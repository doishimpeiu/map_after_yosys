module nngenmod(CLK, RESETN, maxi_awaddr, maxi_awlen, maxi_awsize, maxi_awburst, maxi_awlock, maxi_awcache, maxi_awprot, maxi_awqos, maxi_awuser, maxi_awvalid, maxi_awready, maxi_wdata, maxi_wstrb, maxi_wlast, maxi_wvalid, maxi_wready, maxi_bresp, maxi_bvalid, maxi_bready, maxi_araddr, maxi_arlen, maxi_arsize, maxi_arburst, maxi_arlock, maxi_arcache, maxi_arprot, maxi_arqos, maxi_aruser, maxi_arvalid, maxi_arready, maxi_rdata, maxi_rresp, maxi_rlast, maxi_rvalid, maxi_rready, saxi_awaddr, saxi_awcache, saxi_awprot, saxi_awvalid, saxi_awready, saxi_wdata, saxi_wstrb, saxi_wvalid, saxi_wready, saxi_bresp, saxi_bvalid, saxi_bready, saxi_araddr, saxi_arcache, saxi_arprot, saxi_arvalid, saxi_arready, saxi_rdata, saxi_rresp, saxi_rvalid, saxi_rready);
  input CLK;
  input RESETN;
  input maxi_arready;
  input maxi_awready;
  input [1:0] maxi_bresp;
  input maxi_bvalid;
  input [31:0] maxi_rdata;
  input maxi_rlast;
  input [1:0] maxi_rresp;
  input maxi_rvalid;
  input maxi_wready;
  input [5:0] saxi_araddr;
  input [3:0] saxi_arcache;
  input [2:0] saxi_arprot;
  input saxi_arvalid;
  input [5:0] saxi_awaddr;
  input [3:0] saxi_awcache;
  input [2:0] saxi_awprot;
  input saxi_awvalid;
  input saxi_bready;
  input saxi_rready;
  input [31:0] saxi_wdata;
  input [3:0] saxi_wstrb;
  input saxi_wvalid;
  output [31:0] maxi_araddr;
  output [1:0] maxi_arburst;
  output [3:0] maxi_arcache;
  output [7:0] maxi_arlen;
  output maxi_arlock;
  output [2:0] maxi_arprot;
  output [3:0] maxi_arqos;
  output [2:0] maxi_arsize;
  output [1:0] maxi_aruser;
  output maxi_arvalid;
  output [31:0] maxi_awaddr;
  output [1:0] maxi_awburst;
  output [3:0] maxi_awcache;
  output [7:0] maxi_awlen;
  output maxi_awlock;
  output [2:0] maxi_awprot;
  output [3:0] maxi_awqos;
  output [2:0] maxi_awsize;
  output [1:0] maxi_awuser;
  output maxi_awvalid;
  output maxi_bready;
  output maxi_rready;
  output [31:0] maxi_wdata;
  output maxi_wlast;
  output [3:0] maxi_wstrb;
  output maxi_wvalid;
  output saxi_arready;
  output saxi_awready;
  output [1:0] saxi_bresp;
  output saxi_bvalid;
  output [31:0] saxi_rdata;
  output [1:0] saxi_rresp;
  output saxi_rvalid;
  output saxi_wready;
  wire _00000_;
  wire _00620_;
  wire _01356_;
  wire [31:0] _01468_;
  wire _01646_;
  wire _01657_;
  wire [31:0] _01714_;
  wire [31:0] _01730_;
  wire [31:0] _01732_;
  wire [31:0] _01733_;
  wire _02389_;
  wire _02391_;
  wire _02393_;
  wire _02395_;
  wire _02404_;
  wire _02413_;
  wire _02422_;
  wire _02431_;
  wire _02440_;
  wire _02449_;
  wire _02458_;
  wire _02467_;
  wire _02476_;
  wire _02485_;
  wire _02494_;
  wire _02503_;
  wire _02512_;
  wire _02521_;
  wire _02530_;
  wire _02539_;
  wire _02548_;
  wire _02557_;
  wire _02566_;
  wire _02598_;
  wire _02600_;
  wire _02602_;
  wire _02604_;
  wire _02613_;
  wire _02622_;
  wire _02631_;
  wire _02647_;
  wire _02659_;
  wire [3:0] _02883_;
  wire _03072_;
  wire _03133_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire [31:0] _22041_;
  wire [31:0] _22042_;
  wire [31:0] _22043_;
  wire [31:0] _22044_;
  wire [31:0] _22045_;
  wire [31:0] _22046_;
  wire [31:0] _22047_;
  wire [31:0] _22048_;
  wire [31:0] _22049_;
  wire [31:0] _22050_;
  wire [31:0] _22051_;
  wire [31:0] _22052_;
  wire [31:0] _22053_;
  wire [31:0] _22054_;
  wire [31:0] _22055_;
  wire [31:0] _22056_;
  wire [31:0] _22057_;
  wire [31:0] _22058_;
  wire [31:0] _22059_;
  wire [31:0] _22060_;
  wire [32:0] _22061_;
  wire [32:0] _22062_;
  wire [31:0] _22063_;
  wire [31:0] _22064_;
  wire [32:0] _22065_;
  wire [31:0] _22066_;
  wire [32:0] _22067_;
  wire [31:0] _22068_;
  wire [31:0] _22069_;
  wire [31:0] _22070_;
  wire [31:0] _22071_;
  wire [32:0] _22072_;
  wire [31:0] _22073_;
  wire [31:0] _22074_;
  wire [31:0] _22075_;
  wire [32:0] _22076_;
  wire [31:0] _22077_;
  wire [31:0] _22078_;
  wire [31:0] _22079_;
  wire [31:0] _22080_;
  wire [31:0] _22081_;
  wire [31:0] _22082_;
  wire [31:0] _22083_;
  wire [31:0] _22084_;
  wire [31:0] _22085_;
  wire [31:0] _22086_;
  wire [31:0] _22087_;
  wire [31:0] _22088_;
  wire [31:0] _22089_;
  wire [31:0] _22090_;
  wire [31:0] _22091_;
  wire [31:0] _22092_;
  wire [31:0] _22093_;
  wire [31:0] _22094_;
  wire [31:0] _22095_;
  wire [31:0] _22096_;
  wire [31:0] _22097_;
  wire [31:0] _22098_;
  wire [31:0] _22099_;
  wire [31:0] _22100_;
  wire [31:0] _22101_;
  wire [31:0] _22102_;
  wire [31:0] _22103_;
  wire [31:0] _22104_;
  wire [31:0] _22105_;
  wire [31:0] _22106_;
  wire [31:0] _22107_;
  wire [31:0] _22108_;
  wire [31:0] _22109_;
  wire [31:0] _22110_;
  wire [31:0] _22111_;
  wire [31:0] _22112_;
  wire [31:0] _22113_;
  wire [31:0] _22114_;
  wire [31:0] _22115_;
  wire [31:0] _22116_;
  wire [31:0] _22117_;
  wire [31:0] _22118_;
  wire [31:0] _22119_;
  wire [31:0] _22120_;
  wire [31:0] _22121_;
  wire [31:0] _22122_;
  wire [32:0] _22123_;
  wire [32:0] _22124_;
  wire [31:0] _22125_;
  wire [31:0] _22126_;
  wire [31:0] _22127_;
  wire [31:0] _22128_;
  wire [31:0] _22129_;
  wire [31:0] _22130_;
  wire [31:0] _22131_;
  wire [31:0] _22132_;
  wire [31:0] _22133_;
  wire [31:0] _22134_;
  wire [31:0] _22135_;
  wire [7:0] _22136_;
  wire [7:0] _22137_;
  wire [7:0] _22138_;
  wire [31:0] _22139_;
  wire [31:0] _22140_;
  wire [31:0] _22141_;
  wire [31:0] _22142_;
  wire [31:0] _22143_;
  wire [31:0] _22144_;
  wire [31:0] _22145_;
  wire [31:0] _22146_;
  wire [31:0] _22147_;
  wire [31:0] _22148_;
  wire [31:0] _22149_;
  wire [31:0] _22150_;
  wire [31:0] _22151_;
  wire [31:0] _22152_;
  wire [31:0] _22153_;
  wire [31:0] _22154_;
  wire [31:0] _22155_;
  wire [31:0] _22156_;
  wire [31:0] _22157_;
  wire [31:0] _22158_;
  wire [31:0] _22159_;
  wire [31:0] _22160_;
  wire [31:0] _22161_;
  wire [31:0] _22162_;
  wire [31:0] _22163_;
  wire [31:0] _22164_;
  wire [31:0] _22165_;
  wire [31:0] _22166_;
  wire [31:0] _22167_;
  wire [31:0] _22168_;
  wire [31:0] _22169_;
  wire [31:0] _22170_;
  wire [31:0] _22171_;
  wire [31:0] _22172_;
  wire [31:0] _22173_;
  wire [31:0] _22174_;
  wire [31:0] _22175_;
  wire [31:0] _22176_;
  wire [31:0] _22177_;
  wire [31:0] _22178_;
  wire [31:0] _22179_;
  wire [31:0] _22180_;
  wire [31:0] _22181_;
  wire [31:0] _22182_;
  wire [31:0] _22183_;
  wire [31:0] _22184_;
  wire [31:0] _22185_;
  wire [31:0] _22186_;
  wire [31:0] _22187_;
  wire [31:0] _22188_;
  wire [31:0] _22189_;
  wire [31:0] _22190_;
  wire [31:0] _22191_;
  wire [31:0] _22192_;
  wire [31:0] _22193_;
  wire [31:0] _22194_;
  wire [31:0] _22195_;
  wire [31:0] _22196_;
  wire [31:0] _22197_;
  wire [31:0] _22198_;
  wire [31:0] _22199_;
  wire [31:0] _22200_;
  wire [31:0] _22201_;
  wire [31:0] _22202_;
  wire [31:0] _22203_;
  wire [31:0] _22204_;
  wire [31:0] _22205_;
  wire [31:0] _22206_;
  wire [31:0] _22207_;
  wire [31:0] _22208_;
  wire [31:0] _22209_;
  wire [31:0] _22210_;
  wire [31:0] _22211_;
  wire [31:0] _22212_;
  wire [31:0] _22213_;
  wire [31:0] _22214_;
  wire [31:0] _22215_;
  wire [31:0] _22216_;
  wire [31:0] _22217_;
  wire [31:0] _22218_;
  wire [31:0] _22219_;
  wire [31:0] _22220_;
  wire [31:0] _22221_;
  wire [31:0] _22222_;
  wire [31:0] _22223_;
  wire [31:0] _22224_;
  wire [31:0] _22225_;
  wire [31:0] _22226_;
  wire [31:0] _22227_;
  wire [31:0] _22228_;
  wire [31:0] _22229_;
  wire [31:0] _22230_;
  wire [31:0] _22231_;
  wire [31:0] _22232_;
  wire [31:0] _22233_;
  wire [31:0] _22234_;
  wire [31:0] _22235_;
  wire [31:0] _22236_;
  wire [31:0] _22237_;
  wire [31:0] _22238_;
  wire [31:0] _22239_;
  wire [7:0] _22240_;
  wire [7:0] _22241_;
  wire [7:0] _22242_;
  wire [31:0] _22243_;
  wire [31:0] _22244_;
  wire [31:0] _22245_;
  wire [31:0] _22246_;
  wire [31:0] _22247_;
  wire [31:0] _22248_;
  wire [31:0] _22249_;
  wire [31:0] _22250_;
  wire [31:0] _22251_;
  wire [31:0] _22252_;
  wire [31:0] _22253_;
  wire [31:0] _22254_;
  wire [31:0] _22255_;
  wire [31:0] _22256_;
  wire [31:0] _22257_;
  wire [31:0] _22258_;
  wire [31:0] _22259_;
  wire [31:0] _22260_;
  wire [31:0] _22261_;
  wire [31:0] _22262_;
  wire [31:0] _22263_;
  wire [31:0] _22264_;
  wire [31:0] _22265_;
  wire [31:0] _22266_;
  wire [31:0] _22267_;
  wire [31:0] _22268_;
  wire [31:0] _22269_;
  wire [31:0] _22270_;
  wire [31:0] _22271_;
  wire [31:0] _22272_;
  wire [31:0] _22273_;
  wire [1:0] _22274_;
  wire [31:0] _22275_;
  wire [31:0] _22276_;
  wire [31:0] _22277_;
  wire [31:0] _22278_;
  wire [31:0] _22279_;
  wire [31:0] _22280_;
  wire [31:0] _22281_;
  wire [31:0] _22282_;
  wire [31:0] _22283_;
  wire [31:0] _22284_;
  wire [32:0] _22285_;
  wire [31:0] _22286_;
  wire [31:0] _22287_;
  wire [31:0] _22288_;
  wire [31:0] _22289_;
  wire [31:0] _22290_;
  wire [31:0] _22291_;
  wire [31:0] _22292_;
  wire [31:0] _22293_;
  wire [31:0] _22294_;
  wire [31:0] _22295_;
  wire [31:0] _22296_;
  wire [31:0] _22297_;
  wire [1:0] _22298_;
  wire [31:0] _22299_;
  wire [32:0] _22300_;
  wire [31:0] _22301_;
  wire [31:0] _22302_;
  wire [31:0] _22303_;
  wire [31:0] _22304_;
  wire [31:0] _22305_;
  wire [31:0] _22306_;
  wire [31:0] _22307_;
  wire [31:0] _22308_;
  wire [31:0] _22309_;
  wire [31:0] _22310_;
  wire [31:0] _22311_;
  wire [31:0] _22312_;
  wire [31:0] _22313_;
  wire [31:0] _22314_;
  wire [31:0] _22315_;
  wire [31:0] _22316_;
  wire [31:0] _22317_;
  wire [31:0] _22318_;
  wire [31:0] _22319_;
  wire [31:0] _22320_;
  wire [31:0] _22321_;
  wire [31:0] _22322_;
  wire [31:0] _22323_;
  wire [31:0] _22324_;
  wire [31:0] _22325_;
  wire [31:0] _22326_;
  wire [31:0] _22327_;
  wire [31:0] _22328_;
  wire [31:0] _22329_;
  wire [31:0] _22330_;
  wire [31:0] _22331_;
  wire [31:0] _22332_;
  wire [31:0] _22333_;
  wire [31:0] _22334_;
  wire [31:0] _22335_;
  wire [31:0] _22336_;
  wire [31:0] _22337_;
  wire [31:0] _22338_;
  wire [31:0] _22339_;
  wire [31:0] _22340_;
  wire [31:0] _22341_;
  wire [31:0] _22342_;
  wire [31:0] _22343_;
  wire [31:0] _22344_;
  wire [31:0] _22345_;
  wire [31:0] _22346_;
  wire [31:0] _22347_;
  wire [31:0] _22348_;
  wire [31:0] _22349_;
  wire [31:0] _22350_;
  wire [31:0] _22351_;
  wire [31:0] _22352_;
  wire [31:0] _22353_;
  wire [31:0] _22354_;
  wire [31:0] _22355_;
  wire [31:0] _22356_;
  wire [31:0] _22357_;
  wire [31:0] _22358_;
  wire [31:0] _22359_;
  wire [31:0] _22360_;
  wire [31:0] _22361_;
  wire [31:0] _22362_;
  wire [31:0] _22363_;
  wire [31:0] _22364_;
  wire [31:0] _22365_;
  wire [31:0] _22366_;
  wire [31:0] _22367_;
  wire [31:0] _22368_;
  wire [31:0] _22369_;
  wire [31:0] _22370_;
  wire [31:0] _22371_;
  wire [31:0] _22372_;
  wire [31:0] _22373_;
  wire [31:0] _22374_;
  wire [31:0] _22375_;
  wire [31:0] _22376_;
  wire [31:0] _22377_;
  wire [31:0] _22378_;
  wire [31:0] _22379_;
  wire [31:0] _22380_;
  wire [31:0] _22381_;
  wire [31:0] _22382_;
  wire [31:0] _22383_;
  wire [31:0] _22384_;
  wire [31:0] _22385_;
  wire [31:0] _22386_;
  wire [31:0] _22387_;
  wire [31:0] _22388_;
  wire [31:0] _22389_;
  wire [31:0] _22390_;
  wire [31:0] _22391_;
  wire [31:0] _22392_;
  wire [31:0] _22393_;
  wire [31:0] _22394_;
  wire [31:0] _22395_;
  wire [31:0] _22396_;
  wire [31:0] _22397_;
  wire [31:0] _22398_;
  wire [31:0] _22399_;
  wire [31:0] _22400_;
  wire [31:0] _22401_;
  wire [31:0] _22402_;
  wire [31:0] _22403_;
  wire [31:0] _22404_;
  wire [31:0] _22405_;
  wire [31:0] _22406_;
  wire [31:0] _22407_;
  wire [31:0] _22408_;
  wire [31:0] _22409_;
  wire [31:0] _22410_;
  wire [31:0] _22411_;
  wire [31:0] _22412_;
  wire [31:0] _22413_;
  wire [31:0] _22414_;
  wire [31:0] _22415_;
  wire [31:0] _22416_;
  wire [31:0] _22417_;
  wire [31:0] _22418_;
  wire [31:0] _22419_;
  wire [31:0] _22420_;
  wire [31:0] _22421_;
  wire [31:0] _22422_;
  wire [31:0] _22423_;
  wire [31:0] _22424_;
  wire [31:0] _22425_;
  wire [31:0] _22426_;
  wire [31:0] _22427_;
  wire [31:0] _22428_;
  wire [31:0] _22429_;
  wire [31:0] _22430_;
  wire [31:0] _22431_;
  wire [31:0] _22432_;
  wire [31:0] _22433_;
  wire [31:0] _22434_;
  wire [31:0] _22435_;
  wire [31:0] _22436_;
  wire [31:0] _22437_;
  wire [31:0] _22438_;
  wire [31:0] _22439_;
  wire [31:0] _22440_;
  wire [31:0] _22441_;
  wire [31:0] _22442_;
  wire [31:0] _22443_;
  wire [31:0] _22444_;
  wire [31:0] _22445_;
  wire [31:0] _22446_;
  wire [31:0] _22447_;
  wire [31:0] _22448_;
  wire [31:0] _22449_;
  wire [31:0] _22450_;
  wire [31:0] _22451_;
  wire [31:0] _22452_;
  wire [31:0] _22453_;
  wire [31:0] _22454_;
  wire [31:0] _22455_;
  wire [31:0] _22456_;
  wire [31:0] _22457_;
  wire [31:0] _22458_;
  wire [31:0] _22459_;
  wire [31:0] _22460_;
  wire _22461_;
  wire [31:0] _22462_;
  wire _22463_;
  wire [31:0] _22464_;
  wire [31:0] _22465_;
  wire [31:0] _22466_;
  wire [31:0] _22467_;
  wire [31:0] _22468_;
  wire [31:0] _22469_;
  wire [31:0] _22470_;
  wire _22471_;
  wire [31:0] _22472_;
  wire [31:0] _22473_;
  wire [31:0] _22474_;
  wire [31:0] _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire [31:0] _22500_;
  wire [31:0] _22501_;
  wire [31:0] _22502_;
  wire _22503_;
  wire [31:0] _22504_;
  wire [31:0] _22505_;
  wire [31:0] _22506_;
  wire [31:0] _22507_;
  wire _22508_;
  wire [31:0] _22509_;
  wire [31:0] _22510_;
  wire [31:0] _22511_;
  wire [31:0] _22512_;
  wire [31:0] _22513_;
  wire _22514_;
  wire [31:0] _22515_;
  wire [31:0] _22516_;
  wire [31:0] _22517_;
  wire [31:0] _22518_;
  wire [31:0] _22519_;
  wire _22520_;
  wire [31:0] _22521_;
  wire [31:0] _22522_;
  wire [31:0] _22523_;
  wire [31:0] _22524_;
  wire [31:0] _22525_;
  wire [31:0] _22526_;
  wire [31:0] _22527_;
  wire [31:0] _22528_;
  wire [31:0] _22529_;
  wire [31:0] _22530_;
  wire [31:0] _22531_;
  wire [31:0] _22532_;
  wire [31:0] _22533_;
  wire [31:0] _22534_;
  wire [31:0] _22535_;
  wire [3:0] _22536_;
  wire [31:0] _22537_;
  wire [31:0] _22538_;
  wire [31:0] _22539_;
  wire [31:0] _22540_;
  wire [31:0] _22541_;
  wire [31:0] _22542_;
  wire [31:0] _22543_;
  wire [31:0] _22544_;
  wire [31:0] _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire [31:0] _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire [31:0] _22562_;
  wire [31:0] _22563_;
  wire _22564_;
  wire [31:0] _22565_;
  wire [31:0] _22566_;
  wire _22567_;
  wire [31:0] _22568_;
  wire [31:0] _22569_;
  wire [31:0] _22570_;
  wire [31:0] _22571_;
  wire [31:0] _22572_;
  wire [31:0] _22573_;
  wire [31:0] _22574_;
  wire [31:0] _22575_;
  wire [31:0] _22576_;
  wire [31:0] _22577_;
  wire [31:0] _22578_;
  wire [31:0] _22579_;
  wire [31:0] _22580_;
  wire [31:0] _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire [32:0] _22586_;
  wire [32:0] _22587_;
  wire [32:0] _22588_;
  wire [32:0] _22589_;
  wire [32:0] _22590_;
  wire [32:0] _22591_;
  wire [32:0] _22592_;
  wire [31:0] _22593_;
  wire [31:0] _22594_;
  wire [31:0] _22595_;
  wire [31:0] _22596_;
  wire [31:0] _22597_;
  wire [31:0] _22598_;
  wire [31:0] _22599_;
  wire [31:0] _22600_;
  wire [31:0] _22601_;
  wire [31:0] _22602_;
  wire [31:0] _22603_;
  wire [31:0] _22604_;
  wire [31:0] _22605_;
  wire [31:0] _22606_;
  wire [31:0] _22607_;
  wire [31:0] _22608_;
  wire [31:0] _22609_;
  wire [31:0] _22610_;
  wire [31:0] _22611_;
  wire [31:0] _22612_;
  wire [31:0] _22613_;
  wire [31:0] _22614_;
  wire [31:0] _22615_;
  wire [31:0] _22616_;
  wire [31:0] _22617_;
  wire [31:0] _22618_;
  wire [31:0] _22619_;
  wire [8:0] _22620_;
  wire [31:0] _22621_;
  wire [1:0] _22622_;
  wire [31:0] _22623_;
  wire [31:0] _22624_;
  wire [31:0] _22625_;
  wire [31:0] _22626_;
  wire [31:0] _22627_;
  wire [31:0] _22628_;
  wire [31:0] _22629_;
  wire [31:0] _22630_;
  wire [31:0] _22631_;
  wire [31:0] _22632_;
  wire [31:0] _22633_;
  wire [31:0] _22634_;
  wire [31:0] _22635_;
  wire [31:0] _22636_;
  wire [31:0] _22637_;
  wire [31:0] _22638_;
  wire [31:0] _22639_;
  wire [31:0] _22640_;
  wire [31:0] _22641_;
  wire [31:0] _22642_;
  wire [31:0] _22643_;
  wire [31:0] _22644_;
  wire [31:0] _22645_;
  wire [31:0] _22646_;
  wire [31:0] _22647_;
  wire [31:0] _22648_;
  wire [31:0] _22649_;
  wire [31:0] _22650_;
  wire [31:0] _22651_;
  wire [1:0] _22652_;
  wire [1:0] _22653_;
  wire [31:0] _22654_;
  wire [31:0] _22655_;
  wire [31:0] _22656_;
  wire [31:0] _22657_;
  wire [8:0] _22658_;
  wire [8:0] _22659_;
  wire [8:0] _22660_;
  wire [8:0] _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire [31:0] _22667_;
  wire [31:0] _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire [31:0] _22674_;
  wire [31:0] _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire [31:0] _22681_;
  wire [31:0] _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire [31:0] _22688_;
  wire [31:0] _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire [31:0] _22695_;
  wire [31:0] _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire [31:0] _22702_;
  wire [31:0] _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire [31:0] _22709_;
  wire [31:0] _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire [31:0] _22716_;
  wire [31:0] _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire [31:0] _22727_;
  wire [31:0] _22728_;
  wire [32:0] _22729_;
  wire [32:0] _22730_;
  wire [32:0] _22731_;
  wire [32:0] _22732_;
  wire [32:0] _22733_;
  wire [32:0] _22734_;
  wire [32:0] _22735_;
  wire [31:0] _22736_;
  wire [31:0] _22737_;
  wire [31:0] _22738_;
  wire [31:0] _22739_;
  wire [31:0] _22740_;
  wire [31:0] _22741_;
  wire [31:0] _22742_;
  wire [31:0] _22743_;
  wire [31:0] _22744_;
  wire [31:0] _22745_;
  wire [31:0] _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire [31:0] _22795_;
  wire [31:0] _22796_;
  wire [31:0] _22797_;
  wire _22798_;
  wire [31:0] _22799_;
  wire [31:0] _22800_;
  wire [31:0] _22801_;
  wire [31:0] _22802_;
  wire [31:0] _22803_;
  wire [31:0] _22804_;
  wire [31:0] _22805_;
  wire [31:0] _22806_;
  wire [31:0] _22807_;
  wire [31:0] _22808_;
  wire [31:0] _22809_;
  wire [31:0] _22810_;
  wire [31:0] _22811_;
  wire [31:0] _22812_;
  wire [31:0] _22813_;
  wire [31:0] _22814_;
  wire [31:0] _22815_;
  wire [31:0] _22816_;
  wire [31:0] _22817_;
  wire [31:0] _22818_;
  wire [31:0] _22819_;
  wire [31:0] _22820_;
  wire [1:0] _22821_;
  wire [31:0] _22822_;
  wire [31:0] _22823_;
  wire [31:0] _22824_;
  wire [31:0] _22825_;
  wire [31:0] _22826_;
  wire [31:0] _22827_;
  wire [1:0] _22828_;
  wire [1:0] _22829_;
  wire [31:0] _22830_;
  wire [31:0] _22831_;
  wire [31:0] _22832_;
  wire [31:0] _22833_;
  wire [31:0] _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire [31:0] _22838_;
  wire [31:0] _22839_;
  wire [31:0] _22840_;
  wire [31:0] _22841_;
  wire [31:0] _22842_;
  wire [31:0] _22843_;
  wire [31:0] _22844_;
  wire [31:0] _22845_;
  wire [31:0] _22846_;
  wire [31:0] _22847_;
  wire [31:0] _22848_;
  wire [31:0] _22849_;
  wire [31:0] _22850_;
  wire [31:0] _22851_;
  wire [31:0] _22852_;
  wire [31:0] _22853_;
  wire [31:0] _22854_;
  wire [31:0] _22855_;
  wire [31:0] _22856_;
  wire [31:0] _22857_;
  wire [31:0] _22858_;
  wire [31:0] _22859_;
  wire [31:0] _22860_;
  wire [31:0] _22861_;
  wire [31:0] _22862_;
  wire [31:0] _22863_;
  wire [31:0] _22864_;
  wire [31:0] _22865_;
  wire [31:0] _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire [31:0] _22874_;
  wire _22875_;
  wire [7:0] _22876_;
  wire [31:0] _22877_;
  wire [31:0] _22878_;
  wire [31:0] _22879_;
  wire [31:0] _22880_;
  wire [32:0] _22881_;
  wire [32:0] _22882_;
  wire [32:0] _22883_;
  wire [32:0] _22884_;
  wire [32:0] _22885_;
  wire [32:0] _22886_;
  wire [32:0] _22887_;
  wire [32:0] _22888_;
  wire [32:0] _22889_;
  wire [32:0] _22890_;
  wire [32:0] _22891_;
  wire [32:0] _22892_;
  wire [32:0] _22893_;
  wire [32:0] _22894_;
  wire [32:0] _22895_;
  wire [32:0] _22896_;
  wire [31:0] _22897_;
  wire [31:0] _22898_;
  wire [31:0] _22899_;
  wire [31:0] _22900_;
  wire [32:0] _22901_;
  wire [32:0] _22902_;
  wire [32:0] _22903_;
  wire [32:0] _22904_;
  wire [31:0] _22905_;
  wire [31:0] _22906_;
  wire [31:0] _22907_;
  wire [31:0] _22908_;
  wire [31:0] _22909_;
  wire [31:0] _22910_;
  wire [31:0] _22911_;
  wire [31:0] _22912_;
  wire [31:0] _22913_;
  wire [31:0] _22914_;
  wire [31:0] _22915_;
  wire [31:0] _22916_;
  wire [7:0] _22917_;
  wire [31:0] _22918_;
  wire [31:0] _22919_;
  wire [31:0] _22920_;
  wire [31:0] _22921_;
  wire [32:0] _22922_;
  wire [32:0] _22923_;
  wire [32:0] _22924_;
  wire [32:0] _22925_;
  wire [32:0] _22926_;
  wire [32:0] _22927_;
  wire [32:0] _22928_;
  wire [32:0] _22929_;
  wire [32:0] _22930_;
  wire [32:0] _22931_;
  wire [32:0] _22932_;
  wire [32:0] _22933_;
  wire [32:0] _22934_;
  wire [32:0] _22935_;
  wire [32:0] _22936_;
  wire [32:0] _22937_;
  wire [31:0] _22938_;
  wire [31:0] _22939_;
  wire [31:0] _22940_;
  wire [31:0] _22941_;
  wire [32:0] _22942_;
  wire [32:0] _22943_;
  wire [32:0] _22944_;
  wire [32:0] _22945_;
  wire [31:0] _22946_;
  wire [31:0] _22947_;
  wire [31:0] _22948_;
  wire [31:0] _22949_;
  wire [31:0] _22950_;
  wire [31:0] _22951_;
  wire [31:0] _22952_;
  wire [31:0] _22953_;
  wire [31:0] _22954_;
  wire [31:0] _22955_;
  wire [31:0] _22956_;
  wire [31:0] _22957_;
  wire [3:0] _22958_;
  wire _22959_;
  wire _22960_;
  wire [7:0] _22961_;
  wire [7:0] _22962_;
  wire [7:0] _22963_;
  wire [7:0] _22964_;
  wire [31:0] _22965_;
  wire [31:0] _22966_;
  wire [31:0] _22967_;
  wire [31:0] _22968_;
  wire [32:0] _22969_;
  wire [32:0] _22970_;
  wire [32:0] _22971_;
  wire [32:0] _22972_;
  wire [32:0] _22973_;
  wire [32:0] _22974_;
  wire [32:0] _22975_;
  wire [32:0] _22976_;
  wire [32:0] _22977_;
  wire [32:0] _22978_;
  wire [32:0] _22979_;
  wire [32:0] _22980_;
  wire [32:0] _22981_;
  wire [32:0] _22982_;
  wire [32:0] _22983_;
  wire [32:0] _22984_;
  wire [31:0] _22985_;
  wire [31:0] _22986_;
  wire [31:0] _22987_;
  wire [31:0] _22988_;
  wire [32:0] _22989_;
  wire [32:0] _22990_;
  wire [32:0] _22991_;
  wire [32:0] _22992_;
  wire [31:0] _22993_;
  wire [31:0] _22994_;
  wire [31:0] _22995_;
  wire [31:0] _22996_;
  wire [31:0] _22997_;
  wire [31:0] _22998_;
  wire [31:0] _22999_;
  wire [31:0] _23000_;
  wire [31:0] _23001_;
  wire [31:0] _23002_;
  wire [31:0] _23003_;
  wire [31:0] _23004_;
  wire [31:0] _23005_;
  wire [31:0] _23006_;
  wire [31:0] _23007_;
  wire [31:0] _23008_;
  wire [31:0] _23009_;
  wire [32:0] _23010_;
  wire [32:0] _23011_;
  wire [32:0] _23012_;
  wire [32:0] _23013_;
  wire [32:0] _23014_;
  wire [32:0] _23015_;
  wire [32:0] _23016_;
  wire [32:0] _23017_;
  wire [32:0] _23018_;
  wire [32:0] _23019_;
  wire [32:0] _23020_;
  wire [32:0] _23021_;
  wire [32:0] _23022_;
  wire [32:0] _23023_;
  wire [32:0] _23024_;
  wire [32:0] _23025_;
  wire [31:0] _23026_;
  wire [31:0] _23027_;
  wire [31:0] _23028_;
  wire [31:0] _23029_;
  wire [32:0] _23030_;
  wire [32:0] _23031_;
  wire [32:0] _23032_;
  wire [32:0] _23033_;
  wire [31:0] _23034_;
  wire [31:0] _23035_;
  wire [31:0] _23036_;
  wire [31:0] _23037_;
  wire [31:0] _23038_;
  wire [31:0] _23039_;
  wire [31:0] _23040_;
  wire [31:0] _23041_;
  wire [31:0] _23042_;
  wire [31:0] _23043_;
  wire [31:0] _23044_;
  wire [31:0] _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire [8:0] _23049_;
  wire [7:0] _23050_;
  wire _23051_;
  wire [31:0] _23052_;
  wire [31:0] _23053_;
  wire [7:0] _23054_;
  wire [31:0] _23055_;
  wire [32:0] _23056_;
  wire [32:0] _23057_;
  wire [31:0] _23058_;
  wire [32:0] _23059_;
  wire [31:0] _23060_;
  wire [2:0] _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire [31:0] _23065_;
  wire [7:0] _23066_;
  wire [31:0] _23067_;
  wire [31:0] _23068_;
  wire [2:0] _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire [31:0] _23075_;
  wire [7:0] _23076_;
  wire [31:0] _23077_;
  wire [31:0] _23078_;
  wire [2:0] _23079_;
  wire _23080_;
  wire _23081_;
  wire [3:0] _23082_;
  wire _23083_;
  wire _23084_;
  wire [7:0] _23085_;
  wire _23086_;
  wire [7:0] _23087_;
  wire _23088_;
  wire [7:0] _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire [31:0] _23094_;
  wire [7:0] _23095_;
  wire [31:0] _23096_;
  wire [31:0] _23097_;
  wire [2:0] _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire [31:0] _23104_;
  wire [7:0] _23105_;
  wire [31:0] _23106_;
  wire [31:0] _23107_;
  wire [2:0] _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire [8:0] _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire [31:0] _23122_;
  wire _23123_;
  wire _23124_;
  wire [7:0] _23125_;
  wire [31:0] _23126_;
  wire [31:0] _23127_;
  wire [31:0] _23128_;
  wire [31:0] _23129_;
  wire [32:0] _23130_;
  wire [32:0] _23131_;
  wire [32:0] _23132_;
  wire [32:0] _23133_;
  wire [32:0] _23134_;
  wire [32:0] _23135_;
  wire [32:0] _23136_;
  wire [32:0] _23137_;
  wire [32:0] _23138_;
  wire [32:0] _23139_;
  wire [32:0] _23140_;
  wire [32:0] _23141_;
  wire [32:0] _23142_;
  wire [32:0] _23143_;
  wire [32:0] _23144_;
  wire [32:0] _23145_;
  wire [31:0] _23146_;
  wire [31:0] _23147_;
  wire [31:0] _23148_;
  wire [31:0] _23149_;
  wire [32:0] _23150_;
  wire [32:0] _23151_;
  wire [32:0] _23152_;
  wire [32:0] _23153_;
  wire [31:0] _23154_;
  wire [31:0] _23155_;
  wire [31:0] _23156_;
  wire [31:0] _23157_;
  wire [31:0] _23158_;
  wire [31:0] _23159_;
  wire [31:0] _23160_;
  wire [31:0] _23161_;
  wire [31:0] _23162_;
  wire [31:0] _23163_;
  wire [31:0] _23164_;
  wire [31:0] _23165_;
  wire [3:0] _23166_;
  wire [2:0] _23167_;
  wire [3:0] _23168_;
  wire [31:0] _23169_;
  wire [31:0] _23170_;
  wire [7:0] _23171_;
  wire _23172_;
  wire [31:0] _23173_;
  wire [31:0] _23174_;
  wire [7:0] _23175_;
  wire [31:0] _23176_;
  wire [32:0] _23177_;
  wire [32:0] _23178_;
  wire [31:0] _23179_;
  wire [32:0] _23180_;
  wire [31:0] _23181_;
  wire [2:0] _23182_;
  wire [3:0] _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire [31:0] _23187_;
  wire [7:0] _23188_;
  wire [31:0] _23189_;
  wire [31:0] _23190_;
  wire [2:0] _23191_;
  wire _23192_;
  wire _23193_;
  wire [2:0] _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire [31:0] _23200_;
  wire _23201_;
  wire [7:0] _23202_;
  wire [31:0] _23203_;
  wire [31:0] _23204_;
  wire [31:0] _23205_;
  wire [31:0] _23206_;
  wire [32:0] _23207_;
  wire [32:0] _23208_;
  wire [32:0] _23209_;
  wire [32:0] _23210_;
  wire [32:0] _23211_;
  wire [32:0] _23212_;
  wire [32:0] _23213_;
  wire [32:0] _23214_;
  wire [32:0] _23215_;
  wire [32:0] _23216_;
  wire [32:0] _23217_;
  wire [32:0] _23218_;
  wire [32:0] _23219_;
  wire [32:0] _23220_;
  wire [32:0] _23221_;
  wire [32:0] _23222_;
  wire [31:0] _23223_;
  wire [31:0] _23224_;
  wire [31:0] _23225_;
  wire [31:0] _23226_;
  wire [32:0] _23227_;
  wire [32:0] _23228_;
  wire [32:0] _23229_;
  wire [32:0] _23230_;
  wire [31:0] _23231_;
  wire [31:0] _23232_;
  wire [31:0] _23233_;
  wire [31:0] _23234_;
  wire [31:0] _23235_;
  wire [31:0] _23236_;
  wire [31:0] _23237_;
  wire [31:0] _23238_;
  wire [31:0] _23239_;
  wire [31:0] _23240_;
  wire [31:0] _23241_;
  wire [31:0] _23242_;
  wire [7:0] _23243_;
  wire [31:0] _23244_;
  wire [31:0] _23245_;
  wire [31:0] _23246_;
  wire [31:0] _23247_;
  wire [32:0] _23248_;
  wire [32:0] _23249_;
  wire [32:0] _23250_;
  wire [32:0] _23251_;
  wire [32:0] _23252_;
  wire [32:0] _23253_;
  wire [32:0] _23254_;
  wire [32:0] _23255_;
  wire [32:0] _23256_;
  wire [32:0] _23257_;
  wire [32:0] _23258_;
  wire [32:0] _23259_;
  wire [32:0] _23260_;
  wire [32:0] _23261_;
  wire [32:0] _23262_;
  wire [32:0] _23263_;
  wire [31:0] _23264_;
  wire [31:0] _23265_;
  wire [31:0] _23266_;
  wire [31:0] _23267_;
  wire [32:0] _23268_;
  wire [32:0] _23269_;
  wire [32:0] _23270_;
  wire [32:0] _23271_;
  wire [31:0] _23272_;
  wire [31:0] _23273_;
  wire [31:0] _23274_;
  wire [31:0] _23275_;
  wire [31:0] _23276_;
  wire [31:0] _23277_;
  wire [31:0] _23278_;
  wire [31:0] _23279_;
  wire [31:0] _23280_;
  wire [31:0] _23281_;
  wire [31:0] _23282_;
  wire [31:0] _23283_;
  wire [7:0] _23284_;
  wire [31:0] _23285_;
  wire [31:0] _23286_;
  wire [31:0] _23287_;
  wire [31:0] _23288_;
  wire [32:0] _23289_;
  wire [32:0] _23290_;
  wire [32:0] _23291_;
  wire [32:0] _23292_;
  wire [32:0] _23293_;
  wire [32:0] _23294_;
  wire [32:0] _23295_;
  wire [32:0] _23296_;
  wire [32:0] _23297_;
  wire [32:0] _23298_;
  wire [32:0] _23299_;
  wire [32:0] _23300_;
  wire [32:0] _23301_;
  wire [32:0] _23302_;
  wire [32:0] _23303_;
  wire [32:0] _23304_;
  wire [31:0] _23305_;
  wire [31:0] _23306_;
  wire [31:0] _23307_;
  wire [31:0] _23308_;
  wire [32:0] _23309_;
  wire [32:0] _23310_;
  wire [32:0] _23311_;
  wire [32:0] _23312_;
  wire [31:0] _23313_;
  wire [31:0] _23314_;
  wire [31:0] _23315_;
  wire [31:0] _23316_;
  wire [31:0] _23317_;
  wire [31:0] _23318_;
  wire [31:0] _23319_;
  wire [31:0] _23320_;
  wire [31:0] _23321_;
  wire [31:0] _23322_;
  wire [31:0] _23323_;
  wire [31:0] _23324_;
  wire [7:0] _23325_;
  wire [31:0] _23326_;
  wire [31:0] _23327_;
  wire [31:0] _23328_;
  wire [31:0] _23329_;
  wire [32:0] _23330_;
  wire [32:0] _23331_;
  wire [32:0] _23332_;
  wire [32:0] _23333_;
  wire [32:0] _23334_;
  wire [32:0] _23335_;
  wire [32:0] _23336_;
  wire [32:0] _23337_;
  wire [32:0] _23338_;
  wire [32:0] _23339_;
  wire [32:0] _23340_;
  wire [32:0] _23341_;
  wire [32:0] _23342_;
  wire [32:0] _23343_;
  wire [32:0] _23344_;
  wire [32:0] _23345_;
  wire [31:0] _23346_;
  wire [31:0] _23347_;
  wire [31:0] _23348_;
  wire [31:0] _23349_;
  wire [32:0] _23350_;
  wire [32:0] _23351_;
  wire [32:0] _23352_;
  wire [32:0] _23353_;
  wire [31:0] _23354_;
  wire [31:0] _23355_;
  wire [31:0] _23356_;
  wire [31:0] _23357_;
  wire [31:0] _23358_;
  wire [31:0] _23359_;
  wire [31:0] _23360_;
  wire [31:0] _23361_;
  wire [31:0] _23362_;
  wire [31:0] _23363_;
  wire [31:0] _23364_;
  wire [31:0] _23365_;
  wire [7:0] _23366_;
  wire [31:0] _23367_;
  wire [31:0] _23368_;
  wire [31:0] _23369_;
  wire [31:0] _23370_;
  wire [32:0] _23371_;
  wire [32:0] _23372_;
  wire [32:0] _23373_;
  wire [32:0] _23374_;
  wire [32:0] _23375_;
  wire [32:0] _23376_;
  wire [32:0] _23377_;
  wire [32:0] _23378_;
  wire [32:0] _23379_;
  wire [32:0] _23380_;
  wire [32:0] _23381_;
  wire [32:0] _23382_;
  wire [32:0] _23383_;
  wire [32:0] _23384_;
  wire [32:0] _23385_;
  wire [32:0] _23386_;
  wire [31:0] _23387_;
  wire [31:0] _23388_;
  wire [31:0] _23389_;
  wire [31:0] _23390_;
  wire [32:0] _23391_;
  wire [32:0] _23392_;
  wire [32:0] _23393_;
  wire [32:0] _23394_;
  wire [31:0] _23395_;
  wire [31:0] _23396_;
  wire [31:0] _23397_;
  wire [31:0] _23398_;
  wire [31:0] _23399_;
  wire [31:0] _23400_;
  wire [31:0] _23401_;
  wire [31:0] _23402_;
  wire [31:0] _23403_;
  wire [31:0] _23404_;
  wire [31:0] _23405_;
  wire [31:0] _23406_;
  wire [7:0] _23407_;
  wire [31:0] _23408_;
  wire [31:0] _23409_;
  wire [31:0] _23410_;
  wire [31:0] _23411_;
  wire [32:0] _23412_;
  wire [32:0] _23413_;
  wire [32:0] _23414_;
  wire [32:0] _23415_;
  wire [32:0] _23416_;
  wire [32:0] _23417_;
  wire [32:0] _23418_;
  wire [32:0] _23419_;
  wire [32:0] _23420_;
  wire [32:0] _23421_;
  wire [32:0] _23422_;
  wire [32:0] _23423_;
  wire [32:0] _23424_;
  wire [32:0] _23425_;
  wire [32:0] _23426_;
  wire [32:0] _23427_;
  wire [31:0] _23428_;
  wire [31:0] _23429_;
  wire [31:0] _23430_;
  wire [31:0] _23431_;
  wire [32:0] _23432_;
  wire [32:0] _23433_;
  wire [32:0] _23434_;
  wire [32:0] _23435_;
  wire [31:0] _23436_;
  wire [31:0] _23437_;
  wire [31:0] _23438_;
  wire [31:0] _23439_;
  wire [31:0] _23440_;
  wire [31:0] _23441_;
  wire [31:0] _23442_;
  wire [31:0] _23443_;
  wire [31:0] _23444_;
  wire [31:0] _23445_;
  wire [31:0] _23446_;
  wire [31:0] _23447_;
  wire [7:0] _23448_;
  wire [31:0] _23449_;
  wire [31:0] _23450_;
  wire [31:0] _23451_;
  wire [31:0] _23452_;
  wire [32:0] _23453_;
  wire [32:0] _23454_;
  wire [32:0] _23455_;
  wire [32:0] _23456_;
  wire [32:0] _23457_;
  wire [32:0] _23458_;
  wire [32:0] _23459_;
  wire [32:0] _23460_;
  wire [32:0] _23461_;
  wire [32:0] _23462_;
  wire [32:0] _23463_;
  wire [32:0] _23464_;
  wire [32:0] _23465_;
  wire [32:0] _23466_;
  wire [32:0] _23467_;
  wire [32:0] _23468_;
  wire [31:0] _23469_;
  wire [31:0] _23470_;
  wire [31:0] _23471_;
  wire [31:0] _23472_;
  wire [32:0] _23473_;
  wire [32:0] _23474_;
  wire [32:0] _23475_;
  wire [32:0] _23476_;
  wire [31:0] _23477_;
  wire [31:0] _23478_;
  wire [31:0] _23479_;
  wire [31:0] _23480_;
  wire [31:0] _23481_;
  wire [31:0] _23482_;
  wire [31:0] _23483_;
  wire [31:0] _23484_;
  wire [31:0] _23485_;
  wire [31:0] _23486_;
  wire [31:0] _23487_;
  wire [31:0] _23488_;
  wire [7:0] _23489_;
  wire [31:0] _23490_;
  wire [31:0] _23491_;
  wire [31:0] _23492_;
  wire [31:0] _23493_;
  wire [32:0] _23494_;
  wire [32:0] _23495_;
  wire [32:0] _23496_;
  wire [32:0] _23497_;
  wire [32:0] _23498_;
  wire [32:0] _23499_;
  wire [32:0] _23500_;
  wire [32:0] _23501_;
  wire [32:0] _23502_;
  wire [32:0] _23503_;
  wire [32:0] _23504_;
  wire [32:0] _23505_;
  wire [32:0] _23506_;
  wire [32:0] _23507_;
  wire [32:0] _23508_;
  wire [32:0] _23509_;
  wire [31:0] _23510_;
  wire [31:0] _23511_;
  wire [31:0] _23512_;
  wire [31:0] _23513_;
  wire [32:0] _23514_;
  wire [32:0] _23515_;
  wire [32:0] _23516_;
  wire [32:0] _23517_;
  wire [31:0] _23518_;
  wire [31:0] _23519_;
  wire [31:0] _23520_;
  wire [31:0] _23521_;
  wire [31:0] _23522_;
  wire [31:0] _23523_;
  wire [31:0] _23524_;
  wire [31:0] _23525_;
  wire [31:0] _23526_;
  wire [31:0] _23527_;
  wire [31:0] _23528_;
  wire [31:0] _23529_;
  wire [7:0] _23530_;
  wire [31:0] _23531_;
  wire [31:0] _23532_;
  wire [31:0] _23533_;
  wire [31:0] _23534_;
  wire [32:0] _23535_;
  wire [32:0] _23536_;
  wire [32:0] _23537_;
  wire [32:0] _23538_;
  wire [32:0] _23539_;
  wire [32:0] _23540_;
  wire [32:0] _23541_;
  wire [32:0] _23542_;
  wire [32:0] _23543_;
  wire [32:0] _23544_;
  wire [32:0] _23545_;
  wire [32:0] _23546_;
  wire [32:0] _23547_;
  wire [32:0] _23548_;
  wire [32:0] _23549_;
  wire [32:0] _23550_;
  wire [31:0] _23551_;
  wire [31:0] _23552_;
  wire [31:0] _23553_;
  wire [31:0] _23554_;
  wire [32:0] _23555_;
  wire [32:0] _23556_;
  wire [32:0] _23557_;
  wire [32:0] _23558_;
  wire [31:0] _23559_;
  wire [31:0] _23560_;
  wire [31:0] _23561_;
  wire [31:0] _23562_;
  wire [31:0] _23563_;
  wire [31:0] _23564_;
  wire [31:0] _23565_;
  wire [31:0] _23566_;
  wire [31:0] _23567_;
  wire [31:0] _23568_;
  wire [31:0] _23569_;
  wire [31:0] _23570_;
  wire [7:0] _23571_;
  wire [31:0] _23572_;
  wire [31:0] _23573_;
  wire [31:0] _23574_;
  wire [31:0] _23575_;
  wire [32:0] _23576_;
  wire [32:0] _23577_;
  wire [32:0] _23578_;
  wire [32:0] _23579_;
  wire [32:0] _23580_;
  wire [32:0] _23581_;
  wire [32:0] _23582_;
  wire [32:0] _23583_;
  wire [32:0] _23584_;
  wire [32:0] _23585_;
  wire [32:0] _23586_;
  wire [32:0] _23587_;
  wire [32:0] _23588_;
  wire [32:0] _23589_;
  wire [32:0] _23590_;
  wire [32:0] _23591_;
  wire [31:0] _23592_;
  wire [31:0] _23593_;
  wire [31:0] _23594_;
  wire [31:0] _23595_;
  wire [32:0] _23596_;
  wire [32:0] _23597_;
  wire [32:0] _23598_;
  wire [32:0] _23599_;
  wire [31:0] _23600_;
  wire [31:0] _23601_;
  wire [31:0] _23602_;
  wire [31:0] _23603_;
  wire [31:0] _23604_;
  wire [31:0] _23605_;
  wire [31:0] _23606_;
  wire [31:0] _23607_;
  wire [31:0] _23608_;
  wire [31:0] _23609_;
  wire [31:0] _23610_;
  wire [31:0] _23611_;
  wire [7:0] _23612_;
  wire [31:0] _23613_;
  wire [31:0] _23614_;
  wire [31:0] _23615_;
  wire [31:0] _23616_;
  wire [32:0] _23617_;
  wire [32:0] _23618_;
  wire [32:0] _23619_;
  wire [32:0] _23620_;
  wire [32:0] _23621_;
  wire [32:0] _23622_;
  wire [32:0] _23623_;
  wire [32:0] _23624_;
  wire [32:0] _23625_;
  wire [32:0] _23626_;
  wire [32:0] _23627_;
  wire [32:0] _23628_;
  wire [32:0] _23629_;
  wire [32:0] _23630_;
  wire [32:0] _23631_;
  wire [32:0] _23632_;
  wire [31:0] _23633_;
  wire [31:0] _23634_;
  wire [31:0] _23635_;
  wire [31:0] _23636_;
  wire [32:0] _23637_;
  wire [32:0] _23638_;
  wire [32:0] _23639_;
  wire [32:0] _23640_;
  wire [31:0] _23641_;
  wire [31:0] _23642_;
  wire [31:0] _23643_;
  wire [31:0] _23644_;
  wire [31:0] _23645_;
  wire [31:0] _23646_;
  wire [31:0] _23647_;
  wire [31:0] _23648_;
  wire [31:0] _23649_;
  wire [31:0] _23650_;
  wire [31:0] _23651_;
  wire [31:0] _23652_;
  wire [7:0] _23653_;
  wire [31:0] _23654_;
  wire [31:0] _23655_;
  wire [31:0] _23656_;
  wire [31:0] _23657_;
  wire [32:0] _23658_;
  wire [32:0] _23659_;
  wire [32:0] _23660_;
  wire [32:0] _23661_;
  wire [32:0] _23662_;
  wire [32:0] _23663_;
  wire [32:0] _23664_;
  wire [32:0] _23665_;
  wire [32:0] _23666_;
  wire [32:0] _23667_;
  wire [32:0] _23668_;
  wire [32:0] _23669_;
  wire [32:0] _23670_;
  wire [32:0] _23671_;
  wire [32:0] _23672_;
  wire [32:0] _23673_;
  wire [31:0] _23674_;
  wire [31:0] _23675_;
  wire [31:0] _23676_;
  wire [31:0] _23677_;
  wire [32:0] _23678_;
  wire [32:0] _23679_;
  wire [32:0] _23680_;
  wire [32:0] _23681_;
  wire [31:0] _23682_;
  wire [31:0] _23683_;
  wire [31:0] _23684_;
  wire [31:0] _23685_;
  wire [31:0] _23686_;
  wire [31:0] _23687_;
  wire [31:0] _23688_;
  wire [31:0] _23689_;
  wire [31:0] _23690_;
  wire [31:0] _23691_;
  wire [31:0] _23692_;
  wire [31:0] _23693_;
  wire [7:0] _23694_;
  wire [31:0] _23695_;
  wire [31:0] _23696_;
  wire [31:0] _23697_;
  wire [31:0] _23698_;
  wire [32:0] _23699_;
  wire [32:0] _23700_;
  wire [32:0] _23701_;
  wire [32:0] _23702_;
  wire [32:0] _23703_;
  wire [32:0] _23704_;
  wire [32:0] _23705_;
  wire [32:0] _23706_;
  wire [32:0] _23707_;
  wire [32:0] _23708_;
  wire [32:0] _23709_;
  wire [32:0] _23710_;
  wire [32:0] _23711_;
  wire [32:0] _23712_;
  wire [32:0] _23713_;
  wire [32:0] _23714_;
  wire [31:0] _23715_;
  wire [31:0] _23716_;
  wire [31:0] _23717_;
  wire [31:0] _23718_;
  wire [32:0] _23719_;
  wire [32:0] _23720_;
  wire [32:0] _23721_;
  wire [32:0] _23722_;
  wire [31:0] _23723_;
  wire [31:0] _23724_;
  wire [31:0] _23725_;
  wire [31:0] _23726_;
  wire [31:0] _23727_;
  wire [31:0] _23728_;
  wire [31:0] _23729_;
  wire [31:0] _23730_;
  wire [31:0] _23731_;
  wire [31:0] _23732_;
  wire [31:0] _23733_;
  wire [31:0] _23734_;
  wire [7:0] _23735_;
  wire [31:0] _23736_;
  wire [31:0] _23737_;
  wire [31:0] _23738_;
  wire [31:0] _23739_;
  wire [32:0] _23740_;
  wire [32:0] _23741_;
  wire [32:0] _23742_;
  wire [32:0] _23743_;
  wire [32:0] _23744_;
  wire [32:0] _23745_;
  wire [32:0] _23746_;
  wire [32:0] _23747_;
  wire [32:0] _23748_;
  wire [32:0] _23749_;
  wire [32:0] _23750_;
  wire [32:0] _23751_;
  wire [32:0] _23752_;
  wire [32:0] _23753_;
  wire [32:0] _23754_;
  wire [32:0] _23755_;
  wire [31:0] _23756_;
  wire [31:0] _23757_;
  wire [31:0] _23758_;
  wire [31:0] _23759_;
  wire [32:0] _23760_;
  wire [32:0] _23761_;
  wire [32:0] _23762_;
  wire [32:0] _23763_;
  wire [31:0] _23764_;
  wire [31:0] _23765_;
  wire [31:0] _23766_;
  wire [31:0] _23767_;
  wire [31:0] _23768_;
  wire [31:0] _23769_;
  wire [31:0] _23770_;
  wire [31:0] _23771_;
  wire [31:0] _23772_;
  wire [31:0] _23773_;
  wire [31:0] _23774_;
  wire [31:0] _23775_;
  wire [7:0] _23776_;
  wire [31:0] _23777_;
  wire [31:0] _23778_;
  wire [31:0] _23779_;
  wire [31:0] _23780_;
  wire [32:0] _23781_;
  wire [32:0] _23782_;
  wire [32:0] _23783_;
  wire [32:0] _23784_;
  wire [32:0] _23785_;
  wire [32:0] _23786_;
  wire [32:0] _23787_;
  wire [32:0] _23788_;
  wire [32:0] _23789_;
  wire [32:0] _23790_;
  wire [32:0] _23791_;
  wire [32:0] _23792_;
  wire [32:0] _23793_;
  wire [32:0] _23794_;
  wire [32:0] _23795_;
  wire [32:0] _23796_;
  wire [31:0] _23797_;
  wire [31:0] _23798_;
  wire [31:0] _23799_;
  wire [31:0] _23800_;
  wire [32:0] _23801_;
  wire [32:0] _23802_;
  wire [32:0] _23803_;
  wire [32:0] _23804_;
  wire [31:0] _23805_;
  wire [31:0] _23806_;
  wire [31:0] _23807_;
  wire [31:0] _23808_;
  wire [31:0] _23809_;
  wire [31:0] _23810_;
  wire [31:0] _23811_;
  wire [31:0] _23812_;
  wire [31:0] _23813_;
  wire [31:0] _23814_;
  wire [31:0] _23815_;
  wire [31:0] _23816_;
  wire [7:0] _23817_;
  wire [31:0] _23818_;
  wire [31:0] _23819_;
  wire [31:0] _23820_;
  wire [31:0] _23821_;
  wire [32:0] _23822_;
  wire [32:0] _23823_;
  wire [32:0] _23824_;
  wire [32:0] _23825_;
  wire [32:0] _23826_;
  wire [32:0] _23827_;
  wire [32:0] _23828_;
  wire [32:0] _23829_;
  wire [32:0] _23830_;
  wire [32:0] _23831_;
  wire [32:0] _23832_;
  wire [32:0] _23833_;
  wire [32:0] _23834_;
  wire [32:0] _23835_;
  wire [32:0] _23836_;
  wire [32:0] _23837_;
  wire [31:0] _23838_;
  wire [31:0] _23839_;
  wire [31:0] _23840_;
  wire [31:0] _23841_;
  wire [32:0] _23842_;
  wire [32:0] _23843_;
  wire [32:0] _23844_;
  wire [32:0] _23845_;
  wire [31:0] _23846_;
  wire [31:0] _23847_;
  wire [31:0] _23848_;
  wire [31:0] _23849_;
  wire [31:0] _23850_;
  wire [31:0] _23851_;
  wire [31:0] _23852_;
  wire [31:0] _23853_;
  wire [31:0] _23854_;
  wire [31:0] _23855_;
  wire [31:0] _23856_;
  wire [31:0] _23857_;
  wire [7:0] _23858_;
  wire [31:0] _23859_;
  wire [31:0] _23860_;
  wire [31:0] _23861_;
  wire [31:0] _23862_;
  wire [32:0] _23863_;
  wire [32:0] _23864_;
  wire [32:0] _23865_;
  wire [32:0] _23866_;
  wire [32:0] _23867_;
  wire [32:0] _23868_;
  wire [32:0] _23869_;
  wire [32:0] _23870_;
  wire [32:0] _23871_;
  wire [32:0] _23872_;
  wire [32:0] _23873_;
  wire [32:0] _23874_;
  wire [32:0] _23875_;
  wire [32:0] _23876_;
  wire [32:0] _23877_;
  wire [32:0] _23878_;
  wire [31:0] _23879_;
  wire [31:0] _23880_;
  wire [31:0] _23881_;
  wire [31:0] _23882_;
  wire [32:0] _23883_;
  wire [32:0] _23884_;
  wire [32:0] _23885_;
  wire [32:0] _23886_;
  wire [31:0] _23887_;
  wire [31:0] _23888_;
  wire [31:0] _23889_;
  wire [31:0] _23890_;
  wire [31:0] _23891_;
  wire [31:0] _23892_;
  wire [31:0] _23893_;
  wire [31:0] _23894_;
  wire [31:0] _23895_;
  wire [31:0] _23896_;
  wire [31:0] _23897_;
  wire [31:0] _23898_;
  wire [7:0] _23899_;
  wire [31:0] _23900_;
  wire [31:0] _23901_;
  wire [31:0] _23902_;
  wire [31:0] _23903_;
  wire [32:0] _23904_;
  wire [32:0] _23905_;
  wire [32:0] _23906_;
  wire [32:0] _23907_;
  wire [32:0] _23908_;
  wire [32:0] _23909_;
  wire [32:0] _23910_;
  wire [32:0] _23911_;
  wire [32:0] _23912_;
  wire [32:0] _23913_;
  wire [32:0] _23914_;
  wire [32:0] _23915_;
  wire [32:0] _23916_;
  wire [32:0] _23917_;
  wire [32:0] _23918_;
  wire [32:0] _23919_;
  wire [31:0] _23920_;
  wire [31:0] _23921_;
  wire [31:0] _23922_;
  wire [31:0] _23923_;
  wire [32:0] _23924_;
  wire [32:0] _23925_;
  wire [32:0] _23926_;
  wire [32:0] _23927_;
  wire [31:0] _23928_;
  wire [31:0] _23929_;
  wire [31:0] _23930_;
  wire [31:0] _23931_;
  wire [31:0] _23932_;
  wire [31:0] _23933_;
  wire [31:0] _23934_;
  wire [31:0] _23935_;
  wire [31:0] _23936_;
  wire [31:0] _23937_;
  wire [31:0] _23938_;
  wire [31:0] _23939_;
  wire [3:0] _23940_;
  wire _23941_;
  wire _23942_;
  wire [7:0] _23943_;
  wire [7:0] _23944_;
  wire [7:0] _23945_;
  wire [7:0] _23946_;
  wire [31:0] _23947_;
  wire [31:0] _23948_;
  wire [31:0] _23949_;
  wire [31:0] _23950_;
  wire [32:0] _23951_;
  wire [32:0] _23952_;
  wire [32:0] _23953_;
  wire [32:0] _23954_;
  wire [32:0] _23955_;
  wire [32:0] _23956_;
  wire [32:0] _23957_;
  wire [32:0] _23958_;
  wire [32:0] _23959_;
  wire [32:0] _23960_;
  wire [32:0] _23961_;
  wire [32:0] _23962_;
  wire [32:0] _23963_;
  wire [32:0] _23964_;
  wire [32:0] _23965_;
  wire [32:0] _23966_;
  wire [31:0] _23967_;
  wire [31:0] _23968_;
  wire [31:0] _23969_;
  wire [31:0] _23970_;
  wire [32:0] _23971_;
  wire [32:0] _23972_;
  wire [32:0] _23973_;
  wire [32:0] _23974_;
  wire [31:0] _23975_;
  wire [31:0] _23976_;
  wire [31:0] _23977_;
  wire [31:0] _23978_;
  wire [31:0] _23979_;
  wire [31:0] _23980_;
  wire [31:0] _23981_;
  wire [31:0] _23982_;
  wire [31:0] _23983_;
  wire [31:0] _23984_;
  wire [31:0] _23985_;
  wire [31:0] _23986_;
  wire [31:0] _23987_;
  wire [31:0] _23988_;
  wire [31:0] _23989_;
  wire [31:0] _23990_;
  wire [31:0] _23991_;
  wire [32:0] _23992_;
  wire [32:0] _23993_;
  wire [32:0] _23994_;
  wire [32:0] _23995_;
  wire [32:0] _23996_;
  wire [32:0] _23997_;
  wire [32:0] _23998_;
  wire [32:0] _23999_;
  wire [32:0] _24000_;
  wire [32:0] _24001_;
  wire [32:0] _24002_;
  wire [32:0] _24003_;
  wire [32:0] _24004_;
  wire [32:0] _24005_;
  wire [32:0] _24006_;
  wire [32:0] _24007_;
  wire [31:0] _24008_;
  wire [31:0] _24009_;
  wire [31:0] _24010_;
  wire [31:0] _24011_;
  wire [32:0] _24012_;
  wire [32:0] _24013_;
  wire [32:0] _24014_;
  wire [32:0] _24015_;
  wire [31:0] _24016_;
  wire [31:0] _24017_;
  wire [31:0] _24018_;
  wire [31:0] _24019_;
  wire [31:0] _24020_;
  wire [31:0] _24021_;
  wire [31:0] _24022_;
  wire [31:0] _24023_;
  wire [31:0] _24024_;
  wire [31:0] _24025_;
  wire [31:0] _24026_;
  wire [31:0] _24027_;
  wire [8:0] _24028_;
  wire [1:0] _24029_;
  wire [1:0] _24030_;
  wire [4:0] _24031_;
  wire [7:0] _24032_;
  wire _24033_;
  wire [31:0] _24034_;
  wire [31:0] _24035_;
  wire [7:0] _24036_;
  wire [31:0] _24037_;
  wire [32:0] _24038_;
  wire [32:0] _24039_;
  wire [31:0] _24040_;
  wire [32:0] _24041_;
  wire [31:0] _24042_;
  wire [2:0] _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire [31:0] _24047_;
  wire [7:0] _24048_;
  wire [31:0] _24049_;
  wire [31:0] _24050_;
  wire [2:0] _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire [31:0] _24057_;
  wire [7:0] _24058_;
  wire [31:0] _24059_;
  wire [31:0] _24060_;
  wire [2:0] _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire [31:0] _24067_;
  wire [7:0] _24068_;
  wire [31:0] _24069_;
  wire [31:0] _24070_;
  wire [2:0] _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire [31:0] _24077_;
  wire [7:0] _24078_;
  wire [31:0] _24079_;
  wire [31:0] _24080_;
  wire [2:0] _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire [31:0] _24087_;
  wire [7:0] _24088_;
  wire [31:0] _24089_;
  wire [31:0] _24090_;
  wire [2:0] _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire [31:0] _24097_;
  wire [7:0] _24098_;
  wire [31:0] _24099_;
  wire [31:0] _24100_;
  wire [2:0] _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire [31:0] _24107_;
  wire [7:0] _24108_;
  wire [31:0] _24109_;
  wire [31:0] _24110_;
  wire [2:0] _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire [31:0] _24117_;
  wire [7:0] _24118_;
  wire [31:0] _24119_;
  wire [31:0] _24120_;
  wire [2:0] _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire [31:0] _24127_;
  wire [7:0] _24128_;
  wire [31:0] _24129_;
  wire [31:0] _24130_;
  wire [2:0] _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire [31:0] _24137_;
  wire [7:0] _24138_;
  wire [31:0] _24139_;
  wire [31:0] _24140_;
  wire [2:0] _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire [31:0] _24147_;
  wire [7:0] _24148_;
  wire [31:0] _24149_;
  wire [31:0] _24150_;
  wire [2:0] _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire [31:0] _24157_;
  wire [7:0] _24158_;
  wire [31:0] _24159_;
  wire [31:0] _24160_;
  wire [2:0] _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire [31:0] _24167_;
  wire [7:0] _24168_;
  wire [31:0] _24169_;
  wire [31:0] _24170_;
  wire [2:0] _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire [31:0] _24177_;
  wire [7:0] _24178_;
  wire [31:0] _24179_;
  wire [31:0] _24180_;
  wire [2:0] _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire [31:0] _24187_;
  wire [7:0] _24188_;
  wire [31:0] _24189_;
  wire [31:0] _24190_;
  wire [2:0] _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire [31:0] _24197_;
  wire [7:0] _24198_;
  wire [31:0] _24199_;
  wire [31:0] _24200_;
  wire [2:0] _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire [31:0] _24207_;
  wire [7:0] _24208_;
  wire [31:0] _24209_;
  wire [31:0] _24210_;
  wire [2:0] _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire [31:0] _24217_;
  wire [7:0] _24218_;
  wire [31:0] _24219_;
  wire [31:0] _24220_;
  wire [2:0] _24221_;
  wire _24222_;
  wire _24223_;
  wire [3:0] _24224_;
  wire _24225_;
  wire _24226_;
  wire [7:0] _24227_;
  wire _24228_;
  wire [7:0] _24229_;
  wire _24230_;
  wire [7:0] _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire [31:0] _24236_;
  wire [7:0] _24237_;
  wire [31:0] _24238_;
  wire [31:0] _24239_;
  wire [2:0] _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire [31:0] _24246_;
  wire [7:0] _24247_;
  wire [31:0] _24248_;
  wire [31:0] _24249_;
  wire [2:0] _24250_;
  wire _24251_;
  wire _24252_;
  wire [8:0] _24253_;
  wire [1:0] _24254_;
  wire [1:0] _24255_;
  wire [4:0] _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire [7:0] _24263_;
  wire [7:0] _24264_;
  wire [8:0] _24265_;
  wire [8:0] _24266_;
  wire [31:0] _24267_;
  wire [31:0] _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire [3:0] _24275_;
  wire [7:0] _24276_;
  wire [7:0] _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire [3:0] _24284_;
  wire [7:0] _24285_;
  wire [7:0] _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire [3:0] _24293_;
  wire [7:0] _24294_;
  wire [7:0] _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire [3:0] _24302_;
  wire [7:0] _24303_;
  wire [7:0] _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire [3:0] _24311_;
  wire [7:0] _24312_;
  wire [7:0] _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire [3:0] _24320_;
  wire [7:0] _24321_;
  wire [7:0] _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire [3:0] _24329_;
  wire [7:0] _24330_;
  wire [7:0] _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire [3:0] _24338_;
  wire [7:0] _24339_;
  wire [7:0] _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire [3:0] _24353_;
  wire [3:0] _24354_;
  wire [7:0] _24355_;
  wire [7:0] _24356_;
  wire [7:0] _24357_;
  wire [7:0] _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire [5:0] _24371_;
  wire [5:0] _24372_;
  wire [7:0] _24373_;
  wire [7:0] _24374_;
  wire [31:0] _24375_;
  wire [31:0] _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire [31:0] _24395_;
  wire [31:0] _24396_;
  wire [31:0] _24397_;
  wire [31:0] _24398_;
  wire [31:0] _24399_;
  wire [31:0] _24400_;
  wire [31:0] _24401_;
  wire [31:0] _24402_;
  wire [31:0] _24403_;
  wire _24404_;
  wire _24405_;
  wire [31:0] _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire [31:0] _24423_;
  wire [31:0] _24424_;
  wire [5:0] _24425_;
  wire [5:0] _24426_;
  wire [31:0] _24427_;
  wire [31:0] _24428_;
  wire [32:0] _24429_;
  wire [32:0] _24430_;
  wire [31:0] _24431_;
  wire [31:0] _24432_;
  wire _24433_;
  wire _24434_;
  wire [33:0] _24435_;
  wire [33:0] _24436_;
  wire _24437_;
  wire _24438_;
  wire [31:0] _24439_;
  wire [6:0] _24440_;
  wire [6:0] _24441_;
  wire [6:0] _24442_;
  wire [6:0] _24443_;
  wire [33:0] _24444_;
  wire [33:0] _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire [8:0] _24459_;
  wire [8:0] _24460_;
  wire _24461_;
  wire _24462_;
  wire [7:0] _24463_;
  wire [8:0] _24464_;
  wire [33:0] _24465_;
  wire [33:0] _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire [8:0] _24480_;
  wire [8:0] _24481_;
  wire _24482_;
  wire _24483_;
  wire [7:0] _24484_;
  wire [8:0] _24485_;
  wire [33:0] _24486_;
  wire [33:0] _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire [8:0] _24501_;
  wire [8:0] _24502_;
  wire _24503_;
  wire _24504_;
  wire [7:0] _24505_;
  wire [8:0] _24506_;
  wire _24507_;
  wire _24508_;
  wire [31:0] _24509_;
  wire [33:0] _24510_;
  wire [33:0] _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire [8:0] _24525_;
  wire [8:0] _24526_;
  wire _24527_;
  wire _24528_;
  wire [7:0] _24529_;
  wire [8:0] _24530_;
  wire _24531_;
  wire _24532_;
  wire [7:0] _24533_;
  wire [8:0] _24534_;
  wire [8:0] _24535_;
  wire _24536_;
  wire _24537_;
  wire [7:0] _24538_;
  wire [8:0] _24539_;
  wire [8:0] _24540_;
  wire _24541_;
  wire _24542_;
  wire [7:0] _24543_;
  wire [8:0] _24544_;
  wire [8:0] _24545_;
  wire _24546_;
  wire _24547_;
  wire [7:0] _24548_;
  wire [8:0] _24549_;
  wire [8:0] _24550_;
  wire _24551_;
  wire _24552_;
  wire [7:0] _24553_;
  wire [8:0] _24554_;
  wire [8:0] _24555_;
  wire _24556_;
  wire _24557_;
  wire [7:0] _24558_;
  wire [8:0] _24559_;
  wire [8:0] _24560_;
  wire _24561_;
  wire _24562_;
  wire [7:0] _24563_;
  wire [8:0] _24564_;
  wire [8:0] _24565_;
  wire _24566_;
  wire _24567_;
  wire [7:0] _24568_;
  wire [8:0] _24569_;
  wire [8:0] _24570_;
  wire [1:0] _24571_;
  wire [1:0] _24572_;
  wire [1:0] _24573_;
  wire [8:0] _24574_;
  wire [8:0] _24575_;
  wire [8:0] _24576_;
  wire [8:0] _24577_;
  wire [8:0] _24578_;
  wire [8:0] _24579_;
  wire _24580_;
  wire _24581_;
  wire [33:0] _24582_;
  wire [33:0] _24583_;
  wire [9:0] _24584_;
  wire [9:0] _24585_;
  wire [9:0] _24586_;
  wire _24587_;
  wire _24588_;
  wire [7:0] _24589_;
  wire [8:0] _24590_;
  wire [8:0] _24591_;
  wire [1:0] _24592_;
  wire [1:0] _24593_;
  wire [1:0] _24594_;
  wire [8:0] _24595_;
  wire [8:0] _24596_;
  wire [8:0] _24597_;
  wire [8:0] _24598_;
  wire [8:0] _24599_;
  wire [8:0] _24600_;
  wire _24601_;
  wire _24602_;
  wire [33:0] _24603_;
  wire [33:0] _24604_;
  wire [9:0] _24605_;
  wire [9:0] _24606_;
  wire [9:0] _24607_;
  wire _24608_;
  wire _24609_;
  wire [7:0] _24610_;
  wire [8:0] _24611_;
  wire [8:0] _24612_;
  wire [1:0] _24613_;
  wire [1:0] _24614_;
  wire [1:0] _24615_;
  wire [8:0] _24616_;
  wire [8:0] _24617_;
  wire [8:0] _24618_;
  wire [8:0] _24619_;
  wire [8:0] _24620_;
  wire [8:0] _24621_;
  wire _24622_;
  wire _24623_;
  wire [33:0] _24624_;
  wire [33:0] _24625_;
  wire [9:0] _24626_;
  wire [9:0] _24627_;
  wire [9:0] _24628_;
  wire _24629_;
  wire _24630_;
  wire [7:0] _24631_;
  wire [8:0] _24632_;
  wire [8:0] _24633_;
  wire [1:0] _24634_;
  wire [1:0] _24635_;
  wire [1:0] _24636_;
  wire [8:0] _24637_;
  wire [8:0] _24638_;
  wire [8:0] _24639_;
  wire [8:0] _24640_;
  wire [8:0] _24641_;
  wire [8:0] _24642_;
  wire _24643_;
  wire _24644_;
  wire [33:0] _24645_;
  wire [33:0] _24646_;
  wire [9:0] _24647_;
  wire [9:0] _24648_;
  wire [9:0] _24649_;
  wire _24650_;
  wire _24651_;
  wire [7:0] _24652_;
  wire [8:0] _24653_;
  wire [8:0] _24654_;
  wire _24655_;
  wire _24656_;
  wire [7:0] _24657_;
  wire [8:0] _24658_;
  wire [8:0] _24659_;
  wire _24660_;
  wire _24661_;
  wire [7:0] _24662_;
  wire [8:0] _24663_;
  wire [8:0] _24664_;
  wire _24665_;
  wire _24666_;
  wire [7:0] _24667_;
  wire [8:0] _24668_;
  wire [8:0] _24669_;
  wire _24670_;
  wire _24671_;
  wire [7:0] _24672_;
  wire [8:0] _24673_;
  wire [8:0] _24674_;
  wire _24675_;
  wire _24676_;
  wire [7:0] _24677_;
  wire [8:0] _24678_;
  wire [8:0] _24679_;
  wire _24680_;
  wire _24681_;
  wire [7:0] _24682_;
  wire [8:0] _24683_;
  wire [8:0] _24684_;
  wire _24685_;
  wire _24686_;
  wire [7:0] _24687_;
  wire [8:0] _24688_;
  wire [8:0] _24689_;
  wire _24690_;
  wire _24691_;
  wire [7:0] _24692_;
  wire [8:0] _24693_;
  wire [8:0] _24694_;
  wire [1:0] _24695_;
  wire [1:0] _24696_;
  wire [1:0] _24697_;
  wire [8:0] _24698_;
  wire [8:0] _24699_;
  wire [8:0] _24700_;
  wire [8:0] _24701_;
  wire [8:0] _24702_;
  wire [8:0] _24703_;
  wire _24704_;
  wire _24705_;
  wire [33:0] _24706_;
  wire [33:0] _24707_;
  wire [9:0] _24708_;
  wire [9:0] _24709_;
  wire [9:0] _24710_;
  wire _24711_;
  wire _24712_;
  wire [7:0] _24713_;
  wire [8:0] _24714_;
  wire [8:0] _24715_;
  wire [1:0] _24716_;
  wire [1:0] _24717_;
  wire [1:0] _24718_;
  wire [8:0] _24719_;
  wire [8:0] _24720_;
  wire [8:0] _24721_;
  wire [8:0] _24722_;
  wire [8:0] _24723_;
  wire [8:0] _24724_;
  wire _24725_;
  wire _24726_;
  wire [33:0] _24727_;
  wire [33:0] _24728_;
  wire [9:0] _24729_;
  wire [9:0] _24730_;
  wire [9:0] _24731_;
  wire _24732_;
  wire _24733_;
  wire [7:0] _24734_;
  wire [8:0] _24735_;
  wire [8:0] _24736_;
  wire [1:0] _24737_;
  wire [1:0] _24738_;
  wire [1:0] _24739_;
  wire [8:0] _24740_;
  wire [8:0] _24741_;
  wire [8:0] _24742_;
  wire [8:0] _24743_;
  wire [8:0] _24744_;
  wire [8:0] _24745_;
  wire _24746_;
  wire _24747_;
  wire [33:0] _24748_;
  wire [33:0] _24749_;
  wire [9:0] _24750_;
  wire [9:0] _24751_;
  wire [9:0] _24752_;
  wire _24753_;
  wire _24754_;
  wire [7:0] _24755_;
  wire [8:0] _24756_;
  wire [8:0] _24757_;
  wire [1:0] _24758_;
  wire [1:0] _24759_;
  wire [1:0] _24760_;
  wire [8:0] _24761_;
  wire [8:0] _24762_;
  wire [8:0] _24763_;
  wire [8:0] _24764_;
  wire [8:0] _24765_;
  wire [8:0] _24766_;
  wire _24767_;
  wire _24768_;
  wire [33:0] _24769_;
  wire [33:0] _24770_;
  wire [9:0] _24771_;
  wire [9:0] _24772_;
  wire [9:0] _24773_;
  wire _24774_;
  wire _24775_;
  wire [7:0] _24776_;
  wire [8:0] _24777_;
  wire [8:0] _24778_;
  wire _24779_;
  wire _24780_;
  wire [7:0] _24781_;
  wire [8:0] _24782_;
  wire [8:0] _24783_;
  wire _24784_;
  wire _24785_;
  wire [7:0] _24786_;
  wire [8:0] _24787_;
  wire [8:0] _24788_;
  wire _24789_;
  wire _24790_;
  wire [7:0] _24791_;
  wire [8:0] _24792_;
  wire [8:0] _24793_;
  wire _24794_;
  wire _24795_;
  wire [7:0] _24796_;
  wire [8:0] _24797_;
  wire [8:0] _24798_;
  wire _24799_;
  wire _24800_;
  wire [7:0] _24801_;
  wire [8:0] _24802_;
  wire [8:0] _24803_;
  wire _24804_;
  wire _24805_;
  wire [7:0] _24806_;
  wire [8:0] _24807_;
  wire [8:0] _24808_;
  wire _24809_;
  wire _24810_;
  wire [7:0] _24811_;
  wire [8:0] _24812_;
  wire [8:0] _24813_;
  wire _24814_;
  wire _24815_;
  wire [7:0] _24816_;
  wire [8:0] _24817_;
  wire [8:0] _24818_;
  wire [1:0] _24819_;
  wire [1:0] _24820_;
  wire [1:0] _24821_;
  wire [8:0] _24822_;
  wire [8:0] _24823_;
  wire [8:0] _24824_;
  wire [8:0] _24825_;
  wire [8:0] _24826_;
  wire [8:0] _24827_;
  wire _24828_;
  wire _24829_;
  wire [33:0] _24830_;
  wire [33:0] _24831_;
  wire [9:0] _24832_;
  wire [9:0] _24833_;
  wire [9:0] _24834_;
  wire _24835_;
  wire _24836_;
  wire [7:0] _24837_;
  wire [8:0] _24838_;
  wire [8:0] _24839_;
  wire [1:0] _24840_;
  wire [1:0] _24841_;
  wire [1:0] _24842_;
  wire [8:0] _24843_;
  wire [8:0] _24844_;
  wire [8:0] _24845_;
  wire [8:0] _24846_;
  wire [8:0] _24847_;
  wire [8:0] _24848_;
  wire _24849_;
  wire _24850_;
  wire [33:0] _24851_;
  wire [33:0] _24852_;
  wire [9:0] _24853_;
  wire [9:0] _24854_;
  wire [9:0] _24855_;
  wire _24856_;
  wire _24857_;
  wire [7:0] _24858_;
  wire [8:0] _24859_;
  wire [8:0] _24860_;
  wire [1:0] _24861_;
  wire [1:0] _24862_;
  wire [1:0] _24863_;
  wire [8:0] _24864_;
  wire [8:0] _24865_;
  wire [8:0] _24866_;
  wire [8:0] _24867_;
  wire [8:0] _24868_;
  wire [8:0] _24869_;
  wire _24870_;
  wire _24871_;
  wire [33:0] _24872_;
  wire [33:0] _24873_;
  wire [9:0] _24874_;
  wire [9:0] _24875_;
  wire [9:0] _24876_;
  wire _24877_;
  wire _24878_;
  wire [7:0] _24879_;
  wire [8:0] _24880_;
  wire [8:0] _24881_;
  wire [1:0] _24882_;
  wire [1:0] _24883_;
  wire [1:0] _24884_;
  wire [8:0] _24885_;
  wire [8:0] _24886_;
  wire [8:0] _24887_;
  wire [8:0] _24888_;
  wire [8:0] _24889_;
  wire [8:0] _24890_;
  wire _24891_;
  wire _24892_;
  wire [33:0] _24893_;
  wire [33:0] _24894_;
  wire [9:0] _24895_;
  wire [9:0] _24896_;
  wire [9:0] _24897_;
  wire _24898_;
  wire _24899_;
  wire [7:0] _24900_;
  wire [8:0] _24901_;
  wire [8:0] _24902_;
  wire _24903_;
  wire _24904_;
  wire [7:0] _24905_;
  wire [8:0] _24906_;
  wire [8:0] _24907_;
  wire _24908_;
  wire _24909_;
  wire [7:0] _24910_;
  wire [8:0] _24911_;
  wire [8:0] _24912_;
  wire _24913_;
  wire _24914_;
  wire [7:0] _24915_;
  wire [8:0] _24916_;
  wire [8:0] _24917_;
  wire _24918_;
  wire _24919_;
  wire [7:0] _24920_;
  wire [8:0] _24921_;
  wire [8:0] _24922_;
  wire _24923_;
  wire _24924_;
  wire [7:0] _24925_;
  wire [8:0] _24926_;
  wire [8:0] _24927_;
  wire _24928_;
  wire _24929_;
  wire [7:0] _24930_;
  wire [8:0] _24931_;
  wire [8:0] _24932_;
  wire _24933_;
  wire _24934_;
  wire [7:0] _24935_;
  wire [8:0] _24936_;
  wire [8:0] _24937_;
  wire _24938_;
  wire _24939_;
  wire [7:0] _24940_;
  wire [8:0] _24941_;
  wire [8:0] _24942_;
  wire _24943_;
  wire _24944_;
  wire [7:0] _24945_;
  wire [8:0] _24946_;
  wire [8:0] _24947_;
  wire _24948_;
  wire _24949_;
  wire [7:0] _24950_;
  wire [8:0] _24951_;
  wire [8:0] _24952_;
  wire _24953_;
  wire _24954_;
  wire [7:0] _24955_;
  wire [8:0] _24956_;
  wire [8:0] _24957_;
  wire _24958_;
  wire _24959_;
  wire [7:0] _24960_;
  wire [8:0] _24961_;
  wire [8:0] _24962_;
  wire _24963_;
  wire _24964_;
  wire [7:0] _24965_;
  wire [8:0] _24966_;
  wire [8:0] _24967_;
  wire _24968_;
  wire _24969_;
  wire [7:0] _24970_;
  wire [8:0] _24971_;
  wire [8:0] _24972_;
  wire _24973_;
  wire _24974_;
  wire [7:0] _24975_;
  wire [8:0] _24976_;
  wire [8:0] _24977_;
  wire _24978_;
  wire _24979_;
  wire [7:0] _24980_;
  wire [8:0] _24981_;
  wire [8:0] _24982_;
  wire _24983_;
  wire _24984_;
  wire [7:0] _24985_;
  wire [8:0] _24986_;
  wire [8:0] _24987_;
  wire _24988_;
  wire _24989_;
  wire [7:0] _24990_;
  wire [8:0] _24991_;
  wire [8:0] _24992_;
  wire _24993_;
  wire _24994_;
  wire [7:0] _24995_;
  wire [8:0] _24996_;
  wire [8:0] _24997_;
  wire _24998_;
  wire _24999_;
  wire [7:0] _25000_;
  wire [8:0] _25001_;
  wire [8:0] _25002_;
  wire _25003_;
  wire _25004_;
  wire [7:0] _25005_;
  wire [8:0] _25006_;
  wire [8:0] _25007_;
  wire _25008_;
  wire _25009_;
  wire [7:0] _25010_;
  wire [8:0] _25011_;
  wire [8:0] _25012_;
  wire _25013_;
  wire _25014_;
  wire [7:0] _25015_;
  wire [8:0] _25016_;
  wire [8:0] _25017_;
  wire _25018_;
  wire _25019_;
  wire [7:0] _25020_;
  wire [8:0] _25021_;
  wire [8:0] _25022_;
  wire _25023_;
  wire _25024_;
  wire [7:0] _25025_;
  wire [8:0] _25026_;
  wire [8:0] _25027_;
  wire _25028_;
  wire _25029_;
  wire [7:0] _25030_;
  wire [8:0] _25031_;
  wire [8:0] _25032_;
  wire _25033_;
  wire _25034_;
  wire [7:0] _25035_;
  wire [8:0] _25036_;
  wire [8:0] _25037_;
  wire _25038_;
  wire _25039_;
  wire [7:0] _25040_;
  wire [8:0] _25041_;
  wire [8:0] _25042_;
  wire _25043_;
  wire _25044_;
  wire [33:0] _25045_;
  wire [33:0] _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire [7:0] _25050_;
  wire [7:0] _25051_;
  wire [8:0] _25052_;
  wire [8:0] _25053_;
  wire [8:0] _25054_;
  wire [8:0] _25055_;
  wire [8:0] _25056_;
  wire _25057_;
  wire _25058_;
  wire [33:0] _25059_;
  wire [33:0] _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire [7:0] _25064_;
  wire [7:0] _25065_;
  wire [8:0] _25066_;
  wire [8:0] _25067_;
  wire [8:0] _25068_;
  wire [8:0] _25069_;
  wire [8:0] _25070_;
  wire _25071_;
  wire _25072_;
  wire [33:0] _25073_;
  wire [33:0] _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire [7:0] _25078_;
  wire [7:0] _25079_;
  wire [8:0] _25080_;
  wire [8:0] _25081_;
  wire [8:0] _25082_;
  wire [8:0] _25083_;
  wire [8:0] _25084_;
  wire _25085_;
  wire _25086_;
  wire [33:0] _25087_;
  wire [33:0] _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire [7:0] _25092_;
  wire [7:0] _25093_;
  wire [8:0] _25094_;
  wire [8:0] _25095_;
  wire [8:0] _25096_;
  wire [8:0] _25097_;
  wire [8:0] _25098_;
  wire [33:0] _25099_;
  wire [33:0] _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire [33:0] _25116_;
  wire [33:0] _25117_;
  wire [3:0] _25118_;
  wire [3:0] _25119_;
  wire [3:0] _25120_;
  wire [8:0] _25121_;
  wire [8:0] _25122_;
  wire [8:0] _25123_;
  wire [8:0] _25124_;
  wire [8:0] _25125_;
  wire [8:0] _25126_;
  wire [8:0] _25127_;
  wire [8:0] _25128_;
  wire [8:0] _25129_;
  wire [8:0] _25130_;
  wire [8:0] _25131_;
  wire [8:0] _25132_;
  wire [8:0] _25133_;
  wire [8:0] _25134_;
  wire [8:0] _25135_;
  wire [8:0] _25136_;
  wire [8:0] _25137_;
  wire [8:0] _25138_;
  wire _25139_;
  wire _25140_;
  wire [33:0] _25141_;
  wire [33:0] _25142_;
  wire [9:0] _25143_;
  wire [9:0] _25144_;
  wire [9:0] _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire [7:0] _25149_;
  wire [7:0] _25150_;
  wire [8:0] _25151_;
  wire [8:0] _25152_;
  wire [8:0] _25153_;
  wire [8:0] _25154_;
  wire [8:0] _25155_;
  wire _25156_;
  wire _25157_;
  wire [7:0] _25158_;
  wire [8:0] _25159_;
  wire [8:0] _25160_;
  wire [8:0] _25161_;
  wire [33:0] _25162_;
  wire [33:0] _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire [33:0] _25179_;
  wire [33:0] _25180_;
  wire [3:0] _25181_;
  wire [3:0] _25182_;
  wire [3:0] _25183_;
  wire [8:0] _25184_;
  wire [8:0] _25185_;
  wire [8:0] _25186_;
  wire [8:0] _25187_;
  wire [8:0] _25188_;
  wire [8:0] _25189_;
  wire [8:0] _25190_;
  wire [8:0] _25191_;
  wire [8:0] _25192_;
  wire [8:0] _25193_;
  wire [8:0] _25194_;
  wire [8:0] _25195_;
  wire [8:0] _25196_;
  wire [8:0] _25197_;
  wire [8:0] _25198_;
  wire [8:0] _25199_;
  wire [8:0] _25200_;
  wire [8:0] _25201_;
  wire _25202_;
  wire _25203_;
  wire [33:0] _25204_;
  wire [33:0] _25205_;
  wire [9:0] _25206_;
  wire [9:0] _25207_;
  wire [9:0] _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire [7:0] _25212_;
  wire [7:0] _25213_;
  wire [8:0] _25214_;
  wire [8:0] _25215_;
  wire [8:0] _25216_;
  wire [8:0] _25217_;
  wire [8:0] _25218_;
  wire _25219_;
  wire _25220_;
  wire [7:0] _25221_;
  wire [8:0] _25222_;
  wire [8:0] _25223_;
  wire [8:0] _25224_;
  wire [33:0] _25225_;
  wire [33:0] _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire [33:0] _25242_;
  wire [33:0] _25243_;
  wire [3:0] _25244_;
  wire [3:0] _25245_;
  wire [3:0] _25246_;
  wire [8:0] _25247_;
  wire [8:0] _25248_;
  wire [8:0] _25249_;
  wire [8:0] _25250_;
  wire [8:0] _25251_;
  wire [8:0] _25252_;
  wire [8:0] _25253_;
  wire [8:0] _25254_;
  wire [8:0] _25255_;
  wire [8:0] _25256_;
  wire [8:0] _25257_;
  wire [8:0] _25258_;
  wire [8:0] _25259_;
  wire [8:0] _25260_;
  wire [8:0] _25261_;
  wire [8:0] _25262_;
  wire [8:0] _25263_;
  wire [8:0] _25264_;
  wire _25265_;
  wire _25266_;
  wire [33:0] _25267_;
  wire [33:0] _25268_;
  wire [9:0] _25269_;
  wire [9:0] _25270_;
  wire [9:0] _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire [7:0] _25275_;
  wire [7:0] _25276_;
  wire [8:0] _25277_;
  wire [8:0] _25278_;
  wire [8:0] _25279_;
  wire [8:0] _25280_;
  wire [8:0] _25281_;
  wire _25282_;
  wire _25283_;
  wire [7:0] _25284_;
  wire [8:0] _25285_;
  wire [8:0] _25286_;
  wire [8:0] _25287_;
  wire _25288_;
  wire _25289_;
  wire [31:0] _25290_;
  wire [33:0] _25291_;
  wire [33:0] _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire [33:0] _25308_;
  wire [33:0] _25309_;
  wire [3:0] _25310_;
  wire [3:0] _25311_;
  wire [3:0] _25312_;
  wire [8:0] _25313_;
  wire [8:0] _25314_;
  wire [8:0] _25315_;
  wire [8:0] _25316_;
  wire [8:0] _25317_;
  wire [8:0] _25318_;
  wire [8:0] _25319_;
  wire [8:0] _25320_;
  wire [8:0] _25321_;
  wire [8:0] _25322_;
  wire [8:0] _25323_;
  wire [8:0] _25324_;
  wire [8:0] _25325_;
  wire [8:0] _25326_;
  wire [8:0] _25327_;
  wire [8:0] _25328_;
  wire [8:0] _25329_;
  wire [8:0] _25330_;
  wire _25331_;
  wire _25332_;
  wire [33:0] _25333_;
  wire [33:0] _25334_;
  wire [9:0] _25335_;
  wire [9:0] _25336_;
  wire [9:0] _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire [7:0] _25341_;
  wire [7:0] _25342_;
  wire [8:0] _25343_;
  wire [8:0] _25344_;
  wire [8:0] _25345_;
  wire [8:0] _25346_;
  wire [8:0] _25347_;
  wire _25348_;
  wire _25349_;
  wire [7:0] _25350_;
  wire [8:0] _25351_;
  wire [8:0] _25352_;
  wire [8:0] _25353_;
  wire [33:0] _25354_;
  wire [33:0] _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire [33:0] _25371_;
  wire [33:0] _25372_;
  wire _25373_;
  wire _25374_;
  wire [7:0] _25375_;
  wire [8:0] _25376_;
  wire [8:0] _25377_;
  wire [8:0] _25378_;
  wire [8:0] _25379_;
  wire _25380_;
  wire _25381_;
  wire [7:0] _25382_;
  wire [8:0] _25383_;
  wire [8:0] _25384_;
  wire [8:0] _25385_;
  wire [33:0] _25386_;
  wire [33:0] _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire [33:0] _25403_;
  wire [33:0] _25404_;
  wire _25405_;
  wire _25406_;
  wire [7:0] _25407_;
  wire [8:0] _25408_;
  wire [8:0] _25409_;
  wire [8:0] _25410_;
  wire [8:0] _25411_;
  wire _25412_;
  wire _25413_;
  wire [7:0] _25414_;
  wire [8:0] _25415_;
  wire [8:0] _25416_;
  wire [8:0] _25417_;
  wire [33:0] _25418_;
  wire [33:0] _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire [33:0] _25435_;
  wire [33:0] _25436_;
  wire _25437_;
  wire _25438_;
  wire [7:0] _25439_;
  wire [8:0] _25440_;
  wire [8:0] _25441_;
  wire [8:0] _25442_;
  wire [8:0] _25443_;
  wire _25444_;
  wire _25445_;
  wire [7:0] _25446_;
  wire [8:0] _25447_;
  wire [8:0] _25448_;
  wire [8:0] _25449_;
  wire _25450_;
  wire _25451_;
  wire [31:0] _25452_;
  wire [33:0] _25453_;
  wire [33:0] _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire [33:0] _25470_;
  wire [33:0] _25471_;
  wire _25472_;
  wire _25473_;
  wire [7:0] _25474_;
  wire [8:0] _25475_;
  wire [8:0] _25476_;
  wire [8:0] _25477_;
  wire [8:0] _25478_;
  wire _25479_;
  wire _25480_;
  wire [7:0] _25481_;
  wire [8:0] _25482_;
  wire [8:0] _25483_;
  wire [8:0] _25484_;
  wire _25485_;
  wire _25486_;
  wire [33:0] _25487_;
  wire [33:0] _25488_;
  wire _25489_;
  wire _25490_;
  wire [7:0] _25491_;
  wire [9:0] _25492_;
  wire [9:0] _25493_;
  wire [9:0] _25494_;
  wire _25495_;
  wire _25496_;
  wire [33:0] _25497_;
  wire [33:0] _25498_;
  wire _25499_;
  wire _25500_;
  wire [7:0] _25501_;
  wire [9:0] _25502_;
  wire [9:0] _25503_;
  wire [9:0] _25504_;
  wire _25505_;
  wire _25506_;
  wire [33:0] _25507_;
  wire [33:0] _25508_;
  wire _25509_;
  wire _25510_;
  wire [7:0] _25511_;
  wire [9:0] _25512_;
  wire [9:0] _25513_;
  wire [9:0] _25514_;
  wire _25515_;
  wire _25516_;
  wire [33:0] _25517_;
  wire [33:0] _25518_;
  wire _25519_;
  wire _25520_;
  wire [7:0] _25521_;
  wire [9:0] _25522_;
  wire [9:0] _25523_;
  wire [9:0] _25524_;
  wire [3:0] _25525_;
  wire [3:0] _25526_;
  wire [31:0] _25527_;
  wire [31:0] _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire [5:0] _25532_;
  wire [5:0] _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire [31:0] _25551_;
  wire [31:0] _25552_;
  wire [31:0] _25553_;
  wire [31:0] _25554_;
  wire [31:0] _25555_;
  wire [31:0] _25556_;
  wire [31:0] _25557_;
  wire [31:0] _25558_;
  wire [31:0] _25559_;
  wire [31:0] _25560_;
  wire [31:0] _25561_;
  wire [31:0] _25562_;
  wire [31:0] _25563_;
  wire [31:0] _25564_;
  wire [31:0] _25565_;
  wire [31:0] _25566_;
  wire [31:0] _25567_;
  wire [31:0] _25568_;
  wire [31:0] _25569_;
  wire [31:0] _25570_;
  wire [31:0] _25571_;
  wire [31:0] _25572_;
  wire [31:0] _25573_;
  wire [31:0] _25574_;
  wire [31:0] _25575_;
  wire [31:0] _25576_;
  wire [31:0] _25577_;
  wire [31:0] _25578_;
  wire [31:0] _25579_;
  wire [31:0] _25580_;
  wire [31:0] _25581_;
  wire [31:0] _25582_;
  wire [31:0] _25583_;
  wire [31:0] _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire [31:0] _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire [31:0] _25593_;
  wire _25594_;
  wire _25595_;
  wire [7:0] _25596_;
  wire _25597_;
  wire _25598_;
  wire [7:0] _25599_;
  wire _25600_;
  wire _25601_;
  wire [7:0] _25602_;
  wire _25603_;
  wire _25604_;
  wire [7:0] _25605_;
  wire _25606_;
  wire _25607_;
  wire [7:0] _25608_;
  wire _25609_;
  wire _25610_;
  wire [7:0] _25611_;
  wire _25612_;
  wire _25613_;
  wire [7:0] _25614_;
  wire _25615_;
  wire _25616_;
  wire [7:0] _25617_;
  wire _25618_;
  wire _25619_;
  wire [7:0] _25620_;
  wire _25621_;
  wire _25622_;
  wire [7:0] _25623_;
  wire _25624_;
  wire _25625_;
  wire [7:0] _25626_;
  wire _25627_;
  wire _25628_;
  wire [7:0] _25629_;
  wire _25630_;
  wire _25631_;
  wire [7:0] _25632_;
  wire _25633_;
  wire _25634_;
  wire [7:0] _25635_;
  wire _25636_;
  wire _25637_;
  wire [7:0] _25638_;
  wire _25639_;
  wire _25640_;
  wire [7:0] _25641_;
  wire _25642_;
  wire _25643_;
  wire [7:0] _25644_;
  wire _25645_;
  wire _25646_;
  wire [7:0] _25647_;
  wire _25648_;
  wire _25649_;
  wire [7:0] _25650_;
  wire _25651_;
  wire _25652_;
  wire [7:0] _25653_;
  wire _25654_;
  wire _25655_;
  wire [7:0] _25656_;
  wire _25657_;
  wire _25658_;
  wire [7:0] _25659_;
  wire _25660_;
  wire _25661_;
  wire [7:0] _25662_;
  wire _25663_;
  wire _25664_;
  wire [7:0] _25665_;
  wire _25666_;
  wire _25667_;
  wire [7:0] _25668_;
  wire _25669_;
  wire _25670_;
  wire [7:0] _25671_;
  wire _25672_;
  wire _25673_;
  wire [7:0] _25674_;
  wire _25675_;
  wire _25676_;
  wire [7:0] _25677_;
  wire _25678_;
  wire _25679_;
  wire [7:0] _25680_;
  wire _25681_;
  wire _25682_;
  wire [7:0] _25683_;
  wire _25684_;
  wire _25685_;
  wire [7:0] _25686_;
  wire _25687_;
  wire _25688_;
  wire [7:0] _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire [31:0] _25693_;
  wire [32:0] _25694_;
  wire [31:0] _25695_;
  wire [31:0] _25696_;
  wire [7:0] _25697_;
  wire _25698_;
  wire [31:0] _25699_;
  wire [32:0] _25700_;
  wire [31:0] _25701_;
  wire [31:0] _25702_;
  wire [7:0] _25703_;
  wire _25704_;
  wire [31:0] _25705_;
  wire [32:0] _25706_;
  wire [31:0] _25707_;
  wire [31:0] _25708_;
  wire [7:0] _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire [31:0] _25714_;
  wire [32:0] _25715_;
  wire [31:0] _25716_;
  wire [31:0] _25717_;
  wire [7:0] _25718_;
  wire _25719_;
  wire [31:0] _25720_;
  wire [31:0] _25721_;
  wire [32:0] _25722_;
  wire [32:0] _25723_;
  wire [31:0] _25724_;
  wire [31:0] _25725_;
  wire [31:0] _25726_;
  wire [31:0] _25727_;
  wire [7:0] _25728_;
  wire [7:0] _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire [8:0] _25735_;
  wire [8:0] _25736_;
  wire [8:0] _25737_;
  wire [8:0] _25738_;
  wire [31:0] _25739_;
  wire [32:0] _25740_;
  wire [31:0] _25741_;
  wire [31:0] _25742_;
  wire [7:0] _25743_;
  wire _25744_;
  wire [31:0] _25745_;
  wire [32:0] _25746_;
  wire [31:0] _25747_;
  wire [31:0] _25748_;
  wire [7:0] _25749_;
  wire _25750_;
  wire [31:0] _25751_;
  wire [32:0] _25752_;
  wire [31:0] _25753_;
  wire [31:0] _25754_;
  wire [7:0] _25755_;
  wire _25756_;
  wire [31:0] _25757_;
  wire [32:0] _25758_;
  wire [31:0] _25759_;
  wire [31:0] _25760_;
  wire [7:0] _25761_;
  wire _25762_;
  wire [31:0] _25763_;
  wire [32:0] _25764_;
  wire [31:0] _25765_;
  wire [31:0] _25766_;
  wire [7:0] _25767_;
  wire _25768_;
  wire [31:0] _25769_;
  wire [31:0] _25770_;
  wire [32:0] _25771_;
  wire [32:0] _25772_;
  wire [31:0] _25773_;
  wire [31:0] _25774_;
  wire [31:0] _25775_;
  wire [31:0] _25776_;
  wire [7:0] _25777_;
  wire [7:0] _25778_;
  wire _25779_;
  wire _25780_;
  wire [8:0] _25781_;
  wire [8:0] _25782_;
  wire [31:0] _25783_;
  wire [31:0] _25784_;
  wire [32:0] _25785_;
  wire [32:0] _25786_;
  wire [31:0] _25787_;
  wire [31:0] _25788_;
  wire [31:0] _25789_;
  wire [31:0] _25790_;
  wire [7:0] _25791_;
  wire [7:0] _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire [31:0] _25799_;
  wire [31:0] _25800_;
  wire [31:0] _25801_;
  wire [32:0] _25802_;
  wire [32:0] _25803_;
  wire [32:0] _25804_;
  wire [31:0] _25805_;
  wire [31:0] _25806_;
  wire [31:0] _25807_;
  wire [31:0] _25808_;
  wire [31:0] _25809_;
  wire [31:0] _25810_;
  wire [7:0] _25811_;
  wire [7:0] _25812_;
  wire [7:0] _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire [31:0] _25827_;
  wire [31:0] _25828_;
  wire [31:0] _25829_;
  wire [31:0] _25830_;
  wire [31:0] _25831_;
  wire [31:0] _25832_;
  wire [31:0] _25833_;
  wire [31:0] _25834_;
  wire [31:0] _25835_;
  wire [32:0] _25836_;
  wire [32:0] _25837_;
  wire [32:0] _25838_;
  wire [32:0] _25839_;
  wire [32:0] _25840_;
  wire [32:0] _25841_;
  wire [32:0] _25842_;
  wire [32:0] _25843_;
  wire [32:0] _25844_;
  wire [31:0] _25845_;
  wire [31:0] _25846_;
  wire [31:0] _25847_;
  wire [31:0] _25848_;
  wire [31:0] _25849_;
  wire [31:0] _25850_;
  wire [31:0] _25851_;
  wire [31:0] _25852_;
  wire [31:0] _25853_;
  wire [31:0] _25854_;
  wire [31:0] _25855_;
  wire [31:0] _25856_;
  wire [31:0] _25857_;
  wire [31:0] _25858_;
  wire [31:0] _25859_;
  wire [31:0] _25860_;
  wire [31:0] _25861_;
  wire [31:0] _25862_;
  wire [7:0] _25863_;
  wire [7:0] _25864_;
  wire [7:0] _25865_;
  wire [7:0] _25866_;
  wire [7:0] _25867_;
  wire [7:0] _25868_;
  wire [7:0] _25869_;
  wire [7:0] _25870_;
  wire [7:0] _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire [7:0] _25884_;
  wire [31:0] _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire [3:0] _25899_;
  wire [3:0] _25900_;
  wire [3:0] _25901_;
  wire [31:0] _25902_;
  wire [31:0] _25903_;
  wire [31:0] _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire [7:0] _25909_;
  wire [31:0] _25910_;
  wire [1:0] _25911_;
  wire [65:0] _25912_;
  wire [17:0] _25913_;
  wire [17:0] _25914_;
  wire [17:0] _25915_;
  wire [17:0] _25916_;
  wire [17:0] _25917_;
  wire [17:0] _25918_;
  wire [17:0] _25919_;
  wire [17:0] _25920_;
  wire [17:0] _25921_;
  wire [32:0] _25922_;
  wire [32:0] _25923_;
  wire [31:0] _25924_;
  wire [39:0] _25925_;
  wire [15:0] _25926_;
  wire [15:0] _25927_;
  wire [15:0] _25928_;
  wire [15:0] _25929_;
  wire [15:0] _25930_;
  wire [15:0] _25931_;
  wire [15:0] _25932_;
  wire [15:0] _25933_;
  wire [15:0] _25934_;
  wire [32:0] _25935_;
  wire [31:0] _25936_;
  wire [32:0] _25937_;
  wire [31:0] _25938_;
  wire [31:0] _25939_;
  wire [33:0] _25940_;
  wire [33:0] _25941_;
  wire [33:0] _25942_;
  wire [33:0] _25943_;
  wire [33:0] _25944_;
  wire [33:0] _25945_;
  wire [33:0] _25946_;
  wire [33:0] _25947_;
  wire [33:0] _25948_;
  wire [33:0] _25949_;
  wire [33:0] _25950_;
  wire [33:0] _25951_;
  wire [33:0] _25952_;
  wire [31:0] _25953_;
  wire [31:0] _25954_;
  wire [33:0] _25955_;
  wire [33:0] _25956_;
  wire [33:0] _25957_;
  wire [31:0] _25958_;
  wire [33:0] _25959_;
  wire [33:0] _25960_;
  wire [33:0] _25961_;
  wire [31:0] _25962_;
  wire [33:0] _25963_;
  wire [33:0] _25964_;
  wire [33:0] _25965_;
  wire [31:0] _25966_;
  wire [33:0] _25967_;
  wire [33:0] _25968_;
  wire [33:0] _25969_;
  wire [33:0] _25970_;
  wire [33:0] _25971_;
  wire [33:0] _25972_;
  wire [33:0] _25973_;
  wire [31:0] _25974_;
  wire [31:0] _25975_;
  wire [33:0] _25976_;
  wire [31:0] _25977_;
  wire [33:0] _25978_;
  wire [31:0] _25979_;
  wire [33:0] _25980_;
  wire [31:0] _25981_;
  wire [33:0] _25982_;
  wire [31:0] _25983_;
  wire [31:0] _25984_;
  wire [33:0] _25985_;
  wire [31:0] _25986_;
  wire [33:0] _25987_;
  wire [31:0] _25988_;
  wire [33:0] _25989_;
  wire [31:0] _25990_;
  wire [33:0] _25991_;
  wire [31:0] _25992_;
  wire [31:0] _25993_;
  wire [33:0] _25994_;
  wire [31:0] _25995_;
  wire [33:0] _25996_;
  wire [31:0] _25997_;
  wire [33:0] _25998_;
  wire [31:0] _25999_;
  wire [33:0] _26000_;
  wire [33:0] _26001_;
  wire [33:0] _26002_;
  wire [33:0] _26003_;
  wire [33:0] _26004_;
  wire [33:0] _26005_;
  wire [5:0] _26006_;
  wire [3:0] _26007_;
  wire [3:0] _26008_;
  wire [3:0] _26009_;
  wire [3:0] _26010_;
  wire [3:0] _26011_;
  wire [3:0] _26012_;
  wire [3:0] _26013_;
  wire [3:0] _26014_;
  wire [3:0] _26015_;
  wire [32:0] _26016_;
  wire [32:0] _26017_;
  wire [32:0] _26018_;
  wire [32:0] _26019_;
  wire [32:0] _26020_;
  wire [32:0] _26021_;
  wire [32:0] _26022_;
  wire [32:0] _26023_;
  wire [32:0] _26024_;
  wire [32:0] _26025_;
  wire [32:0] _26026_;
  wire [32:0] _26027_;
  wire [32:0] _26028_;
  wire [32:0] _26029_;
  wire [32:0] _26030_;
  wire [32:0] _26031_;
  wire [32:0] _26032_;
  wire [32:0] _26033_;
  wire [32:0] _26034_;
  wire [32:0] _26035_;
  wire [32:0] _26036_;
  wire [32:0] _26037_;
  wire [32:0] _26038_;
  wire [32:0] _26039_;
  wire [32:0] _26040_;
  wire [32:0] _26041_;
  wire [32:0] _26042_;
  wire [32:0] _26043_;
  wire [32:0] _26044_;
  wire [32:0] _26045_;
  wire [32:0] _26046_;
  wire [32:0] _26047_;
  wire [32:0] _26048_;
  wire [32:0] _26049_;
  wire [32:0] _26050_;
  wire [32:0] _26051_;
  wire [32:0] _26052_;
  wire [32:0] _26053_;
  wire [32:0] _26054_;
  wire [32:0] _26055_;
  wire [32:0] _26056_;
  wire [32:0] _26057_;
  wire [32:0] _26058_;
  wire [32:0] _26059_;
  wire [32:0] _26060_;
  wire [32:0] _26061_;
  wire [32:0] _26062_;
  wire [32:0] _26063_;
  wire [32:0] _26064_;
  wire [32:0] _26065_;
  wire [32:0] _26066_;
  wire [32:0] _26067_;
  wire [32:0] _26068_;
  wire [32:0] _26069_;
  wire [32:0] _26070_;
  wire [32:0] _26071_;
  wire [32:0] _26072_;
  wire [32:0] _26073_;
  wire [32:0] _26074_;
  wire [32:0] _26075_;
  wire [32:0] _26076_;
  wire [32:0] _26077_;
  wire [32:0] _26078_;
  wire [32:0] _26079_;
  wire [32:0] _26080_;
  wire [32:0] _26081_;
  wire [32:0] _26082_;
  wire [32:0] _26083_;
  wire [32:0] _26084_;
  wire [32:0] _26085_;
  wire [32:0] _26086_;
  wire [32:0] _26087_;
  wire [32:0] _26088_;
  wire [32:0] _26089_;
  wire [32:0] _26090_;
  wire [32:0] _26091_;
  wire [32:0] _26092_;
  wire [32:0] _26093_;
  wire [32:0] _26094_;
  wire [32:0] _26095_;
  wire [32:0] _26096_;
  wire [32:0] _26097_;
  wire [32:0] _26098_;
  wire [32:0] _26099_;
  wire [32:0] _26100_;
  wire [32:0] _26101_;
  wire [32:0] _26102_;
  wire [32:0] _26103_;
  wire [32:0] _26104_;
  wire [32:0] _26105_;
  wire [32:0] _26106_;
  wire [32:0] _26107_;
  wire [32:0] _26108_;
  wire [32:0] _26109_;
  wire [32:0] _26110_;
  wire [32:0] _26111_;
  wire [32:0] _26112_;
  wire [32:0] _26113_;
  wire [32:0] _26114_;
  wire [32:0] _26115_;
  wire [32:0] _26116_;
  wire [32:0] _26117_;
  wire [32:0] _26118_;
  wire [32:0] _26119_;
  wire [32:0] _26120_;
  wire [32:0] _26121_;
  wire [32:0] _26122_;
  wire [32:0] _26123_;
  wire [32:0] _26124_;
  wire [32:0] _26125_;
  wire [32:0] _26126_;
  wire [32:0] _26127_;
  wire [32:0] _26128_;
  wire [32:0] _26129_;
  wire [32:0] _26130_;
  wire [32:0] _26131_;
  wire [32:0] _26132_;
  wire [32:0] _26133_;
  wire [32:0] _26134_;
  wire [32:0] _26135_;
  wire [32:0] _26136_;
  wire [32:0] _26137_;
  wire [32:0] _26138_;
  wire [32:0] _26139_;
  wire [32:0] _26140_;
  wire [32:0] _26141_;
  wire [32:0] _26142_;
  wire [32:0] _26143_;
  wire [32:0] _26144_;
  wire [32:0] _26145_;
  wire [32:0] _26146_;
  wire [32:0] _26147_;
  wire [32:0] _26148_;
  wire [32:0] _26149_;
  wire [32:0] _26150_;
  wire [32:0] _26151_;
  wire [32:0] _26152_;
  wire [32:0] _26153_;
  wire [32:0] _26154_;
  wire [32:0] _26155_;
  wire [32:0] _26156_;
  wire [32:0] _26157_;
  wire [32:0] _26158_;
  wire [32:0] _26159_;
  wire [32:0] _26160_;
  wire [32:0] _26161_;
  wire [32:0] _26162_;
  wire [32:0] _26163_;
  wire [32:0] _26164_;
  wire [32:0] _26165_;
  wire [32:0] _26166_;
  wire [32:0] _26167_;
  wire [32:0] _26168_;
  wire [32:0] _26169_;
  wire [32:0] _26170_;
  wire [32:0] _26171_;
  wire [32:0] _26172_;
  wire [32:0] _26173_;
  wire [32:0] _26174_;
  wire [32:0] _26175_;
  wire [32:0] _26176_;
  wire [32:0] _26177_;
  wire [32:0] _26178_;
  wire [32:0] _26179_;
  wire [32:0] _26180_;
  wire [32:0] _26181_;
  wire [32:0] _26182_;
  wire [32:0] _26183_;
  wire [32:0] _26184_;
  wire [32:0] _26185_;
  wire [32:0] _26186_;
  wire [32:0] _26187_;
  wire [32:0] _26188_;
  wire [32:0] _26189_;
  wire [32:0] _26190_;
  wire [32:0] _26191_;
  wire [32:0] _26192_;
  wire [32:0] _26193_;
  wire [32:0] _26194_;
  wire [32:0] _26195_;
  wire [32:0] _26196_;
  wire [32:0] _26197_;
  wire [32:0] _26198_;
  wire [32:0] _26199_;
  wire [32:0] _26200_;
  wire [32:0] _26201_;
  wire [32:0] _26202_;
  wire [32:0] _26203_;
  wire [32:0] _26204_;
  wire [32:0] _26205_;
  wire [32:0] _26206_;
  wire [32:0] _26207_;
  wire [32:0] _26208_;
  wire [32:0] _26209_;
  wire [32:0] _26210_;
  wire [32:0] _26211_;
  wire [32:0] _26212_;
  wire [32:0] _26213_;
  wire [32:0] _26214_;
  wire [32:0] _26215_;
  wire [32:0] _26216_;
  wire [32:0] _26217_;
  wire [32:0] _26218_;
  wire [32:0] _26219_;
  wire [32:0] _26220_;
  wire [32:0] _26221_;
  wire [32:0] _26222_;
  wire [32:0] _26223_;
  wire [32:0] _26224_;
  wire [32:0] _26225_;
  wire [32:0] _26226_;
  wire [32:0] _26227_;
  wire [32:0] _26228_;
  wire [32:0] _26229_;
  wire [32:0] _26230_;
  wire [32:0] _26231_;
  wire [32:0] _26232_;
  wire [32:0] _26233_;
  wire [32:0] _26234_;
  wire [32:0] _26235_;
  wire [32:0] _26236_;
  wire [32:0] _26237_;
  wire [32:0] _26238_;
  wire [32:0] _26239_;
  wire [32:0] _26240_;
  wire [32:0] _26241_;
  wire [32:0] _26242_;
  wire [32:0] _26243_;
  wire [32:0] _26244_;
  wire [32:0] _26245_;
  wire [32:0] _26246_;
  wire [32:0] _26247_;
  wire [32:0] _26248_;
  wire [32:0] _26249_;
  wire [32:0] _26250_;
  wire [32:0] _26251_;
  wire [32:0] _26252_;
  wire [32:0] _26253_;
  wire [32:0] _26254_;
  wire [32:0] _26255_;
  wire [31:0] _26256_;
  wire [32:0] _26257_;
  wire [32:0] _26258_;
  wire [32:0] _26259_;
  wire [32:0] _26260_;
  wire [32:0] _26261_;
  wire [32:0] _26262_;
  wire [32:0] _26263_;
  wire [32:0] _26264_;
  wire [32:0] _26265_;
  wire [32:0] _26266_;
  wire [32:0] _26267_;
  wire [32:0] _26268_;
  wire [32:0] _26269_;
  wire [31:0] _26270_;
  wire [32:0] _26271_;
  wire [32:0] _26272_;
  wire [32:0] _26273_;
  wire [32:0] _26274_;
  wire [32:0] _26275_;
  wire [32:0] _26276_;
  wire [32:0] _26277_;
  wire [32:0] _26278_;
  wire [32:0] _26279_;
  wire [32:0] _26280_;
  wire [32:0] _26281_;
  wire [32:0] _26282_;
  wire [32:0] _26283_;
  wire [32:0] _26284_;
  wire [32:0] _26285_;
  wire [32:0] _26286_;
  wire [32:0] _26287_;
  wire [32:0] _26288_;
  wire [32:0] _26289_;
  wire [32:0] _26290_;
  wire [32:0] _26291_;
  wire [32:0] _26292_;
  wire [32:0] _26293_;
  wire [32:0] _26294_;
  wire [32:0] _26295_;
  wire [32:0] _26296_;
  wire [32:0] _26297_;
  wire [32:0] _26298_;
  wire [32:0] _26299_;
  wire [32:0] _26300_;
  wire [32:0] _26301_;
  wire [32:0] _26302_;
  wire [32:0] _26303_;
  wire [32:0] _26304_;
  wire [32:0] _26305_;
  wire [32:0] _26306_;
  wire [32:0] _26307_;
  wire [32:0] _26308_;
  wire [32:0] _26309_;
  wire [32:0] _26310_;
  wire [32:0] _26311_;
  wire [32:0] _26312_;
  wire [32:0] _26313_;
  wire [32:0] _26314_;
  wire [32:0] _26315_;
  wire [32:0] _26316_;
  wire [32:0] _26317_;
  wire [32:0] _26318_;
  wire [32:0] _26319_;
  wire [31:0] _26320_;
  wire [32:0] _26321_;
  wire [31:0] _26322_;
  wire [32:0] _26323_;
  wire [32:0] _26324_;
  wire [32:0] _26325_;
  wire [1:0] _26326_;
  wire [32:0] _26327_;
  wire [32:0] _26328_;
  wire [32:0] _26329_;
  wire [65:0] _26330_;
  wire [65:0] _26331_;
  wire [65:0] _26332_;
  wire [65:0] _26333_;
  wire [65:0] _26334_;
  wire [65:0] _26335_;
  wire [65:0] _26336_;
  wire [17:0] _26337_;
  wire [17:0] _26338_;
  wire [17:0] _26339_;
  wire [17:0] _26340_;
  wire [17:0] _26341_;
  wire [17:0] _26342_;
  wire [17:0] _26343_;
  wire [17:0] _26344_;
  wire [17:0] _26345_;
  wire [17:0] _26346_;
  wire [17:0] _26347_;
  wire [17:0] _26348_;
  wire [17:0] _26349_;
  wire [17:0] _26350_;
  wire [17:0] _26351_;
  wire [17:0] _26352_;
  wire [17:0] _26353_;
  wire [17:0] _26354_;
  wire [17:0] _26355_;
  wire [17:0] _26356_;
  wire [17:0] _26357_;
  wire [17:0] _26358_;
  wire [17:0] _26359_;
  wire [17:0] _26360_;
  wire [17:0] _26361_;
  wire [17:0] _26362_;
  wire [17:0] _26363_;
  wire [31:0] _26364_;
  wire [31:0] _26365_;
  wire [31:0] _26366_;
  wire [31:0] _26367_;
  wire [31:0] _26368_;
  wire [31:0] _26369_;
  wire [39:0] _26370_;
  wire [39:0] _26371_;
  wire [39:0] _26372_;
  wire [39:0] _26373_;
  wire [39:0] _26374_;
  wire [39:0] _26375_;
  wire [15:0] _26376_;
  wire [15:0] _26377_;
  wire [15:0] _26378_;
  wire [15:0] _26379_;
  wire [15:0] _26380_;
  wire [15:0] _26381_;
  wire [15:0] _26382_;
  wire [15:0] _26383_;
  wire [15:0] _26384_;
  wire [15:0] _26385_;
  wire [15:0] _26386_;
  wire [15:0] _26387_;
  wire [15:0] _26388_;
  wire [15:0] _26389_;
  wire [15:0] _26390_;
  wire [15:0] _26391_;
  wire [15:0] _26392_;
  wire [15:0] _26393_;
  wire [15:0] _26394_;
  wire [15:0] _26395_;
  wire [15:0] _26396_;
  wire [15:0] _26397_;
  wire [15:0] _26398_;
  wire [15:0] _26399_;
  wire [15:0] _26400_;
  wire [15:0] _26401_;
  wire [15:0] _26402_;
  wire [15:0] _26403_;
  wire [15:0] _26404_;
  wire [15:0] _26405_;
  wire [15:0] _26406_;
  wire [15:0] _26407_;
  wire [15:0] _26408_;
  wire [15:0] _26409_;
  wire [15:0] _26410_;
  wire [15:0] _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire [31:0] _26444_;
  wire [31:0] _26445_;
  wire [31:0] _26446_;
  wire [31:0] _26447_;
  wire [31:0] _26448_;
  wire [31:0] _26449_;
  wire [31:0] _26450_;
  wire [31:0] _26451_;
  wire [31:0] _26452_;
  wire [31:0] _26453_;
  wire [31:0] _26454_;
  wire [31:0] _26455_;
  wire [31:0] _26456_;
  wire [31:0] _26457_;
  wire [31:0] _26458_;
  wire [31:0] _26459_;
  wire [31:0] _26460_;
  wire [31:0] _26461_;
  wire [31:0] _26462_;
  wire [31:0] _26463_;
  wire [31:0] _26464_;
  wire [31:0] _26465_;
  wire [31:0] _26466_;
  wire [31:0] _26467_;
  wire [31:0] _26468_;
  wire [31:0] _26469_;
  wire [31:0] _26470_;
  wire [31:0] _26471_;
  wire [31:0] _26472_;
  wire [31:0] _26473_;
  wire [31:0] _26474_;
  wire [31:0] _26475_;
  wire [31:0] _26476_;
  wire [31:0] _26477_;
  wire [31:0] _26478_;
  wire [31:0] _26479_;
  wire [31:0] _26480_;
  wire [31:0] _26481_;
  wire [31:0] _26482_;
  wire [31:0] _26483_;
  wire [31:0] _26484_;
  wire [31:0] _26485_;
  wire [31:0] _26486_;
  wire [31:0] _26487_;
  wire [31:0] _26488_;
  wire [31:0] _26489_;
  wire [31:0] _26490_;
  wire [31:0] _26491_;
  wire [31:0] _26492_;
  wire [31:0] _26493_;
  wire [31:0] _26494_;
  wire [31:0] _26495_;
  wire [31:0] _26496_;
  wire [31:0] _26497_;
  wire [31:0] _26498_;
  wire [31:0] _26499_;
  wire [31:0] _26500_;
  wire [31:0] _26501_;
  wire [31:0] _26502_;
  wire [31:0] _26503_;
  wire [31:0] _26504_;
  wire [31:0] _26505_;
  wire [31:0] _26506_;
  wire [31:0] _26507_;
  wire [31:0] _26508_;
  wire [31:0] _26509_;
  wire [31:0] _26510_;
  wire [32:0] _26511_;
  wire [32:0] _26512_;
  wire [65:0] _26513_;
  wire [39:0] _26514_;
  wire [39:0] _26515_;
  wire [39:0] _26516_;
  wire [31:0] _26517_;
  wire [31:0] _26518_;
  wire [31:0] _26519_;
  wire [31:0] _26520_;
  wire [31:0] _26521_;
  wire [31:0] _26522_;
  wire [31:0] _26523_;
  wire [31:0] _26524_;
  wire [31:0] _26525_;
  wire [31:0] _26526_;
  wire [31:0] _26527_;
  wire [31:0] _26528_;
  wire [31:0] _26529_;
  wire [17:0] _26530_;
  wire [17:0] _26531_;
  wire [17:0] _26532_;
  wire [17:0] _26533_;
  wire [17:0] _26534_;
  wire [17:0] _26535_;
  wire [17:0] _26536_;
  wire [17:0] _26537_;
  wire [17:0] _26538_;
  wire [31:0] _26539_;
  wire [31:0] _26540_;
  wire [31:0] _26541_;
  wire [31:0] _26542_;
  wire [31:0] _26543_;
  wire [31:0] _26544_;
  wire [31:0] _26545_;
  wire [31:0] _26546_;
  wire [31:0] _26547_;
  wire [31:0] _26548_;
  wire [31:0] _26549_;
  wire [31:0] _26550_;
  wire [31:0] _26551_;
  wire [31:0] _26552_;
  wire [31:0] _26553_;
  wire [31:0] _26554_;
  wire [31:0] _26555_;
  wire [31:0] _26556_;
  wire [31:0] _26557_;
  wire [31:0] _26558_;
  wire [31:0] _26559_;
  wire [31:0] _26560_;
  wire [31:0] _26561_;
  wire [31:0] _26562_;
  wire [31:0] _26563_;
  wire [7:0] _26564_;
  wire [7:0] _26565_;
  wire [7:0] _26566_;
  wire [7:0] _26567_;
  wire [7:0] _26568_;
  wire [7:0] _26569_;
  wire [7:0] _26570_;
  wire [7:0] _26571_;
  wire [7:0] _26572_;
  wire [7:0] _26573_;
  wire [7:0] _26574_;
  wire [7:0] _26575_;
  wire [7:0] _26576_;
  wire [7:0] _26577_;
  wire [7:0] _26578_;
  wire [7:0] _26579_;
  wire [7:0] _26580_;
  wire [7:0] _26581_;
  wire [7:0] _26582_;
  wire [7:0] _26583_;
  wire [7:0] _26584_;
  wire [7:0] _26585_;
  wire [7:0] _26586_;
  wire [7:0] _26587_;
  wire [7:0] _26588_;
  wire [7:0] _26589_;
  wire [7:0] _26590_;
  wire [7:0] _26591_;
  wire [7:0] _26592_;
  wire [7:0] _26593_;
  wire [7:0] _26594_;
  wire [7:0] _26595_;
  wire [7:0] _26596_;
  wire [7:0] _26597_;
  wire [7:0] _26598_;
  wire [7:0] _26599_;
  wire [7:0] _26600_;
  wire [7:0] _26601_;
  wire [7:0] _26602_;
  wire [7:0] _26603_;
  wire [7:0] _26604_;
  wire [7:0] _26605_;
  wire [7:0] _26606_;
  wire [7:0] _26607_;
  wire [7:0] _26608_;
  wire [7:0] _26609_;
  wire [7:0] _26610_;
  wire [7:0] _26611_;
  wire [7:0] _26612_;
  wire [7:0] _26613_;
  wire [7:0] _26614_;
  wire [7:0] _26615_;
  wire [7:0] _26616_;
  wire [7:0] _26617_;
  wire [7:0] _26618_;
  wire [7:0] _26619_;
  wire [7:0] _26620_;
  wire [7:0] _26621_;
  wire [7:0] _26622_;
  wire [7:0] _26623_;
  wire [7:0] _26624_;
  wire [7:0] _26625_;
  wire [7:0] _26626_;
  wire [7:0] _26627_;
  wire [31:0] _26628_;
  wire [31:0] _26629_;
  wire [31:0] _26630_;
  wire [8:0] _26631_;
  wire [7:0] _26632_;
  wire [7:0] _26633_;
  wire [7:0] _26634_;
  wire [31:0] _26635_;
  wire [31:0] _26636_;
  wire [31:0] _26637_;
  wire [31:0] _26638_;
  wire [31:0] _26639_;
  wire [31:0] _26640_;
  wire [31:0] _26641_;
  wire [31:0] _26642_;
  wire [31:0] _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire [31:0] _26656_;
  wire [31:0] _26657_;
  wire [31:0] _26658_;
  wire [31:0] _26659_;
  wire [31:0] _26660_;
  wire [31:0] _26661_;
  wire [31:0] _26662_;
  wire [31:0] _26663_;
  wire [31:0] _26664_;
  wire [31:0] _26665_;
  wire [31:0] _26666_;
  wire [31:0] _26667_;
  wire [31:0] _26668_;
  wire [31:0] _26669_;
  wire [31:0] _26670_;
  wire [31:0] _26671_;
  wire [31:0] _26672_;
  wire [31:0] _26673_;
  wire [31:0] _26674_;
  wire [31:0] _26675_;
  wire [31:0] _26676_;
  wire [31:0] _26677_;
  wire [31:0] _26678_;
  wire [31:0] _26679_;
  wire [31:0] _26680_;
  wire [31:0] _26681_;
  wire [31:0] _26682_;
  wire [31:0] _26683_;
  wire [31:0] _26684_;
  wire [31:0] _26685_;
  wire [31:0] _26686_;
  wire [31:0] _26687_;
  wire [31:0] _26688_;
  wire [31:0] _26689_;
  wire [31:0] _26690_;
  wire [31:0] _26691_;
  wire [31:0] _26692_;
  wire [31:0] _26693_;
  wire [31:0] _26694_;
  wire [31:0] _26695_;
  wire [31:0] _26696_;
  wire [31:0] _26697_;
  wire [31:0] _26698_;
  wire [31:0] _26699_;
  wire [31:0] _26700_;
  wire [31:0] _26701_;
  wire [31:0] _26702_;
  wire [31:0] _26703_;
  wire [31:0] _26704_;
  wire [31:0] _26705_;
  wire [31:0] _26706_;
  wire [31:0] _26707_;
  wire [31:0] _26708_;
  wire [31:0] _26709_;
  wire [31:0] _26710_;
  wire [31:0] _26711_;
  wire [31:0] _26712_;
  wire [31:0] _26713_;
  wire [31:0] _26714_;
  wire [31:0] _26715_;
  wire [31:0] _26716_;
  wire [31:0] _26717_;
  wire [31:0] _26718_;
  wire [31:0] _26719_;
  wire [31:0] _26720_;
  wire [31:0] _26721_;
  wire [31:0] _26722_;
  wire [31:0] _26723_;
  wire [31:0] _26724_;
  wire [31:0] _26725_;
  wire [31:0] _26726_;
  wire [31:0] _26727_;
  wire [31:0] _26728_;
  wire [31:0] _26729_;
  wire [31:0] _26730_;
  wire [31:0] _26731_;
  wire [31:0] _26732_;
  wire [31:0] _26733_;
  wire [31:0] _26734_;
  wire [31:0] _26735_;
  wire [31:0] _26736_;
  wire [31:0] _26737_;
  wire [31:0] _26738_;
  wire [31:0] _26739_;
  wire [31:0] _26740_;
  wire [31:0] _26741_;
  wire [31:0] _26742_;
  wire [31:0] _26743_;
  wire [31:0] _26744_;
  wire [31:0] _26745_;
  wire [31:0] _26746_;
  wire [31:0] _26747_;
  wire [31:0] _26748_;
  wire [31:0] _26749_;
  wire [31:0] _26750_;
  wire [31:0] _26751_;
  wire RESETN_inv;
  wire RST;
  wire _RESETN_inv_1;
  wire _RESETN_inv_2;
  wire [7:0] __delay_data_1000;
  wire [7:0] __delay_data_1006;
  wire [7:0] __delay_data_1007;
  wire __delay_data_1008;
  wire __delay_data_1009;
  wire __delay_data_1010;
  wire __delay_data_1011;
  wire __delay_data_1012;
  wire __delay_data_1013;
  wire [7:0] __delay_data_1014;
  wire [7:0] __delay_data_1015;
  wire [7:0] __delay_data_1016;
  wire [7:0] __delay_data_1017;
  wire [7:0] __delay_data_1018;
  wire [7:0] __delay_data_1019;
  wire [7:0] __delay_data_1020;
  wire [7:0] __delay_data_1021;
  wire [7:0] __delay_data_1035;
  wire [7:0] __delay_data_1041;
  wire __delay_data_1042;
  wire __delay_data_1043;
  wire __delay_data_1044;
  wire __delay_data_1045;
  wire __delay_data_1046;
  wire __delay_data_1047;
  wire [7:0] __delay_data_1048;
  wire [7:0] __delay_data_1049;
  wire [7:0] __delay_data_1050;
  wire [7:0] __delay_data_1051;
  wire [7:0] __delay_data_1052;
  wire [7:0] __delay_data_1053;
  wire [7:0] __delay_data_1054;
  wire [7:0] __delay_data_1055;
  wire [7:0] __delay_data_1069;
  wire [7:0] __delay_data_1075;
  wire __delay_data_1076;
  wire __delay_data_1077;
  wire __delay_data_1078;
  wire __delay_data_1079;
  wire __delay_data_1080;
  wire __delay_data_1081;
  wire [7:0] __delay_data_1082;
  wire [7:0] __delay_data_1083;
  wire [7:0] __delay_data_1084;
  wire [7:0] __delay_data_1085;
  wire [7:0] __delay_data_1086;
  wire [7:0] __delay_data_1087;
  wire [7:0] __delay_data_1088;
  wire [7:0] __delay_data_1089;
  wire [7:0] __delay_data_1103;
  wire [7:0] __delay_data_1109;
  wire __delay_data_1110;
  wire __delay_data_1111;
  wire __delay_data_1112;
  wire __delay_data_1113;
  wire __delay_data_1114;
  wire __delay_data_1115;
  wire [7:0] __delay_data_1116;
  wire [7:0] __delay_data_1117;
  wire [7:0] __delay_data_1118;
  wire [7:0] __delay_data_1119;
  wire [7:0] __delay_data_1120;
  wire [7:0] __delay_data_1121;
  wire [7:0] __delay_data_1122;
  wire [7:0] __delay_data_1123;
  wire [7:0] __delay_data_1142;
  wire __delay_data_1143;
  wire __delay_data_1144;
  wire __delay_data_1145;
  wire __delay_data_1146;
  wire __delay_data_1147;
  wire __delay_data_1148;
  wire [7:0] __delay_data_1149;
  wire [7:0] __delay_data_1150;
  wire [7:0] __delay_data_1151;
  wire [7:0] __delay_data_1152;
  wire [7:0] __delay_data_1153;
  wire [7:0] __delay_data_1154;
  wire [7:0] __delay_data_1155;
  wire [7:0] __delay_data_1156;
  wire [7:0] __delay_data_1175;
  wire __delay_data_1176;
  wire __delay_data_1177;
  wire __delay_data_1178;
  wire __delay_data_1179;
  wire __delay_data_1180;
  wire __delay_data_1181;
  wire [7:0] __delay_data_1182;
  wire [7:0] __delay_data_1183;
  wire [7:0] __delay_data_1184;
  wire [7:0] __delay_data_1185;
  wire [7:0] __delay_data_1186;
  wire [7:0] __delay_data_1187;
  wire [7:0] __delay_data_1188;
  wire [7:0] __delay_data_1189;
  wire __delay_data_1196;
  wire __delay_data_1197;
  wire __delay_data_1198;
  wire __delay_data_1199;
  wire __delay_data_1200;
  wire __delay_data_1201;
  wire __delay_data_1202;
  wire __delay_data_1203;
  wire __delay_data_1204;
  wire __delay_data_1205;
  wire __delay_data_1206;
  wire __delay_data_1207;
  wire [7:0] __delay_data_1208;
  wire __delay_data_1209;
  wire __delay_data_1210;
  wire __delay_data_1211;
  wire __delay_data_1212;
  wire __delay_data_1213;
  wire __delay_data_1214;
  wire [7:0] __delay_data_1215;
  wire [7:0] __delay_data_1216;
  wire [7:0] __delay_data_1217;
  wire [7:0] __delay_data_1218;
  wire [7:0] __delay_data_1219;
  wire [7:0] __delay_data_1220;
  wire [7:0] __delay_data_1221;
  wire [7:0] __delay_data_1222;
  wire [7:0] __delay_data_1223;
  wire [7:0] __delay_data_1224;
  wire [7:0] __delay_data_1225;
  wire [7:0] __delay_data_1226;
  wire [7:0] __delay_data_1227;
  wire [7:0] __delay_data_1228;
  wire __delay_data_1229;
  wire [7:0] __delay_data_1230;
  wire [7:0] __delay_data_1231;
  wire [7:0] __delay_data_1232;
  wire [7:0] __delay_data_1233;
  wire [7:0] __delay_data_1234;
  wire [7:0] __delay_data_1235;
  wire [7:0] __delay_data_1236;
  wire [7:0] __delay_data_1237;
  wire [7:0] __delay_data_1238;
  wire [7:0] __delay_data_1239;
  wire [7:0] __delay_data_1240;
  wire [7:0] __delay_data_1241;
  wire [7:0] __delay_data_1242;
  wire [7:0] __delay_data_1243;
  wire [7:0] __delay_data_1244;
  wire [7:0] __delay_data_1245;
  wire [7:0] __delay_data_1246;
  wire [7:0] __delay_data_1247;
  wire [7:0] __delay_data_1248;
  wire [7:0] __delay_data_1249;
  wire [4:0] __delay_data_1250;
  wire [4:0] __delay_data_1251;
  wire [4:0] __delay_data_1252;
  wire [4:0] __delay_data_1253;
  wire [4:0] __delay_data_1254;
  wire [4:0] __delay_data_1255;
  wire [4:0] __delay_data_1256;
  wire [4:0] __delay_data_1257;
  wire [4:0] __delay_data_1258;
  wire [4:0] __delay_data_1259;
  wire [4:0] __delay_data_1260;
  wire [4:0] __delay_data_1261;
  wire [4:0] __delay_data_1262;
  wire [4:0] __delay_data_1263;
  wire [4:0] __delay_data_1264;
  wire [4:0] __delay_data_1265;
  wire [4:0] __delay_data_1266;
  wire [4:0] __delay_data_1267;
  wire [4:0] __delay_data_1268;
  wire [4:0] __delay_data_1269;
  wire [4:0] __delay_data_1270;
  wire [4:0] __delay_data_1271;
  wire [31:0] __delay_data_1272;
  wire [31:0] __delay_data_1273;
  wire [31:0] __delay_data_1274;
  wire [31:0] __delay_data_1275;
  wire [31:0] __delay_data_1276;
  wire [31:0] __delay_data_1277;
  wire [31:0] __delay_data_1278;
  wire [31:0] __delay_data_1279;
  wire [31:0] __delay_data_1280;
  wire [31:0] __delay_data_1281;
  wire [31:0] __delay_data_1282;
  wire [31:0] __delay_data_1283;
  wire [31:0] __delay_data_1284;
  wire [31:0] __delay_data_1285;
  wire [31:0] __delay_data_1286;
  wire [31:0] __delay_data_1287;
  wire [31:0] __delay_data_1288;
  wire [31:0] __delay_data_1289;
  wire [31:0] __delay_data_1290;
  wire [31:0] __delay_data_1291;
  wire [31:0] __delay_data_1292;
  wire [31:0] __delay_data_1293;
  wire [31:0] __delay_data_1294;
  wire [31:0] __delay_data_1295;
  wire [31:0] __delay_data_1296;
  wire [31:0] __delay_data_1297;
  wire [31:0] __delay_data_1298;
  wire [31:0] __delay_data_1299;
  wire [3:0] __delay_data_1300;
  wire [7:0] __delay_data_1301;
  wire [7:0] __delay_data_1302;
  wire [7:0] __delay_data_1303;
  wire [7:0] __delay_data_1304;
  wire [7:0] __delay_data_1305;
  wire [7:0] __delay_data_1306;
  wire [7:0] __delay_data_1307;
  wire [7:0] __delay_data_1308;
  wire [7:0] __delay_data_1309;
  wire [7:0] __delay_data_1310;
  wire [7:0] __delay_data_1311;
  wire [7:0] __delay_data_1312;
  wire [7:0] __delay_data_1313;
  wire [7:0] __delay_data_1314;
  wire [7:0] __delay_data_1315;
  wire [7:0] __delay_data_1316;
  wire [7:0] __delay_data_1317;
  wire [7:0] __delay_data_1318;
  wire [7:0] __delay_data_1319;
  wire [7:0] __delay_data_1320;
  wire [7:0] __delay_data_1321;
  wire [7:0] __delay_data_1322;
  wire [7:0] __delay_data_1323;
  wire [7:0] __delay_data_1324;
  wire [7:0] __delay_data_1325;
  wire [7:0] __delay_data_1326;
  wire [7:0] __delay_data_1327;
  wire [7:0] __delay_data_1328;
  wire [7:0] __delay_data_1329;
  wire [7:0] __delay_data_1330;
  wire [7:0] __delay_data_1331;
  wire [7:0] __delay_data_1332;
  wire [7:0] __delay_data_1333;
  wire [7:0] __delay_data_1334;
  wire [7:0] __delay_data_1335;
  wire [7:0] __delay_data_1336;
  wire [7:0] __delay_data_1337;
  wire [7:0] __delay_data_1338;
  wire [7:0] __delay_data_1339;
  wire [7:0] __delay_data_1340;
  wire [7:0] __delay_data_1341;
  wire [7:0] __delay_data_1342;
  wire [7:0] __delay_data_1343;
  wire [7:0] __delay_data_1344;
  wire [7:0] __delay_data_1345;
  wire [7:0] __delay_data_1346;
  wire [7:0] __delay_data_1347;
  wire [7:0] __delay_data_1348;
  wire [7:0] __delay_data_1349;
  wire [7:0] __delay_data_1350;
  wire [7:0] __delay_data_1351;
  wire [7:0] __delay_data_1352;
  wire [7:0] __delay_data_1353;
  wire [7:0] __delay_data_1354;
  wire [7:0] __delay_data_1355;
  wire [7:0] __delay_data_1356;
  wire [7:0] __delay_data_1357;
  wire [7:0] __delay_data_1358;
  wire __delay_data_1370;
  wire __delay_data_1371;
  wire [3:0] __delay_data_1372;
  wire [7:0] __delay_data_1373;
  wire [7:0] __delay_data_1374;
  wire [2:0] __delay_data_1375;
  wire [2:0] __delay_data_1376;
  wire [2:0] __delay_data_1377;
  wire [7:0] __delay_data_1378;
  wire __delay_data_1379;
  wire __delay_data_1380;
  wire __delay_data_1381;
  wire __delay_data_1382;
  wire [7:0] __delay_data_1383;
  wire [7:0] __delay_data_1384;
  wire [7:0] __delay_data_1385;
  wire [7:0] __delay_data_1386;
  wire [7:0] __delay_data_1387;
  wire [7:0] __delay_data_1388;
  wire __delay_data_1389;
  wire [7:0] __delay_data_1390;
  wire [7:0] __delay_data_1391;
  wire [7:0] __delay_data_1392;
  wire [7:0] __delay_data_1393;
  wire [7:0] __delay_data_1394;
  wire [7:0] __delay_data_1395;
  wire [7:0] __delay_data_1396;
  wire [7:0] __delay_data_1397;
  wire [7:0] __delay_data_1398;
  wire [7:0] __delay_data_1399;
  wire [7:0] __delay_data_1400;
  wire [7:0] __delay_data_1401;
  wire [7:0] __delay_data_1402;
  wire [7:0] __delay_data_1403;
  wire [8:0] __delay_data_1404;
  wire [8:0] __delay_data_1405;
  wire [8:0] __delay_data_1406;
  wire [8:0] __delay_data_1407;
  wire [8:0] __delay_data_1408;
  wire [8:0] __delay_data_1409;
  wire [8:0] __delay_data_1410;
  wire [8:0] __delay_data_1411;
  wire [8:0] __delay_data_1412;
  wire [8:0] __delay_data_1413;
  wire [8:0] __delay_data_1414;
  wire [8:0] __delay_data_1415;
  wire [8:0] __delay_data_1416;
  wire [8:0] __delay_data_1417;
  wire [8:0] __delay_data_1418;
  wire [8:0] __delay_data_1419;
  wire [31:0] __delay_data_1420;
  wire [31:0] __delay_data_1421;
  wire [31:0] __delay_data_1422;
  wire [31:0] __delay_data_1423;
  wire [31:0] __delay_data_1424;
  wire [31:0] __delay_data_1425;
  wire [31:0] __delay_data_1426;
  wire [31:0] __delay_data_1427;
  wire [31:0] __delay_data_1428;
  wire [31:0] __delay_data_1429;
  wire [31:0] __delay_data_1430;
  wire [31:0] __delay_data_1431;
  wire [31:0] __delay_data_1432;
  wire [31:0] __delay_data_1433;
  wire [31:0] __delay_data_1434;
  wire [31:0] __delay_data_1435;
  wire [31:0] __delay_data_1436;
  wire [31:0] __delay_data_1437;
  wire [31:0] __delay_data_1438;
  wire [31:0] __delay_data_1439;
  wire [31:0] __delay_data_1440;
  wire [31:0] __delay_data_1441;
  wire [3:0] __delay_data_1442;
  wire [7:0] __delay_data_1443;
  wire [7:0] __delay_data_1444;
  wire [7:0] __delay_data_1445;
  wire [7:0] __delay_data_1446;
  wire [7:0] __delay_data_1447;
  wire [7:0] __delay_data_1448;
  wire [7:0] __delay_data_1449;
  wire [7:0] __delay_data_1450;
  wire [7:0] __delay_data_1451;
  wire [7:0] __delay_data_1452;
  wire [7:0] __delay_data_1453;
  wire [7:0] __delay_data_1454;
  wire [7:0] __delay_data_1455;
  wire [7:0] __delay_data_1456;
  wire [7:0] __delay_data_1457;
  wire [7:0] __delay_data_1458;
  wire [7:0] __delay_data_1459;
  wire [7:0] __delay_data_1460;
  wire [7:0] __delay_data_1461;
  wire [7:0] __delay_data_1462;
  wire [7:0] __delay_data_1463;
  wire [7:0] __delay_data_1464;
  wire [7:0] __delay_data_1465;
  wire [7:0] __delay_data_1466;
  wire [7:0] __delay_data_1467;
  wire [7:0] __delay_data_1468;
  wire [7:0] __delay_data_1469;
  wire [7:0] __delay_data_1470;
  wire [7:0] __delay_data_1471;
  wire [7:0] __delay_data_1472;
  wire [7:0] __delay_data_1473;
  wire [7:0] __delay_data_1474;
  wire [7:0] __delay_data_1475;
  wire [7:0] __delay_data_1476;
  wire [7:0] __delay_data_1477;
  wire [7:0] __delay_data_1478;
  wire [7:0] __delay_data_1479;
  wire [7:0] __delay_data_1480;
  wire [7:0] __delay_data_1481;
  wire [7:0] __delay_data_1482;
  wire [7:0] __delay_data_1483;
  wire [7:0] __delay_data_1484;
  wire [7:0] __delay_data_1485;
  wire [7:0] __delay_data_1486;
  wire [7:0] __delay_data_1487;
  wire __delay_data_1488;
  wire __delay_data_1489;
  wire __delay_data_1490;
  wire __delay_data_1491;
  wire __delay_data_1492;
  wire __delay_data_1493;
  wire __delay_data_1494;
  wire __delay_data_1495;
  wire __delay_data_1496;
  wire __delay_data_1497;
  wire __delay_data_1498;
  wire __delay_data_573;
  wire [7:0] __delay_data_574;
  wire [7:0] __delay_data_575;
  wire [7:0] __delay_data_576;
  wire [7:0] __delay_data_577;
  wire [7:0] __delay_data_578;
  wire [7:0] __delay_data_579;
  wire [3:0] __delay_data_580;
  wire [3:0] __delay_data_581;
  wire [3:0] __delay_data_582;
  wire [3:0] __delay_data_583;
  wire [3:0] __delay_data_584;
  wire [3:0] __delay_data_585;
  wire [3:0] __delay_data_586;
  wire __delay_data_590;
  wire [7:0] __delay_data_591;
  wire [7:0] __delay_data_592;
  wire [7:0] __delay_data_593;
  wire [7:0] __delay_data_594;
  wire [7:0] __delay_data_595;
  wire [7:0] __delay_data_596;
  wire [3:0] __delay_data_597;
  wire [3:0] __delay_data_598;
  wire [3:0] __delay_data_599;
  wire [3:0] __delay_data_600;
  wire [3:0] __delay_data_601;
  wire [3:0] __delay_data_602;
  wire [3:0] __delay_data_603;
  wire __delay_data_607;
  wire [7:0] __delay_data_608;
  wire [7:0] __delay_data_609;
  wire [7:0] __delay_data_610;
  wire [7:0] __delay_data_611;
  wire [7:0] __delay_data_612;
  wire [7:0] __delay_data_613;
  wire [3:0] __delay_data_614;
  wire [3:0] __delay_data_615;
  wire [3:0] __delay_data_616;
  wire [3:0] __delay_data_617;
  wire [3:0] __delay_data_618;
  wire [3:0] __delay_data_619;
  wire [3:0] __delay_data_620;
  wire __delay_data_624;
  wire [7:0] __delay_data_625;
  wire [7:0] __delay_data_626;
  wire [7:0] __delay_data_627;
  wire [7:0] __delay_data_628;
  wire [7:0] __delay_data_629;
  wire [7:0] __delay_data_630;
  wire [3:0] __delay_data_631;
  wire [3:0] __delay_data_632;
  wire [3:0] __delay_data_633;
  wire [3:0] __delay_data_634;
  wire [3:0] __delay_data_635;
  wire [3:0] __delay_data_636;
  wire [3:0] __delay_data_637;
  wire __delay_data_641;
  wire [7:0] __delay_data_642;
  wire [7:0] __delay_data_643;
  wire [7:0] __delay_data_644;
  wire [7:0] __delay_data_645;
  wire [7:0] __delay_data_646;
  wire [7:0] __delay_data_647;
  wire [3:0] __delay_data_648;
  wire [3:0] __delay_data_649;
  wire [3:0] __delay_data_650;
  wire [3:0] __delay_data_651;
  wire [3:0] __delay_data_652;
  wire [3:0] __delay_data_653;
  wire [3:0] __delay_data_654;
  wire __delay_data_658;
  wire [7:0] __delay_data_659;
  wire [7:0] __delay_data_660;
  wire [7:0] __delay_data_661;
  wire [7:0] __delay_data_662;
  wire [7:0] __delay_data_663;
  wire [7:0] __delay_data_664;
  wire [3:0] __delay_data_665;
  wire [3:0] __delay_data_666;
  wire [3:0] __delay_data_667;
  wire [3:0] __delay_data_668;
  wire [3:0] __delay_data_669;
  wire [3:0] __delay_data_670;
  wire [3:0] __delay_data_671;
  wire __delay_data_675;
  wire [7:0] __delay_data_676;
  wire [7:0] __delay_data_677;
  wire [7:0] __delay_data_678;
  wire [7:0] __delay_data_679;
  wire [7:0] __delay_data_680;
  wire [7:0] __delay_data_681;
  wire [3:0] __delay_data_682;
  wire [3:0] __delay_data_683;
  wire [3:0] __delay_data_684;
  wire [3:0] __delay_data_685;
  wire [3:0] __delay_data_686;
  wire [3:0] __delay_data_687;
  wire [3:0] __delay_data_688;
  wire __delay_data_692;
  wire [7:0] __delay_data_693;
  wire [7:0] __delay_data_694;
  wire [7:0] __delay_data_695;
  wire [7:0] __delay_data_696;
  wire [7:0] __delay_data_697;
  wire [7:0] __delay_data_698;
  wire [3:0] __delay_data_699;
  wire [3:0] __delay_data_700;
  wire [3:0] __delay_data_701;
  wire [3:0] __delay_data_702;
  wire [3:0] __delay_data_703;
  wire [3:0] __delay_data_704;
  wire [3:0] __delay_data_705;
  wire __delay_data_709;
  wire [7:0] __delay_data_710;
  wire [7:0] __delay_data_711;
  wire [7:0] __delay_data_712;
  wire [7:0] __delay_data_713;
  wire [7:0] __delay_data_714;
  wire [7:0] __delay_data_715;
  wire [3:0] __delay_data_716;
  wire [3:0] __delay_data_717;
  wire [3:0] __delay_data_718;
  wire [3:0] __delay_data_719;
  wire [3:0] __delay_data_720;
  wire [3:0] __delay_data_721;
  wire [3:0] __delay_data_722;
  wire __delay_data_728;
  wire [31:0] __delay_data_729;
  wire [31:0] __delay_data_730;
  wire [5:0] __delay_data_731;
  wire [5:0] __delay_data_732;
  wire [5:0] __delay_data_733;
  wire [5:0] __delay_data_734;
  wire __delay_data_735;
  wire __delay_data_736;
  wire __delay_data_737;
  wire __delay_data_738;
  wire [5:0] __delay_data_744;
  wire [5:0] __delay_data_745;
  wire [5:0] __delay_data_746;
  wire [5:0] __delay_data_747;
  wire [39:0] __delay_data_748;
  wire __delay_data_749;
  wire [7:0] __delay_data_868;
  wire __delay_data_869;
  wire [7:0] __delay_data_870;
  wire [7:0] __delay_data_871;
  wire [7:0] __delay_data_874;
  wire [7:0] __delay_data_875;
  wire [7:0] __delay_data_876;
  wire [7:0] __delay_data_877;
  wire [7:0] __delay_data_879;
  wire [7:0] __delay_data_880;
  wire [7:0] __delay_data_883;
  wire [7:0] __delay_data_884;
  wire [7:0] __delay_data_885;
  wire [7:0] __delay_data_886;
  wire [7:0] __delay_data_888;
  wire [7:0] __delay_data_889;
  wire [7:0] __delay_data_892;
  wire [7:0] __delay_data_893;
  wire [7:0] __delay_data_894;
  wire [7:0] __delay_data_902;
  wire [7:0] __delay_data_908;
  wire [7:0] __delay_data_909;
  wire __delay_data_910;
  wire __delay_data_911;
  wire __delay_data_912;
  wire __delay_data_913;
  wire __delay_data_914;
  wire __delay_data_915;
  wire __delay_data_916;
  wire [7:0] __delay_data_917;
  wire [7:0] __delay_data_918;
  wire [7:0] __delay_data_919;
  wire [7:0] __delay_data_920;
  wire [7:0] __delay_data_921;
  wire [7:0] __delay_data_922;
  wire [7:0] __delay_data_923;
  wire [7:0] __delay_data_924;
  wire [7:0] __delay_data_932;
  wire [7:0] __delay_data_935;
  wire [7:0] __delay_data_937;
  wire [7:0] __delay_data_940;
  wire [7:0] __delay_data_942;
  wire [7:0] __delay_data_945;
  wire [7:0] __delay_data_953;
  wire [7:0] __delay_data_959;
  wire [7:0] __delay_data_960;
  wire __delay_data_961;
  wire __delay_data_962;
  wire __delay_data_963;
  wire __delay_data_964;
  wire __delay_data_965;
  wire __delay_data_966;
  wire [7:0] __delay_data_967;
  wire [7:0] __delay_data_968;
  wire [7:0] __delay_data_969;
  wire [7:0] __delay_data_970;
  wire [7:0] __delay_data_971;
  wire [7:0] __delay_data_972;
  wire [7:0] __delay_data_973;
  wire [7:0] __delay_data_974;
  wire [7:0] __delay_data_984;
  wire [7:0] __delay_data_988;
  wire __delay_data_990;
  wire __delay_data_991;
  wire [7:0] __delay_data_992;
  wire __maxi_read_fsm_cond_3_0_1;
  wire __maxi_read_fsm_cond_3_2_1;
  wire __maxi_read_fsm_cond_3_3_1;
  wire __maxi_read_fsm_cond_3_4_1;
  wire __maxi_read_fsm_cond_3_5_1;
  wire __maxi_read_fsm_cond_3_6_1;
  wire __maxi_read_fsm_cond_3_7_1;
  wire __maxi_read_fsm_cond_3_8_1;
  wire __maxi_read_fsm_cond_3_9_1;
  wire __maxi_read_fsm_cond_4_1_1;
  wire __maxi_write_fsm_cond_4_0_1;
  wire [7:0] \__muladd_madd_110.madd._a ;
  wire [7:0] \__muladd_madd_110.madd._b ;
  wire [15:0] \__muladd_madd_110.madd._c ;
  wire [15:0] \__muladd_madd_110.madd._madd ;
  wire [15:0] \__muladd_madd_110.madd._mul ;
  wire [15:0] \__muladd_madd_110.madd._pipe_madd0 ;
  wire [15:0] \__muladd_madd_110.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_125.madd._a ;
  wire [7:0] \__muladd_madd_125.madd._b ;
  wire [15:0] \__muladd_madd_125.madd._c ;
  wire [15:0] \__muladd_madd_125.madd._madd ;
  wire [15:0] \__muladd_madd_125.madd._mul ;
  wire [15:0] \__muladd_madd_125.madd._pipe_madd0 ;
  wire [15:0] \__muladd_madd_125.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_140.madd._a ;
  wire [7:0] \__muladd_madd_140.madd._b ;
  wire [15:0] \__muladd_madd_140.madd._c ;
  wire [15:0] \__muladd_madd_140.madd._madd ;
  wire [15:0] \__muladd_madd_140.madd._mul ;
  wire [15:0] \__muladd_madd_140.madd._pipe_madd0 ;
  wire [15:0] \__muladd_madd_140.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_155.madd._a ;
  wire [7:0] \__muladd_madd_155.madd._b ;
  wire [15:0] \__muladd_madd_155.madd._c ;
  wire [15:0] \__muladd_madd_155.madd._madd ;
  wire [15:0] \__muladd_madd_155.madd._mul ;
  wire [15:0] \__muladd_madd_155.madd._pipe_madd0 ;
  wire [15:0] \__muladd_madd_155.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_170.madd._a ;
  wire [7:0] \__muladd_madd_170.madd._b ;
  wire [15:0] \__muladd_madd_170.madd._c ;
  wire [15:0] \__muladd_madd_170.madd._madd ;
  wire [15:0] \__muladd_madd_170.madd._mul ;
  wire [15:0] \__muladd_madd_170.madd._pipe_madd0 ;
  wire [15:0] \__muladd_madd_170.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_185.madd._a ;
  wire [7:0] \__muladd_madd_185.madd._b ;
  wire [15:0] \__muladd_madd_185.madd._c ;
  wire [15:0] \__muladd_madd_185.madd._madd ;
  wire [15:0] \__muladd_madd_185.madd._mul ;
  wire [15:0] \__muladd_madd_185.madd._pipe_madd0 ;
  wire [15:0] \__muladd_madd_185.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_65.madd._a ;
  wire [7:0] \__muladd_madd_65.madd._b ;
  wire [15:0] \__muladd_madd_65.madd._c ;
  wire [15:0] \__muladd_madd_65.madd._madd ;
  wire [15:0] \__muladd_madd_65.madd._mul ;
  wire [15:0] \__muladd_madd_65.madd._pipe_madd0 ;
  wire [15:0] \__muladd_madd_65.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_80.madd._a ;
  wire [7:0] \__muladd_madd_80.madd._b ;
  wire [15:0] \__muladd_madd_80.madd._c ;
  wire [15:0] \__muladd_madd_80.madd._madd ;
  wire [15:0] \__muladd_madd_80.madd._mul ;
  wire [15:0] \__muladd_madd_80.madd._pipe_madd0 ;
  wire [15:0] \__muladd_madd_80.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_95.madd._a ;
  wire [7:0] \__muladd_madd_95.madd._b ;
  wire [15:0] \__muladd_madd_95.madd._c ;
  wire [15:0] \__muladd_madd_95.madd._madd ;
  wire [15:0] \__muladd_madd_95.madd._mul ;
  wire [15:0] \__muladd_madd_95.madd._pipe_madd0 ;
  wire [15:0] \__muladd_madd_95.madd._pipe_madd1 ;
  wire [15:0] __muladd_madd_odata_reg_110;
  wire [15:0] __muladd_madd_odata_reg_125;
  wire [15:0] __muladd_madd_odata_reg_140;
  wire [15:0] __muladd_madd_odata_reg_155;
  wire [15:0] __muladd_madd_odata_reg_170;
  wire [15:0] __muladd_madd_odata_reg_185;
  wire [15:0] __muladd_madd_odata_reg_65;
  wire [15:0] __muladd_madd_odata_reg_80;
  wire [15:0] __muladd_madd_odata_reg_95;
  wire [31:0] __plusn_data_32;
  wire [31:0] __plusn_data_33;
  wire [31:0] __plusn_data_34;
  wire [31:0] __plusn_data_35;
  wire __reduce_max_13_reduce_reset;
  wire __set_flag_1034_1;
  wire __set_flag_1034_10;
  wire __set_flag_1034_11;
  wire __set_flag_1034_12;
  wire __set_flag_1034_13;
  wire __set_flag_1034_14;
  wire __set_flag_1034_15;
  wire __set_flag_1034_16;
  wire __set_flag_1034_17;
  wire __set_flag_1034_18;
  wire __set_flag_1034_19;
  wire __set_flag_1034_2;
  wire __set_flag_1034_20;
  wire __set_flag_1034_21;
  wire __set_flag_1034_22;
  wire __set_flag_1034_23;
  wire __set_flag_1034_24;
  wire __set_flag_1034_25;
  wire __set_flag_1034_26;
  wire __set_flag_1034_27;
  wire __set_flag_1034_28;
  wire __set_flag_1034_29;
  wire __set_flag_1034_3;
  wire __set_flag_1034_30;
  wire __set_flag_1034_31;
  wire __set_flag_1034_32;
  wire __set_flag_1034_33;
  wire __set_flag_1034_34;
  wire __set_flag_1034_35;
  wire __set_flag_1034_36;
  wire __set_flag_1034_37;
  wire __set_flag_1034_4;
  wire __set_flag_1034_5;
  wire __set_flag_1034_6;
  wire __set_flag_1034_7;
  wire __set_flag_1034_8;
  wire __set_flag_1034_9;
  wire __set_flag_538_1;
  wire __set_flag_538_10;
  wire __set_flag_538_11;
  wire __set_flag_538_12;
  wire __set_flag_538_13;
  wire __set_flag_538_14;
  wire __set_flag_538_15;
  wire __set_flag_538_16;
  wire __set_flag_538_17;
  wire __set_flag_538_18;
  wire __set_flag_538_19;
  wire __set_flag_538_2;
  wire __set_flag_538_20;
  wire __set_flag_538_21;
  wire __set_flag_538_22;
  wire __set_flag_538_23;
  wire __set_flag_538_24;
  wire __set_flag_538_25;
  wire __set_flag_538_26;
  wire __set_flag_538_27;
  wire __set_flag_538_28;
  wire __set_flag_538_29;
  wire __set_flag_538_3;
  wire __set_flag_538_30;
  wire __set_flag_538_31;
  wire __set_flag_538_32;
  wire __set_flag_538_33;
  wire __set_flag_538_34;
  wire __set_flag_538_35;
  wire __set_flag_538_36;
  wire __set_flag_538_37;
  wire __set_flag_538_38;
  wire __set_flag_538_39;
  wire __set_flag_538_4;
  wire __set_flag_538_40;
  wire __set_flag_538_41;
  wire __set_flag_538_42;
  wire __set_flag_538_43;
  wire __set_flag_538_44;
  wire __set_flag_538_45;
  wire __set_flag_538_5;
  wire __set_flag_538_6;
  wire __set_flag_538_7;
  wire __set_flag_538_8;
  wire __set_flag_538_9;
  wire __set_flag_874_1;
  wire __set_flag_874_2;
  wire __set_flag_874_3;
  wire __set_flag_874_4;
  wire __set_flag_874_5;
  wire __set_flag_874_6;
  wire __set_flag_874_7;
  wire __set_flag_874_8;
  wire __set_flag_874_9;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_1;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_10;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_11;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_12;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_13;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_14;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_15;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_16;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_17;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_18;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_19;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_2;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_20;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_21;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_22;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_23;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_24;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_25;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_26;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_27;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_28;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_29;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_3;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_30;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_31;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_32;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_33;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_34;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_35;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_36;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_37;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_38;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_39;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_4;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_40;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_41;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_42;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_43;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_44;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_45;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_5;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_6;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_7;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_8;
  wire [31:0] __stream_conv2d_8_sink_37_sink_offset_0_9;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_1;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_10;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_11;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_12;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_13;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_14;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_15;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_16;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_17;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_18;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_19;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_2;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_20;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_21;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_22;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_23;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_24;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_25;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_26;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_27;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_28;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_29;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_3;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_30;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_31;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_32;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_33;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_34;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_35;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_36;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_37;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_38;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_39;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_4;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_40;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_41;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_42;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_43;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_44;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_45;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_5;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_6;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_7;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_8;
  wire [32:0] __stream_conv2d_8_sink_37_sink_size_1_9;
  wire __stream_conv2d_8_start_1;
  wire __stream_conv2d_8_start_10;
  wire __stream_conv2d_8_start_11;
  wire __stream_conv2d_8_start_12;
  wire __stream_conv2d_8_start_13;
  wire __stream_conv2d_8_start_14;
  wire __stream_conv2d_8_start_15;
  wire __stream_conv2d_8_start_16;
  wire __stream_conv2d_8_start_17;
  wire __stream_conv2d_8_start_18;
  wire __stream_conv2d_8_start_19;
  wire __stream_conv2d_8_start_2;
  wire __stream_conv2d_8_start_20;
  wire __stream_conv2d_8_start_21;
  wire __stream_conv2d_8_start_22;
  wire __stream_conv2d_8_start_23;
  wire __stream_conv2d_8_start_24;
  wire __stream_conv2d_8_start_25;
  wire __stream_conv2d_8_start_26;
  wire __stream_conv2d_8_start_27;
  wire __stream_conv2d_8_start_28;
  wire __stream_conv2d_8_start_29;
  wire __stream_conv2d_8_start_3;
  wire __stream_conv2d_8_start_30;
  wire __stream_conv2d_8_start_31;
  wire __stream_conv2d_8_start_32;
  wire __stream_conv2d_8_start_33;
  wire __stream_conv2d_8_start_34;
  wire __stream_conv2d_8_start_35;
  wire __stream_conv2d_8_start_36;
  wire __stream_conv2d_8_start_37;
  wire __stream_conv2d_8_start_38;
  wire __stream_conv2d_8_start_39;
  wire __stream_conv2d_8_start_4;
  wire __stream_conv2d_8_start_40;
  wire __stream_conv2d_8_start_41;
  wire __stream_conv2d_8_start_42;
  wire __stream_conv2d_8_start_43;
  wire __stream_conv2d_8_start_44;
  wire __stream_conv2d_8_start_45;
  wire __stream_conv2d_8_start_46;
  wire __stream_conv2d_8_start_5;
  wire __stream_conv2d_8_start_6;
  wire __stream_conv2d_8_start_7;
  wire __stream_conv2d_8_start_8;
  wire __stream_conv2d_8_start_9;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_1;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_10;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_11;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_12;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_13;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_14;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_15;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_16;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_17;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_18;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_19;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_2;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_20;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_21;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_22;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_23;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_24;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_25;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_26;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_27;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_28;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_29;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_3;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_30;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_31;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_32;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_33;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_34;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_35;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_36;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_37;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_4;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_5;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_6;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_7;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_8;
  wire [31:0] __stream_matmul_15_sink_21_sink_offset_0_9;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_1;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_10;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_11;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_12;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_13;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_14;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_15;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_16;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_17;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_18;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_19;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_2;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_20;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_21;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_22;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_23;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_24;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_25;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_26;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_27;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_28;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_29;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_3;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_30;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_31;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_32;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_33;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_34;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_35;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_36;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_37;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_4;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_5;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_6;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_7;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_8;
  wire [32:0] __stream_matmul_15_sink_21_sink_size_1_9;
  wire __stream_matmul_15_start_1;
  wire __stream_matmul_15_start_10;
  wire __stream_matmul_15_start_11;
  wire __stream_matmul_15_start_12;
  wire __stream_matmul_15_start_13;
  wire __stream_matmul_15_start_14;
  wire __stream_matmul_15_start_15;
  wire __stream_matmul_15_start_16;
  wire __stream_matmul_15_start_17;
  wire __stream_matmul_15_start_18;
  wire __stream_matmul_15_start_19;
  wire __stream_matmul_15_start_2;
  wire __stream_matmul_15_start_20;
  wire __stream_matmul_15_start_21;
  wire __stream_matmul_15_start_22;
  wire __stream_matmul_15_start_23;
  wire __stream_matmul_15_start_24;
  wire __stream_matmul_15_start_25;
  wire __stream_matmul_15_start_26;
  wire __stream_matmul_15_start_27;
  wire __stream_matmul_15_start_28;
  wire __stream_matmul_15_start_29;
  wire __stream_matmul_15_start_3;
  wire __stream_matmul_15_start_30;
  wire __stream_matmul_15_start_31;
  wire __stream_matmul_15_start_32;
  wire __stream_matmul_15_start_33;
  wire __stream_matmul_15_start_34;
  wire __stream_matmul_15_start_35;
  wire __stream_matmul_15_start_36;
  wire __stream_matmul_15_start_37;
  wire __stream_matmul_15_start_38;
  wire __stream_matmul_15_start_4;
  wire __stream_matmul_15_start_5;
  wire __stream_matmul_15_start_6;
  wire __stream_matmul_15_start_7;
  wire __stream_matmul_15_start_8;
  wire __stream_matmul_15_start_9;
  wire [31:0] __stream_max_pool_serial_9_sink_3_sink_offset_0_1;
  wire [31:0] __stream_max_pool_serial_9_sink_3_sink_offset_0_2;
  wire [31:0] __stream_max_pool_serial_9_sink_3_sink_offset_0_3;
  wire [31:0] __stream_max_pool_serial_9_sink_3_sink_offset_0_4;
  wire [31:0] __stream_max_pool_serial_9_sink_3_sink_offset_0_5;
  wire [31:0] __stream_max_pool_serial_9_sink_3_sink_offset_0_6;
  wire [31:0] __stream_max_pool_serial_9_sink_3_sink_offset_0_7;
  wire [31:0] __stream_max_pool_serial_9_sink_3_sink_offset_0_8;
  wire [31:0] __stream_max_pool_serial_9_sink_3_sink_offset_0_9;
  wire [32:0] __stream_max_pool_serial_9_sink_3_sink_size_1_1;
  wire [32:0] __stream_max_pool_serial_9_sink_3_sink_size_1_2;
  wire [32:0] __stream_max_pool_serial_9_sink_3_sink_size_1_3;
  wire [32:0] __stream_max_pool_serial_9_sink_3_sink_size_1_4;
  wire [32:0] __stream_max_pool_serial_9_sink_3_sink_size_1_5;
  wire [32:0] __stream_max_pool_serial_9_sink_3_sink_size_1_6;
  wire [32:0] __stream_max_pool_serial_9_sink_3_sink_size_1_7;
  wire [32:0] __stream_max_pool_serial_9_sink_3_sink_size_1_8;
  wire [32:0] __stream_max_pool_serial_9_sink_3_sink_size_1_9;
  wire __stream_max_pool_serial_9_start_1;
  wire __stream_max_pool_serial_9_start_10;
  wire __stream_max_pool_serial_9_start_2;
  wire __stream_max_pool_serial_9_start_3;
  wire __stream_max_pool_serial_9_start_4;
  wire __stream_max_pool_serial_9_start_5;
  wire __stream_max_pool_serial_9_start_6;
  wire __stream_max_pool_serial_9_start_7;
  wire __stream_max_pool_serial_9_start_8;
  wire __stream_max_pool_serial_9_start_9;
  wire [15:0] __substreamoutput_data_605;
  wire [15:0] __substreamoutput_data_622;
  wire [15:0] __substreamoutput_data_639;
  wire [15:0] __substreamoutput_data_656;
  wire [15:0] __substreamoutput_data_673;
  wire [15:0] __substreamoutput_data_690;
  wire [15:0] __substreamoutput_data_707;
  wire [15:0] __substreamoutput_data_724;
  wire [31:0] __substreamoutput_data_726;
  wire [31:0] __substreamoutput_data_773;
  wire __substreamoutput_data_774;
  wire [15:0] __substreamoutput_data_856;
  wire [31:0] __substreamoutput_data_858;
  wire [31:0] __substreamoutput_data_861;
  wire __substreamoutput_data_862;
  wire [7:0] __substreamoutput_data_866;
  wire [1:0] __tmp_1015_1;
  wire [1:0] __tmp_1015_2;
  wire [1:0] __tmp_1025_1;
  wire [1:0] __tmp_1025_2;
  wire __tmp_1059_1;
  wire __tmp_1059_10;
  wire __tmp_1059_11;
  wire __tmp_1059_12;
  wire __tmp_1059_13;
  wire __tmp_1059_14;
  wire __tmp_1059_15;
  wire __tmp_1059_16;
  wire __tmp_1059_17;
  wire __tmp_1059_18;
  wire __tmp_1059_19;
  wire __tmp_1059_2;
  wire __tmp_1059_20;
  wire __tmp_1059_21;
  wire __tmp_1059_22;
  wire __tmp_1059_23;
  wire __tmp_1059_24;
  wire __tmp_1059_25;
  wire __tmp_1059_26;
  wire __tmp_1059_27;
  wire __tmp_1059_28;
  wire __tmp_1059_3;
  wire __tmp_1059_4;
  wire __tmp_1059_5;
  wire __tmp_1059_6;
  wire __tmp_1059_7;
  wire __tmp_1059_8;
  wire __tmp_1059_9;
  wire __tmp_1095_1;
  wire __tmp_1095_2;
  wire __tmp_1095_3;
  wire __tmp_1095_4;
  wire __tmp_1095_5;
  wire __tmp_1095_6;
  wire __tmp_1095_7;
  wire __tmp_1095_8;
  wire __tmp_1095_9;
  wire __tmp_1107_10;
  wire __tmp_1107_11;
  wire __tmp_1107_12;
  wire __tmp_1115_35;
  wire __tmp_1115_36;
  wire __tmp_1115_37;
  wire __tmp_1115_38;
  wire __tmp_1117_13;
  wire __tmp_1117_14;
  wire __tmp_1117_15;
  wire __tmp_1117_16;
  wire __tmp_1117_17;
  wire __tmp_1117_18;
  wire __tmp_1117_19;
  wire __tmp_1117_20;
  wire __tmp_1117_21;
  wire __tmp_1117_22;
  wire __tmp_1117_23;
  wire __tmp_1117_24;
  wire __tmp_1117_25;
  wire __tmp_1117_26;
  wire __tmp_1117_27;
  wire __tmp_1117_28;
  wire __tmp_1117_29;
  wire __tmp_1117_30;
  wire __tmp_1117_31;
  wire __tmp_1117_32;
  wire __tmp_1117_33;
  wire __tmp_1117_34;
  wire __tmp_1124_1;
  wire [7:0] __tmp_1125_1;
  wire __tmp_1136_1;
  wire [7:0] __tmp_1137_1;
  wire __tmp_1148_1;
  wire [7:0] __tmp_1149_1;
  wire __tmp_1160_1;
  wire [7:0] __tmp_1161_1;
  wire [1:0] __tmp_339_1;
  wire [1:0] __tmp_339_2;
  wire [1:0] __tmp_359_1;
  wire [1:0] __tmp_359_2;
  wire [1:0] __tmp_369_1;
  wire [1:0] __tmp_369_2;
  wire [1:0] __tmp_379_1;
  wire [1:0] __tmp_379_2;
  wire [1:0] __tmp_389_1;
  wire [1:0] __tmp_389_2;
  wire [1:0] __tmp_399_1;
  wire [1:0] __tmp_399_2;
  wire [1:0] __tmp_409_1;
  wire [1:0] __tmp_409_2;
  wire [1:0] __tmp_419_1;
  wire [1:0] __tmp_419_2;
  wire [1:0] __tmp_429_1;
  wire [1:0] __tmp_429_2;
  wire [1:0] __tmp_439_1;
  wire [1:0] __tmp_439_2;
  wire [1:0] __tmp_449_1;
  wire [1:0] __tmp_449_2;
  wire [1:0] __tmp_459_1;
  wire [1:0] __tmp_459_2;
  wire [1:0] __tmp_469_1;
  wire [1:0] __tmp_469_2;
  wire [1:0] __tmp_479_1;
  wire [1:0] __tmp_479_2;
  wire [1:0] __tmp_489_1;
  wire [1:0] __tmp_489_2;
  wire [1:0] __tmp_499_1;
  wire [1:0] __tmp_499_2;
  wire [1:0] __tmp_509_1;
  wire [1:0] __tmp_509_2;
  wire [1:0] __tmp_519_1;
  wire [1:0] __tmp_519_2;
  wire [1:0] __tmp_529_1;
  wire [1:0] __tmp_529_2;
  wire __tmp_627_1;
  wire __tmp_627_10;
  wire __tmp_627_11;
  wire __tmp_627_12;
  wire __tmp_627_13;
  wire __tmp_627_14;
  wire __tmp_627_15;
  wire __tmp_627_16;
  wire __tmp_627_17;
  wire __tmp_627_18;
  wire __tmp_627_19;
  wire __tmp_627_2;
  wire __tmp_627_20;
  wire __tmp_627_21;
  wire __tmp_627_22;
  wire __tmp_627_23;
  wire __tmp_627_24;
  wire __tmp_627_25;
  wire __tmp_627_26;
  wire __tmp_627_27;
  wire __tmp_627_28;
  wire __tmp_627_29;
  wire __tmp_627_3;
  wire __tmp_627_30;
  wire __tmp_627_31;
  wire __tmp_627_32;
  wire __tmp_627_33;
  wire __tmp_627_34;
  wire __tmp_627_4;
  wire __tmp_627_5;
  wire __tmp_627_6;
  wire __tmp_627_7;
  wire __tmp_627_8;
  wire __tmp_627_9;
  wire __tmp_775_1;
  wire __tmp_775_2;
  wire __tmp_775_3;
  wire __tmp_775_4;
  wire __tmp_775_5;
  wire __tmp_775_6;
  wire __tmp_775_7;
  wire __tmp_775_8;
  wire __tmp_775_9;
  wire __tmp_787_10;
  wire __tmp_787_11;
  wire __tmp_787_12;
  wire __tmp_795_43;
  wire __tmp_795_44;
  wire __tmp_795_45;
  wire __tmp_795_46;
  wire __tmp_797_13;
  wire __tmp_797_14;
  wire __tmp_797_15;
  wire __tmp_797_16;
  wire __tmp_797_17;
  wire __tmp_797_18;
  wire __tmp_797_19;
  wire __tmp_797_20;
  wire __tmp_797_21;
  wire __tmp_797_22;
  wire __tmp_797_23;
  wire __tmp_797_24;
  wire __tmp_797_25;
  wire __tmp_797_26;
  wire __tmp_797_27;
  wire __tmp_797_28;
  wire __tmp_797_29;
  wire __tmp_797_30;
  wire __tmp_797_31;
  wire __tmp_797_32;
  wire __tmp_797_33;
  wire __tmp_797_34;
  wire __tmp_797_35;
  wire __tmp_797_36;
  wire __tmp_797_37;
  wire __tmp_797_38;
  wire __tmp_797_39;
  wire __tmp_797_40;
  wire __tmp_797_41;
  wire __tmp_797_42;
  wire __tmp_804_1;
  wire [7:0] __tmp_805_1;
  wire __tmp_816_1;
  wire [7:0] __tmp_817_1;
  wire __tmp_828_1;
  wire [7:0] __tmp_829_1;
  wire __tmp_840_1;
  wire [7:0] __tmp_841_1;
  wire [1:0] __tmp_865_1;
  wire [1:0] __tmp_865_2;
  wire __tmp_880_8;
  wire __tmp_880_9;
  wire __tmp_884_1;
  wire __tmp_884_2;
  wire __tmp_884_3;
  wire __tmp_884_4;
  wire __tmp_884_5;
  wire __tmp_884_6;
  wire __tmp_884_7;
  wire __tmp_906_10;
  wire __tmp_906_7;
  wire __tmp_906_8;
  wire __tmp_906_9;
  wire __tmp_908_1;
  wire __tmp_908_2;
  wire __tmp_908_3;
  wire __tmp_908_4;
  wire __tmp_908_5;
  wire __tmp_908_6;
  wire __tmp_915_1;
  wire [7:0] __tmp_916_1;
  wire __tmp_927_1;
  wire [7:0] __tmp_928_1;
  wire __tmp_939_1;
  wire [7:0] __tmp_940_1;
  wire __tmp_951_1;
  wire [7:0] __tmp_952_1;
  wire [1:0] __tmp_995_1;
  wire [1:0] __tmp_995_2;
  wire [31:0] __variable_wdata_0;
  wire [5:0] __variable_wdata_1;
  wire [7:0] __variable_wdata_112;
  wire [7:0] __variable_wdata_113;
  wire [3:0] __variable_wdata_114;
  wire [7:0] __variable_wdata_127;
  wire [7:0] __variable_wdata_128;
  wire [3:0] __variable_wdata_129;
  wire [7:0] __variable_wdata_142;
  wire [7:0] __variable_wdata_143;
  wire [3:0] __variable_wdata_144;
  wire [7:0] __variable_wdata_157;
  wire [7:0] __variable_wdata_158;
  wire [3:0] __variable_wdata_159;
  wire [7:0] __variable_wdata_172;
  wire [7:0] __variable_wdata_173;
  wire [3:0] __variable_wdata_174;
  wire [7:0] __variable_wdata_187;
  wire [7:0] __variable_wdata_188;
  wire [4:0] __variable_wdata_194;
  wire [1:0] __variable_wdata_195;
  wire [1:0] __variable_wdata_196;
  wire [8:0] __variable_wdata_197;
  wire [31:0] __variable_wdata_2;
  wire [31:0] __variable_wdata_20;
  wire [31:0] __variable_wdata_210;
  wire [7:0] __variable_wdata_217;
  wire [31:0] __variable_wdata_22;
  wire [7:0] __variable_wdata_224;
  wire [31:0] __variable_wdata_23;
  wire [7:0] __variable_wdata_231;
  wire [7:0] __variable_wdata_238;
  wire [31:0] __variable_wdata_24;
  wire __variable_wdata_244;
  wire __variable_wdata_245;
  wire [3:0] __variable_wdata_246;
  wire [7:0] __variable_wdata_248;
  wire [7:0] __variable_wdata_249;
  wire [31:0] __variable_wdata_25;
  wire [7:0] __variable_wdata_250;
  wire [7:0] __variable_wdata_251;
  wire [7:0] __variable_wdata_252;
  wire [7:0] __variable_wdata_253;
  wire [7:0] __variable_wdata_254;
  wire [7:0] __variable_wdata_255;
  wire [7:0] __variable_wdata_256;
  wire [31:0] __variable_wdata_26;
  wire [31:0] __variable_wdata_27;
  wire [31:0] __variable_wdata_28;
  wire [31:0] __variable_wdata_29;
  wire [31:0] __variable_wdata_30;
  wire [31:0] __variable_wdata_36;
  wire [7:0] __variable_wdata_37;
  wire [5:0] __variable_wdata_38;
  wire [7:0] __variable_wdata_482;
  wire [7:0] __variable_wdata_483;
  wire [7:0] __variable_wdata_484;
  wire [7:0] __variable_wdata_485;
  wire [7:0] __variable_wdata_486;
  wire [7:0] __variable_wdata_487;
  wire [7:0] __variable_wdata_488;
  wire [7:0] __variable_wdata_489;
  wire [7:0] __variable_wdata_490;
  wire [7:0] __variable_wdata_52;
  wire [7:0] __variable_wdata_53;
  wire [3:0] __variable_wdata_54;
  wire [7:0] __variable_wdata_67;
  wire [7:0] __variable_wdata_68;
  wire [3:0] __variable_wdata_69;
  wire [2:0] __variable_wdata_757;
  wire [7:0] __variable_wdata_758;
  wire [3:0] __variable_wdata_759;
  wire [8:0] __variable_wdata_776;
  wire __variable_wdata_777;
  wire __variable_wdata_778;
  wire __variable_wdata_779;
  wire [31:0] __variable_wdata_792;
  wire [7:0] __variable_wdata_799;
  wire [7:0] __variable_wdata_806;
  wire [7:0] __variable_wdata_813;
  wire [7:0] __variable_wdata_82;
  wire [7:0] __variable_wdata_820;
  wire __variable_wdata_826;
  wire __variable_wdata_827;
  wire [3:0] __variable_wdata_828;
  wire [7:0] __variable_wdata_83;
  wire [7:0] __variable_wdata_830;
  wire [3:0] __variable_wdata_84;
  wire [7:0] __variable_wdata_844;
  wire [7:0] __variable_wdata_97;
  wire [7:0] __variable_wdata_98;
  wire [3:0] __variable_wdata_99;
  wire _acc_0_reduce_reset;
  wire [15:0] _cond_data_108;
  wire [31:0] _cond_data_11;
  wire [15:0] _cond_data_123;
  wire [15:0] _cond_data_138;
  wire [15:0] _cond_data_153;
  wire [15:0] _cond_data_168;
  wire [15:0] _cond_data_183;
  wire [31:0] _cond_data_215;
  wire [7:0] _cond_data_222;
  wire [7:0] _cond_data_229;
  wire [7:0] _cond_data_236;
  wire [7:0] _cond_data_243;
  wire [7:0] _cond_data_259;
  wire [7:0] _cond_data_263;
  wire [7:0] _cond_data_266;
  wire [7:0] _cond_data_269;
  wire [7:0] _cond_data_273;
  wire [7:0] _cond_data_276;
  wire [7:0] _cond_data_279;
  wire [7:0] _cond_data_283;
  wire [7:0] _cond_data_286;
  wire [7:0] _cond_data_289;
  wire [7:0] _cond_data_293;
  wire [7:0] _cond_data_296;
  wire [7:0] _cond_data_299;
  wire [7:0] _cond_data_303;
  wire [7:0] _cond_data_306;
  wire [7:0] _cond_data_309;
  wire [7:0] _cond_data_313;
  wire [7:0] _cond_data_316;
  wire [7:0] _cond_data_319;
  wire [7:0] _cond_data_323;
  wire [7:0] _cond_data_326;
  wire [7:0] _cond_data_329;
  wire [7:0] _cond_data_333;
  wire [7:0] _cond_data_336;
  wire [7:0] _cond_data_339;
  wire [7:0] _cond_data_343;
  wire [7:0] _cond_data_346;
  wire [7:0] _cond_data_349;
  wire [7:0] _cond_data_353;
  wire [7:0] _cond_data_356;
  wire [7:0] _cond_data_359;
  wire [7:0] _cond_data_363;
  wire [7:0] _cond_data_366;
  wire [7:0] _cond_data_369;
  wire [7:0] _cond_data_373;
  wire [7:0] _cond_data_376;
  wire [7:0] _cond_data_379;
  wire [7:0] _cond_data_383;
  wire [7:0] _cond_data_386;
  wire [7:0] _cond_data_389;
  wire [7:0] _cond_data_393;
  wire [7:0] _cond_data_396;
  wire [7:0] _cond_data_399;
  wire [7:0] _cond_data_403;
  wire [7:0] _cond_data_406;
  wire [7:0] _cond_data_409;
  wire [7:0] _cond_data_413;
  wire [7:0] _cond_data_416;
  wire [7:0] _cond_data_419;
  wire [7:0] _cond_data_423;
  wire [7:0] _cond_data_426;
  wire [7:0] _cond_data_429;
  wire [39:0] _cond_data_43;
  wire [7:0] _cond_data_433;
  wire [7:0] _cond_data_436;
  wire [39:0] _cond_data_47;
  wire [7:0] _cond_data_51;
  wire [7:0] _cond_data_555;
  wire [7:0] _cond_data_557;
  wire [7:0] _cond_data_559;
  wire [7:0] _cond_data_561;
  wire [7:0] _cond_data_563;
  wire [7:0] _cond_data_565;
  wire [7:0] _cond_data_567;
  wire [7:0] _cond_data_569;
  wire [7:0] _cond_data_571;
  wire [15:0] _cond_data_63;
  wire [7:0] _cond_data_755;
  wire [8:0] _cond_data_771;
  wire [15:0] _cond_data_78;
  wire [31:0] _cond_data_797;
  wire [7:0] _cond_data_804;
  wire [7:0] _cond_data_811;
  wire [7:0] _cond_data_818;
  wire [7:0] _cond_data_825;
  wire [7:0] _cond_data_833;
  wire [7:0] _cond_data_837;
  wire [7:0] _cond_data_853;
  wire [15:0] _cond_data_93;
  wire _control_conv2d_8_cond_14_2_1;
  wire _control_conv2d_8_cond_15_3_1;
  wire _control_conv2d_8_cond_23_4_1;
  wire _control_conv2d_8_cond_24_5_1;
  wire _control_conv2d_8_cond_30_6_1;
  wire _control_conv2d_8_cond_31_7_1;
  wire _control_conv2d_8_cond_37_8_1;
  wire _control_conv2d_8_cond_38_9_1;
  wire _control_conv2d_8_cond_3_0_1;
  wire _control_conv2d_8_cond_48_10_1;
  wire _control_conv2d_8_cond_8_1_1;
  wire _control_matmul_15_cond_14_2_1;
  wire _control_matmul_15_cond_22_3_1;
  wire _control_matmul_15_cond_32_4_1;
  wire _control_matmul_15_cond_3_0_1;
  wire _control_matmul_15_cond_8_1_1;
  wire _control_max_pool_serial_9_cond_11_1_1;
  wire _control_max_pool_serial_9_cond_19_2_1;
  wire _control_max_pool_serial_9_cond_5_0_1;
  wire [3:0] _counter_count_762;
  wire [31:0] _counter_data_762;
  wire [31:0] _d1__maxi_read_fsm;
  wire [31:0] _d1__maxi_write_fsm;
  wire [31:0] _d1_control_conv2d_8;
  wire [31:0] _d1_control_matmul_15;
  wire [31:0] _d1_control_max_pool_serial_9;
  wire [31:0] _dataflow__delay_data_132;
  wire _dataflow__delay_valid_132;
  wire [31:0] _dataflow_cat_data_131;
  wire [31:0] _dataflow_cat_data_74;
  wire [31:0] _dataflow_cat_data_96;
  wire _dataflow_cat_valid_131;
  wire _dataflow_cat_valid_74;
  wire _dataflow_cat_valid_96;
  wire [7:0] _dataflow_slice_data_10;
  wire [7:0] _dataflow_slice_data_100;
  wire [7:0] _dataflow_slice_data_103;
  wire [7:0] _dataflow_slice_data_106;
  wire [7:0] _dataflow_slice_data_109;
  wire [7:0] _dataflow_slice_data_113;
  wire [7:0] _dataflow_slice_data_116;
  wire [7:0] _dataflow_slice_data_119;
  wire [7:0] _dataflow_slice_data_122;
  wire [7:0] _dataflow_slice_data_13;
  wire [7:0] _dataflow_slice_data_17;
  wire [7:0] _dataflow_slice_data_20;
  wire [7:0] _dataflow_slice_data_23;
  wire [7:0] _dataflow_slice_data_26;
  wire [7:0] _dataflow_slice_data_30;
  wire [7:0] _dataflow_slice_data_33;
  wire [7:0] _dataflow_slice_data_36;
  wire [7:0] _dataflow_slice_data_39;
  wire [7:0] _dataflow_slice_data_4;
  wire [7:0] _dataflow_slice_data_43;
  wire [7:0] _dataflow_slice_data_46;
  wire [7:0] _dataflow_slice_data_49;
  wire [7:0] _dataflow_slice_data_52;
  wire [7:0] _dataflow_slice_data_56;
  wire [7:0] _dataflow_slice_data_59;
  wire [7:0] _dataflow_slice_data_62;
  wire [7:0] _dataflow_slice_data_65;
  wire [7:0] _dataflow_slice_data_7;
  wire [7:0] _dataflow_slice_data_78;
  wire [7:0] _dataflow_slice_data_81;
  wire [7:0] _dataflow_slice_data_84;
  wire [7:0] _dataflow_slice_data_87;
  wire _dataflow_slice_valid_10;
  wire _dataflow_slice_valid_100;
  wire _dataflow_slice_valid_103;
  wire _dataflow_slice_valid_106;
  wire _dataflow_slice_valid_109;
  wire _dataflow_slice_valid_113;
  wire _dataflow_slice_valid_116;
  wire _dataflow_slice_valid_119;
  wire _dataflow_slice_valid_122;
  wire _dataflow_slice_valid_13;
  wire _dataflow_slice_valid_17;
  wire _dataflow_slice_valid_20;
  wire _dataflow_slice_valid_23;
  wire _dataflow_slice_valid_26;
  wire _dataflow_slice_valid_30;
  wire _dataflow_slice_valid_33;
  wire _dataflow_slice_valid_36;
  wire _dataflow_slice_valid_39;
  wire _dataflow_slice_valid_4;
  wire _dataflow_slice_valid_43;
  wire _dataflow_slice_valid_46;
  wire _dataflow_slice_valid_49;
  wire _dataflow_slice_valid_52;
  wire _dataflow_slice_valid_56;
  wire _dataflow_slice_valid_59;
  wire _dataflow_slice_valid_62;
  wire _dataflow_slice_valid_65;
  wire _dataflow_slice_valid_7;
  wire _dataflow_slice_valid_78;
  wire _dataflow_slice_valid_81;
  wire _dataflow_slice_valid_84;
  wire _dataflow_slice_valid_87;
  wire _eq_data_337;
  wire _eq_data_341;
  wire _eq_data_344;
  wire _eq_data_427;
  wire _eq_data_431;
  wire _eq_data_434;
  wire _eq_data_831;
  wire _eq_data_835;
  wire _greatereq_data_49;
  wire _greaterthan_data_100;
  wire _greaterthan_data_115;
  wire _greaterthan_data_130;
  wire _greaterthan_data_145;
  wire _greaterthan_data_160;
  wire _greaterthan_data_175;
  wire _greaterthan_data_3;
  wire _greaterthan_data_41;
  wire _greaterthan_data_55;
  wire _greaterthan_data_70;
  wire _greaterthan_data_753;
  wire _greaterthan_data_85;
  wire _lessthan_data_45;
  wire [31:0] _maxi_global_base_addr;
  wire [31:0] _maxi_ram_w32_l128_id0_1_read_global_addr;
  wire [31:0] _maxi_ram_w32_l128_id0_1_read_local_addr;
  wire [31:0] _maxi_ram_w32_l128_id0_1_read_local_stride;
  wire [7:0] _maxi_ram_w32_l128_id0_1_read_op_sel;
  wire [32:0] _maxi_ram_w32_l128_id0_1_read_size;
  wire _maxi_ram_w32_l128_id0_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id0_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id0_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id0_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id0_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id0_1_read_size;
  wire _maxi_ram_w8_l2048_id0_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id0_1_write_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id0_1_write_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id0_1_write_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id0_1_write_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id0_1_write_size;
  wire _maxi_ram_w8_l2048_id0_1_write_start;
  wire [31:0] _maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_size;
  wire _maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_size;
  wire _maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_size;
  wire _maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id19_1_write_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id19_1_write_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id19_1_write_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id19_1_write_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id19_1_write_size;
  wire _maxi_ram_w8_l2048_id19_1_write_start;
  wire [31:0] _maxi_ram_w8_l2048_id1_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id1_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id1_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id1_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id1_1_read_size;
  wire _maxi_ram_w8_l2048_id1_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id1_1_write_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id1_1_write_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id1_1_write_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id1_1_write_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id1_1_write_size;
  wire _maxi_ram_w8_l2048_id1_1_write_start;
  wire [31:0] _maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_size;
  wire _maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id2_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id2_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id2_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id2_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id2_1_read_size;
  wire _maxi_ram_w8_l2048_id2_1_read_start;
  wire [31:0] _maxi_ram_w8_l4096_id0_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l4096_id0_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l4096_id0_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l4096_id0_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l4096_id0_1_read_size;
  wire _maxi_ram_w8_l4096_id0_1_read_start;
  wire [31:0] _maxi_read_cur_global_addr;
  wire [32:0] _maxi_read_cur_size;
  wire [31:0] _maxi_read_fsm;
  wire [31:0] _maxi_read_global_addr;
  wire _maxi_read_idle;
  wire [31:0] _maxi_read_local_addr;
  wire [31:0] _maxi_read_local_stride;
  wire [7:0] _maxi_read_op_sel;
  wire [32:0] _maxi_read_rest_size;
  wire [32:0] _maxi_read_size;
  wire _maxi_read_start;
  wire [31:0] _maxi_write_cur_global_addr;
  wire [32:0] _maxi_write_cur_size;
  wire _maxi_write_data_done;
  wire [31:0] _maxi_write_fsm;
  wire [31:0] _maxi_write_global_addr;
  wire _maxi_write_idle;
  wire [31:0] _maxi_write_local_addr;
  wire [31:0] _maxi_write_local_stride;
  wire [7:0] _maxi_write_op_sel;
  wire [32:0] _maxi_write_rest_size;
  wire [32:0] _maxi_write_size;
  wire _maxi_write_start;
  wire [3:0] _minus_data_102;
  wire [3:0] _minus_data_117;
  wire [3:0] _minus_data_132;
  wire [3:0] _minus_data_147;
  wire [3:0] _minus_data_162;
  wire [3:0] _minus_data_177;
  wire [5:0] _minus_data_5;
  wire [3:0] _minus_data_57;
  wire [3:0] _minus_data_72;
  wire [3:0] _minus_data_87;
  wire [31:0] _plus_data_18;
  wire [7:0] _plus_data_723;
  wire [7:0] _plus_data_739;
  wire [31:0] _plus_data_742;
  wire [7:0] _plus_data_750;
  wire [7:0] _plus_data_855;
  wire [7:0] _plus_data_860;
  wire [31:0] _plus_data_863;
  wire [7:0] _plus_data_865;
  wire _pointer_data_536;
  wire _pointer_data_538;
  wire _pointer_data_540;
  wire _pointer_data_542;
  wire _pointer_data_544;
  wire _pointer_data_546;
  wire _pointer_data_548;
  wire _pointer_data_550;
  wire _pointer_data_552;
  wire _pointer_data_764;
  wire _pointer_data_850;
  wire [32:0] _pulse_count_17;
  wire [8:0] _pulse_count_193;
  wire _pulse_data_17;
  wire _pulse_data_193;
  wire _ram_w32_l128_id0_cond_2_1;
  wire _ram_w32_l128_id0_cond_4_1;
  wire _ram_w8_l2048_id0_0_cond_3_1;
  wire _ram_w8_l2048_id0_1_cond_3_1;
  wire _ram_w8_l2048_id0_2_cond_3_1;
  wire _ram_w8_l2048_id0_3_cond_1_1;
  wire _ram_w8_l2048_id0_3_cond_3_1;
  wire _ram_w8_l2048_id0_3_cond_4_1;
  wire _ram_w8_l2048_id10_0_cond_3_1;
  wire _ram_w8_l2048_id11_0_cond_2_1;
  wire _ram_w8_l2048_id12_0_cond_2_1;
  wire _ram_w8_l2048_id13_0_cond_3_1;
  wire _ram_w8_l2048_id14_0_cond_2_1;
  wire _ram_w8_l2048_id15_0_cond_2_1;
  wire _ram_w8_l2048_id16_0_cond_3_1;
  wire _ram_w8_l2048_id17_0_cond_2_1;
  wire _ram_w8_l2048_id18_0_cond_2_1;
  wire _ram_w8_l2048_id19_0_cond_0_1;
  wire _ram_w8_l2048_id19_1_cond_0_1;
  wire _ram_w8_l2048_id19_2_cond_0_1;
  wire _ram_w8_l2048_id19_3_cond_0_1;
  wire _ram_w8_l2048_id1_0_cond_7_1;
  wire _ram_w8_l2048_id1_1_cond_7_1;
  wire _ram_w8_l2048_id1_2_cond_7_1;
  wire _ram_w8_l2048_id1_3_cond_2_1;
  wire _ram_w8_l2048_id1_3_cond_5_1;
  wire _ram_w8_l2048_id1_3_cond_7_1;
  wire _ram_w8_l2048_id2_3_cond_1_1;
  wire _ram_w8_l2048_id2_3_cond_4_1;
  wire _ram_w8_l2048_id3_3_cond_1_1;
  wire _ram_w8_l2048_id4_3_cond_1_1;
  wire _ram_w8_l2048_id5_3_cond_1_1;
  wire _ram_w8_l2048_id6_3_cond_1_1;
  wire _ram_w8_l2048_id7_3_cond_1_1;
  wire _ram_w8_l2048_id8_3_cond_1_1;
  wire _ram_w8_l2048_id9_0_cond_1_1;
  wire _ram_w8_l2048_id9_2_cond_0_1;
  wire _ram_w8_l4096_id0_3_cond_1_1;
  wire [32:0] _reduceadd_count_15;
  wire [31:0] _reduceadd_data_15;
  wire [8:0] _reducecustom_count_191;
  wire [31:0] _reducecustom_data_191;
  wire _rst_logic_1;
  wire _rst_logic_2;
  wire _saxi_cond_0_1;
  wire _saxi_flag_0;
  wire _saxi_flag_1;
  wire _saxi_flag_10;
  wire _saxi_flag_11;
  wire _saxi_flag_12;
  wire _saxi_flag_13;
  wire _saxi_flag_2;
  wire _saxi_flag_3;
  wire _saxi_flag_4;
  wire _saxi_flag_5;
  wire _saxi_flag_6;
  wire _saxi_flag_7;
  wire _saxi_flag_8;
  wire _saxi_flag_9;
  wire [31:0] _saxi_register_0;
  wire [31:0] _saxi_register_1;
  wire [31:0] _saxi_register_10;
  wire [31:0] _saxi_register_11;
  wire [31:0] _saxi_register_12;
  wire [31:0] _saxi_register_13;
  wire [31:0] _saxi_register_2;
  wire [31:0] _saxi_register_3;
  wire [31:0] _saxi_register_4;
  wire [31:0] _saxi_register_5;
  wire [31:0] _saxi_register_6;
  wire [31:0] _saxi_register_7;
  wire [31:0] _saxi_register_8;
  wire [31:0] _saxi_register_9;
  wire [31:0] _saxi_register_fsm;
  wire [31:0] _saxi_resetval_0;
  wire [31:0] _saxi_resetval_1;
  wire [31:0] _saxi_resetval_10;
  wire [31:0] _saxi_resetval_11;
  wire [31:0] _saxi_resetval_12;
  wire [31:0] _saxi_resetval_13;
  wire [31:0] _saxi_resetval_2;
  wire [31:0] _saxi_resetval_3;
  wire [31:0] _saxi_resetval_4;
  wire [31:0] _saxi_resetval_5;
  wire [31:0] _saxi_resetval_6;
  wire [31:0] _saxi_resetval_7;
  wire [31:0] _saxi_resetval_8;
  wire [31:0] _saxi_resetval_9;
  wire _set_flag_1034;
  wire _set_flag_538;
  wire _set_flag_874;
  wire _set_flag_876;
  wire [17:0] _sll_data_104;
  wire [17:0] _sll_data_119;
  wire [17:0] _sll_data_134;
  wire [17:0] _sll_data_149;
  wire [17:0] _sll_data_164;
  wire [17:0] _sll_data_179;
  wire [17:0] _sll_data_59;
  wire [65:0] _sll_data_7;
  wire [17:0] _sll_data_74;
  wire [17:0] _sll_data_89;
  wire [32:0] _source_stream_conv2d_8_source_19_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_19_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_19_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_19_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_19_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_19_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_19_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_19_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_19_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_19_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_19_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_19_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_19_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_19_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_19_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_19_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_19_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_19_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_19_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_19_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_19_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_19_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_19_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_19_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_20_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_20_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_20_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_20_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_20_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_20_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_20_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_20_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_20_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_20_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_20_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_20_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_20_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_20_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_20_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_20_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_20_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_20_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_20_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_20_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_20_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_20_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_20_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_20_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_21_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_21_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_21_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_21_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_21_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_21_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_21_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_21_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_21_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_21_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_21_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_21_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_21_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_21_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_21_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_21_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_21_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_21_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_21_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_21_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_21_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_21_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_21_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_21_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_22_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_22_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_22_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_22_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_22_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_22_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_22_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_22_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_22_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_22_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_22_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_22_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_22_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_22_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_22_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_22_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_22_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_22_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_22_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_22_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_22_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_22_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_22_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_22_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_23_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_23_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_23_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_23_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_23_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_23_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_23_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_23_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_23_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_23_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_23_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_23_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_23_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_23_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_23_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_23_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_23_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_23_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_23_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_23_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_23_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_23_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_23_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_23_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_24_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_24_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_24_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_24_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_24_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_24_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_24_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_24_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_24_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_24_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_24_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_24_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_24_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_24_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_24_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_24_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_24_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_24_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_24_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_24_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_24_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_24_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_24_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_24_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_25_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_25_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_25_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_25_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_25_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_25_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_25_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_25_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_25_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_25_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_25_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_25_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_25_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_25_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_25_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_25_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_25_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_25_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_25_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_25_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_25_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_25_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_25_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_25_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_26_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_26_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_26_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_26_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_26_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_26_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_26_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_26_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_26_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_26_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_26_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_26_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_26_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_26_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_26_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_26_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_26_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_26_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_26_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_26_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_26_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_26_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_26_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_26_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_27_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_27_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_27_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_27_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_27_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_27_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_27_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_27_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_27_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_27_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_27_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_27_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_27_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_27_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_27_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_27_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_27_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_27_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_27_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_27_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_27_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_27_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_27_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_27_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_28_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_28_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_28_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_28_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_28_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_28_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_28_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_28_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_28_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_28_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_28_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_28_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_28_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_28_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_28_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_28_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_28_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_28_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_28_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_28_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_28_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_28_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_28_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_28_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_29_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_29_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_29_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_29_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_29_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_29_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_29_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_29_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_29_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_29_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_29_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_29_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_29_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_29_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_29_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_29_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_29_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_29_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_29_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_29_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_29_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_29_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_29_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_29_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_30_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_30_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_30_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_30_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_30_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_30_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_30_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_30_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_30_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_30_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_30_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_30_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_30_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_30_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_30_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_30_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_30_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_30_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_30_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_30_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_30_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_30_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_30_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_30_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_31_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_31_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_31_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_31_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_31_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_31_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_31_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_31_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_31_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_31_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_31_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_31_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_31_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_31_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_31_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_31_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_31_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_31_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_31_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_31_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_31_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_31_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_31_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_31_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_32_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_32_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_32_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_32_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_32_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_32_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_32_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_32_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_32_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_32_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_32_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_32_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_32_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_32_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_32_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_32_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_32_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_32_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_32_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_32_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_32_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_32_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_32_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_32_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_33_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_33_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_33_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_33_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_33_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_33_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_33_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_33_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_33_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_33_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_33_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_33_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_33_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_33_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_33_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_33_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_33_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_33_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_33_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_33_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_33_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_33_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_33_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_33_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_34_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_34_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_34_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_34_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_34_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_34_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_34_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_34_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_34_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_34_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_34_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_34_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_34_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_34_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_34_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_34_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_34_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_34_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_34_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_34_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_34_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_34_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_34_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_34_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_35_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_35_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_35_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_35_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_35_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_35_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_35_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_35_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_35_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_35_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_35_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_35_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_35_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_35_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_35_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_35_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_35_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_35_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_35_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_35_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_35_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_35_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_35_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_35_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_36_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_36_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_36_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_36_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_36_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_36_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_36_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_36_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_36_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_36_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_36_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_36_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_36_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_36_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_36_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_36_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_36_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_36_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_36_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_36_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_36_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_36_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_36_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_36_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_6_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_6_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_6_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_6_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_6_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_6_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_6_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_6_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_6_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_6_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_6_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_6_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_6_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_6_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_6_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_6_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_6_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_6_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_6_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_6_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_6_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_6_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_6_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_6_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_8_source_8_pat_count_0;
  wire [32:0] _source_stream_conv2d_8_source_8_pat_count_1;
  wire [32:0] _source_stream_conv2d_8_source_8_pat_count_2;
  wire [32:0] _source_stream_conv2d_8_source_8_pat_count_3;
  wire [31:0] _source_stream_conv2d_8_source_8_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_8_source_8_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_8_source_8_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_8_source_8_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_8_source_8_pat_size_0;
  wire [32:0] _source_stream_conv2d_8_source_8_pat_size_1;
  wire [32:0] _source_stream_conv2d_8_source_8_pat_size_2;
  wire [32:0] _source_stream_conv2d_8_source_8_pat_size_3;
  wire [32:0] _source_stream_conv2d_8_source_8_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_8_source_8_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_8_source_8_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_8_source_8_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_8_source_8_pat_stride_0;
  wire [31:0] _source_stream_conv2d_8_source_8_pat_stride_1;
  wire [31:0] _source_stream_conv2d_8_source_8_pat_stride_2;
  wire [31:0] _source_stream_conv2d_8_source_8_pat_stride_3;
  wire [31:0] _source_stream_conv2d_8_source_8_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_8_source_8_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_8_source_8_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_8_source_8_pat_stride_buf_3;
  wire [32:0] _source_stream_matmul_15_source_19_pat_count_0;
  wire [32:0] _source_stream_matmul_15_source_19_pat_count_1;
  wire [32:0] _source_stream_matmul_15_source_19_pat_count_2;
  wire [32:0] _source_stream_matmul_15_source_19_pat_count_3;
  wire [31:0] _source_stream_matmul_15_source_19_pat_cur_offset_0;
  wire [31:0] _source_stream_matmul_15_source_19_pat_cur_offset_1;
  wire [31:0] _source_stream_matmul_15_source_19_pat_cur_offset_2;
  wire [31:0] _source_stream_matmul_15_source_19_pat_cur_offset_3;
  wire [32:0] _source_stream_matmul_15_source_19_pat_size_0;
  wire [32:0] _source_stream_matmul_15_source_19_pat_size_1;
  wire [32:0] _source_stream_matmul_15_source_19_pat_size_2;
  wire [32:0] _source_stream_matmul_15_source_19_pat_size_3;
  wire [32:0] _source_stream_matmul_15_source_19_pat_size_buf_0;
  wire [32:0] _source_stream_matmul_15_source_19_pat_size_buf_1;
  wire [32:0] _source_stream_matmul_15_source_19_pat_size_buf_2;
  wire [32:0] _source_stream_matmul_15_source_19_pat_size_buf_3;
  wire [31:0] _source_stream_matmul_15_source_19_pat_stride_0;
  wire [31:0] _source_stream_matmul_15_source_19_pat_stride_1;
  wire [31:0] _source_stream_matmul_15_source_19_pat_stride_2;
  wire [31:0] _source_stream_matmul_15_source_19_pat_stride_3;
  wire [31:0] _source_stream_matmul_15_source_19_pat_stride_buf_0;
  wire [31:0] _source_stream_matmul_15_source_19_pat_stride_buf_1;
  wire [31:0] _source_stream_matmul_15_source_19_pat_stride_buf_2;
  wire [31:0] _source_stream_matmul_15_source_19_pat_stride_buf_3;
  wire [32:0] _source_stream_matmul_15_source_20_pat_count_0;
  wire [32:0] _source_stream_matmul_15_source_20_pat_count_1;
  wire [32:0] _source_stream_matmul_15_source_20_pat_count_2;
  wire [32:0] _source_stream_matmul_15_source_20_pat_count_3;
  wire [31:0] _source_stream_matmul_15_source_20_pat_cur_offset_0;
  wire [31:0] _source_stream_matmul_15_source_20_pat_cur_offset_1;
  wire [31:0] _source_stream_matmul_15_source_20_pat_cur_offset_2;
  wire [31:0] _source_stream_matmul_15_source_20_pat_cur_offset_3;
  wire [32:0] _source_stream_matmul_15_source_20_pat_size_0;
  wire [32:0] _source_stream_matmul_15_source_20_pat_size_1;
  wire [32:0] _source_stream_matmul_15_source_20_pat_size_2;
  wire [32:0] _source_stream_matmul_15_source_20_pat_size_3;
  wire [32:0] _source_stream_matmul_15_source_20_pat_size_buf_0;
  wire [32:0] _source_stream_matmul_15_source_20_pat_size_buf_1;
  wire [32:0] _source_stream_matmul_15_source_20_pat_size_buf_2;
  wire [32:0] _source_stream_matmul_15_source_20_pat_size_buf_3;
  wire [31:0] _source_stream_matmul_15_source_20_pat_stride_0;
  wire [31:0] _source_stream_matmul_15_source_20_pat_stride_1;
  wire [31:0] _source_stream_matmul_15_source_20_pat_stride_2;
  wire [31:0] _source_stream_matmul_15_source_20_pat_stride_3;
  wire [31:0] _source_stream_matmul_15_source_20_pat_stride_buf_0;
  wire [31:0] _source_stream_matmul_15_source_20_pat_stride_buf_1;
  wire [31:0] _source_stream_matmul_15_source_20_pat_stride_buf_2;
  wire [31:0] _source_stream_matmul_15_source_20_pat_stride_buf_3;
  wire [32:0] _source_stream_matmul_15_source_6_pat_count_0;
  wire [32:0] _source_stream_matmul_15_source_6_pat_count_1;
  wire [32:0] _source_stream_matmul_15_source_6_pat_count_2;
  wire [32:0] _source_stream_matmul_15_source_6_pat_count_3;
  wire [31:0] _source_stream_matmul_15_source_6_pat_cur_offset_0;
  wire [31:0] _source_stream_matmul_15_source_6_pat_cur_offset_1;
  wire [31:0] _source_stream_matmul_15_source_6_pat_cur_offset_2;
  wire [31:0] _source_stream_matmul_15_source_6_pat_cur_offset_3;
  wire [32:0] _source_stream_matmul_15_source_6_pat_size_0;
  wire [32:0] _source_stream_matmul_15_source_6_pat_size_1;
  wire [32:0] _source_stream_matmul_15_source_6_pat_size_2;
  wire [32:0] _source_stream_matmul_15_source_6_pat_size_3;
  wire [32:0] _source_stream_matmul_15_source_6_pat_size_buf_0;
  wire [32:0] _source_stream_matmul_15_source_6_pat_size_buf_1;
  wire [32:0] _source_stream_matmul_15_source_6_pat_size_buf_2;
  wire [32:0] _source_stream_matmul_15_source_6_pat_size_buf_3;
  wire [31:0] _source_stream_matmul_15_source_6_pat_stride_0;
  wire [31:0] _source_stream_matmul_15_source_6_pat_stride_1;
  wire [31:0] _source_stream_matmul_15_source_6_pat_stride_2;
  wire [31:0] _source_stream_matmul_15_source_6_pat_stride_3;
  wire [31:0] _source_stream_matmul_15_source_6_pat_stride_buf_0;
  wire [31:0] _source_stream_matmul_15_source_6_pat_stride_buf_1;
  wire [31:0] _source_stream_matmul_15_source_6_pat_stride_buf_2;
  wire [31:0] _source_stream_matmul_15_source_6_pat_stride_buf_3;
  wire [32:0] _source_stream_matmul_15_source_8_pat_count_0;
  wire [32:0] _source_stream_matmul_15_source_8_pat_count_1;
  wire [32:0] _source_stream_matmul_15_source_8_pat_count_2;
  wire [32:0] _source_stream_matmul_15_source_8_pat_count_3;
  wire [31:0] _source_stream_matmul_15_source_8_pat_cur_offset_0;
  wire [31:0] _source_stream_matmul_15_source_8_pat_cur_offset_1;
  wire [31:0] _source_stream_matmul_15_source_8_pat_cur_offset_2;
  wire [31:0] _source_stream_matmul_15_source_8_pat_cur_offset_3;
  wire [32:0] _source_stream_matmul_15_source_8_pat_size_0;
  wire [32:0] _source_stream_matmul_15_source_8_pat_size_1;
  wire [32:0] _source_stream_matmul_15_source_8_pat_size_2;
  wire [32:0] _source_stream_matmul_15_source_8_pat_size_3;
  wire [32:0] _source_stream_matmul_15_source_8_pat_size_buf_0;
  wire [32:0] _source_stream_matmul_15_source_8_pat_size_buf_1;
  wire [32:0] _source_stream_matmul_15_source_8_pat_size_buf_2;
  wire [32:0] _source_stream_matmul_15_source_8_pat_size_buf_3;
  wire [31:0] _source_stream_matmul_15_source_8_pat_stride_0;
  wire [31:0] _source_stream_matmul_15_source_8_pat_stride_1;
  wire [31:0] _source_stream_matmul_15_source_8_pat_stride_2;
  wire [31:0] _source_stream_matmul_15_source_8_pat_stride_3;
  wire [31:0] _source_stream_matmul_15_source_8_pat_stride_buf_0;
  wire [31:0] _source_stream_matmul_15_source_8_pat_stride_buf_1;
  wire [31:0] _source_stream_matmul_15_source_8_pat_stride_buf_2;
  wire [31:0] _source_stream_matmul_15_source_8_pat_stride_buf_3;
  wire [32:0] _source_stream_max_pool_serial_9_source_1_pat_count_0;
  wire [32:0] _source_stream_max_pool_serial_9_source_1_pat_count_1;
  wire [32:0] _source_stream_max_pool_serial_9_source_1_pat_count_2;
  wire [32:0] _source_stream_max_pool_serial_9_source_1_pat_count_3;
  wire [31:0] _source_stream_max_pool_serial_9_source_1_pat_cur_offset_0;
  wire [31:0] _source_stream_max_pool_serial_9_source_1_pat_cur_offset_1;
  wire [31:0] _source_stream_max_pool_serial_9_source_1_pat_cur_offset_2;
  wire [31:0] _source_stream_max_pool_serial_9_source_1_pat_cur_offset_3;
  wire [32:0] _source_stream_max_pool_serial_9_source_1_pat_size_0;
  wire [32:0] _source_stream_max_pool_serial_9_source_1_pat_size_1;
  wire [32:0] _source_stream_max_pool_serial_9_source_1_pat_size_2;
  wire [32:0] _source_stream_max_pool_serial_9_source_1_pat_size_3;
  wire [32:0] _source_stream_max_pool_serial_9_source_1_pat_size_buf_0;
  wire [32:0] _source_stream_max_pool_serial_9_source_1_pat_size_buf_1;
  wire [32:0] _source_stream_max_pool_serial_9_source_1_pat_size_buf_2;
  wire [32:0] _source_stream_max_pool_serial_9_source_1_pat_size_buf_3;
  wire [31:0] _source_stream_max_pool_serial_9_source_1_pat_stride_0;
  wire [31:0] _source_stream_max_pool_serial_9_source_1_pat_stride_1;
  wire [31:0] _source_stream_max_pool_serial_9_source_1_pat_stride_2;
  wire [31:0] _source_stream_max_pool_serial_9_source_1_pat_stride_3;
  wire [31:0] _source_stream_max_pool_serial_9_source_1_pat_stride_buf_0;
  wire [31:0] _source_stream_max_pool_serial_9_source_1_pat_stride_buf_1;
  wire [31:0] _source_stream_max_pool_serial_9_source_1_pat_stride_buf_2;
  wire [31:0] _source_stream_max_pool_serial_9_source_1_pat_stride_buf_3;
  wire [15:0] _sra_data_111;
  wire [15:0] _sra_data_126;
  wire [15:0] _sra_data_141;
  wire [15:0] _sra_data_156;
  wire [15:0] _sra_data_171;
  wire [15:0] _sra_data_186;
  wire [31:0] _sra_data_19;
  wire [39:0] _sra_data_40;
  wire [15:0] _sra_data_66;
  wire [15:0] _sra_data_81;
  wire [15:0] _sra_data_96;
  wire [4:0] _stream_conv2d_8_constant_0_next_constant_data;
  wire _stream_conv2d_8_constant_15_next_constant_data;
  wire _stream_conv2d_8_constant_16_next_constant_data;
  wire [3:0] _stream_conv2d_8_constant_17_next_constant_data;
  wire [1:0] _stream_conv2d_8_constant_1_next_constant_data;
  wire [1:0] _stream_conv2d_8_constant_2_next_constant_data;
  wire [8:0] _stream_conv2d_8_constant_3_next_constant_data;
  wire _stream_conv2d_8_done;
  wire _stream_conv2d_8_end_flag;
  wire [31:0] _stream_conv2d_8_fsm;
  wire [32:0] _stream_conv2d_8_sink_37_sink_count;
  wire [31:0] _stream_conv2d_8_sink_37_sink_fsm_20;
  wire [2:0] _stream_conv2d_8_sink_37_sink_mode;
  wire [31:0] _stream_conv2d_8_sink_37_sink_offset;
  wire [7:0] _stream_conv2d_8_sink_37_sink_ram_sel;
  wire [32:0] _stream_conv2d_8_sink_37_sink_size;
  wire [31:0] _stream_conv2d_8_sink_37_sink_stride;
  wire [31:0] _stream_conv2d_8_sink_37_sink_stride_buf;
  wire [31:0] _stream_conv2d_8_sink_37_sink_waddr;
  wire [7:0] _stream_conv2d_8_sink_37_sink_wdata;
  wire _stream_conv2d_8_sink_37_sink_wenable;
  wire _stream_conv2d_8_source_10_idle;
  wire [7:0] _stream_conv2d_8_source_10_source_empty_data;
  wire _stream_conv2d_8_source_12_idle;
  wire [7:0] _stream_conv2d_8_source_12_source_empty_data;
  wire _stream_conv2d_8_source_14_idle;
  wire [7:0] _stream_conv2d_8_source_14_source_empty_data;
  wire _stream_conv2d_8_source_19_idle;
  wire [2:0] _stream_conv2d_8_source_19_source_mode;
  wire [31:0] _stream_conv2d_8_source_19_source_offset;
  wire [31:0] _stream_conv2d_8_source_19_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_19_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_19_source_pat_fsm_2;
  wire [31:0] _stream_conv2d_8_source_19_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_19_source_ram_rdata;
  wire _stream_conv2d_8_source_19_source_ram_renable;
  wire _stream_conv2d_8_source_19_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_19_source_ram_sel;
  wire _stream_conv2d_8_source_20_idle;
  wire [2:0] _stream_conv2d_8_source_20_source_mode;
  wire [31:0] _stream_conv2d_8_source_20_source_offset;
  wire [31:0] _stream_conv2d_8_source_20_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_20_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_20_source_pat_fsm_3;
  wire [31:0] _stream_conv2d_8_source_20_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_20_source_ram_rdata;
  wire _stream_conv2d_8_source_20_source_ram_renable;
  wire _stream_conv2d_8_source_20_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_20_source_ram_sel;
  wire _stream_conv2d_8_source_21_idle;
  wire [2:0] _stream_conv2d_8_source_21_source_mode;
  wire [31:0] _stream_conv2d_8_source_21_source_offset;
  wire [31:0] _stream_conv2d_8_source_21_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_21_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_21_source_pat_fsm_4;
  wire [31:0] _stream_conv2d_8_source_21_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_21_source_ram_rdata;
  wire _stream_conv2d_8_source_21_source_ram_renable;
  wire _stream_conv2d_8_source_21_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_21_source_ram_sel;
  wire _stream_conv2d_8_source_22_idle;
  wire [2:0] _stream_conv2d_8_source_22_source_mode;
  wire [31:0] _stream_conv2d_8_source_22_source_offset;
  wire [31:0] _stream_conv2d_8_source_22_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_22_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_22_source_pat_fsm_5;
  wire [31:0] _stream_conv2d_8_source_22_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_22_source_ram_rdata;
  wire _stream_conv2d_8_source_22_source_ram_renable;
  wire _stream_conv2d_8_source_22_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_22_source_ram_sel;
  wire _stream_conv2d_8_source_23_idle;
  wire [2:0] _stream_conv2d_8_source_23_source_mode;
  wire [31:0] _stream_conv2d_8_source_23_source_offset;
  wire [31:0] _stream_conv2d_8_source_23_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_23_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_23_source_pat_fsm_6;
  wire [31:0] _stream_conv2d_8_source_23_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_23_source_ram_rdata;
  wire _stream_conv2d_8_source_23_source_ram_renable;
  wire _stream_conv2d_8_source_23_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_23_source_ram_sel;
  wire _stream_conv2d_8_source_24_idle;
  wire [2:0] _stream_conv2d_8_source_24_source_mode;
  wire [31:0] _stream_conv2d_8_source_24_source_offset;
  wire [31:0] _stream_conv2d_8_source_24_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_24_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_24_source_pat_fsm_7;
  wire [31:0] _stream_conv2d_8_source_24_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_24_source_ram_rdata;
  wire _stream_conv2d_8_source_24_source_ram_renable;
  wire _stream_conv2d_8_source_24_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_24_source_ram_sel;
  wire _stream_conv2d_8_source_25_idle;
  wire [2:0] _stream_conv2d_8_source_25_source_mode;
  wire [31:0] _stream_conv2d_8_source_25_source_offset;
  wire [31:0] _stream_conv2d_8_source_25_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_25_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_25_source_pat_fsm_8;
  wire [31:0] _stream_conv2d_8_source_25_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_25_source_ram_rdata;
  wire _stream_conv2d_8_source_25_source_ram_renable;
  wire _stream_conv2d_8_source_25_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_25_source_ram_sel;
  wire _stream_conv2d_8_source_26_idle;
  wire [2:0] _stream_conv2d_8_source_26_source_mode;
  wire [31:0] _stream_conv2d_8_source_26_source_offset;
  wire [31:0] _stream_conv2d_8_source_26_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_26_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_26_source_pat_fsm_9;
  wire [31:0] _stream_conv2d_8_source_26_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_26_source_ram_rdata;
  wire _stream_conv2d_8_source_26_source_ram_renable;
  wire _stream_conv2d_8_source_26_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_26_source_ram_sel;
  wire _stream_conv2d_8_source_27_idle;
  wire [2:0] _stream_conv2d_8_source_27_source_mode;
  wire [31:0] _stream_conv2d_8_source_27_source_offset;
  wire [31:0] _stream_conv2d_8_source_27_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_27_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_27_source_pat_fsm_10;
  wire [31:0] _stream_conv2d_8_source_27_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_27_source_ram_rdata;
  wire _stream_conv2d_8_source_27_source_ram_renable;
  wire _stream_conv2d_8_source_27_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_27_source_ram_sel;
  wire _stream_conv2d_8_source_28_idle;
  wire [2:0] _stream_conv2d_8_source_28_source_mode;
  wire [31:0] _stream_conv2d_8_source_28_source_offset;
  wire [31:0] _stream_conv2d_8_source_28_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_28_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_28_source_pat_fsm_11;
  wire [31:0] _stream_conv2d_8_source_28_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_28_source_ram_rdata;
  wire _stream_conv2d_8_source_28_source_ram_renable;
  wire _stream_conv2d_8_source_28_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_28_source_ram_sel;
  wire _stream_conv2d_8_source_29_idle;
  wire [2:0] _stream_conv2d_8_source_29_source_mode;
  wire [31:0] _stream_conv2d_8_source_29_source_offset;
  wire [31:0] _stream_conv2d_8_source_29_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_29_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_29_source_pat_fsm_12;
  wire [31:0] _stream_conv2d_8_source_29_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_29_source_ram_rdata;
  wire _stream_conv2d_8_source_29_source_ram_renable;
  wire _stream_conv2d_8_source_29_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_29_source_ram_sel;
  wire _stream_conv2d_8_source_30_idle;
  wire [2:0] _stream_conv2d_8_source_30_source_mode;
  wire [31:0] _stream_conv2d_8_source_30_source_offset;
  wire [31:0] _stream_conv2d_8_source_30_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_30_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_30_source_pat_fsm_13;
  wire [31:0] _stream_conv2d_8_source_30_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_30_source_ram_rdata;
  wire _stream_conv2d_8_source_30_source_ram_renable;
  wire _stream_conv2d_8_source_30_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_30_source_ram_sel;
  wire _stream_conv2d_8_source_31_idle;
  wire [2:0] _stream_conv2d_8_source_31_source_mode;
  wire [31:0] _stream_conv2d_8_source_31_source_offset;
  wire [31:0] _stream_conv2d_8_source_31_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_31_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_31_source_pat_fsm_14;
  wire [31:0] _stream_conv2d_8_source_31_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_31_source_ram_rdata;
  wire _stream_conv2d_8_source_31_source_ram_renable;
  wire _stream_conv2d_8_source_31_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_31_source_ram_sel;
  wire _stream_conv2d_8_source_32_idle;
  wire [2:0] _stream_conv2d_8_source_32_source_mode;
  wire [31:0] _stream_conv2d_8_source_32_source_offset;
  wire [31:0] _stream_conv2d_8_source_32_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_32_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_32_source_pat_fsm_15;
  wire [31:0] _stream_conv2d_8_source_32_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_32_source_ram_rdata;
  wire _stream_conv2d_8_source_32_source_ram_renable;
  wire _stream_conv2d_8_source_32_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_32_source_ram_sel;
  wire _stream_conv2d_8_source_33_idle;
  wire [2:0] _stream_conv2d_8_source_33_source_mode;
  wire [31:0] _stream_conv2d_8_source_33_source_offset;
  wire [31:0] _stream_conv2d_8_source_33_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_33_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_33_source_pat_fsm_16;
  wire [31:0] _stream_conv2d_8_source_33_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_33_source_ram_rdata;
  wire _stream_conv2d_8_source_33_source_ram_renable;
  wire _stream_conv2d_8_source_33_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_33_source_ram_sel;
  wire _stream_conv2d_8_source_34_idle;
  wire [2:0] _stream_conv2d_8_source_34_source_mode;
  wire [31:0] _stream_conv2d_8_source_34_source_offset;
  wire [31:0] _stream_conv2d_8_source_34_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_34_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_34_source_pat_fsm_17;
  wire [31:0] _stream_conv2d_8_source_34_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_34_source_ram_rdata;
  wire _stream_conv2d_8_source_34_source_ram_renable;
  wire _stream_conv2d_8_source_34_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_34_source_ram_sel;
  wire _stream_conv2d_8_source_35_idle;
  wire [2:0] _stream_conv2d_8_source_35_source_mode;
  wire [31:0] _stream_conv2d_8_source_35_source_offset;
  wire [31:0] _stream_conv2d_8_source_35_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_35_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_35_source_pat_fsm_18;
  wire [31:0] _stream_conv2d_8_source_35_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_35_source_ram_rdata;
  wire _stream_conv2d_8_source_35_source_ram_renable;
  wire _stream_conv2d_8_source_35_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_35_source_ram_sel;
  wire _stream_conv2d_8_source_36_idle;
  wire [2:0] _stream_conv2d_8_source_36_source_mode;
  wire [31:0] _stream_conv2d_8_source_36_source_offset;
  wire [31:0] _stream_conv2d_8_source_36_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_36_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_36_source_pat_fsm_19;
  wire [31:0] _stream_conv2d_8_source_36_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_36_source_ram_rdata;
  wire _stream_conv2d_8_source_36_source_ram_renable;
  wire _stream_conv2d_8_source_36_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_36_source_ram_sel;
  wire _stream_conv2d_8_source_6_idle;
  wire [2:0] _stream_conv2d_8_source_6_source_mode;
  wire [31:0] _stream_conv2d_8_source_6_source_offset;
  wire [31:0] _stream_conv2d_8_source_6_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_6_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_6_source_pat_fsm_0;
  wire [31:0] _stream_conv2d_8_source_6_source_ram_raddr;
  wire [31:0] _stream_conv2d_8_source_6_source_ram_rdata;
  wire _stream_conv2d_8_source_6_source_ram_renable;
  wire _stream_conv2d_8_source_6_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_6_source_ram_sel;
  wire _stream_conv2d_8_source_8_idle;
  wire [2:0] _stream_conv2d_8_source_8_source_mode;
  wire [31:0] _stream_conv2d_8_source_8_source_offset;
  wire [31:0] _stream_conv2d_8_source_8_source_offset_buf;
  wire [31:0] _stream_conv2d_8_source_8_source_pat_all_offset;
  wire [31:0] _stream_conv2d_8_source_8_source_pat_fsm_1;
  wire [31:0] _stream_conv2d_8_source_8_source_ram_raddr;
  wire [7:0] _stream_conv2d_8_source_8_source_ram_rdata;
  wire _stream_conv2d_8_source_8_source_ram_renable;
  wire _stream_conv2d_8_source_8_source_ram_rvalid;
  wire [7:0] _stream_conv2d_8_source_8_source_ram_sel;
  wire _stream_conv2d_8_source_busy;
  wire _stream_conv2d_8_start;
  wire _stream_conv2d_8_start_flag;
  wire _stream_conv2d_8_term_sink;
  wire [8:0] _stream_matmul_15_constant_0_next_constant_data;
  wire _stream_matmul_15_constant_15_next_constant_data;
  wire _stream_matmul_15_constant_16_next_constant_data;
  wire [3:0] _stream_matmul_15_constant_17_next_constant_data;
  wire _stream_matmul_15_constant_1_next_constant_data;
  wire _stream_matmul_15_constant_2_next_constant_data;
  wire _stream_matmul_15_constant_3_next_constant_data;
  wire _stream_matmul_15_done;
  wire _stream_matmul_15_end_flag;
  wire [31:0] _stream_matmul_15_fsm;
  wire [32:0] _stream_matmul_15_sink_21_sink_count;
  wire [31:0] _stream_matmul_15_sink_21_sink_fsm_4;
  wire [2:0] _stream_matmul_15_sink_21_sink_mode;
  wire [31:0] _stream_matmul_15_sink_21_sink_offset;
  wire [7:0] _stream_matmul_15_sink_21_sink_ram_sel;
  wire [32:0] _stream_matmul_15_sink_21_sink_size;
  wire [31:0] _stream_matmul_15_sink_21_sink_stride;
  wire [31:0] _stream_matmul_15_sink_21_sink_stride_buf;
  wire [31:0] _stream_matmul_15_sink_21_sink_waddr;
  wire [7:0] _stream_matmul_15_sink_21_sink_wdata;
  wire _stream_matmul_15_sink_21_sink_wenable;
  wire _stream_matmul_15_source_10_idle;
  wire [7:0] _stream_matmul_15_source_10_source_empty_data;
  wire _stream_matmul_15_source_12_idle;
  wire [7:0] _stream_matmul_15_source_12_source_empty_data;
  wire _stream_matmul_15_source_14_idle;
  wire [7:0] _stream_matmul_15_source_14_source_empty_data;
  wire _stream_matmul_15_source_19_idle;
  wire [2:0] _stream_matmul_15_source_19_source_mode;
  wire [31:0] _stream_matmul_15_source_19_source_offset;
  wire [31:0] _stream_matmul_15_source_19_source_offset_buf;
  wire [31:0] _stream_matmul_15_source_19_source_pat_all_offset;
  wire [31:0] _stream_matmul_15_source_19_source_pat_fsm_2;
  wire [31:0] _stream_matmul_15_source_19_source_ram_raddr;
  wire [7:0] _stream_matmul_15_source_19_source_ram_rdata;
  wire _stream_matmul_15_source_19_source_ram_renable;
  wire _stream_matmul_15_source_19_source_ram_rvalid;
  wire [7:0] _stream_matmul_15_source_19_source_ram_sel;
  wire _stream_matmul_15_source_20_idle;
  wire [2:0] _stream_matmul_15_source_20_source_mode;
  wire [31:0] _stream_matmul_15_source_20_source_offset;
  wire [31:0] _stream_matmul_15_source_20_source_offset_buf;
  wire [31:0] _stream_matmul_15_source_20_source_pat_all_offset;
  wire [31:0] _stream_matmul_15_source_20_source_pat_fsm_3;
  wire [31:0] _stream_matmul_15_source_20_source_ram_raddr;
  wire [7:0] _stream_matmul_15_source_20_source_ram_rdata;
  wire _stream_matmul_15_source_20_source_ram_renable;
  wire _stream_matmul_15_source_20_source_ram_rvalid;
  wire [7:0] _stream_matmul_15_source_20_source_ram_sel;
  wire _stream_matmul_15_source_6_idle;
  wire [2:0] _stream_matmul_15_source_6_source_mode;
  wire [31:0] _stream_matmul_15_source_6_source_offset;
  wire [31:0] _stream_matmul_15_source_6_source_offset_buf;
  wire [31:0] _stream_matmul_15_source_6_source_pat_all_offset;
  wire [31:0] _stream_matmul_15_source_6_source_pat_fsm_0;
  wire [31:0] _stream_matmul_15_source_6_source_ram_raddr;
  wire [31:0] _stream_matmul_15_source_6_source_ram_rdata;
  wire _stream_matmul_15_source_6_source_ram_renable;
  wire _stream_matmul_15_source_6_source_ram_rvalid;
  wire [7:0] _stream_matmul_15_source_6_source_ram_sel;
  wire _stream_matmul_15_source_8_idle;
  wire [2:0] _stream_matmul_15_source_8_source_mode;
  wire [31:0] _stream_matmul_15_source_8_source_offset;
  wire [31:0] _stream_matmul_15_source_8_source_offset_buf;
  wire [31:0] _stream_matmul_15_source_8_source_pat_all_offset;
  wire [31:0] _stream_matmul_15_source_8_source_pat_fsm_1;
  wire [31:0] _stream_matmul_15_source_8_source_ram_raddr;
  wire [7:0] _stream_matmul_15_source_8_source_ram_rdata;
  wire _stream_matmul_15_source_8_source_ram_renable;
  wire _stream_matmul_15_source_8_source_ram_rvalid;
  wire [7:0] _stream_matmul_15_source_8_source_ram_sel;
  wire _stream_matmul_15_source_busy;
  wire _stream_matmul_15_start;
  wire _stream_matmul_15_start_flag;
  wire _stream_matmul_15_term_sink;
  wire [2:0] _stream_max_pool_serial_9_constant_0_next_constant_data;
  wire [3:0] _stream_max_pool_serial_9_constant_2_next_constant_data;
  wire _stream_max_pool_serial_9_end_flag;
  wire [31:0] _stream_max_pool_serial_9_fsm;
  wire _stream_max_pool_serial_9_reduce_reset;
  wire [32:0] _stream_max_pool_serial_9_sink_3_sink_count;
  wire [31:0] _stream_max_pool_serial_9_sink_3_sink_fsm_1;
  wire [2:0] _stream_max_pool_serial_9_sink_3_sink_mode;
  wire [31:0] _stream_max_pool_serial_9_sink_3_sink_offset;
  wire [7:0] _stream_max_pool_serial_9_sink_3_sink_ram_sel;
  wire [32:0] _stream_max_pool_serial_9_sink_3_sink_size;
  wire [31:0] _stream_max_pool_serial_9_sink_3_sink_stride;
  wire [31:0] _stream_max_pool_serial_9_sink_3_sink_stride_buf;
  wire [31:0] _stream_max_pool_serial_9_sink_3_sink_waddr;
  wire [7:0] _stream_max_pool_serial_9_sink_3_sink_wdata;
  wire _stream_max_pool_serial_9_sink_3_sink_wenable;
  wire _stream_max_pool_serial_9_source_1_idle;
  wire [2:0] _stream_max_pool_serial_9_source_1_source_mode;
  wire [31:0] _stream_max_pool_serial_9_source_1_source_offset;
  wire [31:0] _stream_max_pool_serial_9_source_1_source_offset_buf;
  wire [31:0] _stream_max_pool_serial_9_source_1_source_pat_all_offset;
  wire [31:0] _stream_max_pool_serial_9_source_1_source_pat_fsm_0;
  wire [31:0] _stream_max_pool_serial_9_source_1_source_ram_raddr;
  wire [7:0] _stream_max_pool_serial_9_source_1_source_ram_rdata;
  wire _stream_max_pool_serial_9_source_1_source_ram_renable;
  wire _stream_max_pool_serial_9_source_1_source_ram_rvalid;
  wire [7:0] _stream_max_pool_serial_9_source_1_source_ram_sel;
  wire _stream_max_pool_serial_9_source_busy;
  wire _stream_max_pool_serial_9_start;
  wire _stream_max_pool_serial_9_start_flag;
  wire _stream_max_pool_serial_9_term_sink;
  wire _substream__reduce_max_13_size_data_cond_772_43;
  wire _substream__reduce_max_13_x_data_cond_772_42;
  wire _substream_acc_0_rshift_data_cond_727_37;
  wire _substream_acc_0_rshift_data_cond_859_49;
  wire _substream_acc_0_size_data_cond_727_38;
  wire _substream_acc_0_size_data_cond_859_50;
  wire _substream_acc_0_x_data_cond_727_36;
  wire _substream_acc_0_x_data_cond_859_48;
  wire _substream_add_tree_1_var0_data_cond_857_47;
  wire _substream_add_tree_2_var0_data_cond_725_27;
  wire _substream_add_tree_2_var1_data_cond_725_28;
  wire _substream_add_tree_2_var2_data_cond_725_29;
  wire _substream_add_tree_2_var3_data_cond_725_30;
  wire _substream_add_tree_2_var4_data_cond_725_31;
  wire _substream_add_tree_2_var5_data_cond_725_32;
  wire _substream_add_tree_2_var6_data_cond_725_33;
  wire _substream_add_tree_2_var7_data_cond_725_34;
  wire _substream_add_tree_2_var8_data_cond_725_35;
  wire _substream_mul_10_rshift_data_cond_674_20;
  wire _substream_mul_10_x_data_cond_674_18;
  wire _substream_mul_10_y_data_cond_674_19;
  wire _substream_mul_11_rshift_data_cond_691_23;
  wire _substream_mul_11_x_data_cond_691_21;
  wire _substream_mul_11_y_data_cond_691_22;
  wire _substream_mul_12_rshift_data_cond_708_26;
  wire _substream_mul_12_x_data_cond_708_24;
  wire _substream_mul_12_y_data_cond_708_25;
  wire _substream_mul_4_rshift_data_cond_572_2;
  wire _substream_mul_4_rshift_data_cond_854_46;
  wire _substream_mul_4_x_data_cond_572_0;
  wire _substream_mul_4_x_data_cond_854_44;
  wire _substream_mul_4_y_data_cond_572_1;
  wire _substream_mul_4_y_data_cond_854_45;
  wire _substream_mul_5_rshift_data_cond_589_5;
  wire _substream_mul_5_x_data_cond_589_3;
  wire _substream_mul_5_y_data_cond_589_4;
  wire _substream_mul_6_rshift_data_cond_606_8;
  wire _substream_mul_6_x_data_cond_606_6;
  wire _substream_mul_6_y_data_cond_606_7;
  wire _substream_mul_7_rshift_data_cond_623_11;
  wire _substream_mul_7_x_data_cond_623_9;
  wire _substream_mul_7_y_data_cond_623_10;
  wire _substream_mul_8_rshift_data_cond_640_14;
  wire _substream_mul_8_x_data_cond_640_12;
  wire _substream_mul_8_y_data_cond_640_13;
  wire _substream_mul_9_rshift_data_cond_657_17;
  wire _substream_mul_9_x_data_cond_657_15;
  wire _substream_mul_9_y_data_cond_657_16;
  wire _substream_mul_rshift_clip_3_rshift_data_cond_743_41;
  wire _substream_mul_rshift_clip_3_rshift_data_cond_864_53;
  wire _substream_mul_rshift_clip_3_x_data_cond_743_39;
  wire _substream_mul_rshift_clip_3_x_data_cond_864_51;
  wire _substream_mul_rshift_clip_3_y_data_cond_743_40;
  wire _substream_mul_rshift_clip_3_y_data_cond_864_52;
  wire [31:0] \_times_mul_39.mult._a ;
  wire [7:0] \_times_mul_39.mult._b ;
  wire [39:0] \_times_mul_39.mult._mul ;
  wire [39:0] \_times_mul_39.mult._pipe_mul0 ;
  wire [39:0] \_times_mul_39.mult._pipe_mul1 ;
  wire [39:0] _times_mul_odata_reg_39;
  wire [5:0] _tmp_0;
  wire _tmp_1;
  wire [8:0] _tmp_100;
  wire [7:0] _tmp_1000;
  wire _tmp_1003;
  wire [8:0] _tmp_101;
  wire [8:0] _tmp_102;
  wire [7:0] _tmp_1020;
  wire _tmp_1023;
  wire [8:0] _tmp_103;
  wire [7:0] _tmp_1030;
  wire _tmp_1033;
  wire _tmp_1037;
  wire [8:0] _tmp_104;
  wire [8:0] _tmp_105;
  wire [8:0] _tmp_106;
  wire [8:0] _tmp_107;
  wire [8:0] _tmp_108;
  wire [8:0] _tmp_109;
  wire _tmp_1091;
  wire [8:0] _tmp_110;
  wire [8:0] _tmp_111;
  wire _tmp_1119;
  wire [8:0] _tmp_112;
  wire _tmp_1124;
  wire [7:0] _tmp_1125;
  wire _tmp_1126;
  wire _tmp_1127;
  wire _tmp_1128;
  wire _tmp_1129;
  wire [8:0] _tmp_113;
  wire [33:0] _tmp_1130;
  wire _tmp_1131;
  wire _tmp_1136;
  wire [7:0] _tmp_1137;
  wire _tmp_1138;
  wire _tmp_1139;
  wire [8:0] _tmp_114;
  wire _tmp_1140;
  wire _tmp_1141;
  wire [33:0] _tmp_1142;
  wire _tmp_1143;
  wire _tmp_1148;
  wire [7:0] _tmp_1149;
  wire _tmp_1150;
  wire _tmp_1151;
  wire _tmp_1152;
  wire _tmp_1153;
  wire [33:0] _tmp_1154;
  wire _tmp_1155;
  wire _tmp_1160;
  wire [7:0] _tmp_1161;
  wire _tmp_1162;
  wire _tmp_1163;
  wire _tmp_1164;
  wire _tmp_1165;
  wire [33:0] _tmp_1166;
  wire _tmp_1167;
  wire [33:0] _tmp_12;
  wire [3:0] _tmp_124;
  wire [9:0] _tmp_125;
  wire [33:0] _tmp_126;
  wire _tmp_127;
  wire [8:0] _tmp_128;
  wire [8:0] _tmp_129;
  wire _tmp_13;
  wire [8:0] _tmp_130;
  wire [8:0] _tmp_131;
  wire [8:0] _tmp_132;
  wire [8:0] _tmp_133;
  wire [8:0] _tmp_134;
  wire [8:0] _tmp_135;
  wire [8:0] _tmp_136;
  wire [8:0] _tmp_137;
  wire [8:0] _tmp_138;
  wire [8:0] _tmp_139;
  wire [8:0] _tmp_14;
  wire [8:0] _tmp_140;
  wire [8:0] _tmp_141;
  wire [8:0] _tmp_142;
  wire [8:0] _tmp_143;
  wire [8:0] _tmp_144;
  wire [8:0] _tmp_145;
  wire [3:0] _tmp_155;
  wire [9:0] _tmp_161;
  wire [33:0] _tmp_162;
  wire _tmp_163;
  wire [8:0] _tmp_164;
  wire [8:0] _tmp_165;
  wire [8:0] _tmp_166;
  wire [8:0] _tmp_167;
  wire [8:0] _tmp_168;
  wire [8:0] _tmp_169;
  wire [1:0] _tmp_173;
  wire [9:0] _tmp_174;
  wire [33:0] _tmp_175;
  wire _tmp_176;
  wire [8:0] _tmp_177;
  wire [8:0] _tmp_178;
  wire [8:0] _tmp_179;
  wire [8:0] _tmp_180;
  wire [8:0] _tmp_181;
  wire [8:0] _tmp_182;
  wire [1:0] _tmp_186;
  wire [9:0] _tmp_187;
  wire [33:0] _tmp_188;
  wire _tmp_189;
  wire [33:0] _tmp_19;
  wire [8:0] _tmp_190;
  wire [8:0] _tmp_191;
  wire [8:0] _tmp_192;
  wire [8:0] _tmp_193;
  wire [8:0] _tmp_194;
  wire [8:0] _tmp_195;
  wire [1:0] _tmp_199;
  wire _tmp_2;
  wire _tmp_20;
  wire [9:0] _tmp_200;
  wire [33:0] _tmp_201;
  wire _tmp_202;
  wire [8:0] _tmp_203;
  wire [8:0] _tmp_204;
  wire [8:0] _tmp_205;
  wire [8:0] _tmp_206;
  wire [8:0] _tmp_207;
  wire [8:0] _tmp_208;
  wire [33:0] _tmp_21;
  wire [1:0] _tmp_212;
  wire [9:0] _tmp_218;
  wire [33:0] _tmp_219;
  wire _tmp_22;
  wire _tmp_220;
  wire [8:0] _tmp_221;
  wire [8:0] _tmp_222;
  wire [8:0] _tmp_223;
  wire [8:0] _tmp_224;
  wire [8:0] _tmp_225;
  wire [8:0] _tmp_226;
  wire [33:0] _tmp_23;
  wire [1:0] _tmp_230;
  wire [9:0] _tmp_231;
  wire [33:0] _tmp_232;
  wire _tmp_233;
  wire [8:0] _tmp_234;
  wire [8:0] _tmp_235;
  wire [8:0] _tmp_236;
  wire [8:0] _tmp_237;
  wire [8:0] _tmp_238;
  wire [8:0] _tmp_239;
  wire _tmp_24;
  wire [1:0] _tmp_243;
  wire [9:0] _tmp_244;
  wire [33:0] _tmp_245;
  wire _tmp_246;
  wire [8:0] _tmp_247;
  wire [8:0] _tmp_248;
  wire [8:0] _tmp_249;
  wire [33:0] _tmp_25;
  wire [8:0] _tmp_250;
  wire [8:0] _tmp_251;
  wire [8:0] _tmp_252;
  wire [1:0] _tmp_256;
  wire [9:0] _tmp_257;
  wire [33:0] _tmp_258;
  wire _tmp_259;
  wire _tmp_26;
  wire [8:0] _tmp_260;
  wire [8:0] _tmp_261;
  wire [8:0] _tmp_262;
  wire [8:0] _tmp_263;
  wire [8:0] _tmp_264;
  wire [8:0] _tmp_265;
  wire [1:0] _tmp_269;
  wire [9:0] _tmp_275;
  wire [33:0] _tmp_276;
  wire _tmp_277;
  wire [8:0] _tmp_278;
  wire [8:0] _tmp_279;
  wire [8:0] _tmp_280;
  wire [8:0] _tmp_281;
  wire [8:0] _tmp_282;
  wire [8:0] _tmp_283;
  wire [1:0] _tmp_287;
  wire [9:0] _tmp_288;
  wire [33:0] _tmp_289;
  wire _tmp_290;
  wire [8:0] _tmp_291;
  wire [8:0] _tmp_292;
  wire [8:0] _tmp_293;
  wire [8:0] _tmp_294;
  wire [8:0] _tmp_295;
  wire [8:0] _tmp_296;
  wire _tmp_3;
  wire [1:0] _tmp_300;
  wire [9:0] _tmp_301;
  wire [33:0] _tmp_302;
  wire _tmp_303;
  wire [8:0] _tmp_304;
  wire [8:0] _tmp_305;
  wire [8:0] _tmp_306;
  wire [8:0] _tmp_307;
  wire [8:0] _tmp_308;
  wire [8:0] _tmp_309;
  wire [1:0] _tmp_313;
  wire [9:0] _tmp_314;
  wire [33:0] _tmp_315;
  wire _tmp_316;
  wire [8:0] _tmp_317;
  wire [8:0] _tmp_318;
  wire [8:0] _tmp_319;
  wire [9:0] _tmp_32;
  wire [8:0] _tmp_320;
  wire [8:0] _tmp_321;
  wire [8:0] _tmp_322;
  wire [1:0] _tmp_326;
  wire [33:0] _tmp_33;
  wire _tmp_336;
  wire _tmp_34;
  wire [7:0] _tmp_344;
  wire _tmp_347;
  wire [8:0] _tmp_35;
  wire [8:0] _tmp_36;
  wire [7:0] _tmp_364;
  wire _tmp_367;
  wire [8:0] _tmp_37;
  wire [7:0] _tmp_374;
  wire _tmp_377;
  wire [8:0] _tmp_38;
  wire [7:0] _tmp_384;
  wire _tmp_387;
  wire [8:0] _tmp_39;
  wire [7:0] _tmp_394;
  wire _tmp_397;
  wire _tmp_4;
  wire [8:0] _tmp_40;
  wire [7:0] _tmp_404;
  wire _tmp_407;
  wire [8:0] _tmp_41;
  wire [7:0] _tmp_414;
  wire _tmp_417;
  wire [8:0] _tmp_42;
  wire [7:0] _tmp_424;
  wire _tmp_427;
  wire [8:0] _tmp_43;
  wire [7:0] _tmp_434;
  wire _tmp_437;
  wire [8:0] _tmp_44;
  wire [7:0] _tmp_444;
  wire _tmp_447;
  wire [8:0] _tmp_45;
  wire [7:0] _tmp_454;
  wire _tmp_457;
  wire [8:0] _tmp_46;
  wire [7:0] _tmp_464;
  wire _tmp_467;
  wire [8:0] _tmp_47;
  wire [7:0] _tmp_474;
  wire _tmp_477;
  wire [8:0] _tmp_48;
  wire [7:0] _tmp_484;
  wire _tmp_487;
  wire [8:0] _tmp_49;
  wire [7:0] _tmp_494;
  wire _tmp_497;
  wire [3:0] _tmp_5;
  wire [8:0] _tmp_50;
  wire [7:0] _tmp_504;
  wire _tmp_507;
  wire [8:0] _tmp_51;
  wire [7:0] _tmp_514;
  wire _tmp_517;
  wire [8:0] _tmp_52;
  wire [7:0] _tmp_524;
  wire _tmp_527;
  wire [7:0] _tmp_534;
  wire _tmp_537;
  wire _tmp_541;
  wire [31:0] _tmp_6;
  wire [3:0] _tmp_62;
  wire [9:0] _tmp_63;
  wire [33:0] _tmp_64;
  wire _tmp_65;
  wire [8:0] _tmp_66;
  wire [8:0] _tmp_67;
  wire [8:0] _tmp_68;
  wire [8:0] _tmp_69;
  wire _tmp_7;
  wire [8:0] _tmp_70;
  wire [8:0] _tmp_71;
  wire [8:0] _tmp_72;
  wire [8:0] _tmp_73;
  wire [8:0] _tmp_74;
  wire [8:0] _tmp_75;
  wire [8:0] _tmp_76;
  wire [8:0] _tmp_77;
  wire _tmp_771;
  wire [8:0] _tmp_78;
  wire [8:0] _tmp_79;
  wire _tmp_799;
  wire [31:0] _tmp_8;
  wire [8:0] _tmp_80;
  wire _tmp_804;
  wire [7:0] _tmp_805;
  wire _tmp_806;
  wire _tmp_807;
  wire _tmp_808;
  wire _tmp_809;
  wire [8:0] _tmp_81;
  wire [33:0] _tmp_810;
  wire _tmp_811;
  wire _tmp_816;
  wire [7:0] _tmp_817;
  wire _tmp_818;
  wire _tmp_819;
  wire [8:0] _tmp_82;
  wire _tmp_820;
  wire _tmp_821;
  wire [33:0] _tmp_822;
  wire _tmp_823;
  wire _tmp_828;
  wire [7:0] _tmp_829;
  wire [8:0] _tmp_83;
  wire _tmp_830;
  wire _tmp_831;
  wire _tmp_832;
  wire _tmp_833;
  wire [33:0] _tmp_834;
  wire _tmp_835;
  wire _tmp_840;
  wire [7:0] _tmp_841;
  wire _tmp_842;
  wire _tmp_843;
  wire _tmp_844;
  wire _tmp_845;
  wire [33:0] _tmp_846;
  wire [8:0] _tmp_847;
  wire _tmp_848;
  wire [33:0] _tmp_853;
  wire _tmp_854;
  wire [33:0] _tmp_855;
  wire _tmp_856;
  wire [33:0] _tmp_857;
  wire _tmp_858;
  wire [33:0] _tmp_859;
  wire _tmp_860;
  wire [7:0] _tmp_870;
  wire _tmp_873;
  wire _tmp_878;
  wire _tmp_894;
  wire _tmp_910;
  wire _tmp_915;
  wire [7:0] _tmp_916;
  wire _tmp_917;
  wire _tmp_918;
  wire _tmp_919;
  wire _tmp_920;
  wire [33:0] _tmp_921;
  wire _tmp_922;
  wire _tmp_927;
  wire [7:0] _tmp_928;
  wire _tmp_929;
  wire [3:0] _tmp_93;
  wire _tmp_930;
  wire _tmp_931;
  wire _tmp_932;
  wire [33:0] _tmp_933;
  wire _tmp_934;
  wire _tmp_939;
  wire [9:0] _tmp_94;
  wire [7:0] _tmp_940;
  wire _tmp_941;
  wire _tmp_942;
  wire _tmp_943;
  wire _tmp_944;
  wire [33:0] _tmp_945;
  wire _tmp_946;
  wire [33:0] _tmp_95;
  wire _tmp_951;
  wire [7:0] _tmp_952;
  wire _tmp_953;
  wire _tmp_954;
  wire _tmp_955;
  wire _tmp_956;
  wire [33:0] _tmp_957;
  wire _tmp_958;
  wire _tmp_96;
  wire [33:0] _tmp_964;
  wire _tmp_965;
  wire [33:0] _tmp_966;
  wire _tmp_967;
  wire [33:0] _tmp_968;
  wire _tmp_969;
  wire [8:0] _tmp_97;
  wire [33:0] _tmp_970;
  wire _tmp_971;
  wire [33:0] _tmp_975;
  wire _tmp_976;
  wire [33:0] _tmp_977;
  wire _tmp_978;
  wire [33:0] _tmp_979;
  wire [8:0] _tmp_98;
  wire _tmp_980;
  wire [33:0] _tmp_981;
  wire _tmp_982;
  wire [8:0] _tmp_99;
  wire _tmp_992;
  wire [31:0] _wdata_10;
  wire [31:0] _wdata_159;
  wire [31:0] _wdata_17;
  wire [31:0] _wdata_216;
  wire [31:0] _wdata_273;
  wire [31:0] _wdata_30;
  wire [31:0] _wdata_851;
  wire [31:0] _wdata_962;
  wire [31:0] _wdata_973;
  wire _wvalid_11;
  wire _wvalid_160;
  wire _wvalid_18;
  wire _wvalid_217;
  wire _wvalid_274;
  wire _wvalid_31;
  wire _wvalid_852;
  wire _wvalid_963;
  wire _wvalid_974;
  wire axim_flag_1118;
  wire axim_flag_15;
  wire axim_flag_158;
  wire axim_flag_16;
  wire axim_flag_215;
  wire axim_flag_272;
  wire axim_flag_29;
  wire axim_flag_798;
  wire axim_flag_849;
  wire axim_flag_850;
  wire axim_flag_861;
  wire axim_flag_9;
  wire axim_flag_909;
  wire axim_flag_959;
  wire axim_flag_960;
  wire axim_flag_961;
  wire axim_flag_972;
  wire [31:0] control_conv2d_8;
  wire [31:0] control_matmul_15;
  wire [31:0] control_max_pool_serial_9;
  wire [31:0] conv2d_8_act_base_offset;
  wire [31:0] conv2d_8_act_base_offset_bat;
  wire [31:0] conv2d_8_act_base_offset_row;
  wire [31:0] conv2d_8_act_page_comp_offset_0;
  wire [31:0] conv2d_8_act_page_comp_offset_1;
  wire [31:0] conv2d_8_act_page_comp_offset_2;
  wire [31:0] conv2d_8_act_page_comp_offset_buf_0;
  wire [31:0] conv2d_8_act_page_comp_offset_buf_1;
  wire [31:0] conv2d_8_act_page_comp_offset_buf_2;
  wire [31:0] conv2d_8_act_page_dma_offset_0;
  wire [31:0] conv2d_8_act_page_dma_offset_1;
  wire [31:0] conv2d_8_act_page_dma_offset_2;
  wire [31:0] conv2d_8_arg_objaddr_0;
  wire [31:0] conv2d_8_arg_objaddr_1;
  wire [31:0] conv2d_8_arg_objaddr_2;
  wire [31:0] conv2d_8_arg_objaddr_3;
  wire [31:0] conv2d_8_bat_count;
  wire [31:0] conv2d_8_col_count;
  wire [1:0] conv2d_8_col_select;
  wire [31:0] conv2d_8_comp_fsm;
  wire conv2d_8_control_param_index;
  wire conv2d_8_dma_flag_0;
  wire conv2d_8_dma_flag_1;
  wire conv2d_8_dma_flag_2;
  wire conv2d_8_dma_out_mask_0;
  wire conv2d_8_dma_pad_mask_0;
  wire conv2d_8_dma_pad_mask_1;
  wire conv2d_8_dma_pad_mask_2;
  wire [31:0] conv2d_8_filter_base_offset;
  wire [31:0] conv2d_8_filter_page_comp_offset;
  wire [31:0] conv2d_8_filter_page_comp_offset_buf;
  wire [31:0] conv2d_8_filter_page_dma_offset;
  wire [31:0] conv2d_8_mux_act_gaddr_0;
  wire [31:0] conv2d_8_mux_act_gaddr_1;
  wire [31:0] conv2d_8_mux_act_gaddr_2;
  wire conv2d_8_mux_dma_flag_0;
  wire conv2d_8_mux_dma_flag_1;
  wire conv2d_8_mux_dma_flag_2;
  wire conv2d_8_mux_dma_pad_mask_0;
  wire conv2d_8_mux_dma_pad_mask_1;
  wire conv2d_8_mux_dma_pad_mask_2;
  wire conv2d_8_mux_next_dma_flag_0;
  wire conv2d_8_mux_next_dma_flag_1;
  wire conv2d_8_mux_next_dma_flag_2;
  wire [31:0] conv2d_8_next_out_write_size;
  wire [31:0] conv2d_8_next_stream_num_ops;
  wire [31:0] conv2d_8_objaddr;
  wire [31:0] conv2d_8_och_count;
  wire [31:0] conv2d_8_och_count_buf;
  wire [31:0] conv2d_8_out_base_offset;
  wire [31:0] conv2d_8_out_base_offset_bat;
  wire [31:0] conv2d_8_out_base_offset_col;
  wire [31:0] conv2d_8_out_base_offset_och;
  wire [31:0] conv2d_8_out_base_offset_row;
  wire [31:0] conv2d_8_out_base_offset_val;
  wire [31:0] conv2d_8_out_laddr_offset;
  wire conv2d_8_out_page;
  wire [31:0] conv2d_8_out_page_comp_offset;
  wire [31:0] conv2d_8_out_page_comp_offset_buf;
  wire [31:0] conv2d_8_out_page_dma_offset;
  wire [31:0] conv2d_8_out_ram_select;
  wire [31:0] conv2d_8_out_row_count;
  wire [31:0] conv2d_8_prev_bat_count;
  wire [31:0] conv2d_8_prev_och_count;
  wire [31:0] conv2d_8_prev_row_count;
  wire [1:0] conv2d_8_prev_row_select;
  wire [31:0] conv2d_8_row_count;
  wire [31:0] conv2d_8_row_count_buf;
  wire [1:0] conv2d_8_row_select;
  wire [1:0] conv2d_8_row_select_buf;
  wire conv2d_8_skip_comp;
  wire conv2d_8_skip_read_act;
  wire conv2d_8_skip_read_filter;
  wire conv2d_8_skip_write_out;
  wire [31:0] conv2d_8_stream_act_local_0;
  wire [31:0] conv2d_8_stream_act_local_1;
  wire [31:0] conv2d_8_stream_act_local_2;
  wire [31:0] conv2d_8_stream_act_local_3;
  wire [31:0] conv2d_8_stream_act_local_4;
  wire [31:0] conv2d_8_stream_act_local_5;
  wire [31:0] conv2d_8_stream_act_local_6;
  wire [31:0] conv2d_8_stream_act_local_7;
  wire [31:0] conv2d_8_stream_act_local_8;
  wire [31:0] conv2d_8_stream_out_local_col;
  wire conv2d_8_stream_pad_mask_0_0;
  wire conv2d_8_stream_pad_mask_0_1;
  wire conv2d_8_stream_pad_mask_0_2;
  wire conv2d_8_stream_pad_mask_1_0;
  wire conv2d_8_stream_pad_mask_1_1;
  wire conv2d_8_stream_pad_mask_1_2;
  wire conv2d_8_stream_pad_mask_2_0;
  wire conv2d_8_stream_pad_mask_2_1;
  wire conv2d_8_stream_pad_mask_2_2;
  wire [8:0] conv2d_8_stream_pad_masks;
  wire [31:0] conv2d_8_sync_comp_count;
  wire [31:0] conv2d_8_sync_out_count;
  wire conv2d_8_update_filter;
  wire [4:0] cparam_conv2d_8_act_num_row;
  wire [31:0] cparam_conv2d_8_act_offset_values_0;
  wire [31:0] cparam_conv2d_8_act_offset_values_1;
  wire [31:0] cparam_conv2d_8_act_offset_values_2;
  wire [7:0] cparam_conv2d_8_act_read_size;
  wire [6:0] cparam_conv2d_8_act_read_step;
  wire [4:0] cparam_conv2d_8_bias_num;
  wire [1:0] cparam_conv2d_8_col_select_initval;
  wire [3:0] cparam_conv2d_8_cshamt_out_value;
  wire [10:0] cparam_conv2d_8_filter_base_step;
  wire [7:0] cparam_conv2d_8_filter_read_step;
  wire [4:0] cparam_conv2d_8_inc_act_laddr_large;
  wire [4:0] cparam_conv2d_8_inc_sync_out;
  wire [4:0] cparam_conv2d_8_max_col_count;
  wire [6:0] cparam_conv2d_8_och_count_step;
  wire [8:0] cparam_conv2d_8_out_row_step;
  wire cparam_conv2d_8_pad_col_left;
  wire [3:0] cparam_conv2d_8_stream_act_local_large_offset;
  wire [4:0] cparam_conv2d_8_stream_reduce_size;
  wire [4:0] cparam_max_pool_serial_9_act_num_col;
  wire [31:0] cparam_max_pool_serial_9_act_offset_values_1;
  wire [9:0] cparam_max_pool_serial_9_act_row_step;
  wire [5:0] cparam_max_pool_serial_9_inc_act_laddr;
  wire [4:0] cparam_max_pool_serial_9_inc_out_laddr;
  wire [4:0] cparam_max_pool_serial_9_max_col_count;
  wire [7:0] cparam_max_pool_serial_9_out_row_step;
  wire [31:0] main_fsm;
  wire [31:0] matmul_15_act_base_offset;
  wire [31:0] matmul_15_act_base_offset_bat;
  wire [31:0] matmul_15_act_base_offset_row;
  wire [31:0] matmul_15_act_page_comp_offset_0;
  wire [31:0] matmul_15_act_page_comp_offset_buf_0;
  wire [31:0] matmul_15_act_page_dma_offset_0;
  wire [31:0] matmul_15_arg_objaddr_0;
  wire [31:0] matmul_15_arg_objaddr_1;
  wire [31:0] matmul_15_arg_objaddr_2;
  wire [31:0] matmul_15_arg_objaddr_3;
  wire [31:0] matmul_15_bat_count;
  wire [31:0] matmul_15_col_count;
  wire matmul_15_col_select;
  wire [31:0] matmul_15_comp_fsm;
  wire matmul_15_dma_flag_0;
  wire matmul_15_dma_out_mask_0;
  wire matmul_15_dma_pad_mask_0;
  wire [31:0] matmul_15_filter_base_offset;
  wire [31:0] matmul_15_filter_page_comp_offset;
  wire [31:0] matmul_15_filter_page_comp_offset_buf;
  wire [31:0] matmul_15_filter_page_dma_offset;
  wire [31:0] matmul_15_mux_act_gaddr_0;
  wire matmul_15_mux_dma_flag_0;
  wire matmul_15_mux_dma_pad_mask_0;
  wire [31:0] matmul_15_next_out_write_size;
  wire [31:0] matmul_15_next_stream_num_ops;
  wire [31:0] matmul_15_objaddr;
  wire [31:0] matmul_15_och_count;
  wire [31:0] matmul_15_och_count_buf;
  wire [31:0] matmul_15_out_base_offset;
  wire [31:0] matmul_15_out_base_offset_bat;
  wire [31:0] matmul_15_out_base_offset_col;
  wire [31:0] matmul_15_out_base_offset_och;
  wire [31:0] matmul_15_out_base_offset_row;
  wire [31:0] matmul_15_out_base_offset_val;
  wire [31:0] matmul_15_out_laddr_offset;
  wire matmul_15_out_page;
  wire [31:0] matmul_15_out_page_comp_offset;
  wire [31:0] matmul_15_out_page_comp_offset_buf;
  wire [31:0] matmul_15_out_page_dma_offset;
  wire [31:0] matmul_15_out_ram_select;
  wire [31:0] matmul_15_out_row_count;
  wire [31:0] matmul_15_prev_bat_count;
  wire [31:0] matmul_15_prev_och_count;
  wire [31:0] matmul_15_prev_row_count;
  wire matmul_15_prev_row_select;
  wire [31:0] matmul_15_row_count;
  wire [31:0] matmul_15_row_count_buf;
  wire matmul_15_row_select;
  wire matmul_15_row_select_buf;
  wire matmul_15_skip_comp;
  wire matmul_15_skip_read_act;
  wire matmul_15_skip_read_filter;
  wire matmul_15_skip_write_out;
  wire [31:0] matmul_15_stream_act_local_0;
  wire [31:0] matmul_15_stream_out_local_col;
  wire matmul_15_stream_pad_mask_0_0;
  wire matmul_15_stream_pad_masks;
  wire [31:0] matmul_15_sync_comp_count;
  wire [31:0] matmul_15_sync_out_count;
  wire [31:0] max_pool_serial_9_act_base_offset;
  wire [31:0] max_pool_serial_9_act_base_offset_bat;
  wire [31:0] max_pool_serial_9_act_base_offset_row;
  wire max_pool_serial_9_act_page;
  wire [31:0] max_pool_serial_9_act_page_comp_offset;
  wire [31:0] max_pool_serial_9_act_page_comp_offset_buf;
  wire [31:0] max_pool_serial_9_act_page_dma_offset;
  wire [31:0] max_pool_serial_9_arg_objaddr_0;
  wire [31:0] max_pool_serial_9_bat_count;
  wire [31:0] max_pool_serial_9_col_count;
  wire [31:0] max_pool_serial_9_comp_count;
  wire [31:0] max_pool_serial_9_comp_fsm;
  wire max_pool_serial_9_control_param_index;
  wire max_pool_serial_9_dma_pad_mask_0;
  wire max_pool_serial_9_dma_pad_mask_1;
  wire [31:0] max_pool_serial_9_objaddr;
  wire [31:0] max_pool_serial_9_out_base_offset;
  wire [31:0] max_pool_serial_9_out_base_offset_bat;
  wire [31:0] max_pool_serial_9_out_base_offset_row;
  wire [31:0] max_pool_serial_9_out_count;
  wire max_pool_serial_9_out_page;
  wire [31:0] max_pool_serial_9_out_page_comp_offset;
  wire [31:0] max_pool_serial_9_out_page_comp_offset_buf;
  wire [31:0] max_pool_serial_9_out_page_dma_offset;
  wire [31:0] max_pool_serial_9_prev_bat_count;
  wire [31:0] max_pool_serial_9_prev_row_count;
  wire [31:0] max_pool_serial_9_row_count;
  wire [31:0] max_pool_serial_9_row_count_buf;
  wire max_pool_serial_9_skip_comp;
  wire max_pool_serial_9_skip_read_act;
  wire max_pool_serial_9_skip_write_out;
  wire [31:0] max_pool_serial_9_stream_act_local;
  wire [31:0] max_pool_serial_9_stream_out_local;
  wire max_pool_serial_9_stream_pad_mask_0_0;
  wire max_pool_serial_9_stream_pad_mask_0_1;
  wire max_pool_serial_9_stream_pad_mask_1_0;
  wire max_pool_serial_9_stream_pad_mask_1_1;
  wire [3:0] max_pool_serial_9_stream_pad_masks;
  wire [6:0] ram_w32_l128_id0_0_addr;
  wire [31:0] ram_w32_l128_id0_0_rdata;
  wire [6:0] ram_w32_l128_id0_1_addr;
  wire [31:0] ram_w32_l128_id0_1_rdata;
  wire [31:0] ram_w32_l128_id0_1_wdata;
  wire ram_w32_l128_id0_1_wenable;
  wire [8:0] ram_w8_l2048_id0_0_0_addr;
  wire [7:0] ram_w8_l2048_id0_0_0_rdata;
  wire [7:0] ram_w8_l2048_id0_0_0_wdata;
  wire ram_w8_l2048_id0_0_0_wenable;
  wire [8:0] ram_w8_l2048_id0_0_1_addr;
  wire [7:0] ram_w8_l2048_id0_0_1_rdata;
  wire [7:0] ram_w8_l2048_id0_0_1_wdata;
  wire ram_w8_l2048_id0_0_1_wenable;
  wire [8:0] ram_w8_l2048_id0_1_0_addr;
  wire [7:0] ram_w8_l2048_id0_1_0_rdata;
  wire [7:0] ram_w8_l2048_id0_1_0_wdata;
  wire ram_w8_l2048_id0_1_0_wenable;
  wire [8:0] ram_w8_l2048_id0_1_1_addr;
  wire [7:0] ram_w8_l2048_id0_1_1_rdata;
  wire [7:0] ram_w8_l2048_id0_1_1_wdata;
  wire ram_w8_l2048_id0_1_1_wenable;
  wire [8:0] ram_w8_l2048_id0_2_0_addr;
  wire [7:0] ram_w8_l2048_id0_2_0_rdata;
  wire [7:0] ram_w8_l2048_id0_2_0_wdata;
  wire ram_w8_l2048_id0_2_0_wenable;
  wire [8:0] ram_w8_l2048_id0_2_1_addr;
  wire [7:0] ram_w8_l2048_id0_2_1_rdata;
  wire [7:0] ram_w8_l2048_id0_2_1_wdata;
  wire ram_w8_l2048_id0_2_1_wenable;
  wire [8:0] ram_w8_l2048_id0_3_0_addr;
  wire [7:0] ram_w8_l2048_id0_3_0_rdata;
  wire [7:0] ram_w8_l2048_id0_3_0_wdata;
  wire ram_w8_l2048_id0_3_0_wenable;
  wire [8:0] ram_w8_l2048_id0_3_1_addr;
  wire [7:0] ram_w8_l2048_id0_3_1_rdata;
  wire [7:0] ram_w8_l2048_id0_3_1_wdata;
  wire ram_w8_l2048_id0_3_1_wenable;
  wire [8:0] ram_w8_l2048_id10_0_0_addr;
  wire [7:0] ram_w8_l2048_id10_0_0_rdata;
  wire [8:0] ram_w8_l2048_id10_0_1_addr;
  wire [7:0] ram_w8_l2048_id10_0_1_rdata;
  wire [7:0] ram_w8_l2048_id10_0_1_wdata;
  wire ram_w8_l2048_id10_0_1_wenable;
  wire [8:0] ram_w8_l2048_id10_1_0_addr;
  wire [7:0] ram_w8_l2048_id10_1_0_rdata;
  wire [8:0] ram_w8_l2048_id10_1_1_addr;
  wire [7:0] ram_w8_l2048_id10_1_1_rdata;
  wire [7:0] ram_w8_l2048_id10_1_1_wdata;
  wire ram_w8_l2048_id10_1_1_wenable;
  wire [8:0] ram_w8_l2048_id10_2_0_addr;
  wire [7:0] ram_w8_l2048_id10_2_0_rdata;
  wire [8:0] ram_w8_l2048_id10_2_1_addr;
  wire [7:0] ram_w8_l2048_id10_2_1_rdata;
  wire [7:0] ram_w8_l2048_id10_2_1_wdata;
  wire ram_w8_l2048_id10_2_1_wenable;
  wire [8:0] ram_w8_l2048_id10_3_0_addr;
  wire [7:0] ram_w8_l2048_id10_3_0_rdata;
  wire [8:0] ram_w8_l2048_id10_3_1_addr;
  wire [7:0] ram_w8_l2048_id10_3_1_rdata;
  wire [7:0] ram_w8_l2048_id10_3_1_wdata;
  wire ram_w8_l2048_id10_3_1_wenable;
  wire [8:0] ram_w8_l2048_id11_0_0_addr;
  wire [7:0] ram_w8_l2048_id11_0_0_rdata;
  wire [8:0] ram_w8_l2048_id11_0_1_addr;
  wire [7:0] ram_w8_l2048_id11_0_1_rdata;
  wire [7:0] ram_w8_l2048_id11_0_1_wdata;
  wire ram_w8_l2048_id11_0_1_wenable;
  wire [8:0] ram_w8_l2048_id11_1_0_addr;
  wire [7:0] ram_w8_l2048_id11_1_0_rdata;
  wire [8:0] ram_w8_l2048_id11_1_1_addr;
  wire [7:0] ram_w8_l2048_id11_1_1_rdata;
  wire [7:0] ram_w8_l2048_id11_1_1_wdata;
  wire ram_w8_l2048_id11_1_1_wenable;
  wire [8:0] ram_w8_l2048_id11_2_0_addr;
  wire [7:0] ram_w8_l2048_id11_2_0_rdata;
  wire [8:0] ram_w8_l2048_id11_2_1_addr;
  wire [7:0] ram_w8_l2048_id11_2_1_rdata;
  wire [7:0] ram_w8_l2048_id11_2_1_wdata;
  wire ram_w8_l2048_id11_2_1_wenable;
  wire [8:0] ram_w8_l2048_id11_3_0_addr;
  wire [7:0] ram_w8_l2048_id11_3_0_rdata;
  wire [8:0] ram_w8_l2048_id11_3_1_addr;
  wire [7:0] ram_w8_l2048_id11_3_1_rdata;
  wire [7:0] ram_w8_l2048_id11_3_1_wdata;
  wire ram_w8_l2048_id11_3_1_wenable;
  wire [8:0] ram_w8_l2048_id12_0_0_addr;
  wire [7:0] ram_w8_l2048_id12_0_0_rdata;
  wire [8:0] ram_w8_l2048_id12_0_1_addr;
  wire [7:0] ram_w8_l2048_id12_0_1_rdata;
  wire [7:0] ram_w8_l2048_id12_0_1_wdata;
  wire ram_w8_l2048_id12_0_1_wenable;
  wire [8:0] ram_w8_l2048_id12_1_0_addr;
  wire [7:0] ram_w8_l2048_id12_1_0_rdata;
  wire [8:0] ram_w8_l2048_id12_1_1_addr;
  wire [7:0] ram_w8_l2048_id12_1_1_rdata;
  wire [7:0] ram_w8_l2048_id12_1_1_wdata;
  wire ram_w8_l2048_id12_1_1_wenable;
  wire [8:0] ram_w8_l2048_id12_2_0_addr;
  wire [7:0] ram_w8_l2048_id12_2_0_rdata;
  wire [8:0] ram_w8_l2048_id12_2_1_addr;
  wire [7:0] ram_w8_l2048_id12_2_1_rdata;
  wire [7:0] ram_w8_l2048_id12_2_1_wdata;
  wire ram_w8_l2048_id12_2_1_wenable;
  wire [8:0] ram_w8_l2048_id12_3_0_addr;
  wire [7:0] ram_w8_l2048_id12_3_0_rdata;
  wire [8:0] ram_w8_l2048_id12_3_1_addr;
  wire [7:0] ram_w8_l2048_id12_3_1_rdata;
  wire [7:0] ram_w8_l2048_id12_3_1_wdata;
  wire ram_w8_l2048_id12_3_1_wenable;
  wire [8:0] ram_w8_l2048_id13_0_0_addr;
  wire [7:0] ram_w8_l2048_id13_0_0_rdata;
  wire [8:0] ram_w8_l2048_id13_0_1_addr;
  wire [7:0] ram_w8_l2048_id13_0_1_rdata;
  wire [7:0] ram_w8_l2048_id13_0_1_wdata;
  wire ram_w8_l2048_id13_0_1_wenable;
  wire [8:0] ram_w8_l2048_id13_1_0_addr;
  wire [7:0] ram_w8_l2048_id13_1_0_rdata;
  wire [8:0] ram_w8_l2048_id13_1_1_addr;
  wire [7:0] ram_w8_l2048_id13_1_1_rdata;
  wire [7:0] ram_w8_l2048_id13_1_1_wdata;
  wire ram_w8_l2048_id13_1_1_wenable;
  wire [8:0] ram_w8_l2048_id13_2_0_addr;
  wire [7:0] ram_w8_l2048_id13_2_0_rdata;
  wire [8:0] ram_w8_l2048_id13_2_1_addr;
  wire [7:0] ram_w8_l2048_id13_2_1_rdata;
  wire [7:0] ram_w8_l2048_id13_2_1_wdata;
  wire ram_w8_l2048_id13_2_1_wenable;
  wire [8:0] ram_w8_l2048_id13_3_0_addr;
  wire [7:0] ram_w8_l2048_id13_3_0_rdata;
  wire [8:0] ram_w8_l2048_id13_3_1_addr;
  wire [7:0] ram_w8_l2048_id13_3_1_rdata;
  wire [7:0] ram_w8_l2048_id13_3_1_wdata;
  wire ram_w8_l2048_id13_3_1_wenable;
  wire [8:0] ram_w8_l2048_id14_0_0_addr;
  wire [7:0] ram_w8_l2048_id14_0_0_rdata;
  wire [8:0] ram_w8_l2048_id14_0_1_addr;
  wire [7:0] ram_w8_l2048_id14_0_1_rdata;
  wire [7:0] ram_w8_l2048_id14_0_1_wdata;
  wire ram_w8_l2048_id14_0_1_wenable;
  wire [8:0] ram_w8_l2048_id14_1_0_addr;
  wire [7:0] ram_w8_l2048_id14_1_0_rdata;
  wire [8:0] ram_w8_l2048_id14_1_1_addr;
  wire [7:0] ram_w8_l2048_id14_1_1_rdata;
  wire [7:0] ram_w8_l2048_id14_1_1_wdata;
  wire ram_w8_l2048_id14_1_1_wenable;
  wire [8:0] ram_w8_l2048_id14_2_0_addr;
  wire [7:0] ram_w8_l2048_id14_2_0_rdata;
  wire [8:0] ram_w8_l2048_id14_2_1_addr;
  wire [7:0] ram_w8_l2048_id14_2_1_rdata;
  wire [7:0] ram_w8_l2048_id14_2_1_wdata;
  wire ram_w8_l2048_id14_2_1_wenable;
  wire [8:0] ram_w8_l2048_id14_3_0_addr;
  wire [7:0] ram_w8_l2048_id14_3_0_rdata;
  wire [8:0] ram_w8_l2048_id14_3_1_addr;
  wire [7:0] ram_w8_l2048_id14_3_1_rdata;
  wire [7:0] ram_w8_l2048_id14_3_1_wdata;
  wire ram_w8_l2048_id14_3_1_wenable;
  wire [8:0] ram_w8_l2048_id15_0_0_addr;
  wire [7:0] ram_w8_l2048_id15_0_0_rdata;
  wire [8:0] ram_w8_l2048_id15_0_1_addr;
  wire [7:0] ram_w8_l2048_id15_0_1_rdata;
  wire [7:0] ram_w8_l2048_id15_0_1_wdata;
  wire ram_w8_l2048_id15_0_1_wenable;
  wire [8:0] ram_w8_l2048_id15_1_0_addr;
  wire [7:0] ram_w8_l2048_id15_1_0_rdata;
  wire [8:0] ram_w8_l2048_id15_1_1_addr;
  wire [7:0] ram_w8_l2048_id15_1_1_rdata;
  wire [7:0] ram_w8_l2048_id15_1_1_wdata;
  wire ram_w8_l2048_id15_1_1_wenable;
  wire [8:0] ram_w8_l2048_id15_2_0_addr;
  wire [7:0] ram_w8_l2048_id15_2_0_rdata;
  wire [8:0] ram_w8_l2048_id15_2_1_addr;
  wire [7:0] ram_w8_l2048_id15_2_1_rdata;
  wire [7:0] ram_w8_l2048_id15_2_1_wdata;
  wire ram_w8_l2048_id15_2_1_wenable;
  wire [8:0] ram_w8_l2048_id15_3_0_addr;
  wire [7:0] ram_w8_l2048_id15_3_0_rdata;
  wire [8:0] ram_w8_l2048_id15_3_1_addr;
  wire [7:0] ram_w8_l2048_id15_3_1_rdata;
  wire [7:0] ram_w8_l2048_id15_3_1_wdata;
  wire ram_w8_l2048_id15_3_1_wenable;
  wire [8:0] ram_w8_l2048_id16_0_0_addr;
  wire [7:0] ram_w8_l2048_id16_0_0_rdata;
  wire [8:0] ram_w8_l2048_id16_0_1_addr;
  wire [7:0] ram_w8_l2048_id16_0_1_rdata;
  wire [7:0] ram_w8_l2048_id16_0_1_wdata;
  wire ram_w8_l2048_id16_0_1_wenable;
  wire [8:0] ram_w8_l2048_id16_1_0_addr;
  wire [7:0] ram_w8_l2048_id16_1_0_rdata;
  wire [8:0] ram_w8_l2048_id16_1_1_addr;
  wire [7:0] ram_w8_l2048_id16_1_1_rdata;
  wire [7:0] ram_w8_l2048_id16_1_1_wdata;
  wire ram_w8_l2048_id16_1_1_wenable;
  wire [8:0] ram_w8_l2048_id16_2_0_addr;
  wire [7:0] ram_w8_l2048_id16_2_0_rdata;
  wire [8:0] ram_w8_l2048_id16_2_1_addr;
  wire [7:0] ram_w8_l2048_id16_2_1_rdata;
  wire [7:0] ram_w8_l2048_id16_2_1_wdata;
  wire ram_w8_l2048_id16_2_1_wenable;
  wire [8:0] ram_w8_l2048_id16_3_0_addr;
  wire [7:0] ram_w8_l2048_id16_3_0_rdata;
  wire [8:0] ram_w8_l2048_id16_3_1_addr;
  wire [7:0] ram_w8_l2048_id16_3_1_rdata;
  wire [7:0] ram_w8_l2048_id16_3_1_wdata;
  wire ram_w8_l2048_id16_3_1_wenable;
  wire [8:0] ram_w8_l2048_id17_0_0_addr;
  wire [7:0] ram_w8_l2048_id17_0_0_rdata;
  wire [8:0] ram_w8_l2048_id17_0_1_addr;
  wire [7:0] ram_w8_l2048_id17_0_1_rdata;
  wire [7:0] ram_w8_l2048_id17_0_1_wdata;
  wire ram_w8_l2048_id17_0_1_wenable;
  wire [8:0] ram_w8_l2048_id17_1_0_addr;
  wire [7:0] ram_w8_l2048_id17_1_0_rdata;
  wire [8:0] ram_w8_l2048_id17_1_1_addr;
  wire [7:0] ram_w8_l2048_id17_1_1_rdata;
  wire [7:0] ram_w8_l2048_id17_1_1_wdata;
  wire ram_w8_l2048_id17_1_1_wenable;
  wire [8:0] ram_w8_l2048_id17_2_0_addr;
  wire [7:0] ram_w8_l2048_id17_2_0_rdata;
  wire [8:0] ram_w8_l2048_id17_2_1_addr;
  wire [7:0] ram_w8_l2048_id17_2_1_rdata;
  wire [7:0] ram_w8_l2048_id17_2_1_wdata;
  wire ram_w8_l2048_id17_2_1_wenable;
  wire [8:0] ram_w8_l2048_id17_3_0_addr;
  wire [7:0] ram_w8_l2048_id17_3_0_rdata;
  wire [8:0] ram_w8_l2048_id17_3_1_addr;
  wire [7:0] ram_w8_l2048_id17_3_1_rdata;
  wire [7:0] ram_w8_l2048_id17_3_1_wdata;
  wire ram_w8_l2048_id17_3_1_wenable;
  wire [8:0] ram_w8_l2048_id18_0_0_addr;
  wire [7:0] ram_w8_l2048_id18_0_0_rdata;
  wire [8:0] ram_w8_l2048_id18_0_1_addr;
  wire [7:0] ram_w8_l2048_id18_0_1_rdata;
  wire [7:0] ram_w8_l2048_id18_0_1_wdata;
  wire ram_w8_l2048_id18_0_1_wenable;
  wire [8:0] ram_w8_l2048_id18_1_0_addr;
  wire [7:0] ram_w8_l2048_id18_1_0_rdata;
  wire [8:0] ram_w8_l2048_id18_1_1_addr;
  wire [7:0] ram_w8_l2048_id18_1_1_rdata;
  wire [7:0] ram_w8_l2048_id18_1_1_wdata;
  wire ram_w8_l2048_id18_1_1_wenable;
  wire [8:0] ram_w8_l2048_id18_2_0_addr;
  wire [7:0] ram_w8_l2048_id18_2_0_rdata;
  wire [8:0] ram_w8_l2048_id18_2_1_addr;
  wire [7:0] ram_w8_l2048_id18_2_1_rdata;
  wire [7:0] ram_w8_l2048_id18_2_1_wdata;
  wire ram_w8_l2048_id18_2_1_wenable;
  wire [8:0] ram_w8_l2048_id18_3_0_addr;
  wire [7:0] ram_w8_l2048_id18_3_0_rdata;
  wire [8:0] ram_w8_l2048_id18_3_1_addr;
  wire [7:0] ram_w8_l2048_id18_3_1_rdata;
  wire [7:0] ram_w8_l2048_id18_3_1_wdata;
  wire ram_w8_l2048_id18_3_1_wenable;
  wire [8:0] ram_w8_l2048_id19_0_0_addr;
  wire [7:0] ram_w8_l2048_id19_0_0_rdata;
  wire [7:0] ram_w8_l2048_id19_0_0_wdata;
  wire ram_w8_l2048_id19_0_0_wenable;
  wire [8:0] ram_w8_l2048_id19_0_1_addr;
  wire [7:0] ram_w8_l2048_id19_0_1_rdata;
  wire [8:0] ram_w8_l2048_id19_1_0_addr;
  wire [7:0] ram_w8_l2048_id19_1_0_rdata;
  wire [7:0] ram_w8_l2048_id19_1_0_wdata;
  wire ram_w8_l2048_id19_1_0_wenable;
  wire [8:0] ram_w8_l2048_id19_1_1_addr;
  wire [7:0] ram_w8_l2048_id19_1_1_rdata;
  wire [8:0] ram_w8_l2048_id19_2_0_addr;
  wire [7:0] ram_w8_l2048_id19_2_0_rdata;
  wire [7:0] ram_w8_l2048_id19_2_0_wdata;
  wire ram_w8_l2048_id19_2_0_wenable;
  wire [8:0] ram_w8_l2048_id19_2_1_addr;
  wire [7:0] ram_w8_l2048_id19_2_1_rdata;
  wire [8:0] ram_w8_l2048_id19_3_0_addr;
  wire [7:0] ram_w8_l2048_id19_3_0_rdata;
  wire [7:0] ram_w8_l2048_id19_3_0_wdata;
  wire ram_w8_l2048_id19_3_0_wenable;
  wire [8:0] ram_w8_l2048_id19_3_1_addr;
  wire [7:0] ram_w8_l2048_id19_3_1_rdata;
  wire [8:0] ram_w8_l2048_id1_0_0_addr;
  wire [7:0] ram_w8_l2048_id1_0_0_rdata;
  wire [7:0] ram_w8_l2048_id1_0_0_wdata;
  wire ram_w8_l2048_id1_0_0_wenable;
  wire [8:0] ram_w8_l2048_id1_0_1_addr;
  wire [7:0] ram_w8_l2048_id1_0_1_rdata;
  wire [7:0] ram_w8_l2048_id1_0_1_wdata;
  wire ram_w8_l2048_id1_0_1_wenable;
  wire [8:0] ram_w8_l2048_id1_1_0_addr;
  wire [7:0] ram_w8_l2048_id1_1_0_rdata;
  wire [7:0] ram_w8_l2048_id1_1_0_wdata;
  wire ram_w8_l2048_id1_1_0_wenable;
  wire [8:0] ram_w8_l2048_id1_1_1_addr;
  wire [7:0] ram_w8_l2048_id1_1_1_rdata;
  wire [7:0] ram_w8_l2048_id1_1_1_wdata;
  wire ram_w8_l2048_id1_1_1_wenable;
  wire [8:0] ram_w8_l2048_id1_2_0_addr;
  wire [7:0] ram_w8_l2048_id1_2_0_rdata;
  wire [7:0] ram_w8_l2048_id1_2_0_wdata;
  wire ram_w8_l2048_id1_2_0_wenable;
  wire [8:0] ram_w8_l2048_id1_2_1_addr;
  wire [7:0] ram_w8_l2048_id1_2_1_rdata;
  wire [7:0] ram_w8_l2048_id1_2_1_wdata;
  wire ram_w8_l2048_id1_2_1_wenable;
  wire [8:0] ram_w8_l2048_id1_3_0_addr;
  wire [7:0] ram_w8_l2048_id1_3_0_rdata;
  wire [7:0] ram_w8_l2048_id1_3_0_wdata;
  wire ram_w8_l2048_id1_3_0_wenable;
  wire [8:0] ram_w8_l2048_id1_3_1_addr;
  wire [7:0] ram_w8_l2048_id1_3_1_rdata;
  wire [7:0] ram_w8_l2048_id1_3_1_wdata;
  wire ram_w8_l2048_id1_3_1_wenable;
  wire [8:0] ram_w8_l2048_id2_0_0_addr;
  wire [7:0] ram_w8_l2048_id2_0_0_rdata;
  wire [8:0] ram_w8_l2048_id2_0_1_addr;
  wire [7:0] ram_w8_l2048_id2_0_1_rdata;
  wire [7:0] ram_w8_l2048_id2_0_1_wdata;
  wire ram_w8_l2048_id2_0_1_wenable;
  wire [8:0] ram_w8_l2048_id2_1_0_addr;
  wire [7:0] ram_w8_l2048_id2_1_0_rdata;
  wire [8:0] ram_w8_l2048_id2_1_1_addr;
  wire [7:0] ram_w8_l2048_id2_1_1_rdata;
  wire [7:0] ram_w8_l2048_id2_1_1_wdata;
  wire ram_w8_l2048_id2_1_1_wenable;
  wire [8:0] ram_w8_l2048_id2_2_0_addr;
  wire [7:0] ram_w8_l2048_id2_2_0_rdata;
  wire [8:0] ram_w8_l2048_id2_2_1_addr;
  wire [7:0] ram_w8_l2048_id2_2_1_rdata;
  wire [7:0] ram_w8_l2048_id2_2_1_wdata;
  wire ram_w8_l2048_id2_2_1_wenable;
  wire [8:0] ram_w8_l2048_id2_3_0_addr;
  wire [7:0] ram_w8_l2048_id2_3_0_rdata;
  wire [8:0] ram_w8_l2048_id2_3_1_addr;
  wire [7:0] ram_w8_l2048_id2_3_1_rdata;
  wire [7:0] ram_w8_l2048_id2_3_1_wdata;
  wire ram_w8_l2048_id2_3_1_wenable;
  wire [8:0] ram_w8_l2048_id3_0_0_addr;
  wire [7:0] ram_w8_l2048_id3_0_0_rdata;
  wire [8:0] ram_w8_l2048_id3_0_1_addr;
  wire [7:0] ram_w8_l2048_id3_0_1_rdata;
  wire [7:0] ram_w8_l2048_id3_0_1_wdata;
  wire ram_w8_l2048_id3_0_1_wenable;
  wire [8:0] ram_w8_l2048_id3_1_0_addr;
  wire [7:0] ram_w8_l2048_id3_1_0_rdata;
  wire [8:0] ram_w8_l2048_id3_1_1_addr;
  wire [7:0] ram_w8_l2048_id3_1_1_rdata;
  wire [7:0] ram_w8_l2048_id3_1_1_wdata;
  wire ram_w8_l2048_id3_1_1_wenable;
  wire [8:0] ram_w8_l2048_id3_2_0_addr;
  wire [7:0] ram_w8_l2048_id3_2_0_rdata;
  wire [8:0] ram_w8_l2048_id3_2_1_addr;
  wire [7:0] ram_w8_l2048_id3_2_1_rdata;
  wire [7:0] ram_w8_l2048_id3_2_1_wdata;
  wire ram_w8_l2048_id3_2_1_wenable;
  wire [8:0] ram_w8_l2048_id3_3_0_addr;
  wire [7:0] ram_w8_l2048_id3_3_0_rdata;
  wire [8:0] ram_w8_l2048_id3_3_1_addr;
  wire [7:0] ram_w8_l2048_id3_3_1_rdata;
  wire [7:0] ram_w8_l2048_id3_3_1_wdata;
  wire ram_w8_l2048_id3_3_1_wenable;
  wire [8:0] ram_w8_l2048_id4_0_0_addr;
  wire [7:0] ram_w8_l2048_id4_0_0_rdata;
  wire [8:0] ram_w8_l2048_id4_0_1_addr;
  wire [7:0] ram_w8_l2048_id4_0_1_rdata;
  wire [7:0] ram_w8_l2048_id4_0_1_wdata;
  wire ram_w8_l2048_id4_0_1_wenable;
  wire [8:0] ram_w8_l2048_id4_1_0_addr;
  wire [7:0] ram_w8_l2048_id4_1_0_rdata;
  wire [8:0] ram_w8_l2048_id4_1_1_addr;
  wire [7:0] ram_w8_l2048_id4_1_1_rdata;
  wire [7:0] ram_w8_l2048_id4_1_1_wdata;
  wire ram_w8_l2048_id4_1_1_wenable;
  wire [8:0] ram_w8_l2048_id4_2_0_addr;
  wire [7:0] ram_w8_l2048_id4_2_0_rdata;
  wire [8:0] ram_w8_l2048_id4_2_1_addr;
  wire [7:0] ram_w8_l2048_id4_2_1_rdata;
  wire [7:0] ram_w8_l2048_id4_2_1_wdata;
  wire ram_w8_l2048_id4_2_1_wenable;
  wire [8:0] ram_w8_l2048_id4_3_0_addr;
  wire [7:0] ram_w8_l2048_id4_3_0_rdata;
  wire [8:0] ram_w8_l2048_id4_3_1_addr;
  wire [7:0] ram_w8_l2048_id4_3_1_rdata;
  wire [7:0] ram_w8_l2048_id4_3_1_wdata;
  wire ram_w8_l2048_id4_3_1_wenable;
  wire [8:0] ram_w8_l2048_id5_0_0_addr;
  wire [7:0] ram_w8_l2048_id5_0_0_rdata;
  wire [8:0] ram_w8_l2048_id5_0_1_addr;
  wire [7:0] ram_w8_l2048_id5_0_1_rdata;
  wire [7:0] ram_w8_l2048_id5_0_1_wdata;
  wire ram_w8_l2048_id5_0_1_wenable;
  wire [8:0] ram_w8_l2048_id5_1_0_addr;
  wire [7:0] ram_w8_l2048_id5_1_0_rdata;
  wire [8:0] ram_w8_l2048_id5_1_1_addr;
  wire [7:0] ram_w8_l2048_id5_1_1_rdata;
  wire [7:0] ram_w8_l2048_id5_1_1_wdata;
  wire ram_w8_l2048_id5_1_1_wenable;
  wire [8:0] ram_w8_l2048_id5_2_0_addr;
  wire [7:0] ram_w8_l2048_id5_2_0_rdata;
  wire [8:0] ram_w8_l2048_id5_2_1_addr;
  wire [7:0] ram_w8_l2048_id5_2_1_rdata;
  wire [7:0] ram_w8_l2048_id5_2_1_wdata;
  wire ram_w8_l2048_id5_2_1_wenable;
  wire [8:0] ram_w8_l2048_id5_3_0_addr;
  wire [7:0] ram_w8_l2048_id5_3_0_rdata;
  wire [8:0] ram_w8_l2048_id5_3_1_addr;
  wire [7:0] ram_w8_l2048_id5_3_1_rdata;
  wire [7:0] ram_w8_l2048_id5_3_1_wdata;
  wire ram_w8_l2048_id5_3_1_wenable;
  wire [8:0] ram_w8_l2048_id6_0_0_addr;
  wire [7:0] ram_w8_l2048_id6_0_0_rdata;
  wire [8:0] ram_w8_l2048_id6_0_1_addr;
  wire [7:0] ram_w8_l2048_id6_0_1_rdata;
  wire [7:0] ram_w8_l2048_id6_0_1_wdata;
  wire ram_w8_l2048_id6_0_1_wenable;
  wire [8:0] ram_w8_l2048_id6_1_0_addr;
  wire [7:0] ram_w8_l2048_id6_1_0_rdata;
  wire [8:0] ram_w8_l2048_id6_1_1_addr;
  wire [7:0] ram_w8_l2048_id6_1_1_rdata;
  wire [7:0] ram_w8_l2048_id6_1_1_wdata;
  wire ram_w8_l2048_id6_1_1_wenable;
  wire [8:0] ram_w8_l2048_id6_2_0_addr;
  wire [7:0] ram_w8_l2048_id6_2_0_rdata;
  wire [8:0] ram_w8_l2048_id6_2_1_addr;
  wire [7:0] ram_w8_l2048_id6_2_1_rdata;
  wire [7:0] ram_w8_l2048_id6_2_1_wdata;
  wire ram_w8_l2048_id6_2_1_wenable;
  wire [8:0] ram_w8_l2048_id6_3_0_addr;
  wire [7:0] ram_w8_l2048_id6_3_0_rdata;
  wire [8:0] ram_w8_l2048_id6_3_1_addr;
  wire [7:0] ram_w8_l2048_id6_3_1_rdata;
  wire [7:0] ram_w8_l2048_id6_3_1_wdata;
  wire ram_w8_l2048_id6_3_1_wenable;
  wire [8:0] ram_w8_l2048_id7_0_0_addr;
  wire [7:0] ram_w8_l2048_id7_0_0_rdata;
  wire [8:0] ram_w8_l2048_id7_0_1_addr;
  wire [7:0] ram_w8_l2048_id7_0_1_rdata;
  wire [7:0] ram_w8_l2048_id7_0_1_wdata;
  wire ram_w8_l2048_id7_0_1_wenable;
  wire [8:0] ram_w8_l2048_id7_1_0_addr;
  wire [7:0] ram_w8_l2048_id7_1_0_rdata;
  wire [8:0] ram_w8_l2048_id7_1_1_addr;
  wire [7:0] ram_w8_l2048_id7_1_1_rdata;
  wire [7:0] ram_w8_l2048_id7_1_1_wdata;
  wire ram_w8_l2048_id7_1_1_wenable;
  wire [8:0] ram_w8_l2048_id7_2_0_addr;
  wire [7:0] ram_w8_l2048_id7_2_0_rdata;
  wire [8:0] ram_w8_l2048_id7_2_1_addr;
  wire [7:0] ram_w8_l2048_id7_2_1_rdata;
  wire [7:0] ram_w8_l2048_id7_2_1_wdata;
  wire ram_w8_l2048_id7_2_1_wenable;
  wire [8:0] ram_w8_l2048_id7_3_0_addr;
  wire [7:0] ram_w8_l2048_id7_3_0_rdata;
  wire [8:0] ram_w8_l2048_id7_3_1_addr;
  wire [7:0] ram_w8_l2048_id7_3_1_rdata;
  wire [7:0] ram_w8_l2048_id7_3_1_wdata;
  wire ram_w8_l2048_id7_3_1_wenable;
  wire [8:0] ram_w8_l2048_id8_0_0_addr;
  wire [7:0] ram_w8_l2048_id8_0_0_rdata;
  wire [8:0] ram_w8_l2048_id8_0_1_addr;
  wire [7:0] ram_w8_l2048_id8_0_1_rdata;
  wire [7:0] ram_w8_l2048_id8_0_1_wdata;
  wire ram_w8_l2048_id8_0_1_wenable;
  wire [8:0] ram_w8_l2048_id8_1_0_addr;
  wire [7:0] ram_w8_l2048_id8_1_0_rdata;
  wire [8:0] ram_w8_l2048_id8_1_1_addr;
  wire [7:0] ram_w8_l2048_id8_1_1_rdata;
  wire [7:0] ram_w8_l2048_id8_1_1_wdata;
  wire ram_w8_l2048_id8_1_1_wenable;
  wire [8:0] ram_w8_l2048_id8_2_0_addr;
  wire [7:0] ram_w8_l2048_id8_2_0_rdata;
  wire [8:0] ram_w8_l2048_id8_2_1_addr;
  wire [7:0] ram_w8_l2048_id8_2_1_rdata;
  wire [7:0] ram_w8_l2048_id8_2_1_wdata;
  wire ram_w8_l2048_id8_2_1_wenable;
  wire [8:0] ram_w8_l2048_id8_3_0_addr;
  wire [7:0] ram_w8_l2048_id8_3_0_rdata;
  wire [8:0] ram_w8_l2048_id8_3_1_addr;
  wire [7:0] ram_w8_l2048_id8_3_1_rdata;
  wire [7:0] ram_w8_l2048_id8_3_1_wdata;
  wire ram_w8_l2048_id8_3_1_wenable;
  wire [8:0] ram_w8_l2048_id9_0_0_addr;
  wire [7:0] ram_w8_l2048_id9_0_0_rdata;
  wire [8:0] ram_w8_l2048_id9_0_1_addr;
  wire [7:0] ram_w8_l2048_id9_0_1_rdata;
  wire [7:0] ram_w8_l2048_id9_0_1_wdata;
  wire ram_w8_l2048_id9_0_1_wenable;
  wire [8:0] ram_w8_l2048_id9_1_0_addr;
  wire [7:0] ram_w8_l2048_id9_1_0_rdata;
  wire [8:0] ram_w8_l2048_id9_1_1_addr;
  wire [7:0] ram_w8_l2048_id9_1_1_rdata;
  wire [7:0] ram_w8_l2048_id9_1_1_wdata;
  wire ram_w8_l2048_id9_1_1_wenable;
  wire [8:0] ram_w8_l2048_id9_2_0_addr;
  wire [7:0] ram_w8_l2048_id9_2_0_rdata;
  wire [8:0] ram_w8_l2048_id9_2_1_addr;
  wire [7:0] ram_w8_l2048_id9_2_1_rdata;
  wire [7:0] ram_w8_l2048_id9_2_1_wdata;
  wire ram_w8_l2048_id9_2_1_wenable;
  wire [8:0] ram_w8_l2048_id9_3_0_addr;
  wire [7:0] ram_w8_l2048_id9_3_0_rdata;
  wire [8:0] ram_w8_l2048_id9_3_1_addr;
  wire [7:0] ram_w8_l2048_id9_3_1_rdata;
  wire [7:0] ram_w8_l2048_id9_3_1_wdata;
  wire ram_w8_l2048_id9_3_1_wenable;
  wire [9:0] ram_w8_l4096_id0_0_0_addr;
  wire [7:0] ram_w8_l4096_id0_0_0_rdata;
  wire [9:0] ram_w8_l4096_id0_0_1_addr;
  wire [7:0] ram_w8_l4096_id0_0_1_rdata;
  wire [7:0] ram_w8_l4096_id0_0_1_wdata;
  wire ram_w8_l4096_id0_0_1_wenable;
  wire [9:0] ram_w8_l4096_id0_1_0_addr;
  wire [7:0] ram_w8_l4096_id0_1_0_rdata;
  wire [9:0] ram_w8_l4096_id0_1_1_addr;
  wire [7:0] ram_w8_l4096_id0_1_1_rdata;
  wire [7:0] ram_w8_l4096_id0_1_1_wdata;
  wire ram_w8_l4096_id0_1_1_wenable;
  wire [9:0] ram_w8_l4096_id0_2_0_addr;
  wire [7:0] ram_w8_l4096_id0_2_0_rdata;
  wire [9:0] ram_w8_l4096_id0_2_1_addr;
  wire [7:0] ram_w8_l4096_id0_2_1_rdata;
  wire [7:0] ram_w8_l4096_id0_2_1_wdata;
  wire ram_w8_l4096_id0_2_1_wenable;
  wire [9:0] ram_w8_l4096_id0_3_0_addr;
  wire [7:0] ram_w8_l4096_id0_3_0_rdata;
  wire [9:0] ram_w8_l4096_id0_3_1_addr;
  wire [7:0] ram_w8_l4096_id0_3_1_rdata;
  wire [7:0] ram_w8_l4096_id0_3_1_wdata;
  wire ram_w8_l4096_id0_3_1_wenable;
  wire [8:0] req_block_size_156;
  wire [8:0] req_block_size_213;
  wire [8:0] req_block_size_27;
  wire [8:0] req_block_size_270;
  wire rst_logic;
  wire set_req_157;
  wire set_req_214;
  wire set_req_271;
  wire set_req_28;
  assign _22317_[8:0] = _tmp_44;
  assign _22318_[8:0] = _tmp_45;
  assign _22319_[8:0] = _tmp_46;
  assign _22320_[8:0] = _tmp_47;
  assign _22321_[8:0] = _tmp_48;
  assign _22322_[8:0] = _tmp_49;
  assign _22323_[8:0] = _tmp_50;
  assign _22324_[8:0] = _tmp_51;
  assign _22325_[8:0] = _tmp_52;
  assign _22326_[8:0] = _tmp_75;
  assign _22327_[8:0] = _tmp_76;
  assign _22328_[8:0] = _tmp_77;
  assign _22329_[8:0] = _tmp_78;
  assign _22330_[8:0] = _tmp_79;
  assign _22331_[8:0] = _tmp_80;
  assign _22332_[8:0] = _tmp_81;
  assign _22333_[8:0] = _tmp_82;
  assign _22334_[8:0] = _tmp_83;
  assign _22335_[8:0] = _tmp_106;
  assign _22336_[8:0] = _tmp_107;
  assign _22337_[8:0] = _tmp_108;
  assign _22338_[8:0] = _tmp_109;
  assign _22339_[8:0] = _tmp_110;
  assign _22340_[8:0] = _tmp_111;
  assign _22341_[8:0] = _tmp_112;
  assign _22342_[8:0] = _tmp_113;
  assign _22343_[8:0] = _tmp_114;
  assign _22344_[8:0] = _tmp_137;
  assign _22345_[8:0] = _tmp_138;
  assign _22346_[8:0] = _tmp_139;
  assign _22347_[8:0] = _tmp_140;
  assign _22348_[8:0] = _tmp_141;
  assign _22349_[8:0] = _tmp_142;
  assign _22350_[8:0] = _tmp_143;
  assign _22351_[8:0] = _tmp_144;
  assign _22352_[8:0] = _tmp_145;
  assign _22359_[8:0] = _tmp_167;
  assign _22360_[8:0] = _tmp_168;
  assign _22361_[8:0] = _tmp_169;
  assign _22362_[8:0] = _tmp_180;
  assign _22363_[8:0] = _tmp_181;
  assign _22364_[8:0] = _tmp_182;
  assign _22365_[8:0] = _tmp_193;
  assign _22366_[8:0] = _tmp_194;
  assign _22367_[8:0] = _tmp_195;
  assign _22368_[8:0] = _tmp_206;
  assign _22369_[8:0] = _tmp_207;
  assign _22370_[8:0] = _tmp_208;
  assign _22371_[8:0] = _tmp_224;
  assign _22372_[8:0] = _tmp_225;
  assign _22373_[8:0] = _tmp_226;
  assign _22374_[8:0] = _tmp_237;
  assign _22375_[8:0] = _tmp_238;
  assign _22376_[8:0] = _tmp_239;
  assign _22377_[8:0] = _tmp_250;
  assign _22378_[8:0] = _tmp_251;
  assign _22379_[8:0] = _tmp_252;
  assign _22380_[8:0] = _tmp_263;
  assign _22381_[8:0] = _tmp_264;
  assign _22382_[8:0] = _tmp_265;
  assign _22383_[8:0] = _tmp_281;
  assign _22384_[8:0] = _tmp_282;
  assign _22385_[8:0] = _tmp_283;
  assign _22386_[8:0] = _tmp_294;
  assign _22387_[8:0] = _tmp_295;
  assign _22388_[8:0] = _tmp_296;
  assign _22389_[8:0] = _tmp_307;
  assign _22390_[8:0] = _tmp_308;
  assign _22391_[8:0] = _tmp_309;
  assign _22392_[8:0] = _tmp_320;
  assign _22393_[8:0] = _tmp_321;
  assign _22394_[8:0] = _tmp_322;
  assign _25922_[32:31] = 2'h0;
  assign _25923_[32:31] = 2'h0;
  assign _26323_[32:2] = _25922_[30:0];
  assign _26327_[32:2] = _25923_[30:0];
  assign _26330_[15:0] = 16'h0000;
  assign _26331_[31:0] = 0;
  assign _26335_[49:0] = _26330_[65:16];
  assign _26336_[33:0] = _26331_[65:32];
  assign _26365_[30:23] = { _26365_[31], _26365_[31], _26365_[31], _26365_[31], _26365_[31], _26365_[31], _26365_[31], _26365_[31] };
  assign _26369_[31:8] = { _26365_[31], _26365_[22:0] };
  assign _26371_[38:31] = { _26371_[39], _26371_[39], _26371_[39], _26371_[39], _26371_[39], _26371_[39], _26371_[39], _26371_[39] };
  assign _26375_[39:8] = { _26371_[39], _26371_[30:0] };
  assign _26376_[14:7] = { _26376_[15], _26376_[15], _26376_[15], _26376_[15], _26376_[15], _26376_[15], _26376_[15], _26376_[15] };
  assign _26379_[15:8] = { _26376_[15], _26376_[6:0] };
  assign _26380_[14:7] = { _26380_[15], _26380_[15], _26380_[15], _26380_[15], _26380_[15], _26380_[15], _26380_[15], _26380_[15] };
  assign _26383_[15:8] = { _26380_[15], _26380_[6:0] };
  assign _26384_[14:7] = { _26384_[15], _26384_[15], _26384_[15], _26384_[15], _26384_[15], _26384_[15], _26384_[15], _26384_[15] };
  assign _26387_[15:8] = { _26384_[15], _26384_[6:0] };
  assign _26388_[14:7] = { _26388_[15], _26388_[15], _26388_[15], _26388_[15], _26388_[15], _26388_[15], _26388_[15], _26388_[15] };
  assign _26391_[15:8] = { _26388_[15], _26388_[6:0] };
  assign _26392_[14:7] = { _26392_[15], _26392_[15], _26392_[15], _26392_[15], _26392_[15], _26392_[15], _26392_[15], _26392_[15] };
  assign _26395_[15:8] = { _26392_[15], _26392_[6:0] };
  assign _26396_[14:7] = { _26396_[15], _26396_[15], _26396_[15], _26396_[15], _26396_[15], _26396_[15], _26396_[15], _26396_[15] };
  assign _26399_[15:8] = { _26396_[15], _26396_[6:0] };
  assign _26400_[14:7] = { _26400_[15], _26400_[15], _26400_[15], _26400_[15], _26400_[15], _26400_[15], _26400_[15], _26400_[15] };
  assign _26403_[15:8] = { _26400_[15], _26400_[6:0] };
  assign _26404_[14:7] = { _26404_[15], _26404_[15], _26404_[15], _26404_[15], _26404_[15], _26404_[15], _26404_[15], _26404_[15] };
  assign _26407_[15:8] = { _26404_[15], _26404_[6:0] };
  assign _26408_[14:7] = { _26408_[15], _26408_[15], _26408_[15], _26408_[15], _26408_[15], _26408_[15], _26408_[15], _26408_[15] };
  assign _26411_[15:8] = { _26408_[15], _26408_[6:0] };
  assign _26447_[0] = conv2d_8_mux_next_dma_flag_0;
  assign _26449_[0] = conv2d_8_mux_next_dma_flag_1;
  assign _26452_[0] = conv2d_8_mux_next_dma_flag_2;
  assign _26456_[7:0] = _tmp_870;
  assign _26457_[7:0] = _stream_max_pool_serial_9_source_1_source_ram_rdata;
  assign _26458_[0] = _stream_max_pool_serial_9_start_flag;
  assign _26462_[7:0] = _tmp_1000;
  assign _26463_[7:0] = _stream_matmul_15_source_8_source_ram_rdata;
  assign _26467_[7:0] = _tmp_1020;
  assign _26468_[7:0] = _stream_matmul_15_source_19_source_ram_rdata;
  assign _26472_[7:0] = _tmp_1030;
  assign _26473_[7:0] = _stream_matmul_15_source_20_source_ram_rdata;
  assign _26474_[0] = _stream_matmul_15_start_flag;
  assign _26477_[0] = _maxi_write_data_done;
  assign _26510_[0] = _tmp_7;
  assign _26542_[4:0] = cparam_conv2d_8_act_num_row;
  assign _26543_[4:0] = cparam_conv2d_8_bias_num;
  assign _26544_[3:0] = cparam_conv2d_8_cshamt_out_value;
  assign _26545_[4:0] = cparam_conv2d_8_inc_sync_out;
  assign _26546_[0] = cparam_conv2d_8_pad_col_left;
  assign _26547_[4:0] = cparam_conv2d_8_max_col_count;
  assign _26548_[6:0] = cparam_conv2d_8_och_count_step;
  assign _26549_[7:0] = cparam_conv2d_8_act_read_size;
  assign _26550_[4:0] = cparam_conv2d_8_inc_act_laddr_large;
  assign _26551_[6:0] = cparam_conv2d_8_act_read_step;
  assign _26552_[10:0] = cparam_conv2d_8_filter_base_step;
  assign _26553_[7:0] = cparam_conv2d_8_filter_read_step;
  assign _26554_[8:0] = cparam_conv2d_8_out_row_step;
  assign _26555_[4:0] = cparam_conv2d_8_stream_reduce_size;
  assign _26556_[1:0] = cparam_conv2d_8_col_select_initval;
  assign _26557_[3:0] = cparam_conv2d_8_stream_act_local_large_offset;
  assign _26558_[4:0] = cparam_max_pool_serial_9_act_num_col;
  assign _26559_[4:0] = cparam_max_pool_serial_9_max_col_count;
  assign _26560_[9:0] = cparam_max_pool_serial_9_act_row_step;
  assign _26561_[4:0] = cparam_max_pool_serial_9_inc_out_laddr;
  assign _26562_[7:0] = cparam_max_pool_serial_9_out_row_step;
  assign _26563_[5:0] = cparam_max_pool_serial_9_inc_act_laddr;
  assign _26659_[7:0] = _tmp_344;
  assign _26660_[7:0] = _stream_conv2d_8_source_8_source_ram_rdata;
  assign _26664_[7:0] = _tmp_364;
  assign _26665_[7:0] = _stream_conv2d_8_source_19_source_ram_rdata;
  assign _26669_[7:0] = _tmp_374;
  assign _26670_[7:0] = _stream_conv2d_8_source_20_source_ram_rdata;
  assign _26674_[7:0] = _tmp_384;
  assign _26675_[7:0] = _stream_conv2d_8_source_21_source_ram_rdata;
  assign _26679_[7:0] = _tmp_394;
  assign _26680_[7:0] = _stream_conv2d_8_source_22_source_ram_rdata;
  assign _26684_[7:0] = _tmp_404;
  assign _26685_[7:0] = _stream_conv2d_8_source_23_source_ram_rdata;
  assign _26689_[7:0] = _tmp_414;
  assign _26690_[7:0] = _stream_conv2d_8_source_24_source_ram_rdata;
  assign _26694_[7:0] = _tmp_424;
  assign _26695_[7:0] = _stream_conv2d_8_source_25_source_ram_rdata;
  assign _26699_[7:0] = _tmp_434;
  assign _26700_[7:0] = _stream_conv2d_8_source_26_source_ram_rdata;
  assign _26704_[7:0] = _tmp_444;
  assign _26705_[7:0] = _stream_conv2d_8_source_27_source_ram_rdata;
  assign _26709_[7:0] = _tmp_454;
  assign _26710_[7:0] = _stream_conv2d_8_source_28_source_ram_rdata;
  assign _26714_[7:0] = _tmp_464;
  assign _26715_[7:0] = _stream_conv2d_8_source_29_source_ram_rdata;
  assign _26717_[7:0] = _tmp_474;
  assign _26720_[7:0] = _stream_conv2d_8_source_30_source_ram_rdata;
  assign _26724_[7:0] = _tmp_484;
  assign _26725_[7:0] = _stream_conv2d_8_source_31_source_ram_rdata;
  assign _26729_[7:0] = _tmp_494;
  assign _26730_[7:0] = _stream_conv2d_8_source_32_source_ram_rdata;
  assign _26734_[7:0] = _tmp_504;
  assign _26735_[7:0] = _stream_conv2d_8_source_33_source_ram_rdata;
  assign _26739_[7:0] = _tmp_514;
  assign _26740_[7:0] = _stream_conv2d_8_source_34_source_ram_rdata;
  assign _26744_[7:0] = _tmp_524;
  assign _26745_[7:0] = _stream_conv2d_8_source_35_source_ram_rdata;
  assign _26749_[7:0] = _tmp_534;
  assign _26750_[7:0] = _stream_conv2d_8_source_36_source_ram_rdata;
  assign _26751_[0] = _stream_conv2d_8_start_flag;
  assign maxi_arburst = 2'h1;
  assign maxi_arcache = 4'h3;
  assign maxi_arlock = 1'h0;
  assign maxi_arprot = 3'h0;
  assign maxi_arqos = 4'h0;
  assign maxi_arsize = 3'h2;
  assign maxi_aruser = 2'h0;
  assign maxi_awburst = 2'h1;
  assign maxi_awcache = 4'h3;
  assign maxi_awlock = 1'h0;
  assign maxi_awprot = 3'h0;
  assign maxi_awqos = 4'h0;
  assign maxi_awsize = 3'h2;
  assign maxi_awuser = 2'h0;
  assign maxi_bready = 1'h1;
  assign saxi_bresp = 2'h0;
  assign saxi_rresp = 2'h0;
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _26752_ ( .A({ _05055_, _05874_ }), .Y(_21895_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _26753_ ( .A({ control_max_pool_serial_9[1], _05875_, _05885_, control_max_pool_serial_9[0] }), .Y(_05874_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _26754_ ( .A({ _05884_, _05881_, _05876_ }), .Y(_05875_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26755_ ( .A({ _05880_, _05879_, _05878_, _05877_ }), .Y(_05876_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26756_ ( .A(control_max_pool_serial_9[31:28]), .Y(_05877_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26757_ ( .A({ control_max_pool_serial_9[26:25], control_max_pool_serial_9[23], control_max_pool_serial_9[20] }), .Y(_05878_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26758_ ( .A({ control_max_pool_serial_9[11], control_max_pool_serial_9[8:6] }), .Y(_05879_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26759_ ( .A({ control_max_pool_serial_9[19], control_max_pool_serial_9[16], control_max_pool_serial_9[14:13] }), .Y(_05880_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _26760_ ( .A({ _05883_, _05882_, control_max_pool_serial_9[10:9] }), .Y(_05881_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26761_ ( .A({ control_max_pool_serial_9[27], control_max_pool_serial_9[24], control_max_pool_serial_9[22:21] }), .Y(_05882_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26762_ ( .A({ control_max_pool_serial_9[18:17], control_max_pool_serial_9[15], control_max_pool_serial_9[12] }), .Y(_05883_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _26763_ ( .A({ control_max_pool_serial_9[4], control_max_pool_serial_9[5] }), .Y(_05884_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _26764_ ( .A({ control_max_pool_serial_9[2], control_max_pool_serial_9[3] }), .Y(_05885_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _26765_ ( .A({ control_max_pool_serial_9[1], _05886_, _05887_, control_max_pool_serial_9[0] }), .Y(_05055_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _26766_ ( .A({ _05881_, _05876_, control_max_pool_serial_9[4], control_max_pool_serial_9[5] }), .Y(_05886_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _26767_ ( .A(control_max_pool_serial_9[3:2]), .Y(_05887_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _26768_ ( .A({ _05935_, _05888_ }), .Y(_20226_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26769_ ( .A({ _05932_, _05930_, _05923_, _05889_ }), .Y(_05888_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26770_ ( .A({ _05916_, _05911_, _05906_, _05890_ }), .Y(_05889_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26771_ ( .A({ _20546_, _05891_, _20418_, _05902_ }), .Y(_05890_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26772_ ( .A({ _05901_, _05900_, _05897_, _05892_ }), .Y(_05891_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26773_ ( .A({ _05896_, _05895_, _05894_, _05893_ }), .Y(_05892_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26774_ ( .A(control_conv2d_8[23:20]), .Y(_05893_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26775_ ( .A(control_conv2d_8[19:16]), .Y(_05894_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26776_ ( .A(control_conv2d_8[31:28]), .Y(_05895_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26777_ ( .A(control_conv2d_8[27:24]), .Y(_05896_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _26778_ ( .A({ control_conv2d_8[1], _05898_, _05899_, control_conv2d_8[0] }), .Y(_05897_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26779_ ( .A(control_conv2d_8[15:12]), .Y(_05898_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26780_ ( .A(control_conv2d_8[11:8]), .Y(_05899_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _26781_ ( .A(control_conv2d_8[3:2]), .Y(_05900_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _26782_ ( .A({ control_conv2d_8[5], control_conv2d_8[7:6], control_conv2d_8[4] }), .Y(_05901_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26783_ ( .A({ _05901_, _05904_, _05903_, _05892_ }), .Y(_05902_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _26784_ ( .A({ _05899_, _05898_ }), .Y(_05903_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _26785_ ( .A({ control_conv2d_8[3:2], _05905_ }), .Y(_05904_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _26786_ ( .A(control_conv2d_8[1:0]), .Y(_05905_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _26787_ ( .A({ _20194_, _05119_, _05909_, _20290_ }), .Y(_05906_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _26788_ ( .A({ _05908_, _05907_, _05903_, _05892_ }), .Y(_05119_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _26789_ ( .A({ control_conv2d_8[5:4], control_conv2d_8[7:6] }), .Y(_05907_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _26790_ ( .A({ control_conv2d_8[1:0], control_conv2d_8[2], control_conv2d_8[3] }), .Y(_05908_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26791_ ( .A({ _05910_, _05907_, _05903_, _05892_ }), .Y(_05909_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _26792_ ( .A({ control_conv2d_8[2], control_conv2d_8[0], control_conv2d_8[1], control_conv2d_8[3] }), .Y(_05910_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26793_ ( .A({ _20482_, _05912_, _20354_, _05914_ }), .Y(_05911_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26794_ ( .A({ _05901_, _05913_, _05903_, _05892_ }), .Y(_05912_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _26795_ ( .A({ _05905_, control_conv2d_8[2], control_conv2d_8[3] }), .Y(_05913_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26796_ ( .A({ _05915_, _05901_, _05903_, _05892_ }), .Y(_05914_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _26797_ ( .A({ control_conv2d_8[1], control_conv2d_8[2], control_conv2d_8[3], control_conv2d_8[0] }), .Y(_05915_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26798_ ( .A({ _20738_, _05917_, _05919_, _20802_ }), .Y(_05916_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26799_ ( .A({ _05900_, _05918_, _05897_, _05892_ }), .Y(_05917_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _26800_ ( .A({ control_conv2d_8[4], control_conv2d_8[7:5] }), .Y(_05918_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26801_ ( .A({ _05922_, _05920_, _05903_, _05892_ }), .Y(_05919_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _26802_ ( .A({ control_conv2d_8[1:0], _05921_ }), .Y(_05920_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _26803_ ( .A(control_conv2d_8[3:2]), .Y(_05921_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _26804_ ( .A(control_conv2d_8[7:4]), .Y(_05922_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _26805_ ( .A({ _05924_, _05929_, _20834_ }), .Y(_05923_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26806_ ( .A({ _20322_, _05925_, _05927_, _20770_ }), .Y(_05924_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26807_ ( .A({ _05926_, _05901_, _05903_, _05892_ }), .Y(_05925_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26808_ ( .A({ control_conv2d_8[1:0], control_conv2d_8[3:2] }), .Y(_05926_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26809_ ( .A({ _05928_, _05922_, _05903_, _05892_ }), .Y(_05927_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _26810_ ( .A({ control_conv2d_8[2], control_conv2d_8[0], control_conv2d_8[3], control_conv2d_8[1] }), .Y(_05928_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26811_ ( .A({ _05908_, _05922_, _05903_, _05892_ }), .Y(_05929_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _26812_ ( .A({ _20642_, _05931_, _20898_, _05132_ }), .Y(_05930_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26813_ ( .A({ _05918_, _05920_, _05903_, _05892_ }), .Y(_05931_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _26814_ ( .A({ _05900_, _05922_, _05897_, _05892_ }), .Y(_05132_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26815_ ( .A({ _20706_, _05933_, _20386_, _05934_ }), .Y(_05932_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26816_ ( .A({ _05910_, _05918_, _05903_, _05892_ }), .Y(_05933_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26817_ ( .A({ _05901_, _05928_, _05903_, _05892_ }), .Y(_05934_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26818_ ( .A({ _05947_, _05943_, _05940_, _05936_ }), .Y(_05935_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26819_ ( .A({ _20866_, _05937_, _20258_, _05939_ }), .Y(_05936_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26820_ ( .A({ _05938_, _05922_, _05903_, _05892_ }), .Y(_05937_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _26821_ ( .A({ control_conv2d_8[1], control_conv2d_8[2], control_conv2d_8[0], control_conv2d_8[3] }), .Y(_05938_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26822_ ( .A({ _05907_, _05938_, _05903_, _05892_ }), .Y(_05939_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26823_ ( .A({ _20674_, _05941_, _20610_, _05942_ }), .Y(_05940_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26824_ ( .A({ _05918_, _05938_, _05903_, _05892_ }), .Y(_05941_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26825_ ( .A({ _05918_, _05904_, _05903_, _05892_ }), .Y(_05942_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26826_ ( .A({ _20930_, _05944_, _20578_, _05946_ }), .Y(_05943_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26827_ ( .A({ _05900_, _05922_, _05945_, _05892_ }), .Y(_05944_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _26828_ ( .A({ _05905_, _05899_, _05898_ }), .Y(_05945_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26829_ ( .A({ _05928_, _05918_, _05903_, _05892_ }), .Y(_05946_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26830_ ( .A({ _20514_, _05948_, _20450_, _05950_ }), .Y(_05947_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26831_ ( .A({ _05901_, _05949_, _05903_, _05892_ }), .Y(_05948_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _26832_ ( .A({ control_conv2d_8[1:0], _05900_ }), .Y(_05949_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26833_ ( .A({ _05901_, _05951_, _05903_, _05892_ }), .Y(_05950_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _26834_ ( .A({ _05921_, control_conv2d_8[0], control_conv2d_8[1] }), .Y(_05951_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _26835_ ( .A({ _05962_, _05952_ }), .Y(_20225_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26836_ ( .A({ _05961_, _05960_, _05958_, _05953_ }), .Y(_05952_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26837_ ( .A({ _05957_, _05956_, _05955_, _05954_ }), .Y(_05953_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26838_ ( .A({ _20865_, _05937_, _20801_, _05919_ }), .Y(_05954_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26839_ ( .A({ _20449_, _05950_, _20385_, _05934_ }), .Y(_05955_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26840_ ( .A({ _20289_, _05909_, _05914_, _20353_ }), .Y(_05956_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26841_ ( .A({ _20257_, _05939_, _05917_, _20737_ }), .Y(_05957_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _26842_ ( .A({ _05959_, _05931_, _20641_ }), .Y(_05958_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26843_ ( .A({ _20929_, _05944_, _20481_, _05912_ }), .Y(_05959_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26844_ ( .A({ _20513_, _05948_, _20321_, _05925_ }), .Y(_05960_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26845_ ( .A({ _20609_, _05942_, _20417_, _05902_ }), .Y(_05961_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26846_ ( .A({ _05966_, _05965_, _05964_, _05963_ }), .Y(_05962_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26847_ ( .A({ _20545_, _05891_, _05929_, _20833_ }), .Y(_05963_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26848_ ( .A({ _20673_, _05941_, _05933_, _20705_ }), .Y(_05964_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _26849_ ( .A({ _20577_, _05946_, _20897_, _05132_ }), .Y(_05965_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _26850_ ( .A({ _20193_, _05119_, _05927_, _20769_ }), .Y(_05966_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _26851_ ( .A({ _05977_, _05967_ }), .Y(_20223_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26852_ ( .A({ _05976_, _05975_, _05973_, _05968_ }), .Y(_05967_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26853_ ( .A({ _05972_, _05971_, _05970_, _05969_ }), .Y(_05968_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26854_ ( .A({ _20607_, _05942_, _20543_, _05891_ }), .Y(_05969_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _26855_ ( .A({ _20767_, _05927_, _20895_, _05132_ }), .Y(_05970_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26856_ ( .A({ _20415_, _05902_, _05912_, _20479_ }), .Y(_05971_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26857_ ( .A({ _20575_, _05946_, _05933_, _20703_ }), .Y(_05972_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _26858_ ( .A({ _05974_, _05917_, _20735_ }), .Y(_05973_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _26859_ ( .A({ _20191_, _05119_, _05934_, _20383_ }), .Y(_05974_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26860_ ( .A({ _20927_, _05944_, _20799_, _05919_ }), .Y(_05975_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26861_ ( .A({ _20447_, _05950_, _05929_, _20831_ }), .Y(_05976_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26862_ ( .A({ _05981_, _05980_, _05979_, _05978_ }), .Y(_05977_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26863_ ( .A({ _20863_, _05937_, _20255_, _05939_ }), .Y(_05978_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26864_ ( .A({ _20671_, _05941_, _20511_, _05948_ }), .Y(_05979_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26865_ ( .A({ _20287_, _05909_, _05931_, _20639_ }), .Y(_05980_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26866_ ( .A({ _20351_, _05914_, _20319_, _05925_ }), .Y(_05981_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _26867_ ( .A({ _05992_, _05982_ }), .Y(_20222_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26868_ ( .A({ _05991_, _05990_, _05988_, _05983_ }), .Y(_05982_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26869_ ( .A({ _05987_, _05986_, _05985_, _05984_ }), .Y(_05983_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26870_ ( .A({ _20670_, _05941_, _20478_, _05912_ }), .Y(_05984_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26871_ ( .A({ _20926_, _05944_, _20574_, _05946_ }), .Y(_05985_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26872_ ( .A({ _20510_, _05948_, _20414_, _05902_ }), .Y(_05986_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _26873_ ( .A({ _20638_, _05931_, _20894_, _05132_ }), .Y(_05987_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _26874_ ( .A({ _05989_, _05939_, _20254_ }), .Y(_05988_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26875_ ( .A({ _20542_, _05891_, _20382_, _05934_ }), .Y(_05989_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _26876_ ( .A({ _20862_, _05937_, _20190_, _05119_ }), .Y(_05990_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26877_ ( .A({ _20446_, _05950_, _05929_, _20830_ }), .Y(_05991_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26878_ ( .A({ _05996_, _05995_, _05994_, _05993_ }), .Y(_05992_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26879_ ( .A({ _20286_, _05909_, _05919_, _20798_ }), .Y(_05993_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26880_ ( .A({ _20606_, _05942_, _05917_, _20734_ }), .Y(_05994_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26881_ ( .A({ _20766_, _05927_, _20702_, _05933_ }), .Y(_05995_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26882_ ( .A({ _20350_, _05914_, _20318_, _05925_ }), .Y(_05996_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _26883_ ( .A({ _06007_, _05997_ }), .Y(_20221_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26884_ ( .A({ _06006_, _06005_, _06003_, _05998_ }), .Y(_05997_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26885_ ( .A({ _06002_, _06001_, _06000_, _05999_ }), .Y(_05998_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26886_ ( .A({ _20317_, _05925_, _05933_, _20701_ }), .Y(_05999_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26887_ ( .A({ _20573_, _05946_, _05919_, _20797_ }), .Y(_06000_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26888_ ( .A({ _20413_, _05902_, _05931_, _20637_ }), .Y(_06001_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26889_ ( .A({ _20925_, _05944_, _20381_, _05934_ }), .Y(_06002_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _26890_ ( .A({ _06004_, _05132_, _20893_ }), .Y(_06003_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26891_ ( .A({ _20861_, _05937_, _20285_, _05909_ }), .Y(_06004_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _26892_ ( .A({ _20189_, _05119_, _05929_, _20829_ }), .Y(_06005_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26893_ ( .A({ _20253_, _05939_, _05917_, _20733_ }), .Y(_06006_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26894_ ( .A({ _06011_, _06010_, _06009_, _06008_ }), .Y(_06007_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26895_ ( .A({ _20605_, _05942_, _20477_, _05912_ }), .Y(_06008_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26896_ ( .A({ _20445_, _05950_, _20349_, _05914_ }), .Y(_06009_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26897_ ( .A({ _20541_, _05891_, _05927_, _20765_ }), .Y(_06010_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26898_ ( .A({ _20669_, _05941_, _20509_, _05948_ }), .Y(_06011_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _26899_ ( .A({ _05055_, _06012_ }), .Y(_21896_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26900_ ( .A({ control_max_pool_serial_9[1:0], _05885_, _05875_ }), .Y(_06012_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _26901_ ( .A({ _06023_, _06013_ }), .Y(_20219_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26902_ ( .A({ _06022_, _06021_, _06019_, _06014_ }), .Y(_06013_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26903_ ( .A({ _06018_, _06017_, _06016_, _06015_ }), .Y(_06014_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26904_ ( .A({ _20475_, _05912_, _05919_, _20795_ }), .Y(_06015_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26905_ ( .A({ _20283_, _05909_, _05917_, _20731_ }), .Y(_06016_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26906_ ( .A({ _20411_, _05902_, _20315_, _05925_ }), .Y(_06017_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26907_ ( .A({ _20635_, _05931_, _05933_, _20699_ }), .Y(_06018_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _26908_ ( .A({ _06020_, _05132_, _20891_ }), .Y(_06019_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26909_ ( .A({ _20443_, _05950_, _05929_, _20827_ }), .Y(_06020_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _26910_ ( .A({ _20187_, _05119_, _05927_, _20763_ }), .Y(_06021_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26911_ ( .A({ _20571_, _05946_, _20347_, _05914_ }), .Y(_06022_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26912_ ( .A({ _06027_, _06026_, _06025_, _06024_ }), .Y(_06023_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26913_ ( .A({ _20251_, _05939_, _05944_, _20923_ }), .Y(_06024_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26914_ ( .A({ _20507_, _05948_, _05891_, _20539_ }), .Y(_06025_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26915_ ( .A({ _20859_, _05937_, _20667_, _05941_ }), .Y(_06026_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26916_ ( .A({ _20603_, _05942_, _20379_, _05934_ }), .Y(_06027_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _26917_ ( .A({ _06038_, _06028_ }), .Y(_20220_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26918_ ( .A({ _06037_, _06036_, _06034_, _06029_ }), .Y(_06028_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26919_ ( .A({ _06033_, _06032_, _06031_, _06030_ }), .Y(_06029_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26920_ ( .A({ _20540_, _05891_, _20476_, _05912_ }), .Y(_06030_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26921_ ( .A({ _20860_, _05937_, _20700_, _05933_ }), .Y(_06031_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26922_ ( .A({ _20412_, _05902_, _20348_, _05914_ }), .Y(_06032_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26923_ ( .A({ _20796_, _05919_, _05929_, _20828_ }), .Y(_06033_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _26924_ ( .A({ _06035_, _05946_, _20572_ }), .Y(_06034_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26925_ ( .A({ _20316_, _05925_, _05931_, _20636_ }), .Y(_06035_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _26926_ ( .A({ _20188_, _05119_, _05909_, _20284_ }), .Y(_06036_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26927_ ( .A({ _20444_, _05950_, _05927_, _20764_ }), .Y(_06037_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26928_ ( .A({ _06042_, _06041_, _06040_, _06039_ }), .Y(_06038_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26929_ ( .A({ _20252_, _05939_, _05941_, _20668_ }), .Y(_06039_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26930_ ( .A({ _20604_, _05942_, _05917_, _20732_ }), .Y(_06040_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _26931_ ( .A({ _20924_, _05944_, _20892_, _05132_ }), .Y(_06041_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26932_ ( .A({ _20508_, _05948_, _20380_, _05934_ }), .Y(_06042_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _26933_ ( .A({ _06053_, _06043_ }), .Y(_20218_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26934_ ( .A({ _06052_, _06051_, _06049_, _06044_ }), .Y(_06043_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26935_ ( .A({ _06048_, _06047_, _06046_, _06045_ }), .Y(_06044_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26936_ ( .A({ _20442_, _05950_, _20282_, _05909_ }), .Y(_06045_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26937_ ( .A({ _20922_, _05944_, _20634_, _05931_ }), .Y(_06046_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26938_ ( .A({ _20410_, _05902_, _20378_, _05934_ }), .Y(_06047_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26939_ ( .A({ _20858_, _05937_, _20762_, _05927_ }), .Y(_06048_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _26940_ ( .A({ _06050_, _05917_, _20730_ }), .Y(_06049_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26941_ ( .A({ _20506_, _05948_, _05929_, _20826_ }), .Y(_06050_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26942_ ( .A({ _20250_, _05939_, _05941_, _20666_ }), .Y(_06051_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26943_ ( .A({ _20346_, _05914_, _05919_, _20794_ }), .Y(_06052_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26944_ ( .A({ _06057_, _06056_, _06055_, _06054_ }), .Y(_06053_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26945_ ( .A({ _20570_, _05946_, _05933_, _20698_ }), .Y(_06054_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _26946_ ( .A({ _20474_, _05912_, _20890_, _05132_ }), .Y(_06055_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _26947_ ( .A({ _20538_, _05891_, _20186_, _05119_ }), .Y(_06056_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26948_ ( .A({ _20602_, _05942_, _20314_, _05925_ }), .Y(_06057_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _26949_ ( .A({ _06068_, _06058_ }), .Y(_20217_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26950_ ( .A({ _06067_, _06066_, _06064_, _06059_ }), .Y(_06058_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26951_ ( .A({ _06063_, _06062_, _06061_, _06060_ }), .Y(_06059_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26952_ ( .A({ _20921_, _05944_, _20473_, _05912_ }), .Y(_06060_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26953_ ( .A({ _20249_, _05939_, _05927_, _20761_ }), .Y(_06061_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26954_ ( .A({ _20505_, _05948_, _20409_, _05902_ }), .Y(_06062_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26955_ ( .A({ _20537_, _05891_, _05933_, _20697_ }), .Y(_06063_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _26956_ ( .A({ _06065_, _05929_, _20825_ }), .Y(_06064_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26957_ ( .A({ _20665_, _05941_, _20377_, _05934_ }), .Y(_06065_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _26958_ ( .A({ _20185_, _05119_, _05931_, _20633_ }), .Y(_06066_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _26959_ ( .A({ _20441_, _05950_, _20889_, _05132_ }), .Y(_06067_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26960_ ( .A({ _06072_, _06071_, _06070_, _06069_ }), .Y(_06068_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26961_ ( .A({ _20857_, _05937_, _20729_, _05917_ }), .Y(_06069_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26962_ ( .A({ _20601_, _05942_, _20281_, _05909_ }), .Y(_06070_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26963_ ( .A({ _20569_, _05946_, _05919_, _20793_ }), .Y(_06071_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26964_ ( .A({ _20345_, _05914_, _20313_, _05925_ }), .Y(_06072_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _26965_ ( .A({ _05055_, _13919_, _06012_ }), .Y(_13920_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _26966_ ( .A({ _06083_, _06073_ }), .Y(_20216_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26967_ ( .A({ _06082_, _06081_, _06079_, _06074_ }), .Y(_06073_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26968_ ( .A({ _06078_, _06077_, _06076_, _06075_ }), .Y(_06074_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26969_ ( .A({ _20600_, _05942_, _05927_, _20760_ }), .Y(_06075_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _26970_ ( .A({ _20920_, _05944_, _20888_, _05132_ }), .Y(_06076_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26971_ ( .A({ _20472_, _05912_, _20344_, _05914_ }), .Y(_06077_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26972_ ( .A({ _20856_, _05937_, _20792_, _05919_ }), .Y(_06078_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _26973_ ( .A({ _06080_, _05891_, _20536_ }), .Y(_06079_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26974_ ( .A({ _20312_, _05925_, _05933_, _20696_ }), .Y(_06080_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26975_ ( .A({ _20248_, _05939_, _05917_, _20728_ }), .Y(_06081_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26976_ ( .A({ _20280_, _05909_, _05934_, _20376_ }), .Y(_06082_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26977_ ( .A({ _06087_, _06086_, _06085_, _06084_ }), .Y(_06083_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26978_ ( .A({ _20664_, _05941_, _20568_, _05946_ }), .Y(_06084_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26979_ ( .A({ _20408_, _05902_, _05931_, _20632_ }), .Y(_06085_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _26980_ ( .A({ _20184_, _05119_, _05929_, _20824_ }), .Y(_06086_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26981_ ( .A({ _20504_, _05948_, _20440_, _05950_ }), .Y(_06087_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _26982_ ( .A({ _06098_, _06088_ }), .Y(_20215_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26983_ ( .A({ _06097_, _06096_, _06094_, _06089_ }), .Y(_06088_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26984_ ( .A({ _06093_, _06092_, _06091_, _06090_ }), .Y(_06089_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _26985_ ( .A({ _20887_, _05132_, _20695_, _05933_ }), .Y(_06090_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26986_ ( .A({ _20439_, _05950_, _20407_, _05902_ }), .Y(_06091_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26987_ ( .A({ _20311_, _05925_, _05927_, _20759_ }), .Y(_06092_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26988_ ( .A({ _20919_, _05944_, _20823_, _05929_ }), .Y(_06093_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _26989_ ( .A({ _06095_, _05931_, _20631_ }), .Y(_06094_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26990_ ( .A({ _20599_, _05942_, _20279_, _05909_ }), .Y(_06095_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26991_ ( .A({ _20343_, _05914_, _05934_, _20375_ }), .Y(_06096_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26992_ ( .A({ _20503_, _05948_, _20471_, _05912_ }), .Y(_06097_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26993_ ( .A({ _06102_, _06101_, _06100_, _06099_ }), .Y(_06098_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26994_ ( .A({ _20663_, _05941_, _05917_, _20727_ }), .Y(_06099_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26995_ ( .A({ _20855_, _05937_, _20567_, _05946_ }), .Y(_06100_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _26996_ ( .A({ _20247_, _05939_, _05919_, _20791_ }), .Y(_06101_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _26997_ ( .A({ _20535_, _05891_, _20183_, _05119_ }), .Y(_06102_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _26998_ ( .A({ _06113_, _06103_ }), .Y(_20214_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _26999_ ( .A({ _06112_, _06111_, _06109_, _06104_ }), .Y(_06103_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27000_ ( .A({ _06108_, _06107_, _06106_, _06105_ }), .Y(_06104_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27001_ ( .A({ _20278_, _05909_, _05925_, _20310_ }), .Y(_06105_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27002_ ( .A({ _20246_, _05939_, _20182_, _05119_ }), .Y(_06106_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27003_ ( .A({ _20662_, _05941_, _20502_, _05948_ }), .Y(_06107_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27004_ ( .A({ _20438_, _05950_, _05891_, _20534_ }), .Y(_06108_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27005_ ( .A({ _06110_, _05931_, _20630_ }), .Y(_06109_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27006_ ( .A({ _20726_, _05917_, _20886_, _05132_ }), .Y(_06110_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27007_ ( .A({ _20566_, _05946_, _05927_, _20758_ }), .Y(_06111_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27008_ ( .A({ _20918_, _05944_, _20694_, _05933_ }), .Y(_06112_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27009_ ( .A({ _06117_, _06116_, _06115_, _06114_ }), .Y(_06113_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27010_ ( .A({ _20598_, _05942_, _20406_, _05902_ }), .Y(_06114_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27011_ ( .A({ _20342_, _05914_, _05934_, _20374_ }), .Y(_06115_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27012_ ( .A({ _20790_, _05919_, _05929_, _20822_ }), .Y(_06116_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27013_ ( .A({ _20854_, _05937_, _20470_, _05912_ }), .Y(_06117_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27014_ ( .A({ _06128_, _06118_ }), .Y(_20212_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27015_ ( .A({ _06127_, _06126_, _06124_, _06119_ }), .Y(_06118_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27016_ ( .A({ _06123_, _06122_, _06121_, _06120_ }), .Y(_06119_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27017_ ( .A({ _20276_, _05909_, _05925_, _20308_ }), .Y(_06120_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27018_ ( .A({ _20660_, _05941_, _05933_, _20692_ }), .Y(_06121_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27019_ ( .A({ _20564_, _05946_, _20500_, _05948_ }), .Y(_06122_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27020_ ( .A({ _20180_, _05119_, _05934_, _20372_ }), .Y(_06123_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27021_ ( .A({ _06125_, _05919_, _20788_ }), .Y(_06124_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27022_ ( .A({ _20532_, _05891_, _05927_, _20756_ }), .Y(_06125_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27023_ ( .A({ _20244_, _05939_, _05944_, _20916_ }), .Y(_06126_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27024_ ( .A({ _20724_, _05917_, _05929_, _20820_ }), .Y(_06127_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27025_ ( .A({ _06132_, _06131_, _06130_, _06129_ }), .Y(_06128_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27026_ ( .A({ _20404_, _05902_, _05912_, _20468_ }), .Y(_06129_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27027_ ( .A({ _20436_, _05950_, _20340_, _05914_ }), .Y(_06130_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27028_ ( .A({ _20628_, _05931_, _20884_, _05132_ }), .Y(_06131_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27029_ ( .A({ _20852_, _05937_, _20596_, _05942_ }), .Y(_06132_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27030_ ( .A({ _06143_, _06133_ }), .Y(_20211_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27031_ ( .A({ _06142_, _06141_, _06139_, _06134_ }), .Y(_06133_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27032_ ( .A({ _06138_, _06137_, _06136_, _06135_ }), .Y(_06134_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27033_ ( .A({ _20531_, _05891_, _20179_, _05119_ }), .Y(_06135_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27034_ ( .A({ _20307_, _05925_, _05931_, _20627_ }), .Y(_06136_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27035_ ( .A({ _20659_, _05941_, _05944_, _20915_ }), .Y(_06137_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27036_ ( .A({ _20563_, _05946_, _05917_, _20723_ }), .Y(_06138_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27037_ ( .A({ _06140_, _05942_, _20595_ }), .Y(_06139_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27038_ ( .A({ _20467_, _05912_, _20371_, _05934_ }), .Y(_06140_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27039_ ( .A({ _20499_, _05948_, _20403_, _05902_ }), .Y(_06141_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27040_ ( .A({ _20435_, _05950_, _20339_, _05914_ }), .Y(_06142_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27041_ ( .A({ _06147_, _06146_, _06145_, _06144_ }), .Y(_06143_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27042_ ( .A({ _20275_, _05909_, _05929_, _20819_ }), .Y(_06144_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27043_ ( .A({ _20787_, _05919_, _20691_, _05933_ }), .Y(_06145_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27044_ ( .A({ _20755_, _05927_, _20883_, _05132_ }), .Y(_06146_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27045_ ( .A({ _20851_, _05937_, _20243_, _05939_ }), .Y(_06147_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27046_ ( .A({ _06158_, _06148_ }), .Y(_20210_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27047_ ( .A({ _06157_, _06156_, _06154_, _06149_ }), .Y(_06148_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27048_ ( .A({ _06153_, _06152_, _06151_, _06150_ }), .Y(_06149_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27049_ ( .A({ _20914_, _05944_, _20178_, _05119_ }), .Y(_06150_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27050_ ( .A({ _20498_, _05948_, _05927_, _20754_ }), .Y(_06151_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27051_ ( .A({ _20850_, _05937_, _20242_, _05939_ }), .Y(_06152_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27052_ ( .A({ _20658_, _05941_, _05929_, _20818_ }), .Y(_06153_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27053_ ( .A({ _06155_, _05942_, _20594_ }), .Y(_06154_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27054_ ( .A({ _20338_, _05914_, _20306_, _05925_ }), .Y(_06155_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27055_ ( .A({ _20402_, _05902_, _05912_, _20466_ }), .Y(_06156_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27056_ ( .A({ _20434_, _05950_, _20370_, _05934_ }), .Y(_06157_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27057_ ( .A({ _06162_, _06161_, _06160_, _06159_ }), .Y(_06158_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27058_ ( .A({ _20530_, _05891_, _20274_, _05909_ }), .Y(_06159_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27059_ ( .A({ _20626_, _05931_, _20882_, _05132_ }), .Y(_06160_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27060_ ( .A({ _20562_, _05946_, _05919_, _20786_ }), .Y(_06161_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27061_ ( .A({ _20722_, _05917_, _20690_, _05933_ }), .Y(_06162_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27062_ ( .A({ _06173_, _06163_ }), .Y(_20209_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27063_ ( .A({ _06172_, _06171_, _06169_, _06164_ }), .Y(_06163_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27064_ ( .A({ _06168_, _06167_, _06166_, _06165_ }), .Y(_06164_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27065_ ( .A({ _20401_, _05902_, _20881_, _05132_ }), .Y(_06165_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27066_ ( .A({ _20849_, _05937_, _20561_, _05946_ }), .Y(_06166_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27067_ ( .A({ _20465_, _05912_, _20337_, _05914_ }), .Y(_06167_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27068_ ( .A({ _20721_, _05917_, _05929_, _20817_ }), .Y(_06168_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27069_ ( .A({ _06170_, _05927_, _20753_ }), .Y(_06169_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27070_ ( .A({ _20177_, _05119_, _05925_, _20305_ }), .Y(_06170_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27071_ ( .A({ _20241_, _05939_, _05919_, _20785_ }), .Y(_06171_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27072_ ( .A({ _20913_, _05944_, _20433_, _05950_ }), .Y(_06172_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27073_ ( .A({ _06177_, _06176_, _06175_, _06174_ }), .Y(_06173_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27074_ ( .A({ _20273_, _05909_, _05933_, _20689_ }), .Y(_06174_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27075_ ( .A({ _20497_, _05948_, _05931_, _20625_ }), .Y(_06175_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27076_ ( .A({ _20657_, _05941_, _20529_, _05891_ }), .Y(_06176_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27077_ ( .A({ _20593_, _05942_, _20369_, _05934_ }), .Y(_06177_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27078_ ( .A({ _06188_, _06178_ }), .Y(_20208_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27079_ ( .A({ _06187_, _06186_, _06184_, _06179_ }), .Y(_06178_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27080_ ( .A({ _06183_, _06182_, _06181_, _06180_ }), .Y(_06179_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27081_ ( .A({ _20912_, _05944_, _20784_, _05919_ }), .Y(_06180_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27082_ ( .A({ _20592_, _05942_, _20336_, _05914_ }), .Y(_06181_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27083_ ( .A({ _20528_, _05891_, _20368_, _05934_ }), .Y(_06182_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27084_ ( .A({ _20240_, _05939_, _05941_, _20656_ }), .Y(_06183_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27085_ ( .A({ _06185_, _05927_, _20752_ }), .Y(_06184_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27086_ ( .A({ _20464_, _05912_, _05933_, _20688_ }), .Y(_06185_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27087_ ( .A({ _20432_, _05950_, _20304_, _05925_ }), .Y(_06186_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27088_ ( .A({ _20496_, _05948_, _20400_, _05902_ }), .Y(_06187_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27089_ ( .A({ _06192_, _06191_, _06190_, _06189_ }), .Y(_06188_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27090_ ( .A({ _20848_, _05937_, _20272_, _05909_ }), .Y(_06189_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27091_ ( .A({ _20560_, _05946_, _20880_, _05132_ }), .Y(_06190_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27092_ ( .A({ _20176_, _05119_, _05931_, _20624_ }), .Y(_06191_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27093_ ( .A({ _20720_, _05917_, _05929_, _20816_ }), .Y(_06192_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27094_ ( .A({ _06203_, _06193_ }), .Y(_20207_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27095_ ( .A({ _06202_, _06201_, _06199_, _06194_ }), .Y(_06193_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27096_ ( .A({ _06198_, _06197_, _06196_, _06195_ }), .Y(_06194_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27097_ ( .A({ _20495_, _05948_, _05891_, _20527_ }), .Y(_06195_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27098_ ( .A({ _20559_, _05946_, _05929_, _20815_ }), .Y(_06196_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27099_ ( .A({ _20591_, _05942_, _05931_, _20623_ }), .Y(_06197_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27100_ ( .A({ _20719_, _05917_, _20367_, _05934_ }), .Y(_06198_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _27101_ ( .A({ _06200_, _05132_, _20879_ }), .Y(_06199_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27102_ ( .A({ _20271_, _05909_, _05927_, _20751_ }), .Y(_06200_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27103_ ( .A({ _20239_, _05939_, _20175_, _05119_ }), .Y(_06201_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27104_ ( .A({ _20847_, _05937_, _20783_, _05919_ }), .Y(_06202_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27105_ ( .A({ _06207_, _06206_, _06205_, _06204_ }), .Y(_06203_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27106_ ( .A({ _20399_, _05902_, _20303_, _05925_ }), .Y(_06204_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27107_ ( .A({ _20431_, _05950_, _20335_, _05914_ }), .Y(_06205_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27108_ ( .A({ _20911_, _05944_, _20687_, _05933_ }), .Y(_06206_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27109_ ( .A({ _20655_, _05941_, _20463_, _05912_ }), .Y(_06207_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27110_ ( .A({ _06218_, _06208_ }), .Y(_20206_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27111_ ( .A({ _06217_, _06216_, _06214_, _06209_ }), .Y(_06208_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27112_ ( .A({ _06213_, _06212_, _06211_, _06210_ }), .Y(_06209_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27113_ ( .A({ _20270_, _05909_, _05914_, _20334_ }), .Y(_06210_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27114_ ( .A({ _20526_, _05891_, _20174_, _05119_ }), .Y(_06211_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27115_ ( .A({ _20462_, _05912_, _20878_, _05132_ }), .Y(_06212_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27116_ ( .A({ _20846_, _05937_, _20302_, _05925_ }), .Y(_06213_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27117_ ( .A({ _06215_, _05939_, _20238_ }), .Y(_06214_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27118_ ( .A({ _20654_, _05941_, _05919_, _20782_ }), .Y(_06215_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27119_ ( .A({ _20622_, _05931_, _05933_, _20686_ }), .Y(_06216_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27120_ ( .A({ _20558_, _05946_, _05929_, _20814_ }), .Y(_06217_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27121_ ( .A({ _06222_, _06221_, _06220_, _06219_ }), .Y(_06218_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27122_ ( .A({ _20590_, _05942_, _20398_, _05902_ }), .Y(_06219_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27123_ ( .A({ _20430_, _05950_, _20366_, _05934_ }), .Y(_06220_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27124_ ( .A({ _20910_, _05944_, _20750_, _05927_ }), .Y(_06221_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27125_ ( .A({ _20494_, _05948_, _05917_, _20718_ }), .Y(_06222_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27126_ ( .A({ _06233_, _06223_ }), .Y(_20205_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27127_ ( .A({ _06232_, _06231_, _06229_, _06224_ }), .Y(_06223_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27128_ ( .A({ _06228_, _06227_, _06226_, _06225_ }), .Y(_06224_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27129_ ( .A({ _20557_, _05946_, _05929_, _20813_ }), .Y(_06225_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27130_ ( .A({ _20397_, _05902_, _05912_, _20461_ }), .Y(_06226_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27131_ ( .A({ _20909_, _05944_, _20301_, _05925_ }), .Y(_06227_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27132_ ( .A({ _20237_, _05939_, _05891_, _20525_ }), .Y(_06228_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27133_ ( .A({ _06230_, _05919_, _20781_ }), .Y(_06229_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27134_ ( .A({ _20493_, _05948_, _05933_, _20685_ }), .Y(_06230_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27135_ ( .A({ _20429_, _05950_, _20365_, _05934_ }), .Y(_06231_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27136_ ( .A({ _20589_, _05942_, _20333_, _05914_ }), .Y(_06232_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27137_ ( .A({ _06237_, _06236_, _06235_, _06234_ }), .Y(_06233_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27138_ ( .A({ _20845_, _05937_, _20749_, _05927_ }), .Y(_06234_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _27139_ ( .A({ _20173_, _05119_, _20877_, _05132_ }), .Y(_06235_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27140_ ( .A({ _20653_, _05941_, _20621_, _05931_ }), .Y(_06236_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27141_ ( .A({ _20269_, _05909_, _05917_, _20717_ }), .Y(_06237_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27142_ ( .A({ _06248_, _06238_ }), .Y(_20204_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27143_ ( .A({ _06247_, _06246_, _06244_, _06239_ }), .Y(_06238_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27144_ ( .A({ _06243_, _06242_, _06241_, _06240_ }), .Y(_06239_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27145_ ( .A({ _20652_, _05941_, _05927_, _20748_ }), .Y(_06240_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27146_ ( .A({ _20460_, _05912_, _05917_, _20716_ }), .Y(_06241_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27147_ ( .A({ _20524_, _05891_, _05933_, _20684_ }), .Y(_06242_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27148_ ( .A({ _20268_, _05909_, _20876_, _05132_ }), .Y(_06243_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27149_ ( .A({ _06245_, _05948_, _20492_ }), .Y(_06244_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27150_ ( .A({ _20332_, _05914_, _20300_, _05925_ }), .Y(_06245_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27151_ ( .A({ _20588_, _05942_, _20396_, _05902_ }), .Y(_06246_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27152_ ( .A({ _20428_, _05950_, _20364_, _05934_ }), .Y(_06247_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27153_ ( .A({ _06252_, _06251_, _06250_, _06249_ }), .Y(_06248_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27154_ ( .A({ _20236_, _05939_, _05944_, _20908_ }), .Y(_06249_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27155_ ( .A({ _20556_, _05946_, _05929_, _20812_ }), .Y(_06250_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27156_ ( .A({ _20780_, _05919_, _20620_, _05931_ }), .Y(_06251_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27157_ ( .A({ _20844_, _05937_, _20172_, _05119_ }), .Y(_06252_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27158_ ( .A({ _06263_, _06253_ }), .Y(_20203_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27159_ ( .A({ _06262_, _06261_, _06259_, _06254_ }), .Y(_06253_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27160_ ( .A({ _06258_, _06257_, _06256_, _06255_ }), .Y(_06254_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27161_ ( .A({ _20843_, _05937_, _20779_, _05919_ }), .Y(_06255_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27162_ ( .A({ _20491_, _05948_, _05929_, _20811_ }), .Y(_06256_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27163_ ( .A({ _20235_, _05939_, _05927_, _20747_ }), .Y(_06257_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27164_ ( .A({ _20171_, _05119_, _05931_, _20619_ }), .Y(_06258_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27165_ ( .A({ _06260_, _05942_, _20587_ }), .Y(_06259_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27166_ ( .A({ _20299_, _05925_, _05934_, _20363_ }), .Y(_06260_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27167_ ( .A({ _20427_, _05950_, _05912_, _20459_ }), .Y(_06261_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27168_ ( .A({ _20395_, _05902_, _20331_, _05914_ }), .Y(_06262_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27169_ ( .A({ _06267_, _06266_, _06265_, _06264_ }), .Y(_06263_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27170_ ( .A({ _20523_, _05891_, _20267_, _05909_ }), .Y(_06264_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27171_ ( .A({ _20651_, _05941_, _05917_, _20715_ }), .Y(_06265_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27172_ ( .A({ _20907_, _05944_, _20555_, _05946_ }), .Y(_06266_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27173_ ( .A({ _20875_, _05132_, _20683_, _05933_ }), .Y(_06267_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27174_ ( .A({ _06278_, _06268_ }), .Y(_20233_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27175_ ( .A({ _06277_, _06276_, _06274_, _06269_ }), .Y(_06268_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27176_ ( .A({ _06273_, _06272_, _06271_, _06270_ }), .Y(_06269_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27177_ ( .A({ _20681_, _05941_, _20297_, _05909_ }), .Y(_06270_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27178_ ( .A({ _20425_, _05902_, _20329_, _05925_ }), .Y(_06271_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27179_ ( .A({ _20873_, _05937_, _20457_, _05950_ }), .Y(_06272_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27180_ ( .A({ _20809_, _05919_, _20649_, _05931_ }), .Y(_06273_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _27181_ ( .A({ _06275_, _05132_, _20905_ }), .Y(_06274_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27182_ ( .A({ _20585_, _05946_, _20489_, _05912_ }), .Y(_06275_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27183_ ( .A({ _20361_, _05914_, _05934_, _20393_ }), .Y(_06276_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27184_ ( .A({ _20617_, _05942_, _20521_, _05948_ }), .Y(_06277_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27185_ ( .A({ _06282_, _06281_, _06280_, _06279_ }), .Y(_06278_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27186_ ( .A({ _20937_, _05944_, _20745_, _05917_ }), .Y(_06279_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27187_ ( .A({ _20201_, _05119_, _05927_, _20777_ }), .Y(_06280_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27188_ ( .A({ _20265_, _05939_, _05891_, _20553_ }), .Y(_06281_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27189_ ( .A({ _20841_, _05929_, _20713_, _05933_ }), .Y(_06282_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27190_ ( .A({ _06293_, _06283_ }), .Y(_20232_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27191_ ( .A({ _06292_, _06291_, _06289_, _06284_ }), .Y(_06283_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27192_ ( .A({ _06288_, _06287_, _06286_, _06285_ }), .Y(_06284_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27193_ ( .A({ _20936_, _05944_, _20392_, _05934_ }), .Y(_06285_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27194_ ( .A({ _20840_, _05929_, _20648_, _05931_ }), .Y(_06286_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27195_ ( .A({ _20456_, _05950_, _05919_, _20808_ }), .Y(_06287_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27196_ ( .A({ _20296_, _05909_, _05925_, _20328_ }), .Y(_06288_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _27197_ ( .A({ _06290_, _05132_, _20904_ }), .Y(_06289_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27198_ ( .A({ _20680_, _05941_, _05927_, _20776_ }), .Y(_06290_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27199_ ( .A({ _20872_, _05937_, _20264_, _05939_ }), .Y(_06291_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27200_ ( .A({ _20200_, _05119_, _05933_, _20712_ }), .Y(_06292_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27201_ ( .A({ _06297_, _06296_, _06295_, _06294_ }), .Y(_06293_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27202_ ( .A({ _20520_, _05948_, _20360_, _05914_ }), .Y(_06294_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27203_ ( .A({ _20616_, _05942_, _20488_, _05912_ }), .Y(_06295_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27204_ ( .A({ _20552_, _05891_, _05917_, _20744_ }), .Y(_06296_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27205_ ( .A({ _20584_, _05946_, _20424_, _05902_ }), .Y(_06297_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27206_ ( .A({ _06308_, _06298_ }), .Y(_20231_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27207_ ( .A({ _06307_, _06306_, _06304_, _06299_ }), .Y(_06298_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27208_ ( .A({ _06303_, _06302_, _06301_, _06300_ }), .Y(_06299_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27209_ ( .A({ _20487_, _05912_, _05919_, _20807_ }), .Y(_06300_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27210_ ( .A({ _20295_, _05909_, _05927_, _20775_ }), .Y(_06301_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27211_ ( .A({ _20423_, _05902_, _20391_, _05934_ }), .Y(_06302_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27212_ ( .A({ _20839_, _05929_, _20711_, _05933_ }), .Y(_06303_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27213_ ( .A({ _06305_, _05939_, _20263_ }), .Y(_06304_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27214_ ( .A({ _20583_, _05946_, _20359_, _05914_ }), .Y(_06305_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27215_ ( .A({ _20743_, _05917_, _20903_, _05132_ }), .Y(_06306_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27216_ ( .A({ _20199_, _05119_, _05925_, _20327_ }), .Y(_06307_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27217_ ( .A({ _06312_, _06311_, _06310_, _06309_ }), .Y(_06308_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27218_ ( .A({ _20871_, _05937_, _20679_, _05941_ }), .Y(_06309_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27219_ ( .A({ _20615_, _05942_, _20551_, _05891_ }), .Y(_06310_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27220_ ( .A({ _20935_, _05944_, _20647_, _05931_ }), .Y(_06311_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27221_ ( .A({ _20519_, _05948_, _20455_, _05950_ }), .Y(_06312_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27222_ ( .A({ _06323_, _06313_ }), .Y(_20230_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27223_ ( .A({ _06322_, _06321_, _06319_, _06314_ }), .Y(_06313_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27224_ ( .A({ _06318_, _06317_, _06316_, _06315_ }), .Y(_06314_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27225_ ( .A({ _20294_, _05909_, _05925_, _20326_ }), .Y(_06315_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27226_ ( .A({ _20262_, _05939_, _20198_, _05119_ }), .Y(_06316_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27227_ ( .A({ _20486_, _05912_, _05933_, _20710_ }), .Y(_06317_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27228_ ( .A({ _20454_, _05950_, _05891_, _20550_ }), .Y(_06318_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27229_ ( .A({ _06320_, _05931_, _20646_ }), .Y(_06319_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27230_ ( .A({ _20870_, _05937_, _20838_, _05929_ }), .Y(_06320_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27231_ ( .A({ _20678_, _05941_, _05919_, _20806_ }), .Y(_06321_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27232_ ( .A({ _20582_, _05946_, _20902_, _05132_ }), .Y(_06322_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27233_ ( .A({ _06327_, _06326_, _06325_, _06324_ }), .Y(_06323_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27234_ ( .A({ _20614_, _05942_, _20422_, _05902_ }), .Y(_06324_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27235_ ( .A({ _20358_, _05914_, _05934_, _20390_ }), .Y(_06325_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27236_ ( .A({ _20934_, _05944_, _20774_, _05927_ }), .Y(_06326_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27237_ ( .A({ _20518_, _05948_, _05917_, _20742_ }), .Y(_06327_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _27238_ ( .A({ _06345_, _06335_, _06328_ }), .Y(_20229_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27239_ ( .A({ _06334_, _06333_, _06329_ }), .Y(_06328_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _27240_ ( .A({ _06332_, _06330_, _05917_, _20741_ }), .Y(_06329_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _27241_ ( .A({ _06331_, _05908_, _05938_ }), .Y(_06330_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27242_ ( .A({ _05901_, _05903_, _05892_ }), .Y(_06331_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27243_ ( .A({ _20581_, _05946_, _05931_, _20645_ }), .Y(_06332_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27244_ ( .A({ _20933_, _05944_, _20901_, _05132_ }), .Y(_06333_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27245_ ( .A({ _20261_, _05939_, _05927_, _20773_ }), .Y(_06334_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27246_ ( .A({ _06344_, _06343_, _06340_, _06336_ }), .Y(_06335_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27247_ ( .A({ _06337_, _05937_, _20869_ }), .Y(_06336_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _27248_ ( .A({ _06338_, _06339_, _05901_ }), .Y(_06337_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27249_ ( .A({ _05907_, _05913_, _05903_, _05892_ }), .Y(_06338_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27250_ ( .A({ _05921_, _05945_, _05892_ }), .Y(_06339_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27251_ ( .A({ _06341_, _05891_, _20549_ }), .Y(_06340_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27252_ ( .A({ _05926_, _06342_, _06331_, _05910_ }), .Y(_06341_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27253_ ( .A({ _05918_, _05903_, _05892_ }), .Y(_06342_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27254_ ( .A({ _20517_, _05948_, _20357_, _05914_ }), .Y(_06343_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27255_ ( .A({ _20485_, _05912_, _20325_, _05925_ }), .Y(_06344_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27256_ ( .A({ _06359_, _06356_, _06353_, _06346_ }), .Y(_06345_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27257_ ( .A({ _06350_, _06347_ }), .Y(_06346_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _27258_ ( .A({ _05907_, _06348_, _06349_ }), .Y(_06347_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27259_ ( .A({ _05900_, _05945_, _05892_ }), .Y(_06348_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27260_ ( .A({ _05900_, _05897_, _05892_ }), .Y(_06349_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _27261_ ( .A({ _06351_, _06352_, _05949_ }), .Y(_06350_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27262_ ( .A({ _05907_, _05903_, _05892_ }), .Y(_06351_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _27263_ ( .A({ _05900_, control_conv2d_8[0], control_conv2d_8[1] }), .Y(_06352_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27264_ ( .A({ _06355_, _06354_ }), .Y(_06353_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27265_ ( .A({ _20421_, _05902_, _20389_, _05934_ }), .Y(_06354_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27266_ ( .A({ _20677_, _05941_, _20453_, _05950_ }), .Y(_06355_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27267_ ( .A({ _06358_, _06357_ }), .Y(_06356_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27268_ ( .A({ _20805_, _05919_, _05929_, _20837_ }), .Y(_06357_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27269_ ( .A({ _20613_, _05942_, _05933_, _20709_ }), .Y(_06358_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _27270_ ( .A({ _06363_, _06360_, _05119_, _20197_ }), .Y(_06359_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _27271_ ( .A({ _06361_, _06362_, _05909_, _20293_ }), .Y(_06360_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27272_ ( .A({ _05901_, _06352_, _05903_, _05892_ }), .Y(_06361_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27273_ ( .A({ _05901_, _05900_, _05945_, _05892_ }), .Y(_06362_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _27274_ ( .A({ _06364_, _06331_, _05920_ }), .Y(_06363_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27275_ ( .A({ _05921_, _05901_, _05897_, _05892_ }), .Y(_06364_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _27276_ ( .A({ _06382_, _06369_, _06365_ }), .Y(_20228_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _27277_ ( .A({ _06368_, _06366_, _05948_, _20516_ }), .Y(_06365_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27278_ ( .A({ _06367_, _06350_, _06347_ }), .Y(_06366_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _27279_ ( .A({ _05127_, _06342_, _05913_, _05949_ }), .Y(_06367_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27280_ ( .A({ _05926_, _05922_, _05903_, _05892_ }), .Y(_05127_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27281_ ( .A({ _20356_, _05914_, _20324_, _05925_ }), .Y(_06368_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27282_ ( .A({ _06379_, _06376_, _06370_ }), .Y(_06369_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27283_ ( .A({ _06375_, _06373_, _06372_, _06371_ }), .Y(_06370_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27284_ ( .A({ _20548_, _05891_, _05917_, _20740_ }), .Y(_06371_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27285_ ( .A({ _20260_, _05939_, _05933_, _20708_ }), .Y(_06372_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _27286_ ( .A({ _05126_, _06374_, _05937_, _20868_ }), .Y(_06373_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27287_ ( .A({ _05921_, _05918_, _05897_, _05892_ }), .Y(_06374_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27288_ ( .A({ _05908_, _05918_, _05903_, _05892_ }), .Y(_05126_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27289_ ( .A({ _20932_, _05944_, _20452_, _05950_ }), .Y(_06375_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _27290_ ( .A({ _06378_, _06377_, _05902_, _20420_ }), .Y(_06376_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27291_ ( .A({ _20644_, _05931_, _20900_, _05132_ }), .Y(_06377_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _27292_ ( .A({ _06342_, _06348_, _06352_ }), .Y(_06378_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _27293_ ( .A({ _06381_, _06380_, _05919_, _20804_ }), .Y(_06379_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _27294_ ( .A({ _05124_, _06338_, _05119_, _20196_ }), .Y(_06380_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27295_ ( .A({ _05915_, _05918_, _05903_, _05892_ }), .Y(_05124_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _27296_ ( .A({ _06342_, _06339_, _05951_ }), .Y(_06381_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27297_ ( .A({ _06386_, _06385_, _06384_, _06383_ }), .Y(_06382_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27298_ ( .A({ _20676_, _05941_, _05929_, _20836_ }), .Y(_06383_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27299_ ( .A({ _20484_, _05912_, _20388_, _05934_ }), .Y(_06384_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27300_ ( .A({ _20612_, _05942_, _20292_, _05909_ }), .Y(_06385_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27301_ ( .A({ _20580_, _05946_, _05927_, _20772_ }), .Y(_06386_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _27302_ ( .A({ _06405_, _06399_, _06387_ }), .Y(_20227_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27303_ ( .A({ _06398_, _06397_, _06392_, _06388_ }), .Y(_06387_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _27304_ ( .A({ _06390_, _06389_, _05914_, _20355_ }), .Y(_06388_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27305_ ( .A({ _20195_, _05119_, _05925_, _20323_ }), .Y(_06389_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _27306_ ( .A({ _06391_, _05915_, _05904_ }), .Y(_06390_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27307_ ( .A({ _05922_, _05903_, _05892_ }), .Y(_06391_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27308_ ( .A({ _06396_, _06395_, _06394_, _06393_ }), .Y(_06392_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27309_ ( .A({ _20931_, _05944_, _20547_, _05891_ }), .Y(_06393_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27310_ ( .A({ _20675_, _05941_, _05927_, _20771_ }), .Y(_06394_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27311_ ( .A({ _20899_, _05132_, _20707_, _05933_ }), .Y(_06395_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27312_ ( .A({ _20739_, _05917_, _20643_, _05931_ }), .Y(_06396_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27313_ ( .A({ _20867_, _05937_, _20835_, _05929_ }), .Y(_06397_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27314_ ( .A({ _20451_, _05950_, _05919_, _20803_ }), .Y(_06398_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27315_ ( .A({ _06404_, _06363_, _06401_, _06400_ }), .Y(_06399_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _27316_ ( .A({ _05130_, _06381_, _06391_, _05951_ }), .Y(_06400_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27317_ ( .A({ _05922_, _06339_ }), .Y(_05130_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _27318_ ( .A({ _05126_, _05124_, _06403_, _06402_ }), .Y(_06401_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27319_ ( .A({ _05901_, _06339_ }), .Y(_06402_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27320_ ( .A({ _05921_, _05922_, _05897_, _05892_ }), .Y(_06403_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _27321_ ( .A({ _06374_, _06331_, _05908_ }), .Y(_06404_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27322_ ( .A({ _06409_, _06408_, _06407_, _06406_ }), .Y(_06405_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27323_ ( .A({ _20611_, _05942_, _20515_, _05948_ }), .Y(_06406_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27324_ ( .A({ _20419_, _05902_, _20387_, _05934_ }), .Y(_06407_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27325_ ( .A({ _20259_, _05939_, _05946_, _20579_ }), .Y(_06408_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27326_ ( .A({ _20291_, _05909_, _05912_, _20483_ }), .Y(_06409_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27327_ ( .A({ _06430_, _06423_, _06420_, _06410_ }), .Y(_20224_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27328_ ( .A({ _06419_, _06418_, _06416_, _06411_ }), .Y(_06410_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27329_ ( .A({ _06415_, _06414_, _06413_, _06412_ }), .Y(_06411_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27330_ ( .A({ _20320_, _05925_, _05934_, _20384_ }), .Y(_06412_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27331_ ( .A({ _20864_, _05937_, _20800_, _05919_ }), .Y(_06413_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27332_ ( .A({ _20512_, _05948_, _20448_, _05950_ }), .Y(_06414_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27333_ ( .A({ _20480_, _05912_, _20352_, _05914_ }), .Y(_06415_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27334_ ( .A({ _06417_, _05917_, _20736_ }), .Y(_06416_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27335_ ( .A({ _20192_, _05119_, _05927_, _20768_ }), .Y(_06417_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27336_ ( .A({ _20672_, _05941_, _20896_, _05132_ }), .Y(_06418_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27337_ ( .A({ _20928_, _05944_, _20832_, _05929_ }), .Y(_06419_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _27338_ ( .A({ _06390_, _06421_, _05891_, _20544_ }), .Y(_06420_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _27339_ ( .A({ _05124_, _06422_, _06338_ }), .Y(_06421_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27340_ ( .A({ _05949_, _06351_, _05920_, _06331_ }), .Y(_06422_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27341_ ( .A({ _06429_, _06428_, _06424_ }), .Y(_06423_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _27342_ ( .A({ _06427_, _06425_, _05902_, _20416_ }), .Y(_06424_) );
  \$lut  #( .LUT(16'h1fff), .WIDTH(4) ) _27343_ ( .A({ _06426_, _05922_, _05913_, _05910_ }), .Y(_06425_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27344_ ( .A({ _05903_, _05892_ }), .Y(_06426_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27345_ ( .A({ _20608_, _05942_, _05931_, _20640_ }), .Y(_06427_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27346_ ( .A({ _20576_, _05946_, _05933_, _20704_ }), .Y(_06428_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27347_ ( .A({ _20256_, _05939_, _05909_, _20288_ }), .Y(_06429_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27348_ ( .A({ _06431_, _05122_, _05121_ }), .Y(_06430_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27349_ ( .A({ _05938_, _06331_ }), .Y(_05121_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27350_ ( .A({ _05910_, _06331_ }), .Y(_05122_) );
  \$lut  #( .LUT(16'h035f), .WIDTH(4) ) _27351_ ( .A({ _05949_, _06342_, _06391_, _05913_ }), .Y(_06431_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27352_ ( .A({ _06435_, _06434_, _06433_ }), .Y(_06432_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _27353_ ( .A({ _06361_, _06349_, _05907_ }), .Y(_06433_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27354_ ( .A({ _06352_, _06351_, _05910_, _06331_ }), .Y(_06434_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27355_ ( .A({ _20437_, _05950_, _05912_, _20469_ }), .Y(_06435_) );
  \$lut  #( .LUT(16'h01ff), .WIDTH(4) ) _27356_ ( .A({ _06391_, _05910_, _06352_, _05915_ }), .Y(_06436_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27357_ ( .A({ _06442_, _06441_, _06438_ }), .Y(_06437_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _27358_ ( .A({ _06440_, _06439_, _05919_, _20789_ }), .Y(_06438_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27359_ ( .A({ _20277_, _05909_, _05927_, _20757_ }), .Y(_06439_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _27360_ ( .A({ _06364_, _06331_, _05938_ }), .Y(_06440_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27361_ ( .A({ _20181_, _05119_, _05917_, _20725_ }), .Y(_06441_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27362_ ( .A({ _20629_, _05931_, _05933_, _20693_ }), .Y(_06442_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27363_ ( .A({ _06447_, _06446_, _06445_, _06444_ }), .Y(_06443_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27364_ ( .A({ _20405_, _05902_, _20309_, _05925_ }), .Y(_06444_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _27365_ ( .A({ _05124_, _06374_, _05914_, _20341_ }), .Y(_06445_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27366_ ( .A({ _20917_, _05944_, _20501_, _05948_ }), .Y(_06446_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27367_ ( .A({ _20597_, _05942_, _20373_, _05934_ }), .Y(_06447_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _27368_ ( .A({ _06452_, _06451_, _06450_, _06449_ }), .Y(_06448_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27369_ ( .A({ _20533_, _05891_ }), .Y(_06449_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27370_ ( .A({ _20661_, _05941_, _20565_, _05946_ }), .Y(_06450_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27371_ ( .A({ _20853_, _05937_, _20245_, _05939_ }), .Y(_06451_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27372_ ( .A({ _20821_, _05929_, _20885_, _05132_ }), .Y(_06452_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27373_ ( .A({ _06440_, _06390_, _06347_, _06337_ }), .Y(_06453_) );
  \$lut  #( .LUT(16'h44f0), .WIDTH(4) ) _27374_ ( .A({ _05913_, _05130_, _06425_, _06342_ }), .Y(_06454_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27375_ ( .A({ _05918_, _06339_ }), .Y(_05125_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27376_ ( .A({ _06459_, _06458_, _06457_, _06456_ }), .Y(_06455_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27377_ ( .A({ _20234_, _05939_, _05909_, _20266_ }), .Y(_06456_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27378_ ( .A({ _20298_, _05925_, _05934_, _20362_ }), .Y(_06457_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _27379_ ( .A({ _05124_, _06374_, _05929_, _20810_ }), .Y(_06458_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27380_ ( .A({ _20650_, _05941_, _20618_, _05931_ }), .Y(_06459_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27381_ ( .A({ _06464_, _06463_, _06462_, _06461_ }), .Y(_06460_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27382_ ( .A({ _20170_, _05119_, _05912_, _20458_ }), .Y(_06461_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27383_ ( .A({ _20554_, _05946_, _20522_, _05891_ }), .Y(_06462_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27384_ ( .A({ _20490_, _05948_, _20426_, _05950_ }), .Y(_06463_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27385_ ( .A({ _20394_, _05902_, _05917_, _20714_ }), .Y(_06464_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27386_ ( .A({ _06469_, _06468_, _06467_, _06466_ }), .Y(_06465_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27387_ ( .A({ _20586_, _05942_, _05927_, _20746_ }), .Y(_06466_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27388_ ( .A({ _20330_, _05914_, _20874_, _05132_ }), .Y(_06467_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27389_ ( .A({ _20778_, _05919_, _20682_, _05933_ }), .Y(_06468_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27390_ ( .A({ _20842_, _05937_, _05944_, _20906_ }), .Y(_06469_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27391_ ( .A({ _05942_, _05941_, _05939_, _05937_ }), .Y(_06470_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27392_ ( .A({ _06425_, _06390_, _06378_, _06366_ }), .Y(_06471_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27393_ ( .A({ _06478_, _06473_, _06401_, _06400_ }), .Y(_06472_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27394_ ( .A({ _06477_, _06476_, _06475_, _06474_ }), .Y(_06473_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _27395_ ( .A({ _05119_, _05909_, _05902_, _05891_ }), .Y(_06474_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27396_ ( .A({ _05919_, _05917_, _05914_, _05912_ }), .Y(_06475_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27397_ ( .A({ _06338_, _05927_, _05925_, _05929_ }), .Y(_06476_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _27398_ ( .A({ _05132_, _05934_, _05933_, _05931_ }), .Y(_06477_) );
  \$lut  #( .LUT(16'h001f), .WIDTH(4) ) _27399_ ( .A({ _06374_, _06391_, _06352_, _05949_ }), .Y(_06478_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _27400_ ( .A({ _05048_, _06479_ }), .Y(_21894_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _27401_ ( .A({ _06480_, max_pool_serial_9_comp_fsm[2], max_pool_serial_9_comp_fsm[3] }), .Y(_06479_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27402_ ( .A({ max_pool_serial_9_comp_fsm[1:0], _06486_, _06481_ }), .Y(_06480_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27403_ ( .A({ _06485_, _06484_, _06483_, _06482_ }), .Y(_06481_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27404_ ( .A(max_pool_serial_9_comp_fsm[23:20]), .Y(_06482_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27405_ ( .A(max_pool_serial_9_comp_fsm[19:16]), .Y(_06483_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27406_ ( .A(max_pool_serial_9_comp_fsm[31:28]), .Y(_06484_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27407_ ( .A(max_pool_serial_9_comp_fsm[27:24]), .Y(_06485_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27408_ ( .A({ _06489_, _06488_, _06487_ }), .Y(_06486_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27409_ ( .A(max_pool_serial_9_comp_fsm[15:12]), .Y(_06487_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27410_ ( .A(max_pool_serial_9_comp_fsm[7:4]), .Y(_06488_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27411_ ( .A(max_pool_serial_9_comp_fsm[11:8]), .Y(_06489_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _27412_ ( .A({ _06490_, max_pool_serial_9_comp_fsm[0], _06481_, max_pool_serial_9_comp_fsm[1] }), .Y(_05048_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _27413_ ( .A({ _06486_, max_pool_serial_9_comp_fsm[3:2] }), .Y(_06490_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _27414_ ( .A({ _06491_, _21894_ }), .Y(_21893_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _27415_ ( .A({ _06496_, _04898_, _06495_, _06492_ }), .Y(_06491_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27416_ ( .A({ _06494_, _06493_ }), .Y(_06492_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _27417_ ( .A({ _06481_, max_pool_serial_9_comp_fsm[1] }), .Y(_06493_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _27418_ ( .A({ _06486_, max_pool_serial_9_comp_fsm[2], max_pool_serial_9_comp_fsm[3] }), .Y(_06494_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _27419_ ( .A({ _06480_, max_pool_serial_9_comp_fsm[3:2] }), .Y(_06495_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _27420_ ( .A({ _06490_, _06493_, max_pool_serial_9_comp_fsm[0] }), .Y(_04898_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _27421_ ( .A({ _06497_, _06490_, _06494_ }), .Y(_06496_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _27422_ ( .A({ max_pool_serial_9_comp_fsm[1], _06481_, max_pool_serial_9_comp_fsm[0] }), .Y(_06497_) );
  \$lut  #( .LUT(16'h2fff), .WIDTH(4) ) _27423_ ( .A({ _06499_, _06498_, _04898_, _13674_ }), .Y(_13610_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27424_ ( .A({ _06496_, _05048_, _05046_ }), .Y(_06498_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27425_ ( .A({ max_pool_serial_9_comp_fsm[0], _06492_ }), .Y(_05046_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27426_ ( .A({ _13578_, _06479_, _13642_, _06495_ }), .Y(_06499_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27427_ ( .A({ _06500_, _13658_, _06495_ }), .Y(_13626_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27428_ ( .A({ _13594_, _06479_, _13690_, _04898_ }), .Y(_06500_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _27429_ ( .A({ _06496_, _06502_, _05045_, _06501_ }), .Y(_13599_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _27430_ ( .A({ _13663_, _04898_ }), .Y(_06501_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _27431_ ( .A({ _06492_, max_pool_serial_9_comp_fsm[0] }), .Y(_05045_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27432_ ( .A({ _13567_, _06479_, _13631_, _06495_ }), .Y(_06502_) );
  \$lut  #( .LUT(16'h8fff), .WIDTH(4) ) _27433_ ( .A({ _06503_, _06504_, _06495_, _13653_ }), .Y(_13621_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27434_ ( .A({ _13589_, _06479_, _13685_, _04898_ }), .Y(_06503_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _27435_ ( .A({ _06494_, _06497_, _06493_ }), .Y(_06504_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27436_ ( .A({ _06505_, _13592_, _06479_ }), .Y(_13624_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27437_ ( .A({ _13656_, _06495_, _13688_, _04898_ }), .Y(_06505_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27438_ ( .A({ _06506_, _13593_, _06479_ }), .Y(_13625_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27439_ ( .A({ _13657_, _06495_, _13689_, _04898_ }), .Y(_06506_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27440_ ( .A({ _06507_, _13597_, _06479_ }), .Y(_13629_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27441_ ( .A({ _13661_, _06495_, _13693_, _04898_ }), .Y(_06507_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27442_ ( .A({ _06508_, _13595_, _06479_ }), .Y(_13627_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27443_ ( .A({ _13659_, _06495_, _13691_, _04898_ }), .Y(_06508_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27444_ ( .A({ _06509_, _13660_, _06495_ }), .Y(_13628_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27445_ ( .A({ _13596_, _06479_, _13692_, _04898_ }), .Y(_06509_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27446_ ( .A({ _06510_, _13570_, _06479_ }), .Y(_13602_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27447_ ( .A({ _13634_, _06495_, _13666_, _04898_ }), .Y(_06510_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27448_ ( .A({ _06511_, _13662_, _06495_ }), .Y(_13630_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27449_ ( .A({ _13598_, _06479_, _13694_, _04898_ }), .Y(_06511_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27450_ ( .A({ _06512_, _13632_, _06495_ }), .Y(_13600_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27451_ ( .A({ _13568_, _06479_, _13664_, _04898_ }), .Y(_06512_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27452_ ( .A({ _06513_, _13633_, _06495_ }), .Y(_13601_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27453_ ( .A({ _13569_, _06479_, _13665_, _04898_ }), .Y(_06513_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27454_ ( .A({ _06514_, _13571_, _06479_ }), .Y(_13603_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27455_ ( .A({ _13635_, _06495_, _13667_, _04898_ }), .Y(_06514_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27456_ ( .A({ _06515_, _13575_, _06479_ }), .Y(_13607_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27457_ ( .A({ _13639_, _06495_, _13671_, _04898_ }), .Y(_06515_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27458_ ( .A({ _06516_, _13572_, _06479_ }), .Y(_13604_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27459_ ( .A({ _13636_, _06495_, _13668_, _04898_ }), .Y(_06516_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27460_ ( .A({ _06517_, _13637_, _06495_ }), .Y(_13605_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27461_ ( .A({ _13573_, _06479_, _13669_, _04898_ }), .Y(_06517_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27462_ ( .A({ _06518_, _13574_, _06479_ }), .Y(_13606_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27463_ ( .A({ _13638_, _06495_, _13670_, _04898_ }), .Y(_06518_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27464_ ( .A({ _06519_, _13640_, _06495_ }), .Y(_13608_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27465_ ( .A({ _13576_, _06479_, _13672_, _04898_ }), .Y(_06519_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27466_ ( .A({ _06520_, _13641_, _06495_ }), .Y(_13609_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27467_ ( .A({ _13577_, _06479_, _13673_, _04898_ }), .Y(_06520_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27468_ ( .A({ _06521_, _13579_, _06479_ }), .Y(_13611_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27469_ ( .A({ _13643_, _06495_, _13675_, _04898_ }), .Y(_06521_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27470_ ( .A({ _06522_, _13580_, _06479_ }), .Y(_13612_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27471_ ( .A({ _13644_, _06495_, _13676_, _04898_ }), .Y(_06522_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27472_ ( .A({ _06523_, _13581_, _06479_ }), .Y(_13613_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27473_ ( .A({ _13645_, _06495_, _13677_, _04898_ }), .Y(_06523_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27474_ ( .A({ _06524_, _13582_, _06479_ }), .Y(_13614_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27475_ ( .A({ _13646_, _06495_, _13678_, _04898_ }), .Y(_06524_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27476_ ( .A({ _06525_, _13588_, _06479_ }), .Y(_13620_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27477_ ( .A({ _13652_, _06495_, _13684_, _04898_ }), .Y(_06525_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27478_ ( .A({ _06526_, _13583_, _06479_ }), .Y(_13615_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27479_ ( .A({ _13647_, _06495_, _13679_, _04898_ }), .Y(_06526_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27480_ ( .A({ _06527_, _13584_, _06479_ }), .Y(_13616_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27481_ ( .A({ _13648_, _06495_, _13680_, _04898_ }), .Y(_06527_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27482_ ( .A({ _06528_, _13649_, _06495_ }), .Y(_13617_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27483_ ( .A({ _13585_, _06479_, _13681_, _04898_ }), .Y(_06528_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27484_ ( .A({ _06529_, _13650_, _06495_ }), .Y(_13618_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27485_ ( .A({ _13586_, _06479_, _13682_, _04898_ }), .Y(_06529_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27486_ ( .A({ _06530_, _13651_, _06495_ }), .Y(_13619_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27487_ ( .A({ _13587_, _06479_, _13683_, _04898_ }), .Y(_06530_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27488_ ( .A({ _06531_, _13590_, _06479_ }), .Y(_13622_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27489_ ( .A({ _13654_, _06495_, _13686_, _04898_ }), .Y(_06531_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _27490_ ( .A({ _06532_, _13655_, _06495_ }), .Y(_13623_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27491_ ( .A({ _13591_, _06479_, _13687_, _04898_ }), .Y(_06532_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _27492_ ( .A({ _05043_, _06533_ }), .Y(_21892_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27493_ ( .A({ _06542_, _06539_, _06534_ }), .Y(_06533_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27494_ ( .A({ _06538_, _06537_, _06536_, _06535_ }), .Y(_06534_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27495_ ( .A(_stream_max_pool_serial_9_source_1_source_pat_fsm_0[23:20]), .Y(_06535_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27496_ ( .A(_stream_max_pool_serial_9_source_1_source_pat_fsm_0[19:16]), .Y(_06536_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27497_ ( .A(_stream_max_pool_serial_9_source_1_source_pat_fsm_0[31:28]), .Y(_06537_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27498_ ( .A(_stream_max_pool_serial_9_source_1_source_pat_fsm_0[27:24]), .Y(_06538_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27499_ ( .A({ _06541_, _06540_ }), .Y(_06539_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27500_ ( .A(_stream_max_pool_serial_9_source_1_source_pat_fsm_0[15:12]), .Y(_06540_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27501_ ( .A(_stream_max_pool_serial_9_source_1_source_pat_fsm_0[11:8]), .Y(_06541_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _27502_ ( .A({ _06543_, _stream_max_pool_serial_9_source_1_source_pat_fsm_0[3:2], _stream_max_pool_serial_9_source_1_source_pat_fsm_0[0] }), .Y(_06542_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27503_ ( .A(_stream_max_pool_serial_9_source_1_source_pat_fsm_0[7:4]), .Y(_06543_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27504_ ( .A({ _06544_, _06543_, _06539_, _06534_ }), .Y(_05043_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _27505_ ( .A({ _stream_max_pool_serial_9_source_1_source_pat_fsm_0[0], _stream_max_pool_serial_9_source_1_source_pat_fsm_0[3:1] }), .Y(_06544_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27506_ ( .A({ _13562_, _06545_, _13530_, _05043_ }), .Y(_13498_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _27507_ ( .A({ _06533_, _stream_max_pool_serial_9_source_1_source_pat_fsm_0[1] }), .Y(_06545_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27508_ ( .A({ _13535_, _06545_, _13503_, _05043_ }), .Y(_13471_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27509_ ( .A({ _13546_, _06545_, _13514_, _05043_ }), .Y(_13482_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27510_ ( .A({ _13557_, _06545_, _13525_, _05043_ }), .Y(_13493_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27511_ ( .A({ _13560_, _06545_, _13528_, _05043_ }), .Y(_13496_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27512_ ( .A({ _13561_, _06545_, _13529_, _05043_ }), .Y(_13497_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27513_ ( .A({ _13563_, _06545_, _13531_, _05043_ }), .Y(_13499_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27514_ ( .A({ _13564_, _06545_, _13532_, _05043_ }), .Y(_13500_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27515_ ( .A({ _13565_, _06545_, _13533_, _05043_ }), .Y(_13501_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27516_ ( .A({ _13566_, _06545_, _13534_, _05043_ }), .Y(_13502_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27517_ ( .A({ _13536_, _06545_, _13504_, _05043_ }), .Y(_13472_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27518_ ( .A({ _13537_, _06545_, _13505_, _05043_ }), .Y(_13473_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27519_ ( .A({ _13540_, _06545_, _13508_, _05043_ }), .Y(_13476_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27520_ ( .A({ _13538_, _06545_, _13506_, _05043_ }), .Y(_13474_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27521_ ( .A({ _13539_, _06545_, _13507_, _05043_ }), .Y(_13475_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27522_ ( .A({ _13541_, _06545_, _13509_, _05043_ }), .Y(_13477_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27523_ ( .A({ _13542_, _06545_, _13510_, _05043_ }), .Y(_13478_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27524_ ( .A({ _13549_, _06545_, _13517_, _05043_ }), .Y(_13485_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27525_ ( .A({ _13543_, _06545_, _13511_, _05043_ }), .Y(_13479_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27526_ ( .A({ _13544_, _06545_, _13512_, _05043_ }), .Y(_13480_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27527_ ( .A({ _13545_, _06545_, _13513_, _05043_ }), .Y(_13481_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27528_ ( .A({ _13547_, _06545_, _13515_, _05043_ }), .Y(_13483_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27529_ ( .A({ _13551_, _06545_, _13519_, _05043_ }), .Y(_13487_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27530_ ( .A({ _13548_, _06545_, _13516_, _05043_ }), .Y(_13484_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27531_ ( .A({ _13550_, _06545_, _13518_, _05043_ }), .Y(_13486_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27532_ ( .A({ _13552_, _06545_, _13520_, _05043_ }), .Y(_13488_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27533_ ( .A({ _13554_, _06545_, _13522_, _05043_ }), .Y(_13490_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27534_ ( .A({ _13556_, _06545_, _13524_, _05043_ }), .Y(_13492_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27535_ ( .A({ _13553_, _06545_, _13521_, _05043_ }), .Y(_13489_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27536_ ( .A({ _13555_, _06545_, _13523_, _05043_ }), .Y(_13491_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27537_ ( .A({ _13558_, _06545_, _13526_, _05043_ }), .Y(_13494_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _27538_ ( .A({ _13559_, _06545_, _13527_, _05043_ }), .Y(_13495_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27539_ ( .A({ _06554_, _06553_, _06548_, _06546_ }), .Y(_21891_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _27540_ ( .A({ _06547_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[31:29] }), .Y(_06546_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27541_ ( .A(_stream_max_pool_serial_9_sink_3_sink_fsm_1[28:25]), .Y(_06547_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27542_ ( .A({ _06552_, _06551_, _06550_, _06549_ }), .Y(_06548_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27543_ ( .A(_stream_max_pool_serial_9_sink_3_sink_fsm_1[8:5]), .Y(_06549_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27544_ ( .A(_stream_max_pool_serial_9_sink_3_sink_fsm_1[4:1]), .Y(_06550_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27545_ ( .A(_stream_max_pool_serial_9_sink_3_sink_fsm_1[16:13]), .Y(_06551_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27546_ ( .A(_stream_max_pool_serial_9_sink_3_sink_fsm_1[12:9]), .Y(_06552_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27547_ ( .A(_stream_max_pool_serial_9_sink_3_sink_fsm_1[24:21]), .Y(_06553_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27548_ ( .A(_stream_max_pool_serial_9_sink_3_sink_fsm_1[20:17]), .Y(_06554_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27549_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13386_, _13450_ }), .Y(_13418_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27550_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13401_, _13465_ }), .Y(_13433_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27551_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13375_, _13439_ }), .Y(_13407_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27552_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13397_, _13461_ }), .Y(_13429_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27553_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13400_, _13464_ }), .Y(_13432_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27554_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13402_, _13466_ }), .Y(_13434_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27555_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13403_, _13467_ }), .Y(_13435_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27556_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13404_, _13468_ }), .Y(_13436_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27557_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13405_, _13469_ }), .Y(_13437_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27558_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13406_, _13470_ }), .Y(_13438_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27559_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13376_, _13440_ }), .Y(_13408_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27560_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13377_, _13441_ }), .Y(_13409_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27561_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13378_, _13442_ }), .Y(_13410_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27562_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13382_, _13446_ }), .Y(_13414_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27563_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13385_, _13449_ }), .Y(_13417_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27564_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13379_, _13443_ }), .Y(_13411_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27565_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13380_, _13444_ }), .Y(_13412_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27566_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13381_, _13445_ }), .Y(_13413_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27567_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13383_, _13447_ }), .Y(_13415_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27568_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13384_, _13448_ }), .Y(_13416_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27569_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13389_, _13453_ }), .Y(_13421_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27570_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13387_, _13451_ }), .Y(_13419_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27571_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13388_, _13452_ }), .Y(_13420_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27572_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13390_, _13454_ }), .Y(_13422_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27573_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13391_, _13455_ }), .Y(_13423_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27574_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13395_, _13459_ }), .Y(_13427_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27575_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13392_, _13456_ }), .Y(_13424_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27576_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13396_, _13460_ }), .Y(_13428_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27577_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13393_, _13457_ }), .Y(_13425_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27578_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13394_, _13458_ }), .Y(_13426_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27579_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13398_, _13462_ }), .Y(_13430_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27580_ ( .A({ _21891_, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _13399_, _13463_ }), .Y(_13431_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27581_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16455_, _16487_ }), .Y(_16423_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _27582_ ( .A({ _06556_, _06564_, _stream_conv2d_8_source_26_source_pat_fsm_9[1] }), .Y(_06555_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27583_ ( .A({ _06563_, _06562_, _06557_ }), .Y(_06556_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27584_ ( .A({ _06561_, _06560_, _06559_, _06558_ }), .Y(_06557_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27585_ ( .A(_stream_conv2d_8_source_26_source_pat_fsm_9[23:20]), .Y(_06558_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27586_ ( .A(_stream_conv2d_8_source_26_source_pat_fsm_9[19:16]), .Y(_06559_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27587_ ( .A(_stream_conv2d_8_source_26_source_pat_fsm_9[31:28]), .Y(_06560_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27588_ ( .A(_stream_conv2d_8_source_26_source_pat_fsm_9[27:24]), .Y(_06561_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27589_ ( .A(_stream_conv2d_8_source_26_source_pat_fsm_9[15:12]), .Y(_06562_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27590_ ( .A(_stream_conv2d_8_source_26_source_pat_fsm_9[11:8]), .Y(_06563_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _27591_ ( .A({ _06565_, _stream_conv2d_8_source_26_source_pat_fsm_9[3:2] }), .Y(_06564_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27592_ ( .A(_stream_conv2d_8_source_26_source_pat_fsm_9[7:4]), .Y(_06565_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27593_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16454_, _16486_ }), .Y(_16422_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27594_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16450_, _16482_ }), .Y(_16418_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27595_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16439_, _16471_ }), .Y(_16407_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _27596_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16428_, _16460_ }), .Y(_16396_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _27597_ ( .A({ _05080_, _06555_ }), .Y(_21911_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _27598_ ( .A({ _stream_conv2d_8_source_26_source_pat_fsm_9[1], _06556_, _06564_, _stream_conv2d_8_source_26_source_pat_fsm_9[0] }), .Y(_05080_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _27599_ ( .A({ _06584_, _06567_ }), .Y(_06566_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _27600_ ( .A({ _06568_, _06576_, _06573_, control_matmul_15[5] }), .Y(_06567_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27601_ ( .A({ _06572_, _06571_, _06570_, _06569_ }), .Y(_06568_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _27602_ ( .A(control_matmul_15[7:6]), .Y(_06569_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27603_ ( .A(control_matmul_15[19:16]), .Y(_06570_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27604_ ( .A(control_matmul_15[31:28]), .Y(_06571_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27605_ ( .A({ control_matmul_15[26:25], control_matmul_15[23], control_matmul_15[20] }), .Y(_06572_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _27606_ ( .A({ _06574_, _06575_, control_matmul_15[4] }), .Y(_06573_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27607_ ( .A(control_matmul_15[15:12]), .Y(_06574_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27608_ ( .A(control_matmul_15[11:8]), .Y(_06575_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _27609_ ( .A({ control_matmul_15[27], control_matmul_15[24], control_matmul_15[22:21] }), .Y(_06576_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _27610_ ( .A({ control_matmul_15[2], control_matmul_15[3] }), .Y(_06577_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27611_ ( .A({ _06579_, _06567_ }), .Y(_06578_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27612_ ( .A({ control_matmul_15[0], control_matmul_15[1], _06580_ }), .Y(_06579_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _27613_ ( .A({ control_matmul_15[2], control_matmul_15[3] }), .Y(_06580_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27614_ ( .A({ _06582_, _06567_ }), .Y(_06581_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27615_ ( .A({ _06583_, _06580_ }), .Y(_06582_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _27616_ ( .A(control_matmul_15[1:0]), .Y(_06583_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _27617_ ( .A({ _06568_, _06576_, _06585_, control_matmul_15[5] }), .Y(_06584_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27618_ ( .A({ control_matmul_15[4], _06575_, _06574_ }), .Y(_06585_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _27619_ ( .A({ _06577_, control_matmul_15[0], control_matmul_15[1] }), .Y(_06586_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27620_ ( .A({ _06587_, _06567_ }), .Y(_05042_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27621_ ( .A({ _06583_, _06577_ }), .Y(_06587_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27622_ ( .A({ _06589_, _06583_, _06584_ }), .Y(_06588_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27623_ ( .A({ control_matmul_15[2], control_matmul_15[3] }), .Y(_06589_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27624_ ( .A({ _06591_, _06583_, _06567_ }), .Y(_06590_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _27625_ ( .A(control_matmul_15[3:2]), .Y(_06591_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27626_ ( .A({ _06593_, _06567_ }), .Y(_06592_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27627_ ( .A({ control_matmul_15[0], control_matmul_15[1], _06591_ }), .Y(_06593_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27628_ ( .A({ _06595_, _06584_ }), .Y(_06594_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _27629_ ( .A({ control_matmul_15[0], _06580_, control_matmul_15[1] }), .Y(_06595_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27630_ ( .A({ control_matmul_15[0], control_matmul_15[1], _06589_, _06584_ }), .Y(_06596_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27631_ ( .A({ _06597_, _06567_ }), .Y(_05041_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27632_ ( .A({ control_matmul_15[0], control_matmul_15[1], _06577_ }), .Y(_06597_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _27633_ ( .A({ control_matmul_15[0], _06584_, _06577_, control_matmul_15[1] }), .Y(_06598_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27634_ ( .A({ control_matmul_15[0], control_matmul_15[1], _06589_, _06567_ }), .Y(_06599_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _27635_ ( .A({ control_matmul_15[0], _06567_, _06589_, control_matmul_15[1] }), .Y(_06600_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27636_ ( .A({ _06576_, _06602_, _06568_ }), .Y(_06601_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _27637_ ( .A({ control_matmul_15[5], _06574_, _06575_, control_matmul_15[4] }), .Y(_06602_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27638_ ( .A({ _06586_, _06567_ }), .Y(_06603_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27639_ ( .A({ _06605_, _06584_ }), .Y(_06604_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _27640_ ( .A({ _06580_, control_matmul_15[0], control_matmul_15[1] }), .Y(_06605_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _27641_ ( .A({ _06567_, _06605_, _06595_ }), .Y(_06606_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _27642_ ( .A({ _06608_, _05039_, _06584_, _06587_ }), .Y(_06607_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _27643_ ( .A({ _06589_, _06583_, _06567_ }), .Y(_05039_) );
  \$lut  #( .LUT(16'h9fff), .WIDTH(4) ) _27644_ ( .A({ _06583_, _06584_, control_matmul_15[2], control_matmul_15[3] }), .Y(_06608_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27645_ ( .A({ _06610_, _11896_, _12906_ }), .Y(_06609_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27646_ ( .A({ 1'h0, _06611_, _12874_, _06612_ }), .Y(_06610_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27647_ ( .A({ _06576_, _06605_, _06602_, _06568_ }), .Y(_06611_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27648_ ( .A({ _06576_, _06602_, _06582_, _06568_ }), .Y(_06612_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27649_ ( .A({ _06576_, _06602_, _06595_, _06568_ }), .Y(_11896_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27650_ ( .A({ _06576_, _06602_, _06579_, _06568_ }), .Y(_05035_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27651_ ( .A({ _06621_, _06617_, _06615_, _06614_ }), .Y(_06613_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27652_ ( .A({ _13258_, _06578_, _06598_, _13162_ }), .Y(_06614_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27653_ ( .A({ _13194_, _06600_, _06616_, _13002_ }), .Y(_06615_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _27654_ ( .A({ control_matmul_15[0], _06584_, _06589_, control_matmul_15[1] }), .Y(_06616_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _27655_ ( .A({ _06619_, _06618_, _06620_, _13066_ }), .Y(_06617_) );
  \$lut  #( .LUT(16'h6000), .WIDTH(4) ) _27656_ ( .A({ _06577_, _06601_, control_matmul_15[0], control_matmul_15[1] }), .Y(_06618_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _27657_ ( .A({ control_matmul_15[0], _06567_, _06591_, control_matmul_15[1] }), .Y(_06619_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _27658_ ( .A({ control_matmul_15[0], _06584_, _06591_, control_matmul_15[1] }), .Y(_06620_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27659_ ( .A({ _12938_, _06596_, _06622_, _13034_ }), .Y(_06621_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _27660_ ( .A({ _06589_, _06584_, control_matmul_15[0], control_matmul_15[1] }), .Y(_06622_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27661_ ( .A({ _13322_, _05042_, _06592_, _13226_ }), .Y(_06623_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27662_ ( .A({ _13098_, _06594_, _06604_, _13130_ }), .Y(_06624_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27663_ ( .A({ _13290_, _06581_, _06588_, _12970_ }), .Y(_06625_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _27664_ ( .A({ _06637_, _06632_, _06626_ }), .Y(_12831_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27665_ ( .A({ _06631_, _06629_, _06627_, _06607_ }), .Y(_06626_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27666_ ( .A({ _06628_, _06611_, 1'h1 }), .Y(_06627_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27667_ ( .A({ _12895_, _11896_, _06612_, _12863_ }), .Y(_06628_) );
  \$lut  #( .LUT(16'hbf00), .WIDTH(4) ) _27668_ ( .A({ _05040_, _06601_, _06577_, control_matmul_15[0] }), .Y(_06629_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _27669_ ( .A({ _06630_, _06567_ }), .Y(_05040_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _27670_ ( .A({ _06591_, control_matmul_15[0], control_matmul_15[1] }), .Y(_06630_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27671_ ( .A({ _06605_, _06567_, _12799_, _05035_ }), .Y(_06631_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27672_ ( .A({ _06636_, _06635_, _06634_, _06633_ }), .Y(_06632_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27673_ ( .A({ _13215_, _06592_, _06598_, _13151_ }), .Y(_06633_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _27674_ ( .A({ _05038_, _06590_, _06588_, _12959_ }), .Y(_06634_) );
  \$lut  #( .LUT(16'hefff), .WIDTH(4) ) _27675_ ( .A({ _06589_, _06567_, control_matmul_15[0], control_matmul_15[1] }), .Y(_05038_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27676_ ( .A({ _13279_, _06581_, _06594_, _13087_ }), .Y(_06635_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27677_ ( .A({ _13311_, _05042_, _06622_, _13023_ }), .Y(_06636_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27678_ ( .A({ _06642_, _06641_, _06640_, _06638_ }), .Y(_06637_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27679_ ( .A({ _06639_, _06596_, _12927_ }), .Y(_06638_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _27680_ ( .A({ _06584_, _06630_, _06586_ }), .Y(_06639_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27681_ ( .A({ _13119_, _06604_, _06616_, _12991_ }), .Y(_06640_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27682_ ( .A({ _13247_, _06578_, _06620_, _13055_ }), .Y(_06641_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27683_ ( .A({ _13343_, _06603_, _06600_, _13183_ }), .Y(_06642_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27684_ ( .A({ _12890_, _06612_, _12826_, _05035_ }), .Y(_06643_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27685_ ( .A({ _12922_, _11896_, _06611_, 1'h1 }), .Y(_06644_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27686_ ( .A({ _06646_, _06588_, _12986_ }), .Y(_06645_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27687_ ( .A({ _13018_, _06616_, _13082_, _06620_ }), .Y(_06646_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27688_ ( .A({ _06651_, _06650_, _06649_, _06648_ }), .Y(_06647_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27689_ ( .A({ _13242_, _06592_, _13370_, _06603_ }), .Y(_06648_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27690_ ( .A({ _13114_, _06594_, _06596_, _12954_ }), .Y(_06649_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27691_ ( .A({ _13146_, _06604_, _06622_, _13050_ }), .Y(_06650_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27692_ ( .A({ _13306_, _06581_, _06600_, _13210_ }), .Y(_06651_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27693_ ( .A({ _06653_, _11896_, _12917_ }), .Y(_06652_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27694_ ( .A({ _12885_, _06612_, _12821_, _05035_ }), .Y(_06653_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27695_ ( .A({ _06658_, _06657_, _06656_, _06655_ }), .Y(_06654_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27696_ ( .A({ _12981_, _06588_, _06622_, _13045_ }), .Y(_06655_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27697_ ( .A({ _12949_, _06596_, _13013_, _06616_ }), .Y(_06656_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27698_ ( .A({ _06606_, _06581_, _13301_ }), .Y(_06657_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27699_ ( .A({ _13237_, _06592_, _06594_, _13109_ }), .Y(_06658_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _27700_ ( .A({ _06663_, _06662_, _06661_, _06660_ }), .Y(_06659_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27701_ ( .A({ _13141_, _06604_ }), .Y(_06660_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27702_ ( .A({ _13269_, _06578_, _06600_, _13205_ }), .Y(_06661_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27703_ ( .A({ _13173_, _06598_, _06620_, _13077_ }), .Y(_06662_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27704_ ( .A({ _13333_, _05042_, _13365_, _06603_ }), .Y(_06663_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27705_ ( .A({ _06665_, _06611_, 1'h0 }), .Y(_06664_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27706_ ( .A({ _12888_, _06612_, _12824_, _05035_ }), .Y(_06665_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27707_ ( .A({ _06670_, _06669_, _06668_, _06667_ }), .Y(_06666_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27708_ ( .A({ _13304_, _06581_, _06620_, _13080_ }), .Y(_06667_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27709_ ( .A({ _13240_, _06592_, _06616_, _13016_ }), .Y(_06668_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _27710_ ( .A({ _05038_, _06590_, _06594_, _13112_ }), .Y(_06669_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27711_ ( .A({ _13336_, _05042_, _06596_, _12952_ }), .Y(_06670_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _27712_ ( .A({ _06675_, _06674_, _06673_, _06672_ }), .Y(_06671_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27713_ ( .A({ _13208_, _06600_ }), .Y(_06672_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27714_ ( .A({ _13176_, _06598_, _06622_, _13048_ }), .Y(_06673_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27715_ ( .A({ _13272_, _06578_, _06604_, _13144_ }), .Y(_06674_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27716_ ( .A({ _12984_, _06588_, _13368_, _06603_ }), .Y(_06675_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _27717_ ( .A({ _06677_, _06611_, 1'h0 }), .Y(_06676_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27718_ ( .A({ _12889_, _06612_, _12825_, _05035_ }), .Y(_06677_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27719_ ( .A({ _06682_, _06681_, _06680_, _06679_ }), .Y(_06678_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27720_ ( .A({ _12985_, _06588_, _06622_, _13049_ }), .Y(_06679_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27721_ ( .A({ _13113_, _06594_, _06604_, _13145_ }), .Y(_06680_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _27722_ ( .A({ _06639_, _05042_, _13337_ }), .Y(_06681_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27723_ ( .A({ _13305_, _06581_, _06620_, _13081_ }), .Y(_06682_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _27724_ ( .A({ _06687_, _06686_, _06685_, _06684_ }), .Y(_06683_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _27725_ ( .A({ _13369_, _06603_ }), .Y(_06684_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27726_ ( .A({ _13241_, _06592_, _06596_, _12953_ }), .Y(_06685_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27727_ ( .A({ _13209_, _06600_, _06616_, _13017_ }), .Y(_06686_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27728_ ( .A({ _13273_, _06578_, _06598_, _13177_ }), .Y(_06687_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27729_ ( .A({ _06698_, _06697_, _06692_, _06688_ }), .Y(_12859_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27730_ ( .A({ _06691_, _06690_, _06689_ }), .Y(_06688_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27731_ ( .A({ _13307_, _06581_, _06600_, _13211_ }), .Y(_06689_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27732_ ( .A({ 1'h0, _06611_, _12891_, _06612_ }), .Y(_06690_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27733_ ( .A({ _12923_, _11896_, _12827_, _05035_ }), .Y(_06691_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27734_ ( .A({ _06696_, _06695_, _06694_, _06693_ }), .Y(_06692_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27735_ ( .A({ _13243_, _06592_, _06604_, _13147_ }), .Y(_06693_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27736_ ( .A({ _13275_, _06578_, _13371_, _06603_ }), .Y(_06694_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27737_ ( .A({ _12955_, _06596_, _13179_, _06598_ }), .Y(_06695_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27738_ ( .A({ _13339_, _05042_, _06588_, _12987_ }), .Y(_06696_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27739_ ( .A({ _13019_, _06616_, _06622_, _13051_ }), .Y(_06697_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27740_ ( .A({ _13115_, _06594_, _06620_, _13083_ }), .Y(_06698_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27741_ ( .A({ _06709_, _06708_, _06703_, _06699_ }), .Y(_12860_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27742_ ( .A({ _06702_, _06701_, _06700_ }), .Y(_06699_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27743_ ( .A({ _13180_, _06598_, _06604_, _13148_ }), .Y(_06700_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27744_ ( .A({ _12924_, _11896_, _06612_, _12892_ }), .Y(_06701_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27745_ ( .A({ 1'h0, _06611_, _12828_, _05035_ }), .Y(_06702_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27746_ ( .A({ _06707_, _06706_, _06705_, _06704_ }), .Y(_06703_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27747_ ( .A({ _13372_, _06603_, _06600_, _13212_ }), .Y(_06704_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27748_ ( .A({ _13084_, _06620_, _06622_, _13052_ }), .Y(_06705_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27749_ ( .A({ _13340_, _05042_, _06592_, _13244_ }), .Y(_06706_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27750_ ( .A({ _13276_, _06578_, _06616_, _13020_ }), .Y(_06707_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27751_ ( .A({ _12988_, _06588_, _13116_, _06594_ }), .Y(_06708_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27752_ ( .A({ _13308_, _06581_, _06596_, _12956_ }), .Y(_06709_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27753_ ( .A({ _06720_, _06719_, _06714_, _06710_ }), .Y(_12833_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27754_ ( .A({ _06713_, _06712_, _06711_ }), .Y(_06710_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27755_ ( .A({ _13313_, _05042_, _06600_, _13185_ }), .Y(_06711_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27756_ ( .A({ _12897_, _11896_, _06611_, 1'h0 }), .Y(_06712_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27757_ ( .A({ _12865_, _06612_, _12801_, _05035_ }), .Y(_06713_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27758_ ( .A({ _06718_, _06717_, _06716_, _06715_ }), .Y(_06714_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27759_ ( .A({ _13249_, _06578_, _06620_, _13057_ }), .Y(_06715_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27760_ ( .A({ _12929_, _06596_, _13345_, _06603_ }), .Y(_06716_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27761_ ( .A({ _12961_, _06588_, _13217_, _06592_ }), .Y(_06717_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27762_ ( .A({ _13281_, _06581_, _06622_, _13025_ }), .Y(_06718_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27763_ ( .A({ _13153_, _06598_, _06616_, _12993_ }), .Y(_06719_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27764_ ( .A({ _13089_, _06594_, _06604_, _13121_ }), .Y(_06720_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27765_ ( .A({ _06731_, _06730_, _06725_, _06721_ }), .Y(_12861_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27766_ ( .A({ _06724_, _06723_, _06722_ }), .Y(_06721_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27767_ ( .A({ _13181_, _06598_, _06604_, _13149_ }), .Y(_06722_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27768_ ( .A({ _12925_, _11896_, _06612_, _12893_ }), .Y(_06723_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27769_ ( .A({ 1'h0, _06611_, _12829_, _05035_ }), .Y(_06724_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27770_ ( .A({ _06729_, _06728_, _06727_, _06726_ }), .Y(_06725_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27771_ ( .A({ _13373_, _06603_, _06600_, _13213_ }), .Y(_06726_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27772_ ( .A({ _13085_, _06620_, _06622_, _13053_ }), .Y(_06727_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27773_ ( .A({ _13341_, _05042_, _06592_, _13245_ }), .Y(_06728_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27774_ ( .A({ _13277_, _06578_, _06616_, _13021_ }), .Y(_06729_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27775_ ( .A({ _12989_, _06588_, _13117_, _06594_ }), .Y(_06730_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27776_ ( .A({ _13309_, _06581_, _06596_, _12957_ }), .Y(_06731_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27777_ ( .A({ _06742_, _06741_, _06736_, _06732_ }), .Y(_12862_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27778_ ( .A({ _06735_, _06734_, _06733_ }), .Y(_06732_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27779_ ( .A({ _13278_, _06578_, _06600_, _13214_ }), .Y(_06733_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27780_ ( .A({ 1'h0, _06611_, _12830_, _05035_ }), .Y(_06734_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27781_ ( .A({ _12926_, _11896_, _06612_, _12894_ }), .Y(_06735_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27782_ ( .A({ _06740_, _06739_, _06738_, _06737_ }), .Y(_06736_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27783_ ( .A({ _13342_, _05042_, _06604_, _13150_ }), .Y(_06737_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27784_ ( .A({ _13310_, _06581_, _13374_, _06603_ }), .Y(_06738_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27785_ ( .A({ _13182_, _06598_, _06622_, _13054_ }), .Y(_06739_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27786_ ( .A({ _13246_, _06592_, _06620_, _13086_ }), .Y(_06740_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27787_ ( .A({ _13118_, _06594_, _06596_, _12958_ }), .Y(_06741_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27788_ ( .A({ _12990_, _06588_, _13022_, _06616_ }), .Y(_06742_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27789_ ( .A({ _06753_, _06752_, _06747_, _06743_ }), .Y(_12832_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27790_ ( .A({ _06746_, _06745_, _06744_ }), .Y(_06743_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27791_ ( .A({ _13152_, _06598_, _13344_, _06603_ }), .Y(_06744_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27792_ ( .A({ 1'h0, _06611_, _12864_, _06612_ }), .Y(_06745_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27793_ ( .A({ _12896_, _11896_, _12800_, _05035_ }), .Y(_06746_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27794_ ( .A({ _06751_, _06750_, _06749_, _06748_ }), .Y(_06747_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27795_ ( .A({ _13280_, _06581_, _06592_, _13216_ }), .Y(_06748_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27796_ ( .A({ _13248_, _06578_, _13312_, _05042_ }), .Y(_06749_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27797_ ( .A({ _13184_, _06600_, _06620_, _13056_ }), .Y(_06750_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27798_ ( .A({ _13088_, _06594_, _06596_, _12928_ }), .Y(_06751_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27799_ ( .A({ _12992_, _06616_, _06622_, _13024_ }), .Y(_06752_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27800_ ( .A({ _12960_, _06588_, _13120_, _06604_ }), .Y(_06753_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27801_ ( .A({ _06764_, _06763_, _06758_, _06754_ }), .Y(_12834_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27802_ ( .A({ _06757_, _06756_, _06755_ }), .Y(_06754_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27803_ ( .A({ _13090_, _06594_, _13154_, _06598_ }), .Y(_06755_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27804_ ( .A({ _12898_, _11896_, _12802_, _05035_ }), .Y(_06756_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27805_ ( .A({ 1'h0, _06611_, _12866_, _06612_ }), .Y(_06757_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27806_ ( .A({ _06762_, _06761_, _06760_, _06759_ }), .Y(_06758_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27807_ ( .A({ _13250_, _06578_, _13282_, _06581_ }), .Y(_06759_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27808_ ( .A({ _12962_, _06588_, _06596_, _12930_ }), .Y(_06760_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27809_ ( .A({ _13346_, _06603_, _06620_, _13058_ }), .Y(_06761_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27810_ ( .A({ _13218_, _06592_, _06622_, _13026_ }), .Y(_06762_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27811_ ( .A({ _13122_, _06604_, _06616_, _12994_ }), .Y(_06763_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27812_ ( .A({ _13314_, _05042_, _06600_, _13186_ }), .Y(_06764_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27813_ ( .A({ _06775_, _06774_, _06769_, _06765_ }), .Y(_12835_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27814_ ( .A({ _06768_, _06767_, _06766_ }), .Y(_06765_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27815_ ( .A({ _12931_, _06596_, _13059_, _06620_ }), .Y(_06766_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27816_ ( .A({ _12899_, _11896_, _12803_, _05035_ }), .Y(_06767_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27817_ ( .A({ 1'h0, _06611_, _12867_, _06612_ }), .Y(_06768_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27818_ ( .A({ _06773_, _06772_, _06771_, _06770_ }), .Y(_06769_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27819_ ( .A({ _13315_, _05042_, _06592_, _13219_ }), .Y(_06770_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27820_ ( .A({ _13091_, _06594_, _13187_, _06600_ }), .Y(_06771_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27821_ ( .A({ _13283_, _06581_, _06622_, _13027_ }), .Y(_06772_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27822_ ( .A({ _13251_, _06578_, _06616_, _12995_ }), .Y(_06773_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27823_ ( .A({ _12963_, _06588_, _13123_, _06604_ }), .Y(_06774_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27824_ ( .A({ _13155_, _06598_, _13347_, _06603_ }), .Y(_06775_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27825_ ( .A({ _06786_, _06785_, _06780_, _06776_ }), .Y(_12839_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27826_ ( .A({ _06779_, _06778_, _06777_ }), .Y(_06776_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27827_ ( .A({ _13319_, _05042_, _06622_, _13031_ }), .Y(_06777_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27828_ ( .A({ 1'h0, _06611_, _12871_, _06612_ }), .Y(_06778_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27829_ ( .A({ _12903_, _11896_, _12807_, _05035_ }), .Y(_06779_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27830_ ( .A({ _06784_, _06783_, _06782_, _06781_ }), .Y(_06780_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27831_ ( .A({ _12935_, _06596_, _13351_, _06603_ }), .Y(_06781_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27832_ ( .A({ _13287_, _06581_, _06588_, _12967_ }), .Y(_06782_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27833_ ( .A({ _13255_, _06578_, _06600_, _13191_ }), .Y(_06783_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27834_ ( .A({ _13223_, _06592_, _06620_, _13063_ }), .Y(_06784_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27835_ ( .A({ _13095_, _06594_, _06604_, _13127_ }), .Y(_06785_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27836_ ( .A({ _13159_, _06598_, _06616_, _12999_ }), .Y(_06786_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27837_ ( .A({ _06797_, _06796_, _06791_, _06787_ }), .Y(_12844_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27838_ ( .A({ _06790_, _06789_, _06788_ }), .Y(_06787_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27839_ ( .A({ _13228_, _06592_, _06604_, _13132_ }), .Y(_06788_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27840_ ( .A({ _12908_, _11896_, _06611_, 1'h0 }), .Y(_06789_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27841_ ( .A({ _12876_, _06612_, _12812_, _05035_ }), .Y(_06790_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27842_ ( .A({ _06795_, _06794_, _06793_, _06792_ }), .Y(_06791_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27843_ ( .A({ _13292_, _06581_, _13324_, _05042_ }), .Y(_06792_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27844_ ( .A({ _13196_, _06600_, _06616_, _13004_ }), .Y(_06793_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27845_ ( .A({ _12972_, _06588_, _13356_, _06603_ }), .Y(_06794_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27846_ ( .A({ _13260_, _06578_, _06598_, _13164_ }), .Y(_06795_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27847_ ( .A({ _12940_, _06596_, _06622_, _13036_ }), .Y(_06796_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27848_ ( .A({ _13100_, _06594_, _06620_, _13068_ }), .Y(_06797_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27849_ ( .A({ _06808_, _06807_, _06802_, _06798_ }), .Y(_12836_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27850_ ( .A({ _06801_, _06800_, _06799_ }), .Y(_06798_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27851_ ( .A({ _13220_, _06592_, _06622_, _13028_ }), .Y(_06799_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27852_ ( .A({ 1'h0, _06611_, _12868_, _06612_ }), .Y(_06800_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27853_ ( .A({ _12900_, _11896_, _12804_, _05035_ }), .Y(_06801_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27854_ ( .A({ _06806_, _06805_, _06804_, _06803_ }), .Y(_06802_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27855_ ( .A({ _13316_, _05042_, _06596_, _12932_ }), .Y(_06803_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27856_ ( .A({ _13156_, _06598_, _06616_, _12996_ }), .Y(_06804_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27857_ ( .A({ _13252_, _06578_, _06594_, _13092_ }), .Y(_06805_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27858_ ( .A({ _12964_, _06588_, _13124_, _06604_ }), .Y(_06806_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27859_ ( .A({ _13348_, _06603_, _06600_, _13188_ }), .Y(_06807_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27860_ ( .A({ _13284_, _06581_, _06620_, _13060_ }), .Y(_06808_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27861_ ( .A({ _06819_, _06818_, _06813_, _06809_ }), .Y(_12837_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27862_ ( .A({ _06812_, _06811_, _06810_ }), .Y(_06809_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27863_ ( .A({ _13285_, _06581_, _06588_, _12965_ }), .Y(_06810_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27864_ ( .A({ _12901_, _11896_, _06611_, 1'h0 }), .Y(_06811_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27865_ ( .A({ _12869_, _06612_, _12805_, _05035_ }), .Y(_06812_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27866_ ( .A({ _06817_, _06816_, _06815_, _06814_ }), .Y(_06813_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27867_ ( .A({ _13221_, _06592_, _13349_, _06603_ }), .Y(_06814_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27868_ ( .A({ _13189_, _06600_, _06622_, _13029_ }), .Y(_06815_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27869_ ( .A({ _13253_, _06578_, _06604_, _13125_ }), .Y(_06816_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27870_ ( .A({ _13317_, _05042_, _06596_, _12933_ }), .Y(_06817_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27871_ ( .A({ _13093_, _06594_, _13157_, _06598_ }), .Y(_06818_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27872_ ( .A({ _12997_, _06616_, _13061_, _06620_ }), .Y(_06819_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27873_ ( .A({ _06830_, _06829_, _06824_, _06820_ }), .Y(_12838_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27874_ ( .A({ _06823_, _06822_, _06821_ }), .Y(_06820_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27875_ ( .A({ _13094_, _06594_, _06596_, _12934_ }), .Y(_06821_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27876_ ( .A({ _12902_, _11896_, _06611_, 1'h0 }), .Y(_06822_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27877_ ( .A({ _12870_, _06612_, _12806_, _05035_ }), .Y(_06823_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27878_ ( .A({ _06828_, _06827_, _06826_, _06825_ }), .Y(_06824_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27879_ ( .A({ _13318_, _05042_, _06600_, _13190_ }), .Y(_06825_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27880_ ( .A({ _12966_, _06588_, _13062_, _06620_ }), .Y(_06826_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27881_ ( .A({ _13222_, _06592_, _06616_, _12998_ }), .Y(_06827_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27882_ ( .A({ _13126_, _06604_, _06622_, _13030_ }), .Y(_06828_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27883_ ( .A({ _13254_, _06578_, _13350_, _06603_ }), .Y(_06829_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27884_ ( .A({ _13286_, _06581_, _06598_, _13158_ }), .Y(_06830_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27885_ ( .A({ _06841_, _06840_, _06835_, _06831_ }), .Y(_12840_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27886_ ( .A({ _06834_, _06833_, _06832_ }), .Y(_06831_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27887_ ( .A({ _13128_, _06604_, _06616_, _13000_ }), .Y(_06832_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27888_ ( .A({ 1'h0, _06611_, _12872_, _06612_ }), .Y(_06833_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27889_ ( .A({ _12904_, _11896_, _12808_, _05035_ }), .Y(_06834_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27890_ ( .A({ _06839_, _06838_, _06837_, _06836_ }), .Y(_06835_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27891_ ( .A({ _13352_, _06603_, _06620_, _13064_ }), .Y(_06836_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27892_ ( .A({ _13288_, _06581_, _13320_, _05042_ }), .Y(_06837_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27893_ ( .A({ _13192_, _06600_, _06622_, _13032_ }), .Y(_06838_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27894_ ( .A({ _13224_, _06592_, _06598_, _13160_ }), .Y(_06839_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27895_ ( .A({ _13256_, _06578_, _06588_, _12968_ }), .Y(_06840_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27896_ ( .A({ _13096_, _06594_, _06596_, _12936_ }), .Y(_06841_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27897_ ( .A({ _06852_, _06851_, _06846_, _06842_ }), .Y(_12841_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27898_ ( .A({ _06845_, _06844_, _06843_ }), .Y(_06842_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27899_ ( .A({ _13289_, _06581_, _06600_, _13193_ }), .Y(_06843_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27900_ ( .A({ 1'h0, _06611_, _12809_, _05035_ }), .Y(_06844_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27901_ ( .A({ _12905_, _11896_, _06612_, _12873_ }), .Y(_06845_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27902_ ( .A({ _06850_, _06849_, _06848_, _06847_ }), .Y(_06846_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27903_ ( .A({ _13257_, _06578_, _06588_, _12969_ }), .Y(_06847_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27904_ ( .A({ _13321_, _05042_, _06604_, _13129_ }), .Y(_06848_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27905_ ( .A({ _13097_, _06594_, _06622_, _13033_ }), .Y(_06849_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27906_ ( .A({ _12937_, _06596_, _13065_, _06620_ }), .Y(_06850_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27907_ ( .A({ _13353_, _06603_, _06616_, _13001_ }), .Y(_06851_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27908_ ( .A({ _13225_, _06592_, _06598_, _13161_ }), .Y(_06852_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27909_ ( .A({ _06863_, _06862_, _06857_, _06853_ }), .Y(_12843_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27910_ ( .A({ _06856_, _06855_, _06854_ }), .Y(_06853_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27911_ ( .A({ _13259_, _06578_, _06620_, _13067_ }), .Y(_06854_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27912_ ( .A({ 1'h0, _06611_, _12875_, _06612_ }), .Y(_06855_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27913_ ( .A({ _12907_, _11896_, _12811_, _05035_ }), .Y(_06856_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27914_ ( .A({ _06861_, _06860_, _06859_, _06858_ }), .Y(_06857_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27915_ ( .A({ _13323_, _05042_, _13355_, _06603_ }), .Y(_06858_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27916_ ( .A({ _12939_, _06596_, _13195_, _06600_ }), .Y(_06859_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27917_ ( .A({ _12971_, _06588_, _13099_, _06594_ }), .Y(_06860_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27918_ ( .A({ _13163_, _06598_, _06622_, _13035_ }), .Y(_06861_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27919_ ( .A({ _13291_, _06581_, _06592_, _13227_ }), .Y(_06862_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27920_ ( .A({ _13131_, _06604_, _06616_, _13003_ }), .Y(_06863_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27921_ ( .A({ _06874_, _06873_, _06868_, _06864_ }), .Y(_12849_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27922_ ( .A({ _06867_, _06866_, _06865_ }), .Y(_06864_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27923_ ( .A({ _13297_, _06581_, _06600_, _13201_ }), .Y(_06865_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27924_ ( .A({ 1'h0, _06611_, _12881_, _06612_ }), .Y(_06866_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27925_ ( .A({ _12913_, _11896_, _12817_, _05035_ }), .Y(_06867_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27926_ ( .A({ _06872_, _06871_, _06870_, _06869_ }), .Y(_06868_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27927_ ( .A({ _13233_, _06592_, _06604_, _13137_ }), .Y(_06869_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27928_ ( .A({ _13265_, _06578_, _13361_, _06603_ }), .Y(_06870_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27929_ ( .A({ _12945_, _06596_, _13169_, _06598_ }), .Y(_06871_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27930_ ( .A({ _13329_, _05042_, _06588_, _12977_ }), .Y(_06872_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27931_ ( .A({ _13009_, _06616_, _06622_, _13041_ }), .Y(_06873_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27932_ ( .A({ _13105_, _06594_, _06620_, _13073_ }), .Y(_06874_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27933_ ( .A({ _06885_, _06884_, _06879_, _06875_ }), .Y(_12845_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27934_ ( .A({ _06878_, _06877_, _06876_ }), .Y(_06875_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27935_ ( .A({ _12973_, _06588_, _13101_, _06594_ }), .Y(_06876_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27936_ ( .A({ 1'h0, _06611_, _12877_, _06612_ }), .Y(_06877_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27937_ ( .A({ _12909_, _11896_, _12813_, _05035_ }), .Y(_06878_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27938_ ( .A({ _06883_, _06882_, _06881_, _06880_ }), .Y(_06879_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27939_ ( .A({ _13229_, _06592_, _06598_, _13165_ }), .Y(_06880_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27940_ ( .A({ _13325_, _05042_, _06604_, _13133_ }), .Y(_06881_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27941_ ( .A({ _13261_, _06578_, _06620_, _13069_ }), .Y(_06882_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27942_ ( .A({ _13005_, _06616_, _06622_, _13037_ }), .Y(_06883_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27943_ ( .A({ _13293_, _06581_, _06596_, _12941_ }), .Y(_06884_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27944_ ( .A({ _13357_, _06603_, _06600_, _13197_ }), .Y(_06885_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27945_ ( .A({ _06896_, _06895_, _06890_, _06886_ }), .Y(_12854_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27946_ ( .A({ _06889_, _06888_, _06887_ }), .Y(_06886_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27947_ ( .A({ _13174_, _06598_, _06604_, _13142_ }), .Y(_06887_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27948_ ( .A({ _12918_, _11896_, _06612_, _12886_ }), .Y(_06888_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27949_ ( .A({ 1'h0, _06611_, _12822_, _05035_ }), .Y(_06889_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27950_ ( .A({ _06894_, _06893_, _06892_, _06891_ }), .Y(_06890_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27951_ ( .A({ _13366_, _06603_, _06600_, _13206_ }), .Y(_06891_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27952_ ( .A({ _13078_, _06620_, _06622_, _13046_ }), .Y(_06892_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27953_ ( .A({ _13334_, _05042_, _06592_, _13238_ }), .Y(_06893_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27954_ ( .A({ _13270_, _06578_, _06616_, _13014_ }), .Y(_06894_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27955_ ( .A({ _12982_, _06588_, _13110_, _06594_ }), .Y(_06895_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27956_ ( .A({ _13302_, _06581_, _06596_, _12950_ }), .Y(_06896_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27957_ ( .A({ _06907_, _06906_, _06901_, _06897_ }), .Y(_12846_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27958_ ( .A({ _06900_, _06899_, _06898_ }), .Y(_06897_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27959_ ( .A({ _13006_, _06616_, _06622_, _13038_ }), .Y(_06898_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27960_ ( .A({ 1'h0, _06611_, _12814_, _05035_ }), .Y(_06899_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27961_ ( .A({ _12910_, _11896_, _06612_, _12878_ }), .Y(_06900_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27962_ ( .A({ _06905_, _06904_, _06903_, _06902_ }), .Y(_06901_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27963_ ( .A({ _13262_, _06578_, _06600_, _13198_ }), .Y(_06902_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27964_ ( .A({ _13326_, _05042_, _06596_, _12942_ }), .Y(_06903_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27965_ ( .A({ _12974_, _06588_, _13134_, _06604_ }), .Y(_06904_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27966_ ( .A({ _13166_, _06598_, _06620_, _13070_ }), .Y(_06905_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27967_ ( .A({ _13230_, _06592_, _06594_, _13102_ }), .Y(_06906_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27968_ ( .A({ _13294_, _06581_, _13358_, _06603_ }), .Y(_06907_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27969_ ( .A({ _06918_, _06917_, _06912_, _06908_ }), .Y(_12847_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27970_ ( .A({ _06911_, _06910_, _06909_ }), .Y(_06908_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27971_ ( .A({ _13167_, _06598_, _06604_, _13135_ }), .Y(_06909_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27972_ ( .A({ _12911_, _11896_, _06612_, _12879_ }), .Y(_06910_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27973_ ( .A({ 1'h0, _06611_, _12815_, _05035_ }), .Y(_06911_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27974_ ( .A({ _06916_, _06915_, _06914_, _06913_ }), .Y(_06912_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27975_ ( .A({ _13359_, _06603_, _06600_, _13199_ }), .Y(_06913_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27976_ ( .A({ _13071_, _06620_, _06622_, _13039_ }), .Y(_06914_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27977_ ( .A({ _13327_, _05042_, _06592_, _13231_ }), .Y(_06915_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27978_ ( .A({ _13263_, _06578_, _06616_, _13007_ }), .Y(_06916_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27979_ ( .A({ _12975_, _06588_, _13103_, _06594_ }), .Y(_06917_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27980_ ( .A({ _13295_, _06581_, _06596_, _12943_ }), .Y(_06918_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27981_ ( .A({ _06929_, _06928_, _06923_, _06919_ }), .Y(_12848_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27982_ ( .A({ _06922_, _06921_, _06920_ }), .Y(_06919_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27983_ ( .A({ _13328_, _05042_, _06622_, _13040_ }), .Y(_06920_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27984_ ( .A({ 1'h0, _06611_, _12880_, _06612_ }), .Y(_06921_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27985_ ( .A({ _12912_, _11896_, _12816_, _05035_ }), .Y(_06922_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27986_ ( .A({ _06927_, _06926_, _06925_, _06924_ }), .Y(_06923_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27987_ ( .A({ _12944_, _06596_, _13360_, _06603_ }), .Y(_06924_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27988_ ( .A({ _13296_, _06581_, _06588_, _12976_ }), .Y(_06925_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27989_ ( .A({ _13264_, _06578_, _06600_, _13200_ }), .Y(_06926_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27990_ ( .A({ _13232_, _06592_, _06620_, _13072_ }), .Y(_06927_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27991_ ( .A({ _13104_, _06594_, _06604_, _13136_ }), .Y(_06928_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27992_ ( .A({ _13168_, _06598_, _06616_, _13008_ }), .Y(_06929_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _27993_ ( .A({ _06940_, _06939_, _06934_, _06930_ }), .Y(_12850_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _27994_ ( .A({ _06933_, _06932_, _06931_ }), .Y(_06930_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _27995_ ( .A({ _13330_, _05042_, _06622_, _13042_ }), .Y(_06931_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27996_ ( .A({ _12914_, _11896_, _06611_, 1'h0 }), .Y(_06932_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _27997_ ( .A({ _12882_, _06612_, _12818_, _05035_ }), .Y(_06933_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _27998_ ( .A({ _06938_, _06937_, _06936_, _06935_ }), .Y(_06934_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _27999_ ( .A({ _13362_, _06603_, _06604_, _13138_ }), .Y(_06935_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28000_ ( .A({ _13234_, _06592_, _06620_, _13074_ }), .Y(_06936_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28001_ ( .A({ _13298_, _06581_, _06588_, _12978_ }), .Y(_06937_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28002_ ( .A({ _13266_, _06578_, _06616_, _13010_ }), .Y(_06938_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28003_ ( .A({ _13170_, _06598_, _13202_, _06600_ }), .Y(_06939_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28004_ ( .A({ _13106_, _06594_, _06596_, _12946_ }), .Y(_06940_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _28005_ ( .A({ _06951_, _06950_, _06945_, _06941_ }), .Y(_12851_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28006_ ( .A({ _06944_, _06943_, _06942_ }), .Y(_06941_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28007_ ( .A({ _13171_, _06598_, _13363_, _06603_ }), .Y(_06942_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28008_ ( .A({ _12915_, _11896_, _06611_, 1'h0 }), .Y(_06943_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _28009_ ( .A({ _12883_, _06612_, _12819_, _05035_ }), .Y(_06944_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28010_ ( .A({ _06949_, _06948_, _06947_, _06946_ }), .Y(_06945_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28011_ ( .A({ _13299_, _06581_, _06600_, _13203_ }), .Y(_06946_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28012_ ( .A({ _13267_, _06578_, _06616_, _13011_ }), .Y(_06947_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _28013_ ( .A({ _13331_, _05042_, _06620_, _13075_ }), .Y(_06948_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28014_ ( .A({ _13235_, _06592_, _06596_, _12947_ }), .Y(_06949_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28015_ ( .A({ _13107_, _06594_, _06622_, _13043_ }), .Y(_06950_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28016_ ( .A({ _12979_, _06588_, _13139_, _06604_ }), .Y(_06951_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _28017_ ( .A({ _06962_, _06961_, _06956_, _06952_ }), .Y(_12852_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28018_ ( .A({ _06955_, _06954_, _06953_ }), .Y(_06952_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28019_ ( .A({ _12980_, _06588_, _13012_, _06616_ }), .Y(_06953_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28020_ ( .A({ 1'h0, _06611_, _12884_, _06612_ }), .Y(_06954_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _28021_ ( .A({ _12916_, _11896_, _12820_, _05035_ }), .Y(_06955_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28022_ ( .A({ _06960_, _06959_, _06958_, _06957_ }), .Y(_06956_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28023_ ( .A({ _13364_, _06603_, _06604_, _13140_ }), .Y(_06957_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28024_ ( .A({ _13172_, _06598_, _06620_, _13076_ }), .Y(_06958_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _28025_ ( .A({ _13300_, _06581_, _13332_, _05042_ }), .Y(_06959_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28026_ ( .A({ _13268_, _06578_, _06594_, _13108_ }), .Y(_06960_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28027_ ( .A({ _13204_, _06600_, _06622_, _13044_ }), .Y(_06961_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28028_ ( .A({ _13236_, _06592_, _06596_, _12948_ }), .Y(_06962_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _28029_ ( .A({ _06973_, _06972_, _06967_, _06963_ }), .Y(_12855_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28030_ ( .A({ _06966_, _06965_, _06964_ }), .Y(_06963_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28031_ ( .A({ _13239_, _06592_, _06604_, _13143_ }), .Y(_06964_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28032_ ( .A({ _12919_, _11896_, _06611_, 1'h0 }), .Y(_06965_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _28033_ ( .A({ _12887_, _06612_, _12823_, _05035_ }), .Y(_06966_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28034_ ( .A({ _06971_, _06970_, _06969_, _06968_ }), .Y(_06967_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _28035_ ( .A({ _13303_, _06581_, _13335_, _05042_ }), .Y(_06968_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28036_ ( .A({ _13207_, _06600_, _06616_, _13015_ }), .Y(_06969_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28037_ ( .A({ _12983_, _06588_, _13367_, _06603_ }), .Y(_06970_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28038_ ( .A({ _13271_, _06578_, _06598_, _13175_ }), .Y(_06971_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28039_ ( .A({ _12951_, _06596_, _06622_, _13047_ }), .Y(_06972_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _28040_ ( .A({ _13111_, _06594_, _06620_, _13079_ }), .Y(_06973_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28041_ ( .A({ _12760_, _11896_, _06611_, _04373_ }), .Y(_04702_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28042_ ( .A({ _12735_, _11896_, _06611_, _04348_ }), .Y(_04703_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28043_ ( .A({ _12746_, _11896_, _06611_, _04359_ }), .Y(_04704_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28044_ ( .A({ _12757_, _11896_, _06611_, _04370_ }), .Y(_04705_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28045_ ( .A({ _12761_, _11896_, _06611_, _04374_ }), .Y(_04706_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28046_ ( .A({ _12762_, _11896_, _06611_, _04375_ }), .Y(_04707_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28047_ ( .A({ _12763_, _11896_, _06611_, _04376_ }), .Y(_04708_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28048_ ( .A({ _12764_, _11896_, _06611_, _04377_ }), .Y(_04709_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28049_ ( .A({ _12738_, _11896_, _06611_, _04351_ }), .Y(_04710_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28050_ ( .A({ _12765_, _11896_, _06611_, _04378_ }), .Y(_04711_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28051_ ( .A({ _12742_, _11896_, _06611_, _04355_ }), .Y(_04712_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28052_ ( .A({ _12766_, _11896_, _06611_, _04379_ }), .Y(_04713_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28053_ ( .A({ _12736_, _11896_, _06611_, _04349_ }), .Y(_04714_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28054_ ( .A({ _12737_, _11896_, _06611_, _04350_ }), .Y(_04715_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28055_ ( .A({ _12745_, _11896_, _06611_, _04358_ }), .Y(_04716_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28056_ ( .A({ _12739_, _11896_, _06611_, _04352_ }), .Y(_04717_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28057_ ( .A({ _12740_, _11896_, _06611_, _04353_ }), .Y(_04718_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28058_ ( .A({ _12741_, _11896_, _06611_, _04354_ }), .Y(_04719_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28059_ ( .A({ _12743_, _11896_, _06611_, _04356_ }), .Y(_04720_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28060_ ( .A({ _12744_, _11896_, _06611_, _04357_ }), .Y(_04721_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28061_ ( .A({ _12747_, _11896_, _06611_, _04360_ }), .Y(_04722_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28062_ ( .A({ _12750_, _11896_, _06611_, _04363_ }), .Y(_04723_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28063_ ( .A({ _12748_, _11896_, _06611_, _04361_ }), .Y(_04724_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28064_ ( .A({ _12749_, _11896_, _06611_, _04362_ }), .Y(_04725_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28065_ ( .A({ _12752_, _11896_, _06611_, _04365_ }), .Y(_04726_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28066_ ( .A({ _12751_, _11896_, _06611_, _04364_ }), .Y(_04727_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28067_ ( .A({ _12755_, _11896_, _06611_, _04368_ }), .Y(_04728_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28068_ ( .A({ _12753_, _11896_, _06611_, _04366_ }), .Y(_04729_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28069_ ( .A({ _12758_, _11896_, _06611_, _04371_ }), .Y(_04730_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28070_ ( .A({ _12754_, _11896_, _06611_, _04367_ }), .Y(_04731_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28071_ ( .A({ _12756_, _11896_, _06611_, _04369_ }), .Y(_04732_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28072_ ( .A({ _12759_, _11896_, _06611_, _04372_ }), .Y(_04733_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28073_ ( .A({ _05132_, _18550_, _05909_ }), .Y(_18551_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28074_ ( .A({ _05042_, _06611_ }), .Y(_21889_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28075_ ( .A({ _12319_, _11896_, _12351_, _06611_ }), .Y(_04734_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28076_ ( .A({ _12330_, _11896_, _12362_, _06611_ }), .Y(_04735_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28077_ ( .A({ _12341_, _11896_, _12373_, _06611_ }), .Y(_04736_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28078_ ( .A({ _12344_, _11896_, _12376_, _06611_ }), .Y(_04737_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28079_ ( .A({ _12345_, _11896_, _12377_, _06611_ }), .Y(_04738_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28080_ ( .A({ _12346_, _11896_, _12378_, _06611_ }), .Y(_04739_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28081_ ( .A({ _12347_, _11896_, _12379_, _06611_ }), .Y(_04740_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28082_ ( .A({ _12348_, _11896_, _12380_, _06611_ }), .Y(_04741_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28083_ ( .A({ _12349_, _11896_, _12381_, _06611_ }), .Y(_04742_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28084_ ( .A({ _12350_, _11896_, _12382_, _06611_ }), .Y(_04743_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28085_ ( .A({ _12320_, _11896_, _12352_, _06611_ }), .Y(_04744_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28086_ ( .A({ _12321_, _11896_, _12353_, _06611_ }), .Y(_04745_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28087_ ( .A({ _12322_, _11896_, _12354_, _06611_ }), .Y(_04746_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28088_ ( .A({ _12323_, _11896_, _12355_, _06611_ }), .Y(_04747_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28089_ ( .A({ _12324_, _11896_, _12356_, _06611_ }), .Y(_04748_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28090_ ( .A({ _12325_, _11896_, _12357_, _06611_ }), .Y(_04749_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28091_ ( .A({ _12326_, _11896_, _12358_, _06611_ }), .Y(_04750_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28092_ ( .A({ _12327_, _11896_, _12359_, _06611_ }), .Y(_04751_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28093_ ( .A({ _12328_, _11896_, _12360_, _06611_ }), .Y(_04752_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28094_ ( .A({ _12329_, _11896_, _12361_, _06611_ }), .Y(_04753_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28095_ ( .A({ _12331_, _11896_, _12363_, _06611_ }), .Y(_04754_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28096_ ( .A({ _12332_, _11896_, _12364_, _06611_ }), .Y(_04755_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28097_ ( .A({ _12333_, _11896_, _12365_, _06611_ }), .Y(_04756_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28098_ ( .A({ _12334_, _11896_, _12366_, _06611_ }), .Y(_04757_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28099_ ( .A({ _12335_, _11896_, _12367_, _06611_ }), .Y(_04758_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28100_ ( .A({ _12336_, _11896_, _12368_, _06611_ }), .Y(_04759_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28101_ ( .A({ _12337_, _11896_, _12369_, _06611_ }), .Y(_04760_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28102_ ( .A({ _12338_, _11896_, _12370_, _06611_ }), .Y(_04761_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28103_ ( .A({ _12339_, _11896_, _12371_, _06611_ }), .Y(_04762_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28104_ ( .A({ _12340_, _11896_, _12372_, _06611_ }), .Y(_04763_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28105_ ( .A({ _12342_, _11896_, _12374_, _06611_ }), .Y(_04764_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28106_ ( .A({ _12343_, _11896_, _12375_, _06611_ }), .Y(_04765_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28107_ ( .A({ _19388_, _05909_, _06338_, _19420_ }), .Y(_04766_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28108_ ( .A({ _19387_, _05909_, _06338_, _19419_ }), .Y(_04767_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28109_ ( .A({ _19385_, _05909_, _06338_, _19417_ }), .Y(_04768_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28110_ ( .A({ _19384_, _05909_, _06338_, _19416_ }), .Y(_04769_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28111_ ( .A({ _19383_, _05909_, _06338_, _19415_ }), .Y(_04770_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28112_ ( .A({ _19382_, _05909_, _06338_, _19414_ }), .Y(_04771_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28113_ ( .A({ _19381_, _05909_, _06338_, _19413_ }), .Y(_04772_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28114_ ( .A({ _19380_, _05909_, _06338_, _19412_ }), .Y(_04773_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28115_ ( .A({ _19379_, _05909_, _06338_, _19411_ }), .Y(_04774_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28116_ ( .A({ _19378_, _05909_, _06338_, _19410_ }), .Y(_04775_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28117_ ( .A({ _19377_, _05909_, _06338_, _19409_ }), .Y(_04776_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28118_ ( .A({ _19376_, _05909_, _06338_, _19408_ }), .Y(_04777_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28119_ ( .A({ _19374_, _05909_, _06338_, _19406_ }), .Y(_04778_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28120_ ( .A({ _19373_, _05909_, _06338_, _19405_ }), .Y(_04779_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28121_ ( .A({ _19372_, _05909_, _06338_, _19404_ }), .Y(_04780_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28122_ ( .A({ _19371_, _05909_, _06338_, _19403_ }), .Y(_04781_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28123_ ( .A({ _19370_, _05909_, _06338_, _19402_ }), .Y(_04782_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28124_ ( .A({ _19369_, _05909_, _06338_, _19401_ }), .Y(_04783_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28125_ ( .A({ _19368_, _05909_, _06338_, _19400_ }), .Y(_04784_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28126_ ( .A({ _19367_, _05909_, _06338_, _19399_ }), .Y(_04785_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28127_ ( .A({ _19366_, _05909_, _06338_, _19398_ }), .Y(_04786_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28128_ ( .A({ _19365_, _05909_, _06338_, _19397_ }), .Y(_04787_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28129_ ( .A({ _19395_, _05909_, _06338_, _19427_ }), .Y(_04788_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28130_ ( .A({ _19394_, _05909_, _06338_, _19426_ }), .Y(_04789_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28131_ ( .A({ _19393_, _05909_, _06338_, _19425_ }), .Y(_04790_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28132_ ( .A({ _19391_, _05909_, _06338_, _19423_ }), .Y(_04791_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28133_ ( .A({ _19392_, _05909_, _06338_, _19424_ }), .Y(_04792_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28134_ ( .A({ _19390_, _05909_, _06338_, _19422_ }), .Y(_04793_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28135_ ( .A({ _19389_, _05909_, _06338_, _19421_ }), .Y(_04794_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28136_ ( .A({ _19386_, _05909_, _06338_, _19418_ }), .Y(_04795_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28137_ ( .A({ _19375_, _05909_, _06338_, _19407_ }), .Y(_04796_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28138_ ( .A({ _19364_, _05909_, _06338_, _19396_ }), .Y(_04797_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _28139_ ( .A({ _06611_, _04701_ }), .Y(_21888_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28140_ ( .A({ _05042_, _11896_ }), .Y(_04701_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28141_ ( .A({ _11912_, _11896_, _11944_, _06611_ }), .Y(_04798_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28142_ ( .A({ _11901_, _11896_, _11933_, _06611_ }), .Y(_04799_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28143_ ( .A({ _11923_, _11896_, _11955_, _06611_ }), .Y(_04800_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28144_ ( .A({ _11928_, _11896_, _11960_, _06611_ }), .Y(_04801_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28145_ ( .A({ _11926_, _11896_, _11958_, _06611_ }), .Y(_04802_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28146_ ( .A({ _11932_, _11896_, _11964_, _06611_ }), .Y(_04803_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28147_ ( .A({ _11927_, _11896_, _11959_, _06611_ }), .Y(_04804_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28148_ ( .A({ _11929_, _11896_, _11961_, _06611_ }), .Y(_04805_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28149_ ( .A({ _11930_, _11896_, _11962_, _06611_ }), .Y(_04806_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28150_ ( .A({ _11931_, _11896_, _11963_, _06611_ }), .Y(_04807_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28151_ ( .A({ _11902_, _11896_, _11934_, _06611_ }), .Y(_04808_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28152_ ( .A({ _11905_, _11896_, _11937_, _06611_ }), .Y(_04809_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28153_ ( .A({ _11903_, _11896_, _11935_, _06611_ }), .Y(_04810_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28154_ ( .A({ _11909_, _11896_, _11941_, _06611_ }), .Y(_04811_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28155_ ( .A({ _11904_, _11896_, _11936_, _06611_ }), .Y(_04812_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28156_ ( .A({ _11906_, _11896_, _11938_, _06611_ }), .Y(_04813_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28157_ ( .A({ _11907_, _11896_, _11939_, _06611_ }), .Y(_04814_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28158_ ( .A({ _11908_, _11896_, _11940_, _06611_ }), .Y(_04815_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28159_ ( .A({ _11910_, _11896_, _11942_, _06611_ }), .Y(_04816_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28160_ ( .A({ _11914_, _11896_, _11946_, _06611_ }), .Y(_04817_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28161_ ( .A({ _11911_, _11896_, _11943_, _06611_ }), .Y(_04818_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28162_ ( .A({ _11918_, _11896_, _11950_, _06611_ }), .Y(_04819_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28163_ ( .A({ _11913_, _11896_, _11945_, _06611_ }), .Y(_04820_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28164_ ( .A({ _11915_, _11896_, _11947_, _06611_ }), .Y(_04821_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28165_ ( .A({ _11916_, _11896_, _11948_, _06611_ }), .Y(_04822_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28166_ ( .A({ _11917_, _11896_, _11949_, _06611_ }), .Y(_04823_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28167_ ( .A({ _11919_, _11896_, _11951_, _06611_ }), .Y(_04824_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28168_ ( .A({ _11922_, _11896_, _11954_, _06611_ }), .Y(_04825_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28169_ ( .A({ _11920_, _11896_, _11952_, _06611_ }), .Y(_04826_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28170_ ( .A({ _11921_, _11896_, _11953_, _06611_ }), .Y(_04827_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28171_ ( .A({ _11924_, _11896_, _11956_, _06611_ }), .Y(_04828_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28172_ ( .A({ _11925_, _11896_, _11957_, _06611_ }), .Y(_04829_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28173_ ( .A({ _05042_, _11894_, _11896_ }), .Y(_11895_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _28174_ ( .A({ _06988_, _06974_ }), .Y(_21886_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28175_ ( .A({ _05030_, _05028_, _06986_ }), .Y(_06974_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _28176_ ( .A({ _06975_, _06980_, matmul_15_comp_fsm[1] }), .Y(_05030_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _28177_ ( .A({ _06979_, _06976_, matmul_15_comp_fsm[2], matmul_15_comp_fsm[3] }), .Y(_06975_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28178_ ( .A({ _06978_, _06977_ }), .Y(_06976_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28179_ ( .A(matmul_15_comp_fsm[15:12]), .Y(_06977_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28180_ ( .A(matmul_15_comp_fsm[11:8]), .Y(_06978_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28181_ ( .A(matmul_15_comp_fsm[7:4]), .Y(_06979_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28182_ ( .A({ matmul_15_comp_fsm[0], _06981_ }), .Y(_06980_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28183_ ( .A({ _06985_, _06984_, _06983_, _06982_ }), .Y(_06981_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28184_ ( .A(matmul_15_comp_fsm[23:20]), .Y(_06982_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28185_ ( .A(matmul_15_comp_fsm[19:16]), .Y(_06983_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28186_ ( .A(matmul_15_comp_fsm[31:28]), .Y(_06984_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28187_ ( .A(matmul_15_comp_fsm[27:24]), .Y(_06985_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _28188_ ( .A({ matmul_15_comp_fsm[1], _06975_, _06981_, matmul_15_comp_fsm[0] }), .Y(_05028_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28189_ ( .A({ _06980_, _06987_, matmul_15_comp_fsm[1] }), .Y(_06986_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _28190_ ( .A({ matmul_15_comp_fsm[2], _06976_, _06979_, matmul_15_comp_fsm[3] }), .Y(_06987_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _28191_ ( .A({ _04897_, _05027_, _06991_, _06990_ }), .Y(_06988_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _28192_ ( .A({ matmul_15_comp_fsm[1], _06980_, _06975_ }), .Y(_05027_) );
  \$lut  #( .LUT(16'hefff), .WIDTH(4) ) _28193_ ( .A({ _06979_, _06989_, matmul_15_comp_fsm[2], matmul_15_comp_fsm[3] }), .Y(_04897_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _28194_ ( .A({ _06981_, _06976_, matmul_15_comp_fsm[1:0] }), .Y(_06989_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _28195_ ( .A({ matmul_15_comp_fsm[2], _06989_, _06979_, matmul_15_comp_fsm[3] }), .Y(_06990_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _28196_ ( .A({ matmul_15_comp_fsm[1], _06987_, _06981_, matmul_15_comp_fsm[0] }), .Y(_06991_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _28197_ ( .A({ _05027_, _06992_, _06986_ }), .Y(_11820_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _28198_ ( .A({ _11884_, _04897_, _11852_, _06990_ }), .Y(_06992_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28199_ ( .A({ _11892_, _04897_, _11860_, _06990_ }), .Y(_11828_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _28200_ ( .A({ _06993_, _06974_ }), .Y(_11809_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _28201_ ( .A({ _11873_, _04897_, _11841_, _06990_ }), .Y(_06993_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28202_ ( .A({ _06994_, _11830_, _06990_ }), .Y(_11798_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _28203_ ( .A({ _05028_, _04897_, _11862_ }), .Y(_06994_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28204_ ( .A({ _11865_, _04897_, _11833_, _06990_ }), .Y(_11801_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28205_ ( .A({ _11893_, _04897_, _11861_, _06990_ }), .Y(_11829_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28206_ ( .A({ _11891_, _04897_, _11859_, _06990_ }), .Y(_11827_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28207_ ( .A({ _11890_, _04897_, _11858_, _06990_ }), .Y(_11826_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28208_ ( .A({ _11889_, _04897_, _11857_, _06990_ }), .Y(_11825_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28209_ ( .A({ _11888_, _04897_, _11856_, _06990_ }), .Y(_11824_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28210_ ( .A({ _11871_, _04897_, _11839_, _06990_ }), .Y(_11807_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28211_ ( .A({ _11864_, _04897_, _11832_, _06990_ }), .Y(_11800_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28212_ ( .A({ _11870_, _04897_, _11838_, _06990_ }), .Y(_11806_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28213_ ( .A({ _11887_, _04897_, _11855_, _06990_ }), .Y(_11823_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28214_ ( .A({ _11863_, _04897_, _11831_, _06990_ }), .Y(_11799_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28215_ ( .A({ _11872_, _04897_, _11840_, _06990_ }), .Y(_11808_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28216_ ( .A({ _11869_, _04897_, _11837_, _06990_ }), .Y(_11805_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28217_ ( .A({ _11868_, _04897_, _11836_, _06990_ }), .Y(_11804_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28218_ ( .A({ _11867_, _04897_, _11835_, _06990_ }), .Y(_11803_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28219_ ( .A({ _11875_, _04897_, _11843_, _06990_ }), .Y(_11811_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28220_ ( .A({ _11881_, _04897_, _11849_, _06990_ }), .Y(_11817_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28221_ ( .A({ _11866_, _04897_, _11834_, _06990_ }), .Y(_11802_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28222_ ( .A({ _11874_, _04897_, _11842_, _06990_ }), .Y(_11810_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28223_ ( .A({ _11883_, _04897_, _11851_, _06990_ }), .Y(_11819_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28224_ ( .A({ _11882_, _04897_, _11850_, _06990_ }), .Y(_11818_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28225_ ( .A({ _11880_, _04897_, _11848_, _06990_ }), .Y(_11816_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28226_ ( .A({ _11879_, _04897_, _11847_, _06990_ }), .Y(_11815_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28227_ ( .A({ _11877_, _04897_, _11845_, _06990_ }), .Y(_11813_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28228_ ( .A({ _11886_, _04897_, _11854_, _06990_ }), .Y(_11822_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28229_ ( .A({ _11878_, _04897_, _11846_, _06990_ }), .Y(_11814_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28230_ ( .A({ _11876_, _04897_, _11844_, _06990_ }), .Y(_11812_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28231_ ( .A({ _11885_, _04897_, _11853_, _06990_ }), .Y(_11821_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28232_ ( .A({ _05030_, _06991_ }), .Y(_21887_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28233_ ( .A({ _05023_, _06995_ }), .Y(_21885_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28234_ ( .A({ _07004_, _07001_, _06996_ }), .Y(_06995_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28235_ ( .A({ _07000_, _06999_, _06998_, _06997_ }), .Y(_06996_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28236_ ( .A(_stream_matmul_15_source_6_source_pat_fsm_0[23:20]), .Y(_06997_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28237_ ( .A(_stream_matmul_15_source_6_source_pat_fsm_0[19:16]), .Y(_06998_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28238_ ( .A(_stream_matmul_15_source_6_source_pat_fsm_0[31:28]), .Y(_06999_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28239_ ( .A(_stream_matmul_15_source_6_source_pat_fsm_0[27:24]), .Y(_07000_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28240_ ( .A({ _07003_, _07002_ }), .Y(_07001_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28241_ ( .A(_stream_matmul_15_source_6_source_pat_fsm_0[15:12]), .Y(_07002_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28242_ ( .A(_stream_matmul_15_source_6_source_pat_fsm_0[11:8]), .Y(_07003_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _28243_ ( .A({ _07005_, _stream_matmul_15_source_6_source_pat_fsm_0[3:2], _stream_matmul_15_source_6_source_pat_fsm_0[0] }), .Y(_07004_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28244_ ( .A(_stream_matmul_15_source_6_source_pat_fsm_0[7:4]), .Y(_07005_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _28245_ ( .A({ _07006_, _07005_, _07001_, _06996_ }), .Y(_05023_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _28246_ ( .A({ _stream_matmul_15_source_6_source_pat_fsm_0[0], _stream_matmul_15_source_6_source_pat_fsm_0[3:1] }), .Y(_07006_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28247_ ( .A({ _11766_, _07007_, _11734_, _05023_ }), .Y(_11702_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28248_ ( .A({ _06995_, _stream_matmul_15_source_6_source_pat_fsm_0[1] }), .Y(_07007_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28249_ ( .A({ _11777_, _07007_, _11745_, _05023_ }), .Y(_11713_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28250_ ( .A({ _11788_, _07007_, _11756_, _05023_ }), .Y(_11724_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28251_ ( .A({ _11794_, _07007_, _11762_, _05023_ }), .Y(_11730_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28252_ ( .A({ _11791_, _07007_, _11759_, _05023_ }), .Y(_11727_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28253_ ( .A({ _11792_, _07007_, _11760_, _05023_ }), .Y(_11728_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28254_ ( .A({ _11793_, _07007_, _11761_, _05023_ }), .Y(_11729_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28255_ ( .A({ _11767_, _07007_, _11735_, _05023_ }), .Y(_11703_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28256_ ( .A({ _11795_, _07007_, _11763_, _05023_ }), .Y(_11731_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28257_ ( .A({ _11796_, _07007_, _11764_, _05023_ }), .Y(_11732_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28258_ ( .A({ _11797_, _07007_, _11765_, _05023_ }), .Y(_11733_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28259_ ( .A({ _11768_, _07007_, _11736_, _05023_ }), .Y(_11704_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28260_ ( .A({ _11769_, _07007_, _11737_, _05023_ }), .Y(_11705_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28261_ ( .A({ _11770_, _07007_, _11738_, _05023_ }), .Y(_11706_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28262_ ( .A({ _11771_, _07007_, _11739_, _05023_ }), .Y(_11707_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28263_ ( .A({ _11772_, _07007_, _11740_, _05023_ }), .Y(_11708_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28264_ ( .A({ _11776_, _07007_, _11744_, _05023_ }), .Y(_11712_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28265_ ( .A({ _11773_, _07007_, _11741_, _05023_ }), .Y(_11709_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28266_ ( .A({ _11774_, _07007_, _11742_, _05023_ }), .Y(_11710_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28267_ ( .A({ _11775_, _07007_, _11743_, _05023_ }), .Y(_11711_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28268_ ( .A({ _11781_, _07007_, _11749_, _05023_ }), .Y(_11717_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28269_ ( .A({ _11778_, _07007_, _11746_, _05023_ }), .Y(_11714_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28270_ ( .A({ _11779_, _07007_, _11747_, _05023_ }), .Y(_11715_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28271_ ( .A({ _11780_, _07007_, _11748_, _05023_ }), .Y(_11716_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28272_ ( .A({ _11782_, _07007_, _11750_, _05023_ }), .Y(_11718_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28273_ ( .A({ _11783_, _07007_, _11751_, _05023_ }), .Y(_11719_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28274_ ( .A({ _11784_, _07007_, _11752_, _05023_ }), .Y(_11720_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28275_ ( .A({ _11785_, _07007_, _11753_, _05023_ }), .Y(_11721_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28276_ ( .A({ _11786_, _07007_, _11754_, _05023_ }), .Y(_11722_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28277_ ( .A({ _11787_, _07007_, _11755_, _05023_ }), .Y(_11723_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28278_ ( .A({ _11789_, _07007_, _11757_, _05023_ }), .Y(_11725_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28279_ ( .A({ _11790_, _07007_, _11758_, _05023_ }), .Y(_11726_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _28280_ ( .A({ _18227_, _05107_, _18293_, _07019_ }), .Y(_18260_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _28281_ ( .A({ _07008_, _maxi_read_fsm[0], _07017_, _maxi_read_fsm[1] }), .Y(_05107_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28282_ ( .A({ _07014_, _07009_ }), .Y(_07008_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28283_ ( .A({ _07013_, _07012_, _07011_, _07010_ }), .Y(_07009_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28284_ ( .A(_maxi_read_fsm[23:20]), .Y(_07010_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28285_ ( .A(_maxi_read_fsm[19:16]), .Y(_07011_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28286_ ( .A(_maxi_read_fsm[31:28]), .Y(_07012_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28287_ ( .A(_maxi_read_fsm[27:24]), .Y(_07013_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28288_ ( .A({ _07016_, _07015_ }), .Y(_07014_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28289_ ( .A(_maxi_read_fsm[15:12]), .Y(_07015_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28290_ ( .A(_maxi_read_fsm[11:8]), .Y(_07016_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28291_ ( .A({ _07018_, _maxi_read_fsm[2], _maxi_read_fsm[3] }), .Y(_07017_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28292_ ( .A(_maxi_read_fsm[7:4]), .Y(_07018_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _28293_ ( .A({ _07017_, _07008_, _maxi_read_fsm[1:0] }), .Y(_07019_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28294_ ( .A({ _05025_, _07020_ }), .Y(_21884_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28295_ ( .A({ _07021_, _07026_, _stream_matmul_15_source_8_source_pat_fsm_1[0] }), .Y(_07020_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28296_ ( .A({ _07025_, _07024_, _07022_ }), .Y(_07021_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28297_ ( .A({ _07023_, _stream_matmul_15_source_8_source_pat_fsm_1[3:2] }), .Y(_07022_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28298_ ( .A(_stream_matmul_15_source_8_source_pat_fsm_1[7:4]), .Y(_07023_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28299_ ( .A(_stream_matmul_15_source_8_source_pat_fsm_1[15:12]), .Y(_07024_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28300_ ( .A(_stream_matmul_15_source_8_source_pat_fsm_1[11:8]), .Y(_07025_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28301_ ( .A({ _07030_, _07029_, _07028_, _07027_ }), .Y(_07026_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28302_ ( .A(_stream_matmul_15_source_8_source_pat_fsm_1[23:20]), .Y(_07027_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28303_ ( .A(_stream_matmul_15_source_8_source_pat_fsm_1[19:16]), .Y(_07028_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28304_ ( .A(_stream_matmul_15_source_8_source_pat_fsm_1[31:28]), .Y(_07029_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28305_ ( .A(_stream_matmul_15_source_8_source_pat_fsm_1[27:24]), .Y(_07030_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _28306_ ( .A({ _07021_, _stream_matmul_15_source_8_source_pat_fsm_1[0], _07026_, _stream_matmul_15_source_8_source_pat_fsm_1[1] }), .Y(_05025_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28307_ ( .A({ _11670_, _07031_, _11638_, _05025_ }), .Y(_11606_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28308_ ( .A({ _07020_, _stream_matmul_15_source_8_source_pat_fsm_1[1] }), .Y(_07031_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28309_ ( .A({ _11681_, _07031_, _11649_, _05025_ }), .Y(_11617_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28310_ ( .A({ _11692_, _07031_, _11660_, _05025_ }), .Y(_11628_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28311_ ( .A({ _11695_, _07031_, _11663_, _05025_ }), .Y(_11631_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28312_ ( .A({ _11696_, _07031_, _11664_, _05025_ }), .Y(_11632_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28313_ ( .A({ _11697_, _07031_, _11665_, _05025_ }), .Y(_11633_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28314_ ( .A({ _11698_, _07031_, _11666_, _05025_ }), .Y(_11634_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28315_ ( .A({ _11699_, _07031_, _11667_, _05025_ }), .Y(_11635_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28316_ ( .A({ _11700_, _07031_, _11668_, _05025_ }), .Y(_11636_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28317_ ( .A({ _11701_, _07031_, _11669_, _05025_ }), .Y(_11637_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28318_ ( .A({ _11671_, _07031_, _11639_, _05025_ }), .Y(_11607_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28319_ ( .A({ _11672_, _07031_, _11640_, _05025_ }), .Y(_11608_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28320_ ( .A({ _11673_, _07031_, _11641_, _05025_ }), .Y(_11609_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28321_ ( .A({ _11674_, _07031_, _11642_, _05025_ }), .Y(_11610_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28322_ ( .A({ _11675_, _07031_, _11643_, _05025_ }), .Y(_11611_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28323_ ( .A({ _11676_, _07031_, _11644_, _05025_ }), .Y(_11612_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28324_ ( .A({ _11677_, _07031_, _11645_, _05025_ }), .Y(_11613_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28325_ ( .A({ _11678_, _07031_, _11646_, _05025_ }), .Y(_11614_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28326_ ( .A({ _11679_, _07031_, _11647_, _05025_ }), .Y(_11615_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28327_ ( .A({ _11680_, _07031_, _11648_, _05025_ }), .Y(_11616_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28328_ ( .A({ _11682_, _07031_, _11650_, _05025_ }), .Y(_11618_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28329_ ( .A({ _11683_, _07031_, _11651_, _05025_ }), .Y(_11619_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28330_ ( .A({ _11684_, _07031_, _11652_, _05025_ }), .Y(_11620_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28331_ ( .A({ _11685_, _07031_, _11653_, _05025_ }), .Y(_11621_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28332_ ( .A({ _11686_, _07031_, _11654_, _05025_ }), .Y(_11622_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28333_ ( .A({ _11687_, _07031_, _11655_, _05025_ }), .Y(_11623_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28334_ ( .A({ _11688_, _07031_, _11656_, _05025_ }), .Y(_11624_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28335_ ( .A({ _11689_, _07031_, _11657_, _05025_ }), .Y(_11625_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28336_ ( .A({ _11690_, _07031_, _11658_, _05025_ }), .Y(_11626_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28337_ ( .A({ _11691_, _07031_, _11659_, _05025_ }), .Y(_11627_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28338_ ( .A({ _11693_, _07031_, _11661_, _05025_ }), .Y(_11629_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28339_ ( .A({ _11694_, _07031_, _11662_, _05025_ }), .Y(_11630_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28340_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16071_, _16103_ }), .Y(_16039_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28341_ ( .A({ _07033_, _07041_, _stream_conv2d_8_source_30_source_pat_fsm_13[1] }), .Y(_07032_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28342_ ( .A({ _07040_, _07039_, _07034_ }), .Y(_07033_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28343_ ( .A({ _07038_, _07037_, _07036_, _07035_ }), .Y(_07034_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28344_ ( .A(_stream_conv2d_8_source_30_source_pat_fsm_13[23:20]), .Y(_07035_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28345_ ( .A(_stream_conv2d_8_source_30_source_pat_fsm_13[19:16]), .Y(_07036_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28346_ ( .A(_stream_conv2d_8_source_30_source_pat_fsm_13[31:28]), .Y(_07037_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28347_ ( .A(_stream_conv2d_8_source_30_source_pat_fsm_13[27:24]), .Y(_07038_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28348_ ( .A(_stream_conv2d_8_source_30_source_pat_fsm_13[15:12]), .Y(_07039_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28349_ ( .A(_stream_conv2d_8_source_30_source_pat_fsm_13[11:8]), .Y(_07040_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28350_ ( .A({ _07042_, _stream_conv2d_8_source_30_source_pat_fsm_13[3:2] }), .Y(_07041_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28351_ ( .A(_stream_conv2d_8_source_30_source_pat_fsm_13[7:4]), .Y(_07042_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28352_ ( .A({ _05021_, _07043_ }), .Y(_21883_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28353_ ( .A({ _07052_, _07049_, _07044_ }), .Y(_07043_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28354_ ( .A({ _07048_, _07047_, _07046_, _07045_ }), .Y(_07044_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28355_ ( .A(_stream_matmul_15_source_19_source_pat_fsm_2[23:20]), .Y(_07045_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28356_ ( .A(_stream_matmul_15_source_19_source_pat_fsm_2[19:16]), .Y(_07046_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28357_ ( .A(_stream_matmul_15_source_19_source_pat_fsm_2[31:28]), .Y(_07047_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28358_ ( .A(_stream_matmul_15_source_19_source_pat_fsm_2[27:24]), .Y(_07048_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28359_ ( .A({ _07051_, _07050_ }), .Y(_07049_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28360_ ( .A(_stream_matmul_15_source_19_source_pat_fsm_2[15:12]), .Y(_07050_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28361_ ( .A(_stream_matmul_15_source_19_source_pat_fsm_2[11:8]), .Y(_07051_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _28362_ ( .A({ _07053_, _stream_matmul_15_source_19_source_pat_fsm_2[3:2], _stream_matmul_15_source_19_source_pat_fsm_2[0] }), .Y(_07052_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28363_ ( .A(_stream_matmul_15_source_19_source_pat_fsm_2[7:4]), .Y(_07053_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _28364_ ( .A({ _07054_, _07053_, _07049_, _07044_ }), .Y(_05021_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _28365_ ( .A({ _stream_matmul_15_source_19_source_pat_fsm_2[0], _stream_matmul_15_source_19_source_pat_fsm_2[3:1] }), .Y(_07054_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28366_ ( .A({ _11574_, _07055_, _11542_, _05021_ }), .Y(_11510_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28367_ ( .A({ _07043_, _stream_matmul_15_source_19_source_pat_fsm_2[1] }), .Y(_07055_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28368_ ( .A({ _11585_, _07055_, _11553_, _05021_ }), .Y(_11521_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28369_ ( .A({ _11596_, _07055_, _11564_, _05021_ }), .Y(_11532_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28370_ ( .A({ _11599_, _07055_, _11567_, _05021_ }), .Y(_11535_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28371_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17108_, _17140_ }), .Y(_17076_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28372_ ( .A({ _07057_, _07065_, _stream_conv2d_8_source_19_source_pat_fsm_2[1] }), .Y(_07056_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28373_ ( .A({ _07064_, _07063_, _07058_ }), .Y(_07057_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28374_ ( .A({ _07062_, _07061_, _07060_, _07059_ }), .Y(_07058_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28375_ ( .A(_stream_conv2d_8_source_19_source_pat_fsm_2[23:20]), .Y(_07059_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28376_ ( .A(_stream_conv2d_8_source_19_source_pat_fsm_2[19:16]), .Y(_07060_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28377_ ( .A(_stream_conv2d_8_source_19_source_pat_fsm_2[31:28]), .Y(_07061_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28378_ ( .A(_stream_conv2d_8_source_19_source_pat_fsm_2[27:24]), .Y(_07062_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28379_ ( .A(_stream_conv2d_8_source_19_source_pat_fsm_2[15:12]), .Y(_07063_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28380_ ( .A(_stream_conv2d_8_source_19_source_pat_fsm_2[11:8]), .Y(_07064_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28381_ ( .A({ _07066_, _stream_conv2d_8_source_19_source_pat_fsm_2[3:2] }), .Y(_07065_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28382_ ( .A(_stream_conv2d_8_source_19_source_pat_fsm_2[7:4]), .Y(_07066_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28383_ ( .A({ _11600_, _07055_, _11568_, _05021_ }), .Y(_11536_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28384_ ( .A({ _11601_, _07055_, _11569_, _05021_ }), .Y(_11537_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28385_ ( .A({ _11602_, _07055_, _11570_, _05021_ }), .Y(_11538_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28386_ ( .A({ _11603_, _07055_, _11571_, _05021_ }), .Y(_11539_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28387_ ( .A({ _11604_, _07055_, _11572_, _05021_ }), .Y(_11540_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28388_ ( .A({ _11605_, _07055_, _11573_, _05021_ }), .Y(_11541_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28389_ ( .A({ _11575_, _07055_, _11543_, _05021_ }), .Y(_11511_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28390_ ( .A({ _11576_, _07055_, _11544_, _05021_ }), .Y(_11512_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28391_ ( .A({ _11577_, _07055_, _11545_, _05021_ }), .Y(_11513_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28392_ ( .A({ _11578_, _07055_, _11546_, _05021_ }), .Y(_11514_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28393_ ( .A({ _11579_, _07055_, _11547_, _05021_ }), .Y(_11515_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28394_ ( .A({ _11580_, _07055_, _11548_, _05021_ }), .Y(_11516_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28395_ ( .A({ _05071_, _07067_ }), .Y(_21906_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28396_ ( .A({ _07068_, _07073_, _stream_conv2d_8_source_31_source_pat_fsm_14[0] }), .Y(_07067_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28397_ ( .A({ _07072_, _07071_, _07069_ }), .Y(_07068_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28398_ ( .A({ _07070_, _stream_conv2d_8_source_31_source_pat_fsm_14[3:2] }), .Y(_07069_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28399_ ( .A(_stream_conv2d_8_source_31_source_pat_fsm_14[7:4]), .Y(_07070_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28400_ ( .A(_stream_conv2d_8_source_31_source_pat_fsm_14[15:12]), .Y(_07071_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28401_ ( .A(_stream_conv2d_8_source_31_source_pat_fsm_14[11:8]), .Y(_07072_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28402_ ( .A({ _07077_, _07076_, _07075_, _07074_ }), .Y(_07073_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28403_ ( .A(_stream_conv2d_8_source_31_source_pat_fsm_14[23:20]), .Y(_07074_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28404_ ( .A(_stream_conv2d_8_source_31_source_pat_fsm_14[19:16]), .Y(_07075_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28405_ ( .A(_stream_conv2d_8_source_31_source_pat_fsm_14[31:28]), .Y(_07076_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28406_ ( .A(_stream_conv2d_8_source_31_source_pat_fsm_14[27:24]), .Y(_07077_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _28407_ ( .A({ _07068_, _stream_conv2d_8_source_31_source_pat_fsm_14[0], _07073_, _stream_conv2d_8_source_31_source_pat_fsm_14[1] }), .Y(_05071_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28408_ ( .A({ _11581_, _07055_, _11549_, _05021_ }), .Y(_11517_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28409_ ( .A({ _11582_, _07055_, _11550_, _05021_ }), .Y(_11518_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28410_ ( .A({ _11583_, _07055_, _11551_, _05021_ }), .Y(_11519_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28411_ ( .A({ _11584_, _07055_, _11552_, _05021_ }), .Y(_11520_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28412_ ( .A({ _11586_, _07055_, _11554_, _05021_ }), .Y(_11522_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28413_ ( .A({ _11587_, _07055_, _11555_, _05021_ }), .Y(_11523_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28414_ ( .A({ _11588_, _07055_, _11556_, _05021_ }), .Y(_11524_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28415_ ( .A({ _11589_, _07055_, _11557_, _05021_ }), .Y(_11525_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28416_ ( .A({ _11590_, _07055_, _11558_, _05021_ }), .Y(_11526_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28417_ ( .A({ _11591_, _07055_, _11559_, _05021_ }), .Y(_11527_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28418_ ( .A({ _11592_, _07055_, _11560_, _05021_ }), .Y(_11528_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28419_ ( .A({ _11593_, _07055_, _11561_, _05021_ }), .Y(_11529_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28420_ ( .A({ _11594_, _07055_, _11562_, _05021_ }), .Y(_11530_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28421_ ( .A({ _11595_, _07055_, _11563_, _05021_ }), .Y(_11531_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28422_ ( .A({ _11597_, _07055_, _11565_, _05021_ }), .Y(_11533_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28423_ ( .A({ _11598_, _07055_, _11566_, _05021_ }), .Y(_11534_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28424_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16070_, _16102_ }), .Y(_16038_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28425_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17107_, _17139_ }), .Y(_17075_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28426_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16069_, _16101_ }), .Y(_16037_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28427_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16548_, _16580_ }), .Y(_16516_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28428_ ( .A({ _07079_, _07087_, _stream_conv2d_8_source_25_source_pat_fsm_8[1] }), .Y(_07078_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28429_ ( .A({ _07086_, _07085_, _07080_ }), .Y(_07079_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28430_ ( .A({ _07084_, _07083_, _07082_, _07081_ }), .Y(_07080_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28431_ ( .A(_stream_conv2d_8_source_25_source_pat_fsm_8[23:20]), .Y(_07081_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28432_ ( .A(_stream_conv2d_8_source_25_source_pat_fsm_8[19:16]), .Y(_07082_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28433_ ( .A(_stream_conv2d_8_source_25_source_pat_fsm_8[31:28]), .Y(_07083_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28434_ ( .A(_stream_conv2d_8_source_25_source_pat_fsm_8[27:24]), .Y(_07084_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28435_ ( .A(_stream_conv2d_8_source_25_source_pat_fsm_8[15:12]), .Y(_07085_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28436_ ( .A(_stream_conv2d_8_source_25_source_pat_fsm_8[11:8]), .Y(_07086_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28437_ ( .A({ _07088_, _stream_conv2d_8_source_25_source_pat_fsm_8[3:2] }), .Y(_07087_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28438_ ( .A(_stream_conv2d_8_source_25_source_pat_fsm_8[7:4]), .Y(_07088_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28439_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17106_, _17138_ }), .Y(_17074_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28440_ ( .A({ _05020_, _07089_ }), .Y(_21882_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28441_ ( .A({ _07090_, _07095_, _stream_matmul_15_source_20_source_pat_fsm_3[0] }), .Y(_07089_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28442_ ( .A({ _07094_, _07093_, _07091_ }), .Y(_07090_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28443_ ( .A({ _07092_, _stream_matmul_15_source_20_source_pat_fsm_3[3:2] }), .Y(_07091_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28444_ ( .A(_stream_matmul_15_source_20_source_pat_fsm_3[7:4]), .Y(_07092_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28445_ ( .A(_stream_matmul_15_source_20_source_pat_fsm_3[15:12]), .Y(_07093_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28446_ ( .A(_stream_matmul_15_source_20_source_pat_fsm_3[11:8]), .Y(_07094_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28447_ ( .A({ _07099_, _07098_, _07097_, _07096_ }), .Y(_07095_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28448_ ( .A(_stream_matmul_15_source_20_source_pat_fsm_3[23:20]), .Y(_07096_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28449_ ( .A(_stream_matmul_15_source_20_source_pat_fsm_3[19:16]), .Y(_07097_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28450_ ( .A(_stream_matmul_15_source_20_source_pat_fsm_3[31:28]), .Y(_07098_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28451_ ( .A(_stream_matmul_15_source_20_source_pat_fsm_3[27:24]), .Y(_07099_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _28452_ ( .A({ _07090_, _stream_matmul_15_source_20_source_pat_fsm_3[0], _07095_, _stream_matmul_15_source_20_source_pat_fsm_3[1] }), .Y(_05020_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28453_ ( .A({ _11478_, _07100_, _11446_, _05020_ }), .Y(_11414_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28454_ ( .A({ _07089_, _stream_matmul_15_source_20_source_pat_fsm_3[1] }), .Y(_07100_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28455_ ( .A({ _11489_, _07100_, _11457_, _05020_ }), .Y(_11425_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28456_ ( .A({ _11500_, _07100_, _11468_, _05020_ }), .Y(_11436_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28457_ ( .A({ _11503_, _07100_, _11471_, _05020_ }), .Y(_11439_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28458_ ( .A({ _11504_, _07100_, _11472_, _05020_ }), .Y(_11440_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28459_ ( .A({ _11505_, _07100_, _11473_, _05020_ }), .Y(_11441_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28460_ ( .A({ _11506_, _07100_, _11474_, _05020_ }), .Y(_11442_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28461_ ( .A({ _11507_, _07100_, _11475_, _05020_ }), .Y(_11443_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28462_ ( .A({ _11508_, _07100_, _11476_, _05020_ }), .Y(_11444_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28463_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16066_, _16098_ }), .Y(_16034_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28464_ ( .A({ _11509_, _07100_, _11477_, _05020_ }), .Y(_11445_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28465_ ( .A({ _11479_, _07100_, _11447_, _05020_ }), .Y(_11415_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28466_ ( .A({ _11480_, _07100_, _11448_, _05020_ }), .Y(_11416_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28467_ ( .A({ _11481_, _07100_, _11449_, _05020_ }), .Y(_11417_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28468_ ( .A({ _11482_, _07100_, _11450_, _05020_ }), .Y(_11418_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28469_ ( .A({ _11483_, _07100_, _11451_, _05020_ }), .Y(_11419_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28470_ ( .A({ _11484_, _07100_, _11452_, _05020_ }), .Y(_11420_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28471_ ( .A({ _11485_, _07100_, _11453_, _05020_ }), .Y(_11421_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28472_ ( .A({ _11486_, _07100_, _11454_, _05020_ }), .Y(_11422_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28473_ ( .A({ _11487_, _07100_, _11455_, _05020_ }), .Y(_11423_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28474_ ( .A({ _11488_, _07100_, _11456_, _05020_ }), .Y(_11424_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28475_ ( .A({ _11490_, _07100_, _11458_, _05020_ }), .Y(_11426_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28476_ ( .A({ _11491_, _07100_, _11459_, _05020_ }), .Y(_11427_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28477_ ( .A({ _11492_, _07100_, _11460_, _05020_ }), .Y(_11428_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28478_ ( .A({ _11493_, _07100_, _11461_, _05020_ }), .Y(_11429_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28479_ ( .A({ _11494_, _07100_, _11462_, _05020_ }), .Y(_11430_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28480_ ( .A({ _11495_, _07100_, _11463_, _05020_ }), .Y(_11431_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28481_ ( .A({ _11496_, _07100_, _11464_, _05020_ }), .Y(_11432_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28482_ ( .A({ _11497_, _07100_, _11465_, _05020_ }), .Y(_11433_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28483_ ( .A({ _11498_, _07100_, _11466_, _05020_ }), .Y(_11434_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28484_ ( .A({ _11499_, _07100_, _11467_, _05020_ }), .Y(_11435_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28485_ ( .A({ _11501_, _07100_, _11469_, _05020_ }), .Y(_11437_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28486_ ( .A({ _11502_, _07100_, _11470_, _05020_ }), .Y(_11438_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28487_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16547_, _16579_ }), .Y(_16515_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28488_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17105_, _17137_ }), .Y(_17073_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28489_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16545_, _16577_ }), .Y(_16513_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28490_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17103_, _17135_ }), .Y(_17071_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28491_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16544_, _16576_ }), .Y(_16512_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28492_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17102_, _17134_ }), .Y(_17070_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28493_ ( .A({ _07109_, _07108_, _07103_, _07101_ }), .Y(_21881_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _28494_ ( .A({ _07102_, _stream_matmul_15_sink_21_sink_fsm_4[31:29] }), .Y(_07101_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28495_ ( .A(_stream_matmul_15_sink_21_sink_fsm_4[28:25]), .Y(_07102_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28496_ ( .A({ _07107_, _07106_, _07105_, _07104_ }), .Y(_07103_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28497_ ( .A(_stream_matmul_15_sink_21_sink_fsm_4[8:5]), .Y(_07104_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28498_ ( .A(_stream_matmul_15_sink_21_sink_fsm_4[4:1]), .Y(_07105_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28499_ ( .A(_stream_matmul_15_sink_21_sink_fsm_4[16:13]), .Y(_07106_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28500_ ( .A(_stream_matmul_15_sink_21_sink_fsm_4[12:9]), .Y(_07107_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28501_ ( .A(_stream_matmul_15_sink_21_sink_fsm_4[24:21]), .Y(_07108_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28502_ ( .A(_stream_matmul_15_sink_21_sink_fsm_4[20:17]), .Y(_07109_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28503_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11318_, _11382_ }), .Y(_11350_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28504_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11329_, _11393_ }), .Y(_11361_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28505_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11340_, _11404_ }), .Y(_11372_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28506_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11343_, _11407_ }), .Y(_11375_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28507_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11344_, _11408_ }), .Y(_11376_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28508_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11345_, _11409_ }), .Y(_11377_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28509_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11346_, _11410_ }), .Y(_11378_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28510_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11347_, _11411_ }), .Y(_11379_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28511_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11348_, _11412_ }), .Y(_11380_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28512_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11349_, _11413_ }), .Y(_11381_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28513_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11319_, _11383_ }), .Y(_11351_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28514_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11320_, _11384_ }), .Y(_11352_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28515_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11321_, _11385_ }), .Y(_11353_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28516_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11322_, _11386_ }), .Y(_11354_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28517_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11323_, _11387_ }), .Y(_11355_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28518_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11324_, _11388_ }), .Y(_11356_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28519_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11325_, _11389_ }), .Y(_11357_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28520_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11326_, _11390_ }), .Y(_11358_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28521_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11327_, _11391_ }), .Y(_11359_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28522_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11328_, _11392_ }), .Y(_11360_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28523_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11330_, _11394_ }), .Y(_11362_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28524_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11331_, _11395_ }), .Y(_11363_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28525_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11332_, _11396_ }), .Y(_11364_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28526_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11333_, _11397_ }), .Y(_11365_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28527_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16543_, _16575_ }), .Y(_16511_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28528_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11334_, _11398_ }), .Y(_11366_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28529_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11335_, _11399_ }), .Y(_11367_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28530_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11336_, _11400_ }), .Y(_11368_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28531_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11337_, _11401_ }), .Y(_11369_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28532_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11338_, _11402_ }), .Y(_11370_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28533_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11339_, _11403_ }), .Y(_11371_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28534_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11341_, _11405_ }), .Y(_11373_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28535_ ( .A({ _21881_, _stream_matmul_15_sink_21_sink_fsm_4[0], _11342_, _11406_ }), .Y(_11374_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28536_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17101_, _17133_ }), .Y(_17069_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28537_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16542_, _16574_ }), .Y(_16510_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28538_ ( .A({ _07110_, _17380_, _07122_ }), .Y(_17412_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28539_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17444_, _17476_ }), .Y(_07110_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28540_ ( .A({ _07112_, _07119_, conv2d_8_comp_fsm[3] }), .Y(_07111_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _28541_ ( .A({ _07118_, _07113_, conv2d_8_comp_fsm[1:0] }), .Y(_07112_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28542_ ( .A({ _07117_, _07116_, _07115_, _07114_ }), .Y(_07113_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28543_ ( .A(conv2d_8_comp_fsm[23:20]), .Y(_07114_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28544_ ( .A(conv2d_8_comp_fsm[19:16]), .Y(_07115_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28545_ ( .A(conv2d_8_comp_fsm[31:28]), .Y(_07116_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28546_ ( .A(conv2d_8_comp_fsm[27:24]), .Y(_07117_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28547_ ( .A(conv2d_8_comp_fsm[7:4]), .Y(_07118_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28548_ ( .A({ _07121_, _07120_ }), .Y(_07119_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28549_ ( .A(conv2d_8_comp_fsm[15:12]), .Y(_07120_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28550_ ( .A(conv2d_8_comp_fsm[11:8]), .Y(_07121_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28551_ ( .A({ _07124_, _07123_ }), .Y(_07122_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _28552_ ( .A({ conv2d_8_comp_fsm[1], _07119_, _07113_, conv2d_8_comp_fsm[0] }), .Y(_07123_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28553_ ( .A({ conv2d_8_comp_fsm[2], _07118_, conv2d_8_comp_fsm[3] }), .Y(_07124_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28554_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17131_, _17163_ }), .Y(_17099_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28555_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16541_, _16573_ }), .Y(_16509_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28556_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17130_, _17162_ }), .Y(_17098_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28557_ ( .A({ _07125_, _17379_, _07122_ }), .Y(_17411_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28558_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17443_, _17475_ }), .Y(_07125_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28559_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16540_, _16572_ }), .Y(_16508_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28560_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17129_, _17161_ }), .Y(_17097_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28561_ ( .A({ _07126_, _17377_, _07122_ }), .Y(_17409_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28562_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17441_, _17473_ }), .Y(_07126_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28563_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16356_, _16388_ }), .Y(_16324_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28564_ ( .A({ _07128_, _07136_, _stream_conv2d_8_source_27_source_pat_fsm_10[1] }), .Y(_07127_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28565_ ( .A({ _07135_, _07134_, _07129_ }), .Y(_07128_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28566_ ( .A({ _07133_, _07132_, _07131_, _07130_ }), .Y(_07129_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28567_ ( .A(_stream_conv2d_8_source_27_source_pat_fsm_10[23:20]), .Y(_07130_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28568_ ( .A(_stream_conv2d_8_source_27_source_pat_fsm_10[19:16]), .Y(_07131_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28569_ ( .A(_stream_conv2d_8_source_27_source_pat_fsm_10[31:28]), .Y(_07132_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28570_ ( .A(_stream_conv2d_8_source_27_source_pat_fsm_10[27:24]), .Y(_07133_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28571_ ( .A(_stream_conv2d_8_source_27_source_pat_fsm_10[15:12]), .Y(_07134_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28572_ ( .A(_stream_conv2d_8_source_27_source_pat_fsm_10[11:8]), .Y(_07135_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28573_ ( .A({ _07137_, _stream_conv2d_8_source_27_source_pat_fsm_10[3:2] }), .Y(_07136_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28574_ ( .A(_stream_conv2d_8_source_27_source_pat_fsm_10[7:4]), .Y(_07137_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28575_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16538_, _16570_ }), .Y(_16506_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28576_ ( .A({ _07138_, _17376_, _07122_ }), .Y(_17408_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28577_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17440_, _17472_ }), .Y(_07138_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28578_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17128_, _17160_ }), .Y(_17096_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28579_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16536_, _16568_ }), .Y(_16504_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28580_ ( .A({ _07139_, _17375_, _07122_ }), .Y(_17407_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28581_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17439_, _17471_ }), .Y(_07139_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28582_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17127_, _17159_ }), .Y(_17095_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28583_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16534_, _16566_ }), .Y(_16502_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28584_ ( .A({ _07140_, _17374_, _07122_ }), .Y(_17406_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28585_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17438_, _17470_ }), .Y(_07140_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28586_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17126_, _17158_ }), .Y(_17094_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28587_ ( .A({ _07141_, _17373_, _07122_ }), .Y(_17405_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28588_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17437_, _17469_ }), .Y(_07141_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28589_ ( .A({ _07142_, _17372_, _07122_ }), .Y(_17404_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28590_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17436_, _17468_ }), .Y(_07142_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28591_ ( .A({ _07143_, _17371_, _07122_ }), .Y(_17403_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28592_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17435_, _17467_ }), .Y(_07143_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28593_ ( .A({ _05102_, _07122_ }), .Y(_21922_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _28594_ ( .A({ _07144_, _07145_, conv2d_8_comp_fsm[1] }), .Y(_05102_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28595_ ( .A({ conv2d_8_comp_fsm[0], _07113_, _07119_ }), .Y(_07144_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28596_ ( .A({ _07118_, conv2d_8_comp_fsm[2], conv2d_8_comp_fsm[3] }), .Y(_07145_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28597_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16055_, _16087_ }), .Y(_16023_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28598_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16355_, _16387_ }), .Y(_16323_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28599_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16533_, _16565_ }), .Y(_16501_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28600_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17122_, _17154_ }), .Y(_17090_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28601_ ( .A({ _07146_, _17370_, _07122_ }), .Y(_17402_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28602_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17434_, _17466_ }), .Y(_07146_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28603_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16044_, _16076_ }), .Y(_16012_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28604_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16353_, _16385_ }), .Y(_16321_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28605_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16532_, _16564_ }), .Y(_16500_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28606_ ( .A({ _07147_, _17369_, _07122_ }), .Y(_17401_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28607_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17433_, _17465_ }), .Y(_07147_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28608_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17111_, _17143_ }), .Y(_17079_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28609_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16164_, _16196_ }), .Y(_16132_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28610_ ( .A({ _07149_, _07157_, _stream_conv2d_8_source_29_source_pat_fsm_12[1] }), .Y(_07148_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28611_ ( .A({ _07156_, _07155_, _07150_ }), .Y(_07149_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28612_ ( .A({ _07154_, _07153_, _07152_, _07151_ }), .Y(_07150_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28613_ ( .A(_stream_conv2d_8_source_29_source_pat_fsm_12[23:20]), .Y(_07151_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28614_ ( .A(_stream_conv2d_8_source_29_source_pat_fsm_12[19:16]), .Y(_07152_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28615_ ( .A(_stream_conv2d_8_source_29_source_pat_fsm_12[31:28]), .Y(_07153_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28616_ ( .A(_stream_conv2d_8_source_29_source_pat_fsm_12[27:24]), .Y(_07154_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28617_ ( .A(_stream_conv2d_8_source_29_source_pat_fsm_12[15:12]), .Y(_07155_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28618_ ( .A(_stream_conv2d_8_source_29_source_pat_fsm_12[11:8]), .Y(_07156_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28619_ ( .A({ _07158_, _stream_conv2d_8_source_29_source_pat_fsm_12[3:2] }), .Y(_07157_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28620_ ( .A(_stream_conv2d_8_source_29_source_pat_fsm_12[7:4]), .Y(_07158_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28621_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16352_, _16384_ }), .Y(_16320_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28622_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16531_, _16563_ }), .Y(_16499_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28623_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17100_, _17132_ }), .Y(_17068_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28624_ ( .A({ _07159_, _17368_, _07122_ }), .Y(_17400_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28625_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17432_, _17464_ }), .Y(_07159_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28626_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16351_, _16383_ }), .Y(_16319_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28627_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16530_, _16562_ }), .Y(_16498_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28628_ ( .A({ _07160_, _17366_, _07122_ }), .Y(_17398_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28629_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17430_, _17462_ }), .Y(_07160_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28630_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16350_, _16382_ }), .Y(_16318_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28631_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16529_, _16561_ }), .Y(_16497_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28632_ ( .A({ _07161_, _17365_, _07122_ }), .Y(_17397_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28633_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17429_, _17461_ }), .Y(_07161_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28634_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16349_, _16381_ }), .Y(_16317_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28635_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16528_, _16560_ }), .Y(_16496_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28636_ ( .A({ _07162_, _17364_, _07122_ }), .Y(_17396_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28637_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17428_, _17460_ }), .Y(_07162_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28638_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16348_, _16380_ }), .Y(_16316_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28639_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16527_, _16559_ }), .Y(_16495_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28640_ ( .A({ _07163_, _17363_, _07122_ }), .Y(_17395_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28641_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17427_, _17459_ }), .Y(_07163_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28642_ ( .A({ _05094_, _07056_ }), .Y(_21918_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _28643_ ( .A({ _stream_conv2d_8_source_19_source_pat_fsm_2[1], _07057_, _07065_, _stream_conv2d_8_source_19_source_pat_fsm_2[0] }), .Y(_05094_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28644_ ( .A({ _07164_, _17362_, _07122_ }), .Y(_17394_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28645_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17426_, _17458_ }), .Y(_07164_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28646_ ( .A({ _07165_, _17361_, _07122_ }), .Y(_17393_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28647_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17425_, _17457_ }), .Y(_07165_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28648_ ( .A({ _07166_, _17360_, _07122_ }), .Y(_17392_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28649_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17424_, _17456_ }), .Y(_07166_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28650_ ( .A({ _07167_, _17359_, _07122_ }), .Y(_17391_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28651_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17423_, _17455_ }), .Y(_07167_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28652_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16163_, _16195_ }), .Y(_16131_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28653_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16347_, _16379_ }), .Y(_16315_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28654_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16526_, _16558_ }), .Y(_16494_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28655_ ( .A({ _07168_, _17358_, _07122_ }), .Y(_17390_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28656_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17422_, _17454_ }), .Y(_07168_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _28657_ ( .A({ _07177_, _07176_, _07171_, _07169_ }), .Y(_05232_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _28658_ ( .A({ _07170_, matmul_15_och_count[31:29] }), .Y(_07169_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28659_ ( .A(matmul_15_och_count[28:25]), .Y(_07170_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28660_ ( .A({ _07175_, _07174_, _07173_, _07172_ }), .Y(_07171_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28661_ ( .A(matmul_15_och_count[16:13]), .Y(_07172_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28662_ ( .A(matmul_15_och_count[12:9]), .Y(_07173_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28663_ ( .A(matmul_15_och_count[8:5]), .Y(_07174_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _28664_ ( .A({ matmul_15_och_count[4:3], matmul_15_och_count[1], matmul_15_och_count[2] }), .Y(_07175_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28665_ ( .A(matmul_15_och_count[24:21]), .Y(_07176_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28666_ ( .A(matmul_15_och_count[20:17]), .Y(_07177_) );
  \$lut  #( .LUT(16'hf2ff), .WIDTH(4) ) _28667_ ( .A({ _07223_, _07200_, _07178_, _07220_ }), .Y(_05248_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _28668_ ( .A({ _07197_, _07194_, _07191_, _07179_ }), .Y(_07178_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _28669_ ( .A({ _07186_, _07190_, _07180_, _07189_ }), .Y(_07179_) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _28670_ ( .A({ matmul_15_sync_comp_count[5], _07181_, _07185_, _04343_ }), .Y(_07180_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _28671_ ( .A({ _07184_, _04341_, matmul_15_sync_comp_count[3], _07182_ }), .Y(_07181_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _28672_ ( .A({ _04338_, matmul_15_sync_comp_count[2], _07183_ }), .Y(_07182_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _28673_ ( .A({ _04316_, matmul_15_sync_comp_count[0], matmul_15_sync_comp_count[1], _04327_ }), .Y(_07183_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28674_ ( .A({ matmul_15_sync_comp_count[4], _04342_ }), .Y(_07184_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28675_ ( .A({ _04342_, matmul_15_sync_comp_count[4] }), .Y(_07185_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _28676_ ( .A({ _07188_, _07187_, _04345_, matmul_15_sync_comp_count[7] }), .Y(_07186_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28677_ ( .A({ matmul_15_sync_comp_count[11], _04318_, matmul_15_sync_comp_count[10], _04317_ }), .Y(_07187_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28678_ ( .A({ matmul_15_sync_comp_count[9], _04347_, matmul_15_sync_comp_count[8], _04346_ }), .Y(_07188_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28679_ ( .A({ _04344_, matmul_15_sync_comp_count[6] }), .Y(_07189_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _28680_ ( .A({ matmul_15_sync_comp_count[6], _04344_, matmul_15_sync_comp_count[7], _04345_ }), .Y(_07190_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _28681_ ( .A({ _07192_, _07187_, _07193_ }), .Y(_07191_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28682_ ( .A({ matmul_15_sync_comp_count[10], matmul_15_sync_comp_count[11], _04317_, _04318_ }), .Y(_07192_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28683_ ( .A({ matmul_15_sync_comp_count[8], matmul_15_sync_comp_count[9], _04346_, _04347_ }), .Y(_07193_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28684_ ( .A({ _07196_, _07195_ }), .Y(_07194_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28685_ ( .A({ matmul_15_sync_comp_count[15], _04322_, matmul_15_sync_comp_count[14], _04321_ }), .Y(_07195_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28686_ ( .A({ matmul_15_sync_comp_count[13], _04320_, matmul_15_sync_comp_count[12], _04319_ }), .Y(_07196_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _28687_ ( .A({ _07199_, _07195_, _07198_ }), .Y(_07197_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28688_ ( .A({ matmul_15_sync_comp_count[12], matmul_15_sync_comp_count[13], _04319_, _04320_ }), .Y(_07198_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _28689_ ( .A({ matmul_15_sync_comp_count[14], matmul_15_sync_comp_count[15], _04321_, _04322_ }), .Y(_07199_) );
  \$lut  #( .LUT(16'hf400), .WIDTH(4) ) _28690_ ( .A({ _07215_, _07219_, _07218_, _07201_ }), .Y(_07200_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _28691_ ( .A({ _07214_, _07202_, _07213_ }), .Y(_07201_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _28692_ ( .A({ _07207_, _07203_, _07209_ }), .Y(_07202_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _28693_ ( .A({ _07206_, _07204_, _04328_, matmul_15_sync_comp_count[20] }), .Y(_07203_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _28694_ ( .A({ _07205_, _04329_, matmul_15_sync_comp_count[21] }), .Y(_07204_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28695_ ( .A({ matmul_15_sync_comp_count[23], _04331_, matmul_15_sync_comp_count[22], _04330_ }), .Y(_07205_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _28696_ ( .A({ matmul_15_sync_comp_count[20], _04328_, matmul_15_sync_comp_count[21], _04329_ }), .Y(_07206_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _28697_ ( .A({ _07208_, _07204_, _07206_ }), .Y(_07207_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _28698_ ( .A({ matmul_15_sync_comp_count[22], matmul_15_sync_comp_count[23], _04330_, _04331_ }), .Y(_07208_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _28699_ ( .A({ _07211_, _07210_, _07212_ }), .Y(_07209_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28700_ ( .A({ matmul_15_sync_comp_count[19], _04326_, matmul_15_sync_comp_count[18], _04325_ }), .Y(_07210_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28701_ ( .A({ matmul_15_sync_comp_count[18], matmul_15_sync_comp_count[19], _04325_, _04326_ }), .Y(_07211_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28702_ ( .A({ matmul_15_sync_comp_count[16], matmul_15_sync_comp_count[17], _04323_, _04324_ }), .Y(_07212_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28703_ ( .A({ matmul_15_sync_comp_count[25], _04333_, matmul_15_sync_comp_count[24], _04332_ }), .Y(_07213_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28704_ ( .A({ matmul_15_sync_comp_count[24], matmul_15_sync_comp_count[25], _04332_, _04333_ }), .Y(_07214_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28705_ ( .A({ _07217_, _07216_ }), .Y(_07215_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28706_ ( .A({ matmul_15_sync_comp_count[31], _04340_, matmul_15_sync_comp_count[30], _04339_ }), .Y(_07216_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28707_ ( .A({ matmul_15_sync_comp_count[29], _04337_, matmul_15_sync_comp_count[28], _04336_ }), .Y(_07217_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28708_ ( .A({ matmul_15_sync_comp_count[27], _04335_, matmul_15_sync_comp_count[26], _04334_ }), .Y(_07218_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28709_ ( .A({ matmul_15_sync_comp_count[26], matmul_15_sync_comp_count[27], _04334_, _04335_ }), .Y(_07219_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28710_ ( .A({ _07222_, _07213_, _07221_ }), .Y(_07220_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28711_ ( .A({ _07210_, _07218_, _07215_, _07203_ }), .Y(_07221_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28712_ ( .A({ matmul_15_sync_comp_count[17], _04324_, matmul_15_sync_comp_count[16], _04323_ }), .Y(_07222_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28713_ ( .A({ _07226_, _07224_ }), .Y(_07223_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _28714_ ( .A({ _07216_, matmul_15_sync_comp_count[29], _04337_, _07225_ }), .Y(_07224_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28715_ ( .A({ matmul_15_sync_comp_count[28], _04336_ }), .Y(_07225_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _28716_ ( .A({ matmul_15_sync_comp_count[30], matmul_15_sync_comp_count[31], _04339_, _04340_ }), .Y(_07226_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28717_ ( .A({ _07227_, _17357_, _07122_ }), .Y(_17389_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28718_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17421_, _17453_ }), .Y(_07227_) );
  \$lut  #( .LUT(16'h0bff), .WIDTH(4) ) _28719_ ( .A({ _07232_, _07228_, cparam_max_pool_serial_9_max_col_count[4], max_pool_serial_9_col_count[4] }), .Y(_05247_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _28720_ ( .A({ _07231_, cparam_max_pool_serial_9_max_col_count[3], max_pool_serial_9_col_count[3], _07229_ }), .Y(_07228_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _28721_ ( .A({ cparam_max_pool_serial_9_max_col_count[2], max_pool_serial_9_col_count[2], _07230_ }), .Y(_07229_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28722_ ( .A({ cparam_max_pool_serial_9_max_col_count[0], cparam_max_pool_serial_9_max_col_count[1], max_pool_serial_9_col_count[0], max_pool_serial_9_col_count[1] }), .Y(_07230_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28723_ ( .A({ max_pool_serial_9_col_count[4], cparam_max_pool_serial_9_max_col_count[4] }), .Y(_07231_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28724_ ( .A({ _07240_, _07239_, _07238_, _07233_ }), .Y(_07232_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28725_ ( .A({ _07237_, _07236_, _07235_, _07234_ }), .Y(_07233_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _28726_ ( .A({ max_pool_serial_9_col_count[28], max_pool_serial_9_col_count[25], max_pool_serial_9_col_count[22] }), .Y(_07234_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28727_ ( .A({ max_pool_serial_9_col_count[19], max_pool_serial_9_col_count[17], max_pool_serial_9_col_count[15], max_pool_serial_9_col_count[12] }), .Y(_07235_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28728_ ( .A({ max_pool_serial_9_col_count[29], max_pool_serial_9_col_count[27], max_pool_serial_9_col_count[24], max_pool_serial_9_col_count[18] }), .Y(_07236_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28729_ ( .A({ max_pool_serial_9_col_count[11], max_pool_serial_9_col_count[8], max_pool_serial_9_col_count[6:5] }), .Y(_07237_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28730_ ( .A({ max_pool_serial_9_col_count[21], max_pool_serial_9_col_count[16], max_pool_serial_9_col_count[14:13] }), .Y(_07238_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28731_ ( .A({ max_pool_serial_9_col_count[30], max_pool_serial_9_col_count[26], max_pool_serial_9_col_count[23], max_pool_serial_9_col_count[20] }), .Y(_07239_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28732_ ( .A({ max_pool_serial_9_col_count[10:9], max_pool_serial_9_col_count[7], max_pool_serial_9_col_count[31] }), .Y(_07240_) );
  \$lut  #( .LUT(16'h8eff), .WIDTH(4) ) _28733_ ( .A({ _07244_, cparam_max_pool_serial_9_max_col_count[4], max_pool_serial_9_row_count[4], _07241_ }), .Y(_05246_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _28734_ ( .A({ max_pool_serial_9_row_count[3], cparam_max_pool_serial_9_max_col_count[3], _07242_ }), .Y(_07241_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _28735_ ( .A({ max_pool_serial_9_row_count[2], cparam_max_pool_serial_9_max_col_count[2], _07243_ }), .Y(_07242_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _28736_ ( .A({ cparam_max_pool_serial_9_max_col_count[0], cparam_max_pool_serial_9_max_col_count[1], max_pool_serial_9_row_count[0], max_pool_serial_9_row_count[1] }), .Y(_07243_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28737_ ( .A({ _07252_, _07251_, _07250_, _07245_ }), .Y(_07244_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28738_ ( .A({ _07249_, _07248_, _07247_, _07246_ }), .Y(_07245_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28739_ ( .A({ max_pool_serial_9_row_count[15:14], max_pool_serial_9_row_count[12:11] }), .Y(_07246_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28740_ ( .A({ max_pool_serial_9_row_count[10], max_pool_serial_9_row_count[8:6] }), .Y(_07247_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28741_ ( .A({ max_pool_serial_9_row_count[29:28], max_pool_serial_9_row_count[26], max_pool_serial_9_row_count[24] }), .Y(_07248_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28742_ ( .A({ max_pool_serial_9_row_count[22], max_pool_serial_9_row_count[20], max_pool_serial_9_row_count[18], max_pool_serial_9_row_count[16] }), .Y(_07249_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _28743_ ( .A({ max_pool_serial_9_row_count[27], max_pool_serial_9_row_count[25], max_pool_serial_9_row_count[23] }), .Y(_07250_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28744_ ( .A({ max_pool_serial_9_row_count[21], max_pool_serial_9_row_count[19], max_pool_serial_9_row_count[17], max_pool_serial_9_row_count[13] }), .Y(_07251_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28745_ ( .A({ max_pool_serial_9_row_count[9], max_pool_serial_9_row_count[5], max_pool_serial_9_row_count[31:30] }), .Y(_07252_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _28746_ ( .A({ _07274_, _07298_, _07300_, _07253_ }), .Y(_05245_) );
  \$lut  #( .LUT(16'hef00), .WIDTH(4) ) _28747_ ( .A({ _07270_, _07273_, _07254_, _07268_ }), .Y(_07253_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _28748_ ( .A({ _07263_, _07267_, _07255_, _07266_ }), .Y(_07254_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _28749_ ( .A({ _07256_, _04311_, max_pool_serial_9_comp_count[5] }), .Y(_07255_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _28750_ ( .A({ _07262_, _07261_, _07257_, _07260_ }), .Y(_07256_) );
  \$lut  #( .LUT(16'hddd4), .WIDTH(4) ) _28751_ ( .A({ _07259_, _07258_, max_pool_serial_9_comp_count[2], _04306_ }), .Y(_07257_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _28752_ ( .A({ _04284_, max_pool_serial_9_comp_count[0], _04295_, max_pool_serial_9_comp_count[1] }), .Y(_07258_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28753_ ( .A({ max_pool_serial_9_comp_count[1], _04295_ }), .Y(_07259_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28754_ ( .A({ _04309_, max_pool_serial_9_comp_count[3] }), .Y(_07260_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _28755_ ( .A({ max_pool_serial_9_comp_count[3], _04309_, max_pool_serial_9_comp_count[4], _04310_ }), .Y(_07261_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _28756_ ( .A({ _04310_, max_pool_serial_9_comp_count[4], _04311_, max_pool_serial_9_comp_count[5] }), .Y(_07262_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _28757_ ( .A({ _07265_, _07264_, _04313_, max_pool_serial_9_comp_count[7] }), .Y(_07263_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28758_ ( .A({ max_pool_serial_9_comp_count[11], _04286_, max_pool_serial_9_comp_count[10], _04285_ }), .Y(_07264_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28759_ ( .A({ max_pool_serial_9_comp_count[9], _04315_, max_pool_serial_9_comp_count[8], _04314_ }), .Y(_07265_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28760_ ( .A({ _04312_, max_pool_serial_9_comp_count[6] }), .Y(_07266_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _28761_ ( .A({ max_pool_serial_9_comp_count[6], _04312_, max_pool_serial_9_comp_count[7], _04313_ }), .Y(_07267_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28762_ ( .A({ _07269_, _07264_ }), .Y(_07268_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28763_ ( .A({ max_pool_serial_9_comp_count[8], max_pool_serial_9_comp_count[9], _04314_, _04315_ }), .Y(_07269_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28764_ ( .A({ _07272_, _07271_ }), .Y(_07270_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28765_ ( .A({ max_pool_serial_9_comp_count[15], _04290_, max_pool_serial_9_comp_count[14], _04289_ }), .Y(_07271_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28766_ ( .A({ max_pool_serial_9_comp_count[13], _04288_, max_pool_serial_9_comp_count[12], _04287_ }), .Y(_07272_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _28767_ ( .A({ max_pool_serial_9_comp_count[10], max_pool_serial_9_comp_count[11], _04285_, _04286_ }), .Y(_07273_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _28768_ ( .A({ _07296_, _07286_, _07275_, _07294_ }), .Y(_07274_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _28769_ ( .A({ _07276_, _07278_, _07280_ }), .Y(_07275_) );
  \$lut  #( .LUT(16'h001f), .WIDTH(4) ) _28770_ ( .A({ _07285_, _07277_, _07284_, _07281_ }), .Y(_07276_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _28771_ ( .A({ _07280_, _07278_, _04296_, max_pool_serial_9_comp_count[20] }), .Y(_07277_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _28772_ ( .A({ _07279_, _04297_, max_pool_serial_9_comp_count[21] }), .Y(_07278_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28773_ ( .A({ max_pool_serial_9_comp_count[23], _04299_, max_pool_serial_9_comp_count[22], _04298_ }), .Y(_07279_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _28774_ ( .A({ max_pool_serial_9_comp_count[20], _04296_, max_pool_serial_9_comp_count[21], _04297_ }), .Y(_07280_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _28775_ ( .A({ _07282_, max_pool_serial_9_comp_count[17], _04292_, _07283_ }), .Y(_07281_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28776_ ( .A({ max_pool_serial_9_comp_count[19], _04294_, max_pool_serial_9_comp_count[18], _04293_ }), .Y(_07282_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28777_ ( .A({ max_pool_serial_9_comp_count[16], _04291_ }), .Y(_07283_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28778_ ( .A({ max_pool_serial_9_comp_count[18], max_pool_serial_9_comp_count[19], _04293_, _04294_ }), .Y(_07284_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28779_ ( .A({ max_pool_serial_9_comp_count[22], max_pool_serial_9_comp_count[23], _04298_, _04299_ }), .Y(_07285_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _28780_ ( .A({ _07287_, _07291_, _07293_, _07292_ }), .Y(_07286_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _28781_ ( .A({ _07290_, _07288_, _04304_, max_pool_serial_9_comp_count[28] }), .Y(_07287_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _28782_ ( .A({ _07289_, _04305_, max_pool_serial_9_comp_count[29] }), .Y(_07288_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28783_ ( .A({ max_pool_serial_9_comp_count[31], _04308_, max_pool_serial_9_comp_count[30], _04307_ }), .Y(_07289_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _28784_ ( .A({ max_pool_serial_9_comp_count[28], _04304_, max_pool_serial_9_comp_count[29], _04305_ }), .Y(_07290_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28785_ ( .A({ max_pool_serial_9_comp_count[26], max_pool_serial_9_comp_count[27], _04302_, _04303_ }), .Y(_07291_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28786_ ( .A({ max_pool_serial_9_comp_count[27], _04303_, max_pool_serial_9_comp_count[26], _04302_ }), .Y(_07292_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28787_ ( .A({ max_pool_serial_9_comp_count[24], max_pool_serial_9_comp_count[25], _04300_, _04301_ }), .Y(_07293_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28788_ ( .A({ _07295_, _07292_, _07287_ }), .Y(_07294_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28789_ ( .A({ max_pool_serial_9_comp_count[25], _04301_, max_pool_serial_9_comp_count[24], _04300_ }), .Y(_07295_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _28790_ ( .A({ _07297_, _07288_, _07290_ }), .Y(_07296_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28791_ ( .A({ max_pool_serial_9_comp_count[30], max_pool_serial_9_comp_count[31], _04307_, _04308_ }), .Y(_07297_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28792_ ( .A({ _07299_, _07282_, _07277_, _07294_ }), .Y(_07298_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _28793_ ( .A({ max_pool_serial_9_comp_count[17], _04292_, max_pool_serial_9_comp_count[16], _04291_ }), .Y(_07299_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _28794_ ( .A({ _07301_, _07271_, _07302_ }), .Y(_07300_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28795_ ( .A({ max_pool_serial_9_comp_count[14], max_pool_serial_9_comp_count[15], _04289_, _04290_ }), .Y(_07301_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _28796_ ( .A({ max_pool_serial_9_comp_count[12], max_pool_serial_9_comp_count[13], _04287_, _04288_ }), .Y(_07302_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _28797_ ( .A({ _07308_, _07303_ }), .Y(_05244_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28798_ ( .A({ _07307_, _07306_, _07305_, _07304_ }), .Y(_07303_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28799_ ( .A({ _04262_, _04261_, _04260_, _04259_ }), .Y(_07304_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28800_ ( .A({ _04258_, _04257_, _04256_, _04255_ }), .Y(_07305_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28801_ ( .A({ _04276_, _04275_, _04273_, _04272_ }), .Y(_07306_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28802_ ( .A({ _04270_, _04269_, _04267_, _04264_ }), .Y(_07307_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28803_ ( .A({ _04271_, _04268_, _04266_, _04265_ }), .Y(_07308_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _28804_ ( .A({ _07309_, _07318_, _07315_, _maxi_write_rest_size[8] }), .Y(_05263_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28805_ ( .A({ _07314_, _07310_ }), .Y(_07309_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _28806_ ( .A({ _07313_, _07311_, _maxi_write_rest_size[20:19] }), .Y(_07310_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _28807_ ( .A({ _07312_, _maxi_write_rest_size[32:30] }), .Y(_07311_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28808_ ( .A({ _maxi_write_rest_size[28:27], _maxi_write_rest_size[25], _maxi_write_rest_size[22] }), .Y(_07312_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28809_ ( .A({ _maxi_write_rest_size[21], _maxi_write_rest_size[18:16] }), .Y(_07313_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28810_ ( .A({ _maxi_write_rest_size[29], _maxi_write_rest_size[26], _maxi_write_rest_size[24:23] }), .Y(_07314_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28811_ ( .A({ _07317_, _07316_ }), .Y(_07315_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28812_ ( .A(_maxi_write_rest_size[7:4]), .Y(_07316_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28813_ ( .A(_maxi_write_rest_size[3:0]), .Y(_07317_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _28814_ ( .A({ _07319_, _maxi_write_rest_size[14], _maxi_write_rest_size[11:10] }), .Y(_07318_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28815_ ( .A({ _maxi_write_rest_size[15], _maxi_write_rest_size[13:12], _maxi_write_rest_size[9] }), .Y(_07319_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28816_ ( .A({ _07320_, _17387_, _07122_ }), .Y(_17419_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28817_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17451_, _17483_ }), .Y(_07320_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28818_ ( .A({ _07321_, _17386_, _07122_ }), .Y(_17418_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28819_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17450_, _17482_ }), .Y(_07321_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28820_ ( .A({ _18414_, _07019_, _18350_, maxi_rready }), .Y(_18382_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28821_ ( .A({ _maxi_read_fsm[1:0], _07017_, _07008_ }), .Y(maxi_rready) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28822_ ( .A({ _07322_, _17385_, _07122_ }), .Y(_17417_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28823_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17449_, _17481_ }), .Y(_07322_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28824_ ( .A({ _18413_, _07019_, _18349_, maxi_rready }), .Y(_18381_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28825_ ( .A({ _07323_, _17384_, _07122_ }), .Y(_17416_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28826_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17448_, _17480_ }), .Y(_07323_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28827_ ( .A({ _18411_, _07019_, _18347_, maxi_rready }), .Y(_18379_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28828_ ( .A({ _07324_, _17383_, _07122_ }), .Y(_17415_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28829_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17447_, _17479_ }), .Y(_07324_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28830_ ( .A({ _18410_, _07019_, _18346_, maxi_rready }), .Y(_18378_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28831_ ( .A({ _07325_, _17382_, _07122_ }), .Y(_17414_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28832_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17446_, _17478_ }), .Y(_07325_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _28833_ ( .A({ _07326_, _17381_, _07122_ }), .Y(_17413_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _28834_ ( .A({ _07111_, conv2d_8_comp_fsm[2], _17445_, _17477_ }), .Y(_07326_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28835_ ( .A({ _18409_, _07019_, _18345_, maxi_rready }), .Y(_18377_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28836_ ( .A({ _18408_, _07019_, _18344_, maxi_rready }), .Y(_18376_) );
  \$lut  #( .LUT(16'h8fff), .WIDTH(4) ) _28837_ ( .A({ _07327_, _07329_, _07328_, _17442_ }), .Y(_17410_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _28838_ ( .A({ _17474_, _04899_, _17378_, _07122_ }), .Y(_07327_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28839_ ( .A({ _07111_, conv2d_8_comp_fsm[2] }), .Y(_04899_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _28840_ ( .A({ conv2d_8_comp_fsm[2], _07111_ }), .Y(_07328_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28841_ ( .A({ _05101_, _07330_ }), .Y(_07329_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28842_ ( .A({ _07144_, _07124_, conv2d_8_comp_fsm[1] }), .Y(_07330_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _28843_ ( .A({ conv2d_8_comp_fsm[1], _07145_, _07144_ }), .Y(_05101_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28844_ ( .A({ _18406_, _07019_, _18342_, maxi_rready }), .Y(_18374_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28845_ ( .A({ _18407_, _07019_, _18343_, maxi_rready }), .Y(_18375_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _28846_ ( .A({ _05100_, _05102_, _07332_, _07331_ }), .Y(_17399_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _28847_ ( .A({ _07330_, _07328_, _17431_ }), .Y(_07331_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _28848_ ( .A({ _17463_, _04899_, _17367_, _07122_ }), .Y(_07332_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _28849_ ( .A({ _07145_, _07123_ }), .Y(_05100_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28850_ ( .A({ _18405_, _07019_, _18341_, maxi_rready }), .Y(_18373_) );
  \$lut  #( .LUT(16'h8fff), .WIDTH(4) ) _28851_ ( .A({ _07333_, _05100_, _07328_, _17420_ }), .Y(_17388_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _28852_ ( .A({ _17452_, _04899_, _17356_, _07122_ }), .Y(_07333_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28853_ ( .A({ _18404_, _07019_, _18340_, maxi_rready }), .Y(_18372_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28854_ ( .A({ _18403_, _07019_, _18339_, maxi_rready }), .Y(_18371_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28855_ ( .A({ _18402_, _07019_, _18338_, maxi_rready }), .Y(_18370_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28856_ ( .A({ _18400_, _07019_, _18336_, maxi_rready }), .Y(_18368_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28857_ ( .A({ _18399_, _07019_, _18335_, maxi_rready }), .Y(_18367_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28858_ ( .A({ _18398_, _07019_, _18334_, maxi_rready }), .Y(_18366_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28859_ ( .A({ _18397_, _07019_, _18333_, maxi_rready }), .Y(_18365_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28860_ ( .A({ _15989_, _07334_, _15957_, _05071_ }), .Y(_15925_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _28861_ ( .A({ _07067_, _stream_conv2d_8_source_31_source_pat_fsm_14[1] }), .Y(_07334_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28862_ ( .A({ _16000_, _07334_, _15968_, _05071_ }), .Y(_15936_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28863_ ( .A({ _16010_, _07334_, _15978_, _05071_ }), .Y(_15946_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28864_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16161_, _16193_ }), .Y(_16129_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28865_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16346_, _16378_ }), .Y(_16314_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28866_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16525_, _16557_ }), .Y(_16493_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28867_ ( .A({ _18396_, _07019_, _18332_, maxi_rready }), .Y(_18364_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28868_ ( .A({ _15999_, _07334_, _15967_, _05071_ }), .Y(_15935_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28869_ ( .A({ _15988_, _07334_, _15956_, _05071_ }), .Y(_15924_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28870_ ( .A({ _16009_, _07334_, _15977_, _05071_ }), .Y(_15945_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28871_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16160_, _16192_ }), .Y(_16128_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28872_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16345_, _16377_ }), .Y(_16313_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28873_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16555_, _16587_ }), .Y(_16523_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28874_ ( .A({ _18395_, _07019_, _18331_, maxi_rready }), .Y(_18363_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28875_ ( .A({ _16008_, _07334_, _15976_, _05071_ }), .Y(_15944_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28876_ ( .A({ _15998_, _07334_, _15966_, _05071_ }), .Y(_15934_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28877_ ( .A({ _15987_, _07334_, _15955_, _05071_ }), .Y(_15923_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28878_ ( .A({ _05072_, _07032_ }), .Y(_21907_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _28879_ ( .A({ _stream_conv2d_8_source_30_source_pat_fsm_13[1], _07033_, _07041_, _stream_conv2d_8_source_30_source_pat_fsm_13[0] }), .Y(_05072_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28880_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16068_, _16100_ }), .Y(_16036_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28881_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16159_, _16191_ }), .Y(_16127_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28882_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16344_, _16376_ }), .Y(_16312_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28883_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16554_, _16586_ }), .Y(_16522_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28884_ ( .A({ _18394_, _07019_, _18330_, maxi_rready }), .Y(_18362_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28885_ ( .A({ _15986_, _07334_, _15954_, _05071_ }), .Y(_15922_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28886_ ( .A({ _15997_, _07334_, _15965_, _05071_ }), .Y(_15933_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _28887_ ( .A({ _16007_, _07334_, _15975_, _05071_ }), .Y(_15943_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28888_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16067_, _16099_ }), .Y(_16035_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28889_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16158_, _16190_ }), .Y(_16126_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28890_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16342_, _16374_ }), .Y(_16310_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28891_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16553_, _16585_ }), .Y(_16521_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28892_ ( .A({ _18393_, _07019_, _18329_, maxi_rready }), .Y(_18361_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28893_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16065_, _16097_ }), .Y(_16033_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28894_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16157_, _16189_ }), .Y(_16125_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28895_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16341_, _16373_ }), .Y(_16309_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28896_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16552_, _16584_ }), .Y(_16520_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28897_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17028_, _17060_ }), .Y(_16996_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28898_ ( .A({ _07336_, _07344_, _stream_conv2d_8_source_20_source_pat_fsm_3[1] }), .Y(_07335_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28899_ ( .A({ _07343_, _07342_, _07337_ }), .Y(_07336_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28900_ ( .A({ _07341_, _07340_, _07339_, _07338_ }), .Y(_07337_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28901_ ( .A(_stream_conv2d_8_source_20_source_pat_fsm_3[23:20]), .Y(_07338_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28902_ ( .A(_stream_conv2d_8_source_20_source_pat_fsm_3[19:16]), .Y(_07339_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28903_ ( .A(_stream_conv2d_8_source_20_source_pat_fsm_3[31:28]), .Y(_07340_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28904_ ( .A(_stream_conv2d_8_source_20_source_pat_fsm_3[27:24]), .Y(_07341_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28905_ ( .A(_stream_conv2d_8_source_20_source_pat_fsm_3[15:12]), .Y(_07342_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28906_ ( .A(_stream_conv2d_8_source_20_source_pat_fsm_3[11:8]), .Y(_07343_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28907_ ( .A({ _07345_, _stream_conv2d_8_source_20_source_pat_fsm_3[3:2] }), .Y(_07344_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28908_ ( .A(_stream_conv2d_8_source_20_source_pat_fsm_3[7:4]), .Y(_07345_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28909_ ( .A({ _18392_, _07019_, _18328_, maxi_rready }), .Y(_18360_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28910_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16064_, _16096_ }), .Y(_16032_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28911_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16156_, _16188_ }), .Y(_16124_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28912_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16340_, _16372_ }), .Y(_16308_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28913_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16551_, _16583_ }), .Y(_16519_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28914_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17027_, _17059_ }), .Y(_16995_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28915_ ( .A({ _18391_, _07019_, _18327_, maxi_rready }), .Y(_18359_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28916_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16063_, _16095_ }), .Y(_16031_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28917_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16155_, _16187_ }), .Y(_16123_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28918_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16339_, _16371_ }), .Y(_16307_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28919_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16550_, _16582_ }), .Y(_16518_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28920_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17025_, _17057_ }), .Y(_16993_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _28921_ ( .A({ _05100_, _05102_, _07346_ }), .Y(_21921_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28922_ ( .A({ _07329_, _07111_, _07122_ }), .Y(_07346_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28923_ ( .A({ _18421_, _07019_, _18357_, maxi_rready }), .Y(_18389_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28924_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16154_, _16186_ }), .Y(_16122_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28925_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16338_, _16370_ }), .Y(_16306_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28926_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16549_, _16581_ }), .Y(_16517_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28927_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17024_, _17056_ }), .Y(_16992_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28928_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16153_, _16185_ }), .Y(_16121_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28929_ ( .A({ _18420_, _07019_, _18356_, maxi_rready }), .Y(_18388_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28930_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16337_, _16369_ }), .Y(_16305_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28931_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16546_, _16578_ }), .Y(_16514_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28932_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17023_, _17055_ }), .Y(_16991_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28933_ ( .A({ _18419_, _07019_, _18355_, maxi_rready }), .Y(_18387_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28934_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16152_, _16184_ }), .Y(_16120_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28935_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16336_, _16368_ }), .Y(_16304_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28936_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16535_, _16567_ }), .Y(_16503_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28937_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17022_, _17054_ }), .Y(_16990_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28938_ ( .A({ _18418_, _07019_, _18354_, maxi_rready }), .Y(_18386_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28939_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16150_, _16182_ }), .Y(_16118_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28940_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16335_, _16367_ }), .Y(_16303_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28941_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16524_, _16556_ }), .Y(_16492_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28942_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17021_, _17053_ }), .Y(_16989_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28943_ ( .A({ _18417_, _07019_, _18353_, maxi_rready }), .Y(_18385_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28944_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16334_, _16366_ }), .Y(_16302_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28945_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17020_, _17052_ }), .Y(_16988_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28946_ ( .A({ _18416_, _07019_, _18352_, maxi_rready }), .Y(_18384_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28947_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16333_, _16365_ }), .Y(_16301_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28948_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17019_, _17051_ }), .Y(_16987_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28949_ ( .A({ _18415_, _07019_, _18351_, maxi_rready }), .Y(_18383_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28950_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16363_, _16395_ }), .Y(_16331_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28951_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17018_, _17050_ }), .Y(_16986_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28952_ ( .A({ _18412_, _07019_, _18348_, maxi_rready }), .Y(_18380_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28953_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16362_, _16394_ }), .Y(_16330_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28954_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17017_, _17049_ }), .Y(_16985_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28955_ ( .A({ _18401_, _07019_, _18337_, maxi_rready }), .Y(_18369_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28956_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16361_, _16393_ }), .Y(_16329_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28957_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17016_, _17048_ }), .Y(_16984_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _28958_ ( .A({ _18390_, _07019_, _18326_, maxi_rready }), .Y(_18358_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28959_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16360_, _16392_ }), .Y(_16328_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28960_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17014_, _17046_ }), .Y(_16982_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28961_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16359_, _16391_ }), .Y(_16327_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28962_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17013_, _17045_ }), .Y(_16981_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28963_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16358_, _16390_ }), .Y(_16326_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28964_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17012_, _17044_ }), .Y(_16980_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28965_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16357_, _16389_ }), .Y(_16325_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28966_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17011_, _17043_ }), .Y(_16979_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _28967_ ( .A({ maxi_rready, _07019_ }), .Y(_21923_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28968_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17009_, _17041_ }), .Y(_16977_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28969_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17007_, _17039_ }), .Y(_16975_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28970_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17006_, _17038_ }), .Y(_16974_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28971_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17005_, _17037_ }), .Y(_16973_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28972_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17035_, _17067_ }), .Y(_17003_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28973_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17034_, _17066_ }), .Y(_17002_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28974_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17033_, _17065_ }), .Y(_17001_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28975_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17032_, _17064_ }), .Y(_17000_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28976_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17031_, _17063_ }), .Y(_16999_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28977_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17030_, _17062_ }), .Y(_16998_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28978_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17029_, _17061_ }), .Y(_16997_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28979_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17026_, _17058_ }), .Y(_16994_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28980_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17004_, _17036_ }), .Y(_16972_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28981_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16932_, _16964_ }), .Y(_16900_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _28982_ ( .A({ _07348_, _07356_, _stream_conv2d_8_source_21_source_pat_fsm_4[1] }), .Y(_07347_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _28983_ ( .A({ _07355_, _07354_, _07349_ }), .Y(_07348_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _28984_ ( .A({ _07353_, _07352_, _07351_, _07350_ }), .Y(_07349_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28985_ ( .A(_stream_conv2d_8_source_21_source_pat_fsm_4[23:20]), .Y(_07350_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28986_ ( .A(_stream_conv2d_8_source_21_source_pat_fsm_4[19:16]), .Y(_07351_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28987_ ( .A(_stream_conv2d_8_source_21_source_pat_fsm_4[31:28]), .Y(_07352_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28988_ ( .A(_stream_conv2d_8_source_21_source_pat_fsm_4[27:24]), .Y(_07353_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28989_ ( .A(_stream_conv2d_8_source_21_source_pat_fsm_4[15:12]), .Y(_07354_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28990_ ( .A(_stream_conv2d_8_source_21_source_pat_fsm_4[11:8]), .Y(_07355_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _28991_ ( .A({ _07357_, _stream_conv2d_8_source_21_source_pat_fsm_4[3:2] }), .Y(_07356_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _28992_ ( .A(_stream_conv2d_8_source_21_source_pat_fsm_4[7:4]), .Y(_07357_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28993_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16931_, _16963_ }), .Y(_16899_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28994_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16929_, _16961_ }), .Y(_16897_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _28995_ ( .A({ _05092_, _07335_ }), .Y(_21917_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _28996_ ( .A({ _stream_conv2d_8_source_20_source_pat_fsm_3[1], _07336_, _07344_, _stream_conv2d_8_source_20_source_pat_fsm_3[0] }), .Y(_05092_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28997_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16928_, _16960_ }), .Y(_16896_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28998_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16927_, _16959_ }), .Y(_16895_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _28999_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16926_, _16958_ }), .Y(_16894_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29000_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16925_, _16957_ }), .Y(_16893_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29001_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16924_, _16956_ }), .Y(_16892_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29002_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16921_, _16953_ }), .Y(_16889_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29003_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16920_, _16952_ }), .Y(_16888_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29004_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16918_, _16950_ }), .Y(_16886_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29005_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16917_, _16949_ }), .Y(_16885_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29006_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16916_, _16948_ }), .Y(_16884_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29007_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16062_, _16094_ }), .Y(_16030_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29008_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16149_, _16181_ }), .Y(_16117_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29009_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16354_, _16386_ }), .Y(_16322_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29010_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16915_, _16947_ }), .Y(_16883_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29011_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16061_, _16093_ }), .Y(_16029_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29012_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16148_, _16180_ }), .Y(_16116_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29013_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16343_, _16375_ }), .Y(_16311_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29014_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16644_, _16676_ }), .Y(_16612_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29015_ ( .A({ _07359_, _07367_, _stream_conv2d_8_source_24_source_pat_fsm_7[1] }), .Y(_07358_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29016_ ( .A({ _07366_, _07365_, _07360_ }), .Y(_07359_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29017_ ( .A({ _07364_, _07363_, _07362_, _07361_ }), .Y(_07360_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29018_ ( .A(_stream_conv2d_8_source_24_source_pat_fsm_7[23:20]), .Y(_07361_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29019_ ( .A(_stream_conv2d_8_source_24_source_pat_fsm_7[19:16]), .Y(_07362_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29020_ ( .A(_stream_conv2d_8_source_24_source_pat_fsm_7[31:28]), .Y(_07363_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29021_ ( .A(_stream_conv2d_8_source_24_source_pat_fsm_7[27:24]), .Y(_07364_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29022_ ( .A(_stream_conv2d_8_source_24_source_pat_fsm_7[15:12]), .Y(_07365_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29023_ ( .A(_stream_conv2d_8_source_24_source_pat_fsm_7[11:8]), .Y(_07366_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29024_ ( .A({ _07368_, _stream_conv2d_8_source_24_source_pat_fsm_7[3:2] }), .Y(_07367_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29025_ ( .A(_stream_conv2d_8_source_24_source_pat_fsm_7[7:4]), .Y(_07368_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29026_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16914_, _16946_ }), .Y(_16882_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29027_ ( .A({ _17573_, _07122_, _17637_, _05102_ }), .Y(_17605_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29028_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16060_, _16092_ }), .Y(_16028_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29029_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16147_, _16179_ }), .Y(_16115_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29030_ ( .A({ _07127_, _stream_conv2d_8_source_27_source_pat_fsm_10[0], _16332_, _16364_ }), .Y(_16300_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29031_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16641_, _16673_ }), .Y(_16609_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29032_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16913_, _16945_ }), .Y(_16881_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29033_ ( .A({ _17572_, _07122_, _17636_, _05102_ }), .Y(_17604_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29034_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16146_, _16178_ }), .Y(_16114_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29035_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16640_, _16672_ }), .Y(_16608_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29036_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16912_, _16944_ }), .Y(_16880_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29037_ ( .A({ _17570_, _07122_, _17634_, _05102_ }), .Y(_17602_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29038_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16145_, _16177_ }), .Y(_16113_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29039_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16639_, _16671_ }), .Y(_16607_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29040_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16911_, _16943_ }), .Y(_16879_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29041_ ( .A({ _17569_, _07122_, _17633_, _05102_ }), .Y(_17601_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29042_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16144_, _16176_ }), .Y(_16112_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29043_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16638_, _16670_ }), .Y(_16606_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29044_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16909_, _16941_ }), .Y(_16877_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29045_ ( .A({ _17568_, _07122_, _17632_, _05102_ }), .Y(_17600_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29046_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16143_, _16175_ }), .Y(_16111_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29047_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16637_, _16669_ }), .Y(_16605_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29048_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16939_, _16971_ }), .Y(_16907_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29049_ ( .A({ _17567_, _07122_, _17631_, _05102_ }), .Y(_17599_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29050_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16142_, _16174_ }), .Y(_16110_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29051_ ( .A({ _05078_, _07127_ }), .Y(_21910_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29052_ ( .A({ _stream_conv2d_8_source_27_source_pat_fsm_10[1], _07128_, _07136_, _stream_conv2d_8_source_27_source_pat_fsm_10[0] }), .Y(_05078_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29053_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16636_, _16668_ }), .Y(_16604_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29054_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16938_, _16970_ }), .Y(_16906_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29055_ ( .A({ _17566_, _07122_, _17630_, _05102_ }), .Y(_17598_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29056_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16141_, _16173_ }), .Y(_16109_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29057_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16635_, _16667_ }), .Y(_16603_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29058_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16937_, _16969_ }), .Y(_16905_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29059_ ( .A({ _17565_, _07122_, _17629_, _05102_ }), .Y(_17597_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29060_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16171_, _16203_ }), .Y(_16139_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29061_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16634_, _16666_ }), .Y(_16602_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29062_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16936_, _16968_ }), .Y(_16904_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29063_ ( .A({ _17564_, _07122_, _17628_, _05102_ }), .Y(_17596_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29064_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16170_, _16202_ }), .Y(_16138_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29065_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16633_, _16665_ }), .Y(_16601_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29066_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16935_, _16967_ }), .Y(_16903_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29067_ ( .A({ _17563_, _07122_, _17627_, _05102_ }), .Y(_17595_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29068_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16169_, _16201_ }), .Y(_16137_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29069_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16632_, _16664_ }), .Y(_16600_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29070_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16934_, _16966_ }), .Y(_16902_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29071_ ( .A({ _17562_, _07122_, _17626_, _05102_ }), .Y(_17594_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29072_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16168_, _16200_ }), .Y(_16136_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29073_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16630_, _16662_ }), .Y(_16598_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29074_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16933_, _16965_ }), .Y(_16901_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29075_ ( .A({ _17561_, _07122_, _17625_, _05102_ }), .Y(_17593_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29076_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16167_, _16199_ }), .Y(_16135_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29077_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16629_, _16661_ }), .Y(_16597_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29078_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16930_, _16962_ }), .Y(_16898_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29079_ ( .A({ _17559_, _07122_, _17623_, _05102_ }), .Y(_17591_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29080_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16166_, _16198_ }), .Y(_16134_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29081_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16627_, _16659_ }), .Y(_16595_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29082_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16919_, _16951_ }), .Y(_16887_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29083_ ( .A({ _17558_, _07122_, _17622_, _05102_ }), .Y(_17590_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29084_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16626_, _16658_ }), .Y(_16594_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29085_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16836_, _16868_ }), .Y(_16804_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29086_ ( .A({ _07370_, _07378_, _stream_conv2d_8_source_22_source_pat_fsm_5[1] }), .Y(_07369_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29087_ ( .A({ _07377_, _07376_, _07371_ }), .Y(_07370_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29088_ ( .A({ _07375_, _07374_, _07373_, _07372_ }), .Y(_07371_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29089_ ( .A(_stream_conv2d_8_source_22_source_pat_fsm_5[23:20]), .Y(_07372_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29090_ ( .A(_stream_conv2d_8_source_22_source_pat_fsm_5[19:16]), .Y(_07373_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29091_ ( .A(_stream_conv2d_8_source_22_source_pat_fsm_5[31:28]), .Y(_07374_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29092_ ( .A(_stream_conv2d_8_source_22_source_pat_fsm_5[27:24]), .Y(_07375_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29093_ ( .A(_stream_conv2d_8_source_22_source_pat_fsm_5[15:12]), .Y(_07376_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29094_ ( .A(_stream_conv2d_8_source_22_source_pat_fsm_5[11:8]), .Y(_07377_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29095_ ( .A({ _07379_, _stream_conv2d_8_source_22_source_pat_fsm_5[3:2] }), .Y(_07378_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29096_ ( .A(_stream_conv2d_8_source_22_source_pat_fsm_5[7:4]), .Y(_07379_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29097_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16908_, _16940_ }), .Y(_16876_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29098_ ( .A({ _17557_, _07122_, _17621_, _05102_ }), .Y(_17589_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29099_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16625_, _16657_ }), .Y(_16593_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29100_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16833_, _16865_ }), .Y(_16801_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29101_ ( .A({ _17556_, _07122_, _17620_, _05102_ }), .Y(_17588_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29102_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16624_, _16656_ }), .Y(_16592_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29103_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16832_, _16864_ }), .Y(_16800_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29104_ ( .A({ _17555_, _07122_, _17619_, _05102_ }), .Y(_17587_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29105_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16623_, _16655_ }), .Y(_16591_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29106_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16831_, _16863_ }), .Y(_16799_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29107_ ( .A({ _17554_, _07122_, _17618_, _05102_ }), .Y(_17586_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29108_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16622_, _16654_ }), .Y(_16590_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29109_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16830_, _16862_ }), .Y(_16798_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29110_ ( .A({ _05090_, _07347_ }), .Y(_21916_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29111_ ( .A({ _stream_conv2d_8_source_21_source_pat_fsm_4[1], _07348_, _07356_, _stream_conv2d_8_source_21_source_pat_fsm_4[0] }), .Y(_05090_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29112_ ( .A({ _17553_, _07122_, _17617_, _05102_ }), .Y(_17585_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29113_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16621_, _16653_ }), .Y(_16589_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29114_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16829_, _16861_ }), .Y(_16797_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29115_ ( .A({ _17552_, _07122_, _17616_, _05102_ }), .Y(_17584_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29116_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16651_, _16683_ }), .Y(_16619_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29117_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16828_, _16860_ }), .Y(_16796_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29118_ ( .A({ _17551_, _07122_, _17615_, _05102_ }), .Y(_17583_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29119_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16650_, _16682_ }), .Y(_16618_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29120_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16827_, _16859_ }), .Y(_16795_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29121_ ( .A({ _17550_, _07122_, _17614_, _05102_ }), .Y(_17582_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29122_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16649_, _16681_ }), .Y(_16617_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29123_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16826_, _16858_ }), .Y(_16794_) );
  \$lut  #( .LUT(16'h4dff), .WIDTH(4) ) _29124_ ( .A({ _07383_, cparam_conv2d_8_max_col_count[4], conv2d_8_col_count[4], _07380_ }), .Y(_05242_) );
  \$lut  #( .LUT(8'h71), .WIDTH(3) ) _29125_ ( .A({ cparam_conv2d_8_max_col_count[3], conv2d_8_col_count[3], _07381_ }), .Y(_07380_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _29126_ ( .A({ conv2d_8_col_count[2], cparam_conv2d_8_max_col_count[2], _07382_ }), .Y(_07381_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _29127_ ( .A({ cparam_conv2d_8_max_col_count[0], cparam_conv2d_8_max_col_count[1], conv2d_8_col_count[0], conv2d_8_col_count[1] }), .Y(_07382_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29128_ ( .A({ _07391_, _07390_, _07389_, _07384_ }), .Y(_07383_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29129_ ( .A({ _07388_, _07387_, _07386_, _07385_ }), .Y(_07384_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29130_ ( .A({ conv2d_8_col_count[20], conv2d_8_col_count[17:16], conv2d_8_col_count[13] }), .Y(_07385_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29131_ ( .A(conv2d_8_col_count[10:7]), .Y(_07386_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29132_ ( .A({ conv2d_8_col_count[5], conv2d_8_col_count[31:29] }), .Y(_07387_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29133_ ( .A({ conv2d_8_col_count[28], conv2d_8_col_count[25:23] }), .Y(_07388_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _29134_ ( .A({ conv2d_8_col_count[27:26], conv2d_8_col_count[22] }), .Y(_07389_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29135_ ( .A({ conv2d_8_col_count[21], conv2d_8_col_count[19:18], conv2d_8_col_count[15] }), .Y(_07390_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29136_ ( .A({ conv2d_8_col_count[14], conv2d_8_col_count[12:11], conv2d_8_col_count[6] }), .Y(_07391_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29137_ ( .A({ _17580_, _07122_, _17644_, _05102_ }), .Y(_17612_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29138_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16648_, _16680_ }), .Y(_16616_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29139_ ( .A({ _07397_, _07392_ }), .Y(_05243_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29140_ ( .A({ _07396_, _07395_, _07394_, _07393_ }), .Y(_07392_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29141_ ( .A({ _04202_, _04201_, _04200_, _04199_ }), .Y(_07393_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29142_ ( .A({ _04197_, _04196_, _04195_, _04194_ }), .Y(_07394_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29143_ ( .A({ _04211_, _04210_, _04208_, _04207_ }), .Y(_07395_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29144_ ( .A({ _04206_, _04205_, _04204_, _04203_ }), .Y(_07396_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29145_ ( .A({ _07401_, _07400_, _07399_, _07398_ }), .Y(_07397_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _29146_ ( .A({ _04212_, _04209_, _04187_, _04198_ }), .Y(_07398_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29147_ ( .A({ _04216_, _04215_, _04214_, _04213_ }), .Y(_07399_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29148_ ( .A({ _04193_, _04192_, _04191_, _04190_ }), .Y(_07400_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29149_ ( .A({ _04189_, _04188_, _04218_, _04217_ }), .Y(_07401_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29150_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16825_, _16857_ }), .Y(_16793_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29151_ ( .A({ _17579_, _07122_, _17643_, _05102_ }), .Y(_17611_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29152_ ( .A({ _17991_, _07122_, _17637_, _05102_ }), .Y(_18023_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29153_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16647_, _16679_ }), .Y(_16615_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29154_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16824_, _16856_ }), .Y(_16792_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29155_ ( .A({ _17578_, _07122_, _17642_, _05102_ }), .Y(_17610_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29156_ ( .A({ _17990_, _07122_, _17636_, _05102_ }), .Y(_18022_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29157_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16646_, _16678_ }), .Y(_16614_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29158_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16822_, _16854_ }), .Y(_16790_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29159_ ( .A({ _17577_, _07122_, _17641_, _05102_ }), .Y(_17609_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29160_ ( .A({ _17988_, _07122_, _17634_, _05102_ }), .Y(_18020_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29161_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16645_, _16677_ }), .Y(_16613_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29162_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16821_, _16853_ }), .Y(_16789_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29163_ ( .A({ _17576_, _07122_, _17640_, _05102_ }), .Y(_17608_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29164_ ( .A({ _17987_, _07122_, _17633_, _05102_ }), .Y(_18019_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29165_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16642_, _16674_ }), .Y(_16610_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29166_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16820_, _16852_ }), .Y(_16788_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29167_ ( .A({ _17575_, _07122_, _17639_, _05102_ }), .Y(_17607_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29168_ ( .A({ _17986_, _07122_, _17632_, _05102_ }), .Y(_18018_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29169_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16631_, _16663_ }), .Y(_16599_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29170_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16819_, _16851_ }), .Y(_16787_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29171_ ( .A({ _17574_, _07122_, _17638_, _05102_ }), .Y(_17606_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29172_ ( .A({ _17985_, _07122_, _17631_, _05102_ }), .Y(_18017_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29173_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16620_, _16652_ }), .Y(_16588_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29174_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16818_, _16850_ }), .Y(_16786_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29175_ ( .A({ _17571_, _07122_, _17635_, _05102_ }), .Y(_17603_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29176_ ( .A({ _17984_, _07122_, _17630_, _05102_ }), .Y(_18016_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29177_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16817_, _16849_ }), .Y(_16785_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29178_ ( .A({ _17560_, _07122_, _17624_, _05102_ }), .Y(_17592_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29179_ ( .A({ _17983_, _07122_, _17629_, _05102_ }), .Y(_18015_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29180_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16816_, _16848_ }), .Y(_16784_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29181_ ( .A({ _17549_, _07122_, _17613_, _05102_ }), .Y(_17581_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29182_ ( .A({ _17982_, _07122_, _17628_, _05102_ }), .Y(_18014_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29183_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16815_, _16847_ }), .Y(_16783_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29184_ ( .A({ _17981_, _07122_, _17627_, _05102_ }), .Y(_18013_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29185_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16814_, _16846_ }), .Y(_16782_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29186_ ( .A({ _17980_, _07122_, _17626_, _05102_ }), .Y(_18012_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29187_ ( .A({ _05084_, _07358_ }), .Y(_21913_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29188_ ( .A({ _stream_conv2d_8_source_24_source_pat_fsm_7[1], _07359_, _07367_, _stream_conv2d_8_source_24_source_pat_fsm_7[0] }), .Y(_05084_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29189_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16813_, _16845_ }), .Y(_16781_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29190_ ( .A({ _17979_, _07122_, _17625_, _05102_ }), .Y(_18011_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29191_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16843_, _16875_ }), .Y(_16811_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29192_ ( .A({ _17977_, _07122_, _17623_, _05102_ }), .Y(_18009_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29193_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16842_, _16874_ }), .Y(_16810_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29194_ ( .A({ _17976_, _07122_, _17622_, _05102_ }), .Y(_18008_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29195_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16841_, _16873_ }), .Y(_16809_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29196_ ( .A({ _17975_, _07122_, _17621_, _05102_ }), .Y(_18007_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29197_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16840_, _16872_ }), .Y(_16808_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29198_ ( .A({ _17974_, _07122_, _17620_, _05102_ }), .Y(_18006_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29199_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16740_, _16772_ }), .Y(_16708_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29200_ ( .A({ _07403_, _07411_, _stream_conv2d_8_source_23_source_pat_fsm_6[1] }), .Y(_07402_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29201_ ( .A({ _07410_, _07409_, _07404_ }), .Y(_07403_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29202_ ( .A({ _07408_, _07407_, _07406_, _07405_ }), .Y(_07404_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29203_ ( .A(_stream_conv2d_8_source_23_source_pat_fsm_6[23:20]), .Y(_07405_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29204_ ( .A(_stream_conv2d_8_source_23_source_pat_fsm_6[19:16]), .Y(_07406_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29205_ ( .A(_stream_conv2d_8_source_23_source_pat_fsm_6[31:28]), .Y(_07407_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29206_ ( .A(_stream_conv2d_8_source_23_source_pat_fsm_6[27:24]), .Y(_07408_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29207_ ( .A(_stream_conv2d_8_source_23_source_pat_fsm_6[15:12]), .Y(_07409_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29208_ ( .A(_stream_conv2d_8_source_23_source_pat_fsm_6[11:8]), .Y(_07410_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29209_ ( .A({ _07412_, _stream_conv2d_8_source_23_source_pat_fsm_6[3:2] }), .Y(_07411_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29210_ ( .A(_stream_conv2d_8_source_23_source_pat_fsm_6[7:4]), .Y(_07412_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29211_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16838_, _16870_ }), .Y(_16806_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29212_ ( .A({ _17973_, _07122_, _17619_, _05102_ }), .Y(_18005_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29213_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16739_, _16771_ }), .Y(_16707_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29214_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16837_, _16869_ }), .Y(_16805_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29215_ ( .A({ _07418_, _07413_ }), .Y(_05241_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29216_ ( .A({ _07417_, _07416_, _07415_, _07414_ }), .Y(_07413_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29217_ ( .A({ _04165_, _04164_, _04163_, _04162_ }), .Y(_07414_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29218_ ( .A({ _04161_, _04160_, _04159_, _04158_ }), .Y(_07415_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29219_ ( .A({ _04179_, _04178_, _04176_, _04175_ }), .Y(_07416_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29220_ ( .A({ _04173_, _04172_, _04170_, _04167_ }), .Y(_07417_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29221_ ( .A({ _04174_, _04171_, _04169_, _04168_ }), .Y(_07418_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29222_ ( .A({ _17972_, _07122_, _17618_, _05102_ }), .Y(_18004_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29223_ ( .A({ _17971_, _07122_, _17617_, _05102_ }), .Y(_18003_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _29224_ ( .A({ _07419_, _07428_, _07425_, _maxi_read_rest_size[8] }), .Y(_05262_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29225_ ( .A({ _07424_, _07420_ }), .Y(_07419_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _29226_ ( .A({ _07423_, _07421_, _maxi_read_rest_size[20:19] }), .Y(_07420_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29227_ ( .A({ _07422_, _maxi_read_rest_size[32:30] }), .Y(_07421_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29228_ ( .A({ _maxi_read_rest_size[28:27], _maxi_read_rest_size[25], _maxi_read_rest_size[22] }), .Y(_07422_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29229_ ( .A({ _maxi_read_rest_size[21], _maxi_read_rest_size[18:16] }), .Y(_07423_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29230_ ( .A({ _maxi_read_rest_size[29], _maxi_read_rest_size[26], _maxi_read_rest_size[24:23] }), .Y(_07424_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29231_ ( .A({ _07427_, _07426_ }), .Y(_07425_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29232_ ( .A(_maxi_read_rest_size[7:4]), .Y(_07426_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29233_ ( .A(_maxi_read_rest_size[3:0]), .Y(_07427_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29234_ ( .A({ _07429_, _maxi_read_rest_size[14], _maxi_read_rest_size[11:10] }), .Y(_07428_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29235_ ( .A({ _maxi_read_rest_size[15], _maxi_read_rest_size[13:12], _maxi_read_rest_size[9] }), .Y(_07429_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29236_ ( .A({ _15995_, _07334_, _15963_, _05071_ }), .Y(_15931_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _29237_ ( .A({ _07440_, _07432_, _11212_ }), .Y(conv2d_8_update_filter) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _29238_ ( .A({ cparam_conv2d_8_max_col_count[2], conv2d_8_row_count[2], _07431_ }), .Y(_07430_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29239_ ( .A({ cparam_conv2d_8_max_col_count[0], cparam_conv2d_8_max_col_count[1], conv2d_8_row_count[0], conv2d_8_row_count[1] }), .Y(_07431_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29240_ ( .A({ _07439_, _07438_, _07433_ }), .Y(_07432_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29241_ ( .A({ _07437_, _07436_, _07435_, _07434_ }), .Y(_07433_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29242_ ( .A(conv2d_8_row_count[23:20]), .Y(_07434_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29243_ ( .A(conv2d_8_row_count[19:16]), .Y(_07435_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29244_ ( .A({ conv2d_8_row_count[27], conv2d_8_row_count[31:29] }), .Y(_07436_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29245_ ( .A({ conv2d_8_row_count[28], conv2d_8_row_count[26:24] }), .Y(_07437_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29246_ ( .A(conv2d_8_row_count[15:12]), .Y(_07438_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29247_ ( .A(conv2d_8_row_count[11:8]), .Y(_07439_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _29248_ ( .A(conv2d_8_row_count[7:5]), .Y(_07440_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29249_ ( .A({ _15984_, _07334_, _15952_, _05071_ }), .Y(_15920_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29250_ ( .A({ _16002_, _07334_, _15970_, _05071_ }), .Y(_15938_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29251_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16165_, _16197_ }), .Y(_16133_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29252_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16260_, _16292_ }), .Y(_16228_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29253_ ( .A({ _07442_, _07450_, _stream_conv2d_8_source_28_source_pat_fsm_11[1] }), .Y(_07441_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29254_ ( .A({ _07449_, _07448_, _07443_ }), .Y(_07442_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29255_ ( .A({ _07447_, _07446_, _07445_, _07444_ }), .Y(_07443_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29256_ ( .A(_stream_conv2d_8_source_28_source_pat_fsm_11[23:20]), .Y(_07444_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29257_ ( .A(_stream_conv2d_8_source_28_source_pat_fsm_11[19:16]), .Y(_07445_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29258_ ( .A(_stream_conv2d_8_source_28_source_pat_fsm_11[31:28]), .Y(_07446_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29259_ ( .A(_stream_conv2d_8_source_28_source_pat_fsm_11[27:24]), .Y(_07447_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29260_ ( .A(_stream_conv2d_8_source_28_source_pat_fsm_11[15:12]), .Y(_07448_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29261_ ( .A(_stream_conv2d_8_source_28_source_pat_fsm_11[11:8]), .Y(_07449_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29262_ ( .A({ _07451_, _stream_conv2d_8_source_28_source_pat_fsm_11[3:2] }), .Y(_07450_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29263_ ( .A(_stream_conv2d_8_source_28_source_pat_fsm_11[7:4]), .Y(_07451_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29264_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16737_, _16769_ }), .Y(_16705_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29265_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16834_, _16866_ }), .Y(_16802_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29266_ ( .A({ _17970_, _07122_, _17616_, _05102_ }), .Y(_18002_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29267_ ( .A({ _07457_, _07452_ }), .Y(_05240_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29268_ ( .A({ _07456_, _07455_, _07454_, _07453_ }), .Y(_07452_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29269_ ( .A({ _04009_, _04008_, _04007_, _04006_ }), .Y(_07453_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29270_ ( .A({ _04004_, _04003_, _04002_, _04001_ }), .Y(_07454_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29271_ ( .A({ _04018_, _04017_, _04015_, _04014_ }), .Y(_07455_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29272_ ( .A({ _04013_, _04012_, _04011_, _04010_ }), .Y(_07456_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29273_ ( .A({ _07461_, _07460_, _07459_, _07458_ }), .Y(_07457_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _29274_ ( .A({ _04019_, _04016_, _03994_, _04005_ }), .Y(_07458_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29275_ ( .A({ _04023_, _04022_, _04021_, _04020_ }), .Y(_07459_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29276_ ( .A({ _04000_, _03999_, _03998_, _03997_ }), .Y(_07460_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29277_ ( .A({ _03996_, _03995_, _04025_, _04024_ }), .Y(_07461_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _29278_ ( .A({ _07483_, _07480_, _07476_, _07463_ }), .Y(_07462_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _29279_ ( .A({ _07471_, _07475_, _07464_, _07474_ }), .Y(_07463_) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _29280_ ( .A({ conv2d_8_sync_comp_count[5], _07465_, _07470_, _03925_ }), .Y(_07464_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _29281_ ( .A({ _07466_, _07469_, _07468_, _07467_ }), .Y(_07465_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29282_ ( .A({ conv2d_8_sync_comp_count[3], _03923_, conv2d_8_sync_comp_count[4], _03924_ }), .Y(_07466_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29283_ ( .A({ conv2d_8_sync_comp_count[2], _03920_ }), .Y(_07467_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _29284_ ( .A({ _03898_, conv2d_8_sync_comp_count[0], conv2d_8_sync_comp_count[1], _03909_ }), .Y(_07468_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29285_ ( .A({ _03920_, conv2d_8_sync_comp_count[2], _03923_, conv2d_8_sync_comp_count[3] }), .Y(_07469_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29286_ ( .A({ _03924_, conv2d_8_sync_comp_count[4] }), .Y(_07470_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _29287_ ( .A({ _07473_, _07472_, _03927_, conv2d_8_sync_comp_count[7] }), .Y(_07471_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29288_ ( .A({ conv2d_8_sync_comp_count[11], _03900_, conv2d_8_sync_comp_count[10], _03899_ }), .Y(_07472_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29289_ ( .A({ conv2d_8_sync_comp_count[9], _03929_, conv2d_8_sync_comp_count[8], _03928_ }), .Y(_07473_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29290_ ( .A({ _03926_, conv2d_8_sync_comp_count[6] }), .Y(_07474_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29291_ ( .A({ conv2d_8_sync_comp_count[6], _03926_, conv2d_8_sync_comp_count[7], _03927_ }), .Y(_07475_) );
  \$lut  #( .LUT(16'h0071), .WIDTH(4) ) _29292_ ( .A({ _07477_, _03900_, conv2d_8_sync_comp_count[11], _07479_ }), .Y(_07476_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _29293_ ( .A({ _07472_, conv2d_8_sync_comp_count[9], _03929_, _07478_ }), .Y(_07477_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29294_ ( .A({ conv2d_8_sync_comp_count[8], _03928_ }), .Y(_07478_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29295_ ( .A({ conv2d_8_sync_comp_count[10], _03899_ }), .Y(_07479_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29296_ ( .A({ _07482_, _07481_ }), .Y(_07480_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29297_ ( .A({ conv2d_8_sync_comp_count[15], _03904_, conv2d_8_sync_comp_count[14], _03903_ }), .Y(_07481_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29298_ ( .A({ conv2d_8_sync_comp_count[13], _03902_, conv2d_8_sync_comp_count[12], _03901_ }), .Y(_07482_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _29299_ ( .A({ _07485_, _07481_, _07484_ }), .Y(_07483_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29300_ ( .A({ conv2d_8_sync_comp_count[12], conv2d_8_sync_comp_count[13], _03901_, _03902_ }), .Y(_07484_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29301_ ( .A({ conv2d_8_sync_comp_count[14], conv2d_8_sync_comp_count[15], _03903_, _03904_ }), .Y(_07485_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29302_ ( .A({ _07493_, _07487_ }), .Y(_07486_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29303_ ( .A({ _07492_, _07488_ }), .Y(_07487_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _29304_ ( .A({ _07491_, _07489_, _03910_, conv2d_8_sync_comp_count[20] }), .Y(_07488_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _29305_ ( .A({ _07490_, _03911_, conv2d_8_sync_comp_count[21] }), .Y(_07489_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29306_ ( .A({ conv2d_8_sync_comp_count[23], _03913_, conv2d_8_sync_comp_count[22], _03912_ }), .Y(_07490_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29307_ ( .A({ conv2d_8_sync_comp_count[20], _03910_, conv2d_8_sync_comp_count[21], _03911_ }), .Y(_07491_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29308_ ( .A({ conv2d_8_sync_comp_count[19], _03908_, conv2d_8_sync_comp_count[18], _03907_ }), .Y(_07492_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29309_ ( .A({ conv2d_8_sync_comp_count[17], _03906_, conv2d_8_sync_comp_count[16], _03905_ }), .Y(_07493_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _29310_ ( .A({ _07497_, _07495_, _07487_, _07499_ }), .Y(_07494_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29311_ ( .A({ _07488_, _07496_ }), .Y(_07495_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _29312_ ( .A({ conv2d_8_sync_comp_count[18], conv2d_8_sync_comp_count[19], _03907_, _03908_ }), .Y(_07496_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _29313_ ( .A({ _07498_, _07489_, _07491_ }), .Y(_07497_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _29314_ ( .A({ conv2d_8_sync_comp_count[22], conv2d_8_sync_comp_count[23], _03912_, _03913_ }), .Y(_07498_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29315_ ( .A({ conv2d_8_sync_comp_count[16], conv2d_8_sync_comp_count[17], _03905_, _03906_ }), .Y(_07499_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29316_ ( .A({ _07504_, _07501_ }), .Y(_07500_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29317_ ( .A({ _07503_, _07502_ }), .Y(_07501_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29318_ ( .A({ conv2d_8_sync_comp_count[31], _03922_, conv2d_8_sync_comp_count[30], _03921_ }), .Y(_07502_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29319_ ( .A({ conv2d_8_sync_comp_count[29], _03919_, conv2d_8_sync_comp_count[28], _03918_ }), .Y(_07503_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29320_ ( .A({ conv2d_8_sync_comp_count[27], _03917_, conv2d_8_sync_comp_count[26], _03916_ }), .Y(_07504_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29321_ ( .A({ conv2d_8_sync_comp_count[25], _03915_, conv2d_8_sync_comp_count[24], _03914_ }), .Y(_07505_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _29322_ ( .A({ _07510_, _07507_, _07501_, _07509_ }), .Y(_07506_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _29323_ ( .A({ _07502_, conv2d_8_sync_comp_count[29], _03919_, _07508_ }), .Y(_07507_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29324_ ( .A({ conv2d_8_sync_comp_count[28], _03918_ }), .Y(_07508_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29325_ ( .A({ conv2d_8_sync_comp_count[26], conv2d_8_sync_comp_count[27], _03916_, _03917_ }), .Y(_07509_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _29326_ ( .A({ conv2d_8_sync_comp_count[30], conv2d_8_sync_comp_count[31], _03921_, _03922_ }), .Y(_07510_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29327_ ( .A({ conv2d_8_sync_comp_count[24], conv2d_8_sync_comp_count[25], _03914_, _03915_ }), .Y(_07511_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29328_ ( .A({ _07524_, _07523_, _07521_, _07512_ }), .Y(_05238_) );
  \$lut  #( .LUT(16'hf400), .WIDTH(4) ) _29329_ ( .A({ _07516_, _07513_, _counter_count_762[3], _21867_ }), .Y(_07512_) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _29330_ ( .A({ _21864_, _07514_, _07515_, _counter_count_762[2] }), .Y(_07513_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29331_ ( .A({ _21842_, _counter_count_762[0], _21853_, _counter_count_762[1] }), .Y(_07514_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29332_ ( .A({ _counter_count_762[1], _21853_ }), .Y(_07515_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29333_ ( .A({ _07520_, _07519_, _07518_, _07517_ }), .Y(_07516_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29334_ ( .A({ _21857_, _21854_, _21851_, _21850_ }), .Y(_07517_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29335_ ( .A({ _21865_, _21863_, _21861_, _21858_ }), .Y(_07518_) );
  \$lut  #( .LUT(16'h000d), .WIDTH(4) ) _29336_ ( .A({ _21870_, _21869_, _counter_count_762[3], _21867_ }), .Y(_07519_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29337_ ( .A({ _21848_, _21845_, _21843_, _21873_ }), .Y(_07520_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29338_ ( .A({ _07522_, _21871_, _21868_ }), .Y(_07521_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29339_ ( .A({ _21847_, _21846_, _21844_, _21872_ }), .Y(_07522_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29340_ ( .A({ _21856_, _21855_, _21852_, _21849_ }), .Y(_07523_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29341_ ( .A({ _21866_, _21862_, _21860_, _21859_ }), .Y(_07524_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29342_ ( .A({ _17969_, _07122_, _17615_, _05102_ }), .Y(_18001_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29343_ ( .A({ _17968_, _07122_, _17614_, _05102_ }), .Y(_18000_) );
  \$lut  #( .LUT(8'h71), .WIDTH(3) ) _29344_ ( .A({ _21835_, _pulse_count_193[3], _07526_ }), .Y(_07525_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _29345_ ( .A({ _pulse_count_193[2], _21832_, _07527_ }), .Y(_07526_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _29346_ ( .A({ _21810_, _pulse_count_193[0], _pulse_count_193[1], _21821_ }), .Y(_07527_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29347_ ( .A({ _21839_, _pulse_count_193[7] }), .Y(_07528_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29348_ ( .A({ _pulse_count_193[7], _21839_, _pulse_count_193[6], _21838_ }), .Y(_07529_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29349_ ( .A({ _07533_, _07531_ }), .Y(_07530_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29350_ ( .A({ _07532_, _21833_, _21825_, _21823_ }), .Y(_07531_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29351_ ( .A({ _21817_, _21814_, _21831_, _21826_ }), .Y(_07532_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29352_ ( .A({ _07537_, _07536_, _07535_, _07534_ }), .Y(_07533_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29353_ ( .A({ _21824_, _21820_, _21819_, _21816_ }), .Y(_07534_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29354_ ( .A({ _21815_, _21813_, _21812_, _21841_ }), .Y(_07535_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29355_ ( .A({ _21818_, _21811_, _21828_, _21827_ }), .Y(_07536_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29356_ ( .A({ _21834_, _21830_, _21829_, _21822_ }), .Y(_07537_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29357_ ( .A({ _17998_, _07122_, _17644_, _05102_ }), .Y(_18030_) );
  \$lut  #( .LUT(8'h71), .WIDTH(3) ) _29358_ ( .A({ _21837_, _reducecustom_count_191[5], _07539_ }), .Y(_07538_) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _29359_ ( .A({ _21836_, _07540_, _07543_, _reducecustom_count_191[4] }), .Y(_07539_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _29360_ ( .A({ _07542_, _reducecustom_count_191[2], _21832_, _07541_ }), .Y(_07540_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _29361_ ( .A({ _21810_, _21821_, _reducecustom_count_191[0], _reducecustom_count_191[1] }), .Y(_07541_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29362_ ( .A({ _21835_, _reducecustom_count_191[3] }), .Y(_07542_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29363_ ( .A({ _reducecustom_count_191[3], _21835_ }), .Y(_07543_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29364_ ( .A({ _17996_, _07122_, _17642_, _05102_ }), .Y(_18028_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29365_ ( .A({ _17995_, _07122_, _17641_, _05102_ }), .Y(_18027_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29366_ ( .A({ _17994_, _07122_, _17640_, _05102_ }), .Y(_18026_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29367_ ( .A({ _17993_, _07122_, _17639_, _05102_ }), .Y(_18025_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29368_ ( .A({ _17992_, _07122_, _17638_, _05102_ }), .Y(_18024_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29369_ ( .A({ _17989_, _07122_, _17635_, _05102_ }), .Y(_18021_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29370_ ( .A({ _17978_, _07122_, _17624_, _05102_ }), .Y(_18010_) );
  \$lut  #( .LUT(16'h004f), .WIDTH(4) ) _29371_ ( .A({ _07588_, _07561_, _07586_, _07544_ }), .Y(_05234_) );
  \$lut  #( .LUT(16'hbf00), .WIDTH(4) ) _29372_ ( .A({ _07556_, _07560_, _07557_, _07545_ }), .Y(_07544_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _29373_ ( .A({ _07555_, _07550_, _11298_, _07553_ }), .Y(_07545_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29374_ ( .A({ _21799_, _pulse_count_17[2], _21803_, _pulse_count_17[3] }), .Y(_07546_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29375_ ( .A({ _pulse_count_17[3], _21803_, _pulse_count_17[4], _21804_ }), .Y(_07547_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29376_ ( .A({ _21804_, _pulse_count_17[4], _21805_, _pulse_count_17[5] }), .Y(_07548_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29377_ ( .A({ _pulse_count_17[5], _21805_, _pulse_count_17[6], _21806_ }), .Y(_07549_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _29378_ ( .A({ _07552_, _07551_, _21809_, _pulse_count_17[9] }), .Y(_07550_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29379_ ( .A({ _pulse_count_17[8], _21808_, _pulse_count_17[9], _21809_ }), .Y(_07551_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29380_ ( .A({ _pulse_count_17[11], _21779_, _pulse_count_17[10], _21778_ }), .Y(_07552_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29381_ ( .A({ _07554_, _07552_, _07551_ }), .Y(_07553_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29382_ ( .A({ _21808_, _pulse_count_17[8], _21809_, _pulse_count_17[9] }), .Y(_07554_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _29383_ ( .A({ _pulse_count_17[10], _pulse_count_17[11], _21778_, _21779_ }), .Y(_07555_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _29384_ ( .A({ _07558_, _07557_, _07559_ }), .Y(_07556_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29385_ ( .A({ _pulse_count_17[15], _21783_, _pulse_count_17[14], _21782_ }), .Y(_07557_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29386_ ( .A({ _pulse_count_17[14], _pulse_count_17[15], _21782_, _21783_ }), .Y(_07558_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29387_ ( .A({ _pulse_count_17[12], _pulse_count_17[13], _21780_, _21781_ }), .Y(_07559_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29388_ ( .A({ _pulse_count_17[13], _21781_, _pulse_count_17[12], _21780_ }), .Y(_07560_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _29389_ ( .A({ _07562_, _07575_, _07585_ }), .Y(_07561_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _29390_ ( .A({ _07571_, _07563_, _07566_, _07574_ }), .Y(_07562_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _29391_ ( .A({ _07564_, _07569_, _07570_, _07565_ }), .Y(_07563_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _29392_ ( .A({ _07568_, _07565_, _21794_, _pulse_count_17[25] }), .Y(_07564_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29393_ ( .A({ _07567_, _07566_ }), .Y(_07565_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29394_ ( .A({ _pulse_count_17[31], _21801_, _pulse_count_17[30], _21800_ }), .Y(_07566_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29395_ ( .A({ _pulse_count_17[29], _21798_, _pulse_count_17[28], _21797_ }), .Y(_07567_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29396_ ( .A({ _pulse_count_17[27], _21796_, _pulse_count_17[26], _21795_ }), .Y(_07568_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29397_ ( .A({ _pulse_count_17[24], _21793_, _pulse_count_17[25], _21794_ }), .Y(_07569_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29398_ ( .A({ _pulse_count_17[26], _pulse_count_17[27], _21795_, _21796_ }), .Y(_07570_) );
  \$lut  #( .LUT(16'h0071), .WIDTH(4) ) _29399_ ( .A({ _07573_, _21801_, _pulse_count_17[31], _07572_ }), .Y(_07571_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29400_ ( .A({ _pulse_count_17[30], _21800_ }), .Y(_07572_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29401_ ( .A({ _pulse_count_17[32], _21802_ }), .Y(_07573_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29402_ ( .A({ _pulse_count_17[28], _pulse_count_17[29], _21797_, _21798_ }), .Y(_07574_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _29403_ ( .A({ _07584_, _07576_, _07578_, _07580_ }), .Y(_07575_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _29404_ ( .A({ _07577_, _07581_, _07583_, _07582_ }), .Y(_07576_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _29405_ ( .A({ _07580_, _07578_, _21789_, _pulse_count_17[20] }), .Y(_07577_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _29406_ ( .A({ _07579_, _pulse_count_17[22], _21791_ }), .Y(_07578_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _29407_ ( .A({ _pulse_count_17[23], _21792_, _21790_, _pulse_count_17[21] }), .Y(_07579_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29408_ ( .A({ _pulse_count_17[20], _21789_, _pulse_count_17[21], _21790_ }), .Y(_07580_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29409_ ( .A({ _pulse_count_17[18], _pulse_count_17[19], _21786_, _21787_ }), .Y(_07581_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29410_ ( .A({ _pulse_count_17[19], _21787_, _pulse_count_17[18], _21786_ }), .Y(_07582_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29411_ ( .A({ _pulse_count_17[16], _pulse_count_17[17], _21784_, _21785_ }), .Y(_07583_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _29412_ ( .A({ _pulse_count_17[22], _pulse_count_17[23], _21791_, _21792_ }), .Y(_07584_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _29413_ ( .A({ _07569_, _07564_, _21793_, _pulse_count_17[24] }), .Y(_07585_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29414_ ( .A({ _07587_, _07582_, _07577_, _07585_ }), .Y(_07586_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29415_ ( .A({ _pulse_count_17[17], _21785_, _pulse_count_17[16], _21784_ }), .Y(_07587_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29416_ ( .A({ _21802_, _pulse_count_17[32] }), .Y(_07588_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29417_ ( .A({ _17967_, _07122_, _17613_, _05102_ }), .Y(_17999_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _29418_ ( .A({ _07623_, _07612_, _07632_, _07590_ }), .Y(_07589_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _29419_ ( .A({ _07608_, _07605_, _07611_, _07591_ }), .Y(_07590_) );
  \$lut  #( .LUT(16'hffb0), .WIDTH(4) ) _29420_ ( .A({ _07602_, _11220_, _07604_, _07592_ }), .Y(_07591_) );
  \$lut  #( .LUT(16'h00f4), .WIDTH(4) ) _29421_ ( .A({ _07598_, _07599_, _07600_, _07593_ }), .Y(_07592_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _29422_ ( .A({ _07597_, _07596_, _07594_, _07595_ }), .Y(_07593_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29423_ ( .A({ _reduceadd_count_15[2], _21799_ }), .Y(_07594_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _29424_ ( .A({ _21777_, _21788_, _reduceadd_count_15[0], _reduceadd_count_15[1] }), .Y(_07595_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29425_ ( .A({ _21799_, _reduceadd_count_15[2], _21803_, _reduceadd_count_15[3] }), .Y(_07596_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29426_ ( .A({ _reduceadd_count_15[3], _21803_, _reduceadd_count_15[4], _21804_ }), .Y(_07597_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29427_ ( .A({ _21806_, _reduceadd_count_15[6] }), .Y(_07598_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29428_ ( .A({ _reduceadd_count_15[5], _21805_ }), .Y(_07599_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29429_ ( .A({ _21804_, _reduceadd_count_15[4], _21805_, _reduceadd_count_15[5] }), .Y(_07600_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29430_ ( .A({ _21779_, _reduceadd_count_15[11], _21778_, _reduceadd_count_15[10] }), .Y(_07601_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29431_ ( .A({ _07601_, _07603_ }), .Y(_07602_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _29432_ ( .A({ _reduceadd_count_15[8], _21808_, _21809_, _reduceadd_count_15[9] }), .Y(_07603_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29433_ ( .A({ _reduceadd_count_15[6], _21806_, _reduceadd_count_15[7], _21807_ }), .Y(_07604_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29434_ ( .A({ _07607_, _07606_ }), .Y(_07605_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29435_ ( .A({ _21783_, _reduceadd_count_15[15], _21782_, _reduceadd_count_15[14] }), .Y(_07606_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29436_ ( .A({ _21781_, _reduceadd_count_15[13], _21780_, _reduceadd_count_15[12] }), .Y(_07607_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _29437_ ( .A({ _07610_, _07606_, _07609_ }), .Y(_07608_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _29438_ ( .A({ _reduceadd_count_15[12], _21780_, _21781_, _reduceadd_count_15[13] }), .Y(_07609_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _29439_ ( .A({ _reduceadd_count_15[14], _21782_, _21783_, _reduceadd_count_15[15] }), .Y(_07610_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _29440_ ( .A({ _reduceadd_count_15[10], _21778_, _21779_, _reduceadd_count_15[11] }), .Y(_07611_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _29441_ ( .A({ _07622_, _07620_, _07613_ }), .Y(_07612_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _29442_ ( .A({ _07614_, _07619_, _07617_, _07618_ }), .Y(_07613_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29443_ ( .A({ _07616_, _07615_ }), .Y(_07614_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29444_ ( .A({ _21792_, _reduceadd_count_15[23], _21791_, _reduceadd_count_15[22] }), .Y(_07615_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29445_ ( .A({ _21790_, _reduceadd_count_15[21], _21789_, _reduceadd_count_15[20] }), .Y(_07616_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29446_ ( .A({ _21787_, _reduceadd_count_15[19], _21786_, _reduceadd_count_15[18] }), .Y(_07617_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _29447_ ( .A({ _reduceadd_count_15[16], _21784_, _21785_, _reduceadd_count_15[17] }), .Y(_07618_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _29448_ ( .A({ _reduceadd_count_15[18], _21786_, _21787_, _reduceadd_count_15[19] }), .Y(_07619_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _29449_ ( .A({ _07615_, _reduceadd_count_15[21], _21790_, _07621_ }), .Y(_07620_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29450_ ( .A({ _reduceadd_count_15[20], _21789_ }), .Y(_07621_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _29451_ ( .A({ _reduceadd_count_15[22], _21791_, _21792_, _reduceadd_count_15[23] }), .Y(_07622_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29452_ ( .A({ _07630_, _07628_, _07624_ }), .Y(_07623_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _29453_ ( .A({ _07627_, _07625_, _reduceadd_count_15[28], _21797_ }), .Y(_07624_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _29454_ ( .A({ _07626_, _21801_, _reduceadd_count_15[31] }), .Y(_07625_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _29455_ ( .A({ _21800_, _reduceadd_count_15[30], _21798_, _reduceadd_count_15[29] }), .Y(_07626_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29456_ ( .A({ _reduceadd_count_15[28], _21797_, _reduceadd_count_15[29], _21798_ }), .Y(_07627_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _29457_ ( .A({ _07629_, _reduceadd_count_15[24], _21793_ }), .Y(_07628_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29458_ ( .A({ _reduceadd_count_15[24], _21793_, _reduceadd_count_15[25], _21794_ }), .Y(_07629_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _29459_ ( .A({ _07631_, _21795_, _reduceadd_count_15[26] }), .Y(_07630_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _29460_ ( .A({ _21796_, _reduceadd_count_15[27], _21794_, _reduceadd_count_15[25] }), .Y(_07631_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29461_ ( .A({ _07633_, _07617_, _07614_ }), .Y(_07632_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29462_ ( .A({ _21785_, _reduceadd_count_15[17], _21784_, _reduceadd_count_15[16] }), .Y(_07633_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _29463_ ( .A({ _07635_, _07630_, _07629_ }), .Y(_07634_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _29464_ ( .A({ _reduceadd_count_15[26], _21795_, _21796_, _reduceadd_count_15[27] }), .Y(_07635_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _29465_ ( .A({ _reduceadd_count_15[30], _21800_, _reduceadd_count_15[31], _21801_ }), .Y(_07636_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29466_ ( .A({ _07637_, _18539_, _07019_ }), .Y(_18443_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29467_ ( .A({ _18475_, maxi_rready, _18507_, _07638_ }), .Y(_07637_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29468_ ( .A({ _07017_, _07639_ }), .Y(_07638_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _29469_ ( .A({ _maxi_read_fsm[1], _07009_, _07014_, _maxi_read_fsm[0] }), .Y(_07639_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29470_ ( .A({ _07640_, _18542_, _07019_ }), .Y(_18446_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29471_ ( .A({ _18478_, maxi_rready, _18510_, _07638_ }), .Y(_07640_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29472_ ( .A({ _07641_, _18541_, _07019_ }), .Y(_18445_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29473_ ( .A({ _18477_, maxi_rready, _18509_, _07638_ }), .Y(_07641_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29474_ ( .A({ _07642_, _18536_, _07019_ }), .Y(_18440_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29475_ ( .A({ _18472_, maxi_rready, _18504_, _07638_ }), .Y(_07642_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29476_ ( .A({ _07643_, _18538_, _07019_ }), .Y(_18442_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29477_ ( .A({ _18474_, maxi_rready, _18506_, _07638_ }), .Y(_07643_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29478_ ( .A({ _07644_, _18537_, _07019_ }), .Y(_18441_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29479_ ( .A({ _18473_, maxi_rready, _18505_, _07638_ }), .Y(_07644_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29480_ ( .A({ _07645_, _18533_, _07019_ }), .Y(_18437_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29481_ ( .A({ _18469_, maxi_rready, _18501_, _07638_ }), .Y(_07645_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29482_ ( .A({ _07646_, _18535_, _07019_ }), .Y(_18439_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29483_ ( .A({ _18471_, maxi_rready, _18503_, _07638_ }), .Y(_07646_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29484_ ( .A({ _07647_, _18534_, _07019_ }), .Y(_18438_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29485_ ( .A({ _18470_, maxi_rready, _18502_, _07638_ }), .Y(_07647_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29486_ ( .A({ _07648_, _18530_, _07019_ }), .Y(_18434_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29487_ ( .A({ _18466_, maxi_rready, _18498_, _07638_ }), .Y(_07648_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29488_ ( .A({ _07649_, _18532_, _07019_ }), .Y(_18436_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29489_ ( .A({ _18468_, maxi_rready, _18500_, _07638_ }), .Y(_07649_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29490_ ( .A({ _07650_, _18531_, _07019_ }), .Y(_18435_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29491_ ( .A({ _18467_, maxi_rready, _18499_, _07638_ }), .Y(_07650_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29492_ ( .A({ _07651_, _18526_, _07019_ }), .Y(_18430_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29493_ ( .A({ _18462_, maxi_rready, _18494_, _07638_ }), .Y(_07651_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29494_ ( .A({ _07652_, _18528_, _07019_ }), .Y(_18432_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29495_ ( .A({ _18464_, maxi_rready, _18496_, _07638_ }), .Y(_07652_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29496_ ( .A({ _07653_, _18527_, _07019_ }), .Y(_18431_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29497_ ( .A({ _18463_, maxi_rready, _18495_, _07638_ }), .Y(_07653_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29498_ ( .A({ _07654_, _18523_, _07019_ }), .Y(_18427_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29499_ ( .A({ _18459_, maxi_rready, _18491_, _07638_ }), .Y(_07654_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29500_ ( .A({ _07655_, _18525_, _07019_ }), .Y(_18429_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29501_ ( .A({ _18461_, maxi_rready, _18493_, _07638_ }), .Y(_07655_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29502_ ( .A({ _07656_, _18524_, _07019_ }), .Y(_18428_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29503_ ( .A({ _18460_, maxi_rready, _18492_, _07638_ }), .Y(_07656_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29504_ ( .A({ _07657_, _18520_, _07019_ }), .Y(_18424_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29505_ ( .A({ _18456_, maxi_rready, _18488_, _07638_ }), .Y(_07657_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29506_ ( .A({ _07658_, _18522_, _07019_ }), .Y(_18426_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29507_ ( .A({ _18458_, maxi_rready, _18490_, _07638_ }), .Y(_07658_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29508_ ( .A({ _07659_, _18521_, _07019_ }), .Y(_18425_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29509_ ( .A({ _18457_, maxi_rready, _18489_, _07638_ }), .Y(_07659_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29510_ ( .A({ _07660_, _18548_, _07019_ }), .Y(_18452_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29511_ ( .A({ _18484_, maxi_rready, _18516_, _07638_ }), .Y(_07660_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29512_ ( .A({ _07661_, _18519_, _07019_ }), .Y(_18423_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29513_ ( .A({ _18455_, maxi_rready, _18487_, _07638_ }), .Y(_07661_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29514_ ( .A({ _07662_, _18549_, _07019_ }), .Y(_18453_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29515_ ( .A({ _18485_, maxi_rready, _18517_, _07638_ }), .Y(_07662_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29516_ ( .A({ _07663_, _18545_, _07019_ }), .Y(_18449_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29517_ ( .A({ _18481_, maxi_rready, _18513_, _07638_ }), .Y(_07663_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29518_ ( .A({ _07664_, _18547_, _07019_ }), .Y(_18451_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29519_ ( .A({ _18483_, maxi_rready, _18515_, _07638_ }), .Y(_07664_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29520_ ( .A({ _07665_, _18546_, _07019_ }), .Y(_18450_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29521_ ( .A({ _18482_, maxi_rready, _18514_, _07638_ }), .Y(_07665_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29522_ ( .A({ _07666_, _18540_, _07019_ }), .Y(_18444_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _29523_ ( .A({ _07667_, _07638_, _18508_ }), .Y(_07666_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _29524_ ( .A({ _05105_, maxi_rready, _18476_ }), .Y(_07667_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _29525_ ( .A({ _07008_, _07668_, _maxi_read_fsm[0] }), .Y(_05105_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _29526_ ( .A({ _maxi_read_fsm[2], _07018_, _maxi_read_fsm[1], _maxi_read_fsm[3] }), .Y(_07668_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29527_ ( .A({ _07669_, _18544_, _07019_ }), .Y(_18448_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29528_ ( .A({ _18480_, maxi_rready, _18512_, _07638_ }), .Y(_07669_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29529_ ( .A({ _07670_, _18543_, _07019_ }), .Y(_18447_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29530_ ( .A({ _18479_, maxi_rready, _18511_, _07638_ }), .Y(_07670_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29531_ ( .A({ _07671_, _18529_, _07019_ }), .Y(_18433_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _29532_ ( .A({ _07672_, maxi_rready, _18465_ }), .Y(_07671_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _29533_ ( .A({ _05107_, _07638_, _18497_ }), .Y(_07672_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29534_ ( .A({ _07673_, _18518_, _07019_ }), .Y(_18422_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _29535_ ( .A({ _07674_, maxi_rready, _18454_ }), .Y(_07673_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _29536_ ( .A({ _05105_, _07638_, _18486_ }), .Y(_07674_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29537_ ( .A({ _05107_, _07019_ }), .Y(_04830_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29538_ ( .A({ _07675_, _21923_ }), .Y(_21924_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _29539_ ( .A({ _05107_, _07638_, _07008_, _07668_ }), .Y(_07675_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29540_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16923_, _16955_ }), .Y(_16891_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29541_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16736_, _16768_ }), .Y(_16704_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29542_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16823_, _16855_ }), .Y(_16791_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29543_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16733_, _16765_ }), .Y(_16701_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29544_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16732_, _16764_ }), .Y(_16700_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29545_ ( .A({ _05067_, _07676_ }), .Y(_21904_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29546_ ( .A({ _07677_, _07682_, _stream_conv2d_8_source_33_source_pat_fsm_16[0] }), .Y(_07676_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29547_ ( .A({ _07681_, _07680_, _07678_ }), .Y(_07677_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29548_ ( .A({ _07679_, _stream_conv2d_8_source_33_source_pat_fsm_16[3:2] }), .Y(_07678_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29549_ ( .A(_stream_conv2d_8_source_33_source_pat_fsm_16[7:4]), .Y(_07679_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29550_ ( .A(_stream_conv2d_8_source_33_source_pat_fsm_16[15:12]), .Y(_07680_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29551_ ( .A(_stream_conv2d_8_source_33_source_pat_fsm_16[11:8]), .Y(_07681_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29552_ ( .A({ _07686_, _07685_, _07684_, _07683_ }), .Y(_07682_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29553_ ( .A(_stream_conv2d_8_source_33_source_pat_fsm_16[23:20]), .Y(_07683_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29554_ ( .A(_stream_conv2d_8_source_33_source_pat_fsm_16[19:16]), .Y(_07684_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29555_ ( .A(_stream_conv2d_8_source_33_source_pat_fsm_16[31:28]), .Y(_07685_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29556_ ( .A(_stream_conv2d_8_source_33_source_pat_fsm_16[27:24]), .Y(_07686_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29557_ ( .A({ _07677_, _stream_conv2d_8_source_33_source_pat_fsm_16[0], _07682_, _stream_conv2d_8_source_33_source_pat_fsm_16[1] }), .Y(_05067_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29558_ ( .A({ _15788_, _07687_, _15756_, _05067_ }), .Y(_15724_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29559_ ( .A({ _07676_, _stream_conv2d_8_source_33_source_pat_fsm_16[1] }), .Y(_07687_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29560_ ( .A({ _15799_, _07687_, _15767_, _05067_ }), .Y(_15735_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29561_ ( .A({ _15810_, _07687_, _15778_, _05067_ }), .Y(_15746_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29562_ ( .A({ _15813_, _07687_, _15781_, _05067_ }), .Y(_15749_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29563_ ( .A({ _15814_, _07687_, _15782_, _05067_ }), .Y(_15750_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29564_ ( .A({ _15815_, _07687_, _15783_, _05067_ }), .Y(_15751_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29565_ ( .A({ _15816_, _07687_, _15784_, _05067_ }), .Y(_15752_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29566_ ( .A({ _15817_, _07687_, _15785_, _05067_ }), .Y(_15753_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29567_ ( .A({ _15818_, _07687_, _15786_, _05067_ }), .Y(_15754_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29568_ ( .A({ _15819_, _07687_, _15787_, _05067_ }), .Y(_15755_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29569_ ( .A({ _15789_, _07687_, _15757_, _05067_ }), .Y(_15725_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29570_ ( .A({ _15790_, _07687_, _15758_, _05067_ }), .Y(_15726_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29571_ ( .A({ _15791_, _07687_, _15759_, _05067_ }), .Y(_15727_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29572_ ( .A({ _15792_, _07687_, _15760_, _05067_ }), .Y(_15728_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29573_ ( .A({ _15793_, _07687_, _15761_, _05067_ }), .Y(_15729_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29574_ ( .A({ _15794_, _07687_, _15762_, _05067_ }), .Y(_15730_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29575_ ( .A({ _15795_, _07687_, _15763_, _05067_ }), .Y(_15731_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29576_ ( .A({ _15796_, _07687_, _15764_, _05067_ }), .Y(_15732_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29577_ ( .A({ _15797_, _07687_, _15765_, _05067_ }), .Y(_15733_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29578_ ( .A({ _15798_, _07687_, _15766_, _05067_ }), .Y(_15734_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29579_ ( .A({ _15800_, _07687_, _15768_, _05067_ }), .Y(_15736_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29580_ ( .A({ _15801_, _07687_, _15769_, _05067_ }), .Y(_15737_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29581_ ( .A({ _15802_, _07687_, _15770_, _05067_ }), .Y(_15738_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29582_ ( .A({ _15803_, _07687_, _15771_, _05067_ }), .Y(_15739_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29583_ ( .A({ _15804_, _07687_, _15772_, _05067_ }), .Y(_15740_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29584_ ( .A({ _15805_, _07687_, _15773_, _05067_ }), .Y(_15741_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29585_ ( .A({ _05082_, _07078_ }), .Y(_21912_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29586_ ( .A({ _stream_conv2d_8_source_25_source_pat_fsm_8[1], _07079_, _07087_, _stream_conv2d_8_source_25_source_pat_fsm_8[0] }), .Y(_05082_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29587_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17010_, _17042_ }), .Y(_16978_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29588_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17015_, _17047_ }), .Y(_16983_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29589_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16922_, _16954_ }), .Y(_16890_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29590_ ( .A({ _15806_, _07687_, _15774_, _05067_ }), .Y(_15742_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29591_ ( .A({ _15807_, _07687_, _15775_, _05067_ }), .Y(_15743_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29592_ ( .A({ _15808_, _07687_, _15776_, _05067_ }), .Y(_15744_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29593_ ( .A({ _15809_, _07687_, _15777_, _05067_ }), .Y(_15745_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29594_ ( .A({ _15811_, _07687_, _15779_, _05067_ }), .Y(_15747_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29595_ ( .A({ _15812_, _07687_, _15780_, _05067_ }), .Y(_15748_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29596_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16735_, _16767_ }), .Y(_16703_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29597_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16812_, _16844_ }), .Y(_16780_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29598_ ( .A({ _07335_, _stream_conv2d_8_source_20_source_pat_fsm_3[0], _17008_, _17040_ }), .Y(_16976_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29599_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16741_, _16773_ }), .Y(_16709_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29600_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17124_, _17156_ }), .Y(_17092_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29601_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17104_, _17136_ }), .Y(_17072_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29602_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16539_, _16571_ }), .Y(_16507_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29603_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17125_, _17157_ }), .Y(_17093_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29604_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16643_, _16675_ }), .Y(_16611_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29605_ ( .A({ _07347_, _stream_conv2d_8_source_21_source_pat_fsm_4[0], _16910_, _16942_ }), .Y(_16878_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29606_ ( .A({ _07358_, _stream_conv2d_8_source_24_source_pat_fsm_7[0], _16628_, _16660_ }), .Y(_16596_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29607_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16835_, _16867_ }), .Y(_16803_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29608_ ( .A({ _07369_, _stream_conv2d_8_source_22_source_pat_fsm_5[0], _16839_, _16871_ }), .Y(_16807_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29609_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16734_, _16766_ }), .Y(_16702_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29610_ ( .A({ _07078_, _stream_conv2d_8_source_25_source_pat_fsm_8[0], _16537_, _16569_ }), .Y(_16505_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29611_ ( .A({ _05066_, _07688_ }), .Y(_21903_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29612_ ( .A({ _07689_, _07694_, _stream_conv2d_8_source_34_source_pat_fsm_17[0] }), .Y(_07688_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29613_ ( .A({ _07693_, _07692_, _07690_ }), .Y(_07689_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29614_ ( .A({ _07691_, _stream_conv2d_8_source_34_source_pat_fsm_17[3:2] }), .Y(_07690_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29615_ ( .A(_stream_conv2d_8_source_34_source_pat_fsm_17[7:4]), .Y(_07691_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29616_ ( .A(_stream_conv2d_8_source_34_source_pat_fsm_17[15:12]), .Y(_07692_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29617_ ( .A(_stream_conv2d_8_source_34_source_pat_fsm_17[11:8]), .Y(_07693_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29618_ ( .A({ _07698_, _07697_, _07696_, _07695_ }), .Y(_07694_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29619_ ( .A(_stream_conv2d_8_source_34_source_pat_fsm_17[23:20]), .Y(_07695_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29620_ ( .A(_stream_conv2d_8_source_34_source_pat_fsm_17[19:16]), .Y(_07696_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29621_ ( .A(_stream_conv2d_8_source_34_source_pat_fsm_17[31:28]), .Y(_07697_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29622_ ( .A(_stream_conv2d_8_source_34_source_pat_fsm_17[27:24]), .Y(_07698_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29623_ ( .A({ _07689_, _stream_conv2d_8_source_34_source_pat_fsm_17[0], _07694_, _stream_conv2d_8_source_34_source_pat_fsm_17[1] }), .Y(_05066_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29624_ ( .A({ _15692_, _07699_, _15660_, _05066_ }), .Y(_15628_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29625_ ( .A({ _07688_, _stream_conv2d_8_source_34_source_pat_fsm_17[1] }), .Y(_07699_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29626_ ( .A({ _15703_, _07699_, _15671_, _05066_ }), .Y(_15639_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29627_ ( .A({ _15714_, _07699_, _15682_, _05066_ }), .Y(_15650_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29628_ ( .A({ _15717_, _07699_, _15685_, _05066_ }), .Y(_15653_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29629_ ( .A({ _15718_, _07699_, _15686_, _05066_ }), .Y(_15654_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29630_ ( .A({ _15719_, _07699_, _15687_, _05066_ }), .Y(_15655_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29631_ ( .A({ _15720_, _07699_, _15688_, _05066_ }), .Y(_15656_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29632_ ( .A({ _15721_, _07699_, _15689_, _05066_ }), .Y(_15657_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29633_ ( .A({ _15722_, _07699_, _15690_, _05066_ }), .Y(_15658_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29634_ ( .A({ _15723_, _07699_, _15691_, _05066_ }), .Y(_15659_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29635_ ( .A({ _15693_, _07699_, _15661_, _05066_ }), .Y(_15629_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29636_ ( .A({ _15694_, _07699_, _15662_, _05066_ }), .Y(_15630_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29637_ ( .A({ _15695_, _07699_, _15663_, _05066_ }), .Y(_15631_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29638_ ( .A({ _15696_, _07699_, _15664_, _05066_ }), .Y(_15632_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29639_ ( .A({ _15697_, _07699_, _15665_, _05066_ }), .Y(_15633_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29640_ ( .A({ _15698_, _07699_, _15666_, _05066_ }), .Y(_15634_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29641_ ( .A({ _15699_, _07699_, _15667_, _05066_ }), .Y(_15635_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29642_ ( .A({ _15700_, _07699_, _15668_, _05066_ }), .Y(_15636_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29643_ ( .A({ _15701_, _07699_, _15669_, _05066_ }), .Y(_15637_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29644_ ( .A({ _15702_, _07699_, _15670_, _05066_ }), .Y(_15638_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29645_ ( .A({ _15704_, _07699_, _15672_, _05066_ }), .Y(_15640_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29646_ ( .A({ _15705_, _07699_, _15673_, _05066_ }), .Y(_15641_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29647_ ( .A({ _15706_, _07699_, _15674_, _05066_ }), .Y(_15642_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29648_ ( .A({ _15707_, _07699_, _15675_, _05066_ }), .Y(_15643_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29649_ ( .A({ _15708_, _07699_, _15676_, _05066_ }), .Y(_15644_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29650_ ( .A({ _15709_, _07699_, _15677_, _05066_ }), .Y(_15645_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29651_ ( .A({ _15710_, _07699_, _15678_, _05066_ }), .Y(_15646_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29652_ ( .A({ _15711_, _07699_, _15679_, _05066_ }), .Y(_15647_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29653_ ( .A({ _15712_, _07699_, _15680_, _05066_ }), .Y(_15648_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29654_ ( .A({ _15713_, _07699_, _15681_, _05066_ }), .Y(_15649_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29655_ ( .A({ _15715_, _07699_, _15683_, _05066_ }), .Y(_15651_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29656_ ( .A({ _15716_, _07699_, _15684_, _05066_ }), .Y(_15652_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29657_ ( .A({ _17799_, _07122_, _17637_, _05102_ }), .Y(_17831_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29658_ ( .A({ _17776_, _07122_, _17614_, _05102_ }), .Y(_17808_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29659_ ( .A({ _17997_, _07122_, _17643_, _05102_ }), .Y(_18029_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29660_ ( .A({ _07705_, _07700_ }), .Y(matmul_15_dma_out_mask_0) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29661_ ( .A({ _07704_, _07703_, _07702_, _07701_ }), .Y(_07700_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29662_ ( .A(matmul_15_out_row_count[23:20]), .Y(_07701_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29663_ ( .A(matmul_15_out_row_count[19:16]), .Y(_07702_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29664_ ( .A(matmul_15_out_row_count[31:28]), .Y(_07703_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29665_ ( .A(matmul_15_out_row_count[27:24]), .Y(_07704_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29666_ ( .A({ _07709_, _07708_, _07707_, _07706_ }), .Y(_07705_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29667_ ( .A(matmul_15_out_row_count[7:4]), .Y(_07706_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29668_ ( .A(matmul_15_out_row_count[3:0]), .Y(_07707_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29669_ ( .A(matmul_15_out_row_count[15:12]), .Y(_07708_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29670_ ( .A(matmul_15_out_row_count[11:8]), .Y(_07709_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29671_ ( .A({ _07715_, _07710_ }), .Y(matmul_15_dma_pad_mask_0) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29672_ ( .A({ _07714_, _07713_, _07712_, _07711_ }), .Y(_07710_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29673_ ( .A(matmul_15_row_count[31:28]), .Y(_07711_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29674_ ( .A(matmul_15_row_count[27:24]), .Y(_07712_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29675_ ( .A(matmul_15_row_count[23:20]), .Y(_07713_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29676_ ( .A(matmul_15_row_count[19:16]), .Y(_07714_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29677_ ( .A({ _07719_, _07718_, _07717_, _07716_ }), .Y(_07715_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29678_ ( .A(matmul_15_row_count[7:4]), .Y(_07716_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29679_ ( .A(matmul_15_row_count[3:0]), .Y(_07717_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29680_ ( .A(matmul_15_row_count[15:12]), .Y(_07718_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29681_ ( .A(matmul_15_row_count[11:8]), .Y(_07719_) );
  \$lut  #( .LUT(16'h4dff), .WIDTH(4) ) _29682_ ( .A({ _07244_, cparam_max_pool_serial_9_act_num_col[4], max_pool_serial_9_row_count[4], _07720_ }), .Y(max_pool_serial_9_dma_pad_mask_0) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _29683_ ( .A({ cparam_max_pool_serial_9_act_num_col[3], max_pool_serial_9_row_count[3], _07721_ }), .Y(_07720_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _29684_ ( .A({ cparam_max_pool_serial_9_act_num_col[2], max_pool_serial_9_row_count[2], _07722_ }), .Y(_07721_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29685_ ( .A({ cparam_max_pool_serial_9_act_num_col[0], cparam_max_pool_serial_9_act_num_col[1], max_pool_serial_9_row_count[0], max_pool_serial_9_row_count[1] }), .Y(_07722_) );
  \$lut  #( .LUT(16'h2fff), .WIDTH(4) ) _29686_ ( .A({ _07726_, _07730_, _07723_, _07735_ }), .Y(max_pool_serial_9_dma_pad_mask_1) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _29687_ ( .A({ _07724_, cparam_max_pool_serial_9_act_num_col[3], _03571_ }), .Y(_07723_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _29688_ ( .A({ _03568_, cparam_max_pool_serial_9_act_num_col[2], _07725_ }), .Y(_07724_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _29689_ ( .A({ cparam_max_pool_serial_9_act_num_col[0], _03546_, _03557_, cparam_max_pool_serial_9_act_num_col[1] }), .Y(_07725_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _29690_ ( .A({ _07729_, _07727_, _03576_, _03573_ }), .Y(_07726_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29691_ ( .A({ _07728_, _03569_, _03565_, _03564_ }), .Y(_07727_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29692_ ( .A({ _03561_, _03560_, _03558_, _03554_ }), .Y(_07728_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29693_ ( .A({ _03552_, _03551_, _03549_, _03577_ }), .Y(_07729_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29694_ ( .A({ _07734_, _07733_, _07732_, _07731_ }), .Y(_07730_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29695_ ( .A({ _03562_, _03559_, _03556_, _03555_ }), .Y(_07731_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29696_ ( .A({ _03570_, _03567_, _03566_, _03563_ }), .Y(_07732_) );
  \$lut  #( .LUT(16'h000d), .WIDTH(4) ) _29697_ ( .A({ _03575_, _03574_, cparam_max_pool_serial_9_act_num_col[4], _03572_ }), .Y(_07733_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29698_ ( .A({ _03553_, _03550_, _03548_, _03547_ }), .Y(_07734_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _29699_ ( .A({ cparam_max_pool_serial_9_act_num_col[3], _03571_, cparam_max_pool_serial_9_act_num_col[4], _03572_ }), .Y(_07735_) );
  \$lut  #( .LUT(16'hf4ff), .WIDTH(4) ) _29700_ ( .A({ _07741_, _07736_, conv2d_8_out_row_count[4], cparam_conv2d_8_inc_sync_out[4] }), .Y(conv2d_8_dma_out_mask_0) );
  \$lut  #( .LUT(16'h000d), .WIDTH(4) ) _29701_ ( .A({ _07740_, _07737_, conv2d_8_out_row_count[4], cparam_conv2d_8_inc_sync_out[4] }), .Y(_07736_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _29702_ ( .A({ _07739_, cparam_conv2d_8_inc_sync_out[1], conv2d_8_out_row_count[1], _07738_ }), .Y(_07737_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29703_ ( .A({ cparam_conv2d_8_inc_sync_out[0], conv2d_8_out_row_count[0] }), .Y(_07738_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _29704_ ( .A({ cparam_conv2d_8_inc_sync_out[3], conv2d_8_out_row_count[3], cparam_conv2d_8_inc_sync_out[2], conv2d_8_out_row_count[2] }), .Y(_07739_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _29705_ ( .A({ cparam_conv2d_8_inc_sync_out[2], cparam_conv2d_8_inc_sync_out[3], conv2d_8_out_row_count[2], conv2d_8_out_row_count[3] }), .Y(_07740_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29706_ ( .A({ _07749_, _07748_, _07744_, _07742_ }), .Y(_07741_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29707_ ( .A({ _07743_, conv2d_8_out_row_count[31:29] }), .Y(_07742_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29708_ ( .A({ conv2d_8_out_row_count[27:26], conv2d_8_out_row_count[24], conv2d_8_out_row_count[21] }), .Y(_07743_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29709_ ( .A({ _07747_, _07746_, _07745_ }), .Y(_07744_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29710_ ( .A({ conv2d_8_out_row_count[28], conv2d_8_out_row_count[25], conv2d_8_out_row_count[23:22] }), .Y(_07745_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29711_ ( .A({ conv2d_8_out_row_count[12], conv2d_8_out_row_count[9], conv2d_8_out_row_count[7:6] }), .Y(_07746_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29712_ ( .A({ conv2d_8_out_row_count[19:18], conv2d_8_out_row_count[16], conv2d_8_out_row_count[13] }), .Y(_07747_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29713_ ( .A({ conv2d_8_out_row_count[11:10], conv2d_8_out_row_count[8], conv2d_8_out_row_count[5] }), .Y(_07748_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29714_ ( .A({ conv2d_8_out_row_count[20], conv2d_8_out_row_count[17], conv2d_8_out_row_count[15:14] }), .Y(_07749_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29715_ ( .A({ _18159_, _07122_, cparam_conv2d_8_col_select_initval[0], _05102_ }), .Y(_18161_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29716_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17292_, _17324_ }), .Y(_17260_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29717_ ( .A({ _07751_, _07759_, _stream_conv2d_8_source_6_source_pat_fsm_0[1] }), .Y(_07750_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29718_ ( .A({ _07758_, _07757_, _07752_ }), .Y(_07751_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29719_ ( .A({ _07756_, _07755_, _07754_, _07753_ }), .Y(_07752_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29720_ ( .A(_stream_conv2d_8_source_6_source_pat_fsm_0[23:20]), .Y(_07753_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29721_ ( .A(_stream_conv2d_8_source_6_source_pat_fsm_0[19:16]), .Y(_07754_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29722_ ( .A(_stream_conv2d_8_source_6_source_pat_fsm_0[31:28]), .Y(_07755_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29723_ ( .A(_stream_conv2d_8_source_6_source_pat_fsm_0[27:24]), .Y(_07756_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29724_ ( .A(_stream_conv2d_8_source_6_source_pat_fsm_0[15:12]), .Y(_07757_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29725_ ( .A(_stream_conv2d_8_source_6_source_pat_fsm_0[11:8]), .Y(_07758_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29726_ ( .A({ _07760_, _stream_conv2d_8_source_6_source_pat_fsm_0[3:2] }), .Y(_07759_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29727_ ( .A(_stream_conv2d_8_source_6_source_pat_fsm_0[7:4]), .Y(_07760_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29728_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16729_, _16761_ }), .Y(_16697_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29729_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16257_, _16289_ }), .Y(_16225_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29730_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16151_, _16183_ }), .Y(_16119_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29731_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16058_, _16090_ }), .Y(_16026_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29732_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16727_, _16759_ }), .Y(_16695_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29733_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16256_, _16288_ }), .Y(_16224_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29734_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16255_, _16287_ }), .Y(_16223_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29735_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16140_, _16172_ }), .Y(_16108_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29736_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16254_, _16286_ }), .Y(_16222_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29737_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16252_, _16284_ }), .Y(_16220_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29738_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16452_, _16484_ }), .Y(_16420_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29739_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16248_, _16280_ }), .Y(_16216_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29740_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16447_, _16479_ }), .Y(_16415_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29741_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16244_, _16276_ }), .Y(_16212_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29742_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16057_, _16089_ }), .Y(_16025_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29743_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16444_, _16476_ }), .Y(_16412_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29744_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16241_, _16273_ }), .Y(_16209_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29745_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16056_, _16088_ }), .Y(_16024_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29746_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16435_, _16467_ }), .Y(_16403_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29747_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16434_, _16466_ }), .Y(_16402_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29748_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16264_, _16296_ }), .Y(_16232_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29749_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16433_, _16465_ }), .Y(_16401_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29750_ ( .A({ _17795_, _07122_, _17633_, _05102_ }), .Y(_17827_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29751_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16432_, _16464_ }), .Y(_16400_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29752_ ( .A({ _17789_, _07122_, _17627_, _05102_ }), .Y(_17821_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29753_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16431_, _16463_ }), .Y(_16399_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29754_ ( .A({ _17782_, _07122_, _17620_, _05102_ }), .Y(_17814_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29755_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17219_, _17251_ }), .Y(_17187_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29756_ ( .A({ _07762_, _07770_, _stream_conv2d_8_source_8_source_pat_fsm_1[1] }), .Y(_07761_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29757_ ( .A({ _07769_, _07768_, _07763_ }), .Y(_07762_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29758_ ( .A({ _07767_, _07766_, _07765_, _07764_ }), .Y(_07763_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29759_ ( .A(_stream_conv2d_8_source_8_source_pat_fsm_1[23:20]), .Y(_07764_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29760_ ( .A(_stream_conv2d_8_source_8_source_pat_fsm_1[19:16]), .Y(_07765_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29761_ ( .A(_stream_conv2d_8_source_8_source_pat_fsm_1[31:28]), .Y(_07766_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29762_ ( .A(_stream_conv2d_8_source_8_source_pat_fsm_1[27:24]), .Y(_07767_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29763_ ( .A(_stream_conv2d_8_source_8_source_pat_fsm_1[15:12]), .Y(_07768_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29764_ ( .A(_stream_conv2d_8_source_8_source_pat_fsm_1[11:8]), .Y(_07769_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29765_ ( .A({ _07771_, _stream_conv2d_8_source_8_source_pat_fsm_1[3:2] }), .Y(_07770_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29766_ ( .A(_stream_conv2d_8_source_8_source_pat_fsm_1[7:4]), .Y(_07771_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29767_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16430_, _16462_ }), .Y(_16398_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29768_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16263_, _16295_ }), .Y(_16231_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29769_ ( .A({ _17806_, _07122_, _17644_, _05102_ }), .Y(_17838_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29770_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17213_, _17245_ }), .Y(_17181_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29771_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16429_, _16461_ }), .Y(_16397_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29772_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16262_, _16294_ }), .Y(_16230_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29773_ ( .A({ _17800_, _07122_, _17638_, _05102_ }), .Y(_17832_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29774_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17206_, _17238_ }), .Y(_17174_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29775_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16459_, _16491_ }), .Y(_16427_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29776_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16261_, _16293_ }), .Y(_16229_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29777_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17202_, _17234_ }), .Y(_17170_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29778_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16457_, _16489_ }), .Y(_16425_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29779_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16236_, _16268_ }), .Y(_16204_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29780_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16051_, _16083_ }), .Y(_16019_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29781_ ( .A({ _16005_, _07334_, _15973_, _05071_ }), .Y(_15941_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29782_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17198_, _17230_ }), .Y(_17166_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29783_ ( .A({ _05076_, _07441_ }), .Y(_21909_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29784_ ( .A({ _stream_conv2d_8_source_28_source_pat_fsm_11[1], _07442_, _07450_, _stream_conv2d_8_source_28_source_pat_fsm_11[0] }), .Y(_05076_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29785_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16050_, _16082_ }), .Y(_16018_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29786_ ( .A({ _15991_, _07334_, _15959_, _05071_ }), .Y(_15927_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29787_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17225_, _17257_ }), .Y(_17193_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29788_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16049_, _16081_ }), .Y(_16017_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29789_ ( .A({ _15980_, _07334_, _15948_, _05071_ }), .Y(_15916_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29790_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17207_, _17239_ }), .Y(_17175_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29791_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16047_, _16079_ }), .Y(_16015_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29792_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17316_, _17348_ }), .Y(_17284_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29793_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17315_, _17347_ }), .Y(_17283_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29794_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17313_, _17345_ }), .Y(_17281_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29795_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17312_, _17344_ }), .Y(_17280_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29796_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17311_, _17343_ }), .Y(_17279_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29797_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17310_, _17342_ }), .Y(_17278_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29798_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17309_, _17341_ }), .Y(_17277_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29799_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17308_, _17340_ }), .Y(_17276_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29800_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17307_, _17339_ }), .Y(_17275_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29801_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17306_, _17338_ }), .Y(_17274_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29802_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17305_, _17337_ }), .Y(_17273_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29803_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17304_, _17336_ }), .Y(_17272_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29804_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17302_, _17334_ }), .Y(_17270_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29805_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17301_, _17333_ }), .Y(_17269_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29806_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17300_, _17332_ }), .Y(_17268_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29807_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17299_, _17331_ }), .Y(_17267_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29808_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17298_, _17330_ }), .Y(_17266_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29809_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17297_, _17329_ }), .Y(_17265_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29810_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17296_, _17328_ }), .Y(_17264_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29811_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17295_, _17327_ }), .Y(_17263_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29812_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17294_, _17326_ }), .Y(_17262_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29813_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17293_, _17325_ }), .Y(_17261_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29814_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17323_, _17355_ }), .Y(_17291_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29815_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17322_, _17354_ }), .Y(_17290_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29816_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17321_, _17353_ }), .Y(_17289_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29817_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17320_, _17352_ }), .Y(_17288_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29818_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17319_, _17351_ }), .Y(_17287_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29819_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17318_, _17350_ }), .Y(_17286_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29820_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17317_, _17349_ }), .Y(_17285_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29821_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17314_, _17346_ }), .Y(_17282_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29822_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16731_, _16763_ }), .Y(_16699_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29823_ ( .A({ _07750_, _stream_conv2d_8_source_6_source_pat_fsm_0[0], _17303_, _17335_ }), .Y(_17271_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29824_ ( .A({ _05088_, _07369_ }), .Y(_21915_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29825_ ( .A({ _stream_conv2d_8_source_22_source_pat_fsm_5[1], _07370_, _07378_, _stream_conv2d_8_source_22_source_pat_fsm_5[0] }), .Y(_05088_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29826_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16730_, _16762_ }), .Y(_16698_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29827_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16259_, _16291_ }), .Y(_16227_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29828_ ( .A({ _07148_, _stream_conv2d_8_source_29_source_pat_fsm_12[0], _16162_, _16194_ }), .Y(_16130_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29829_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16059_, _16091_ }), .Y(_16027_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29830_ ( .A({ _16006_, _07334_, _15974_, _05071_ }), .Y(_15942_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29831_ ( .A({ _15985_, _07334_, _15953_, _05071_ }), .Y(_15921_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29832_ ( .A({ _15996_, _07334_, _15964_, _05071_ }), .Y(_15932_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29833_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16728_, _16760_ }), .Y(_16696_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29834_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16726_, _16758_ }), .Y(_16694_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29835_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16725_, _16757_ }), .Y(_16693_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29836_ ( .A({ _05098_, _07750_ }), .Y(_21920_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29837_ ( .A({ _stream_conv2d_8_source_6_source_pat_fsm_0[1], _07751_, _07759_, _stream_conv2d_8_source_6_source_pat_fsm_0[0] }), .Y(_05098_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29838_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16724_, _16756_ }), .Y(_16692_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29839_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16723_, _16755_ }), .Y(_16691_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29840_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16722_, _16754_ }), .Y(_16690_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29841_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16721_, _16753_ }), .Y(_16689_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29842_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16720_, _16752_ }), .Y(_16688_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29843_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16719_, _16751_ }), .Y(_16687_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29844_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16718_, _16750_ }), .Y(_16686_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29845_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16717_, _16749_ }), .Y(_16685_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29846_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16747_, _16779_ }), .Y(_16715_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29847_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16746_, _16778_ }), .Y(_16714_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29848_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16745_, _16777_ }), .Y(_16713_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29849_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16744_, _16776_ }), .Y(_16712_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29850_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16743_, _16775_ }), .Y(_16711_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29851_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16742_, _16774_ }), .Y(_16710_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29852_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16738_, _16770_ }), .Y(_16706_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29853_ ( .A({ _07402_, _stream_conv2d_8_source_23_source_pat_fsm_6[0], _16716_, _16748_ }), .Y(_16684_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29854_ ( .A({ _05086_, _07402_ }), .Y(_21914_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29855_ ( .A({ _stream_conv2d_8_source_23_source_pat_fsm_6[1], _07403_, _07411_, _stream_conv2d_8_source_23_source_pat_fsm_6[0] }), .Y(_05086_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29856_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16253_, _16285_ }), .Y(_16221_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29857_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16251_, _16283_ }), .Y(_16219_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29858_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16250_, _16282_ }), .Y(_16218_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29859_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16451_, _16483_ }), .Y(_16419_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29860_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16249_, _16281_ }), .Y(_16217_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29861_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16449_, _16481_ }), .Y(_16417_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29862_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16246_, _16278_ }), .Y(_16214_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29863_ ( .A({ _05074_, _07148_ }), .Y(_21908_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29864_ ( .A({ _stream_conv2d_8_source_29_source_pat_fsm_12[1], _07149_, _07157_, _stream_conv2d_8_source_29_source_pat_fsm_12[0] }), .Y(_05074_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29865_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16448_, _16480_ }), .Y(_16416_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29866_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16245_, _16277_ }), .Y(_16213_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29867_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16446_, _16478_ }), .Y(_16414_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29868_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16243_, _16275_ }), .Y(_16211_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29869_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16445_, _16477_ }), .Y(_16413_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29870_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16242_, _16274_ }), .Y(_16210_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29871_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16443_, _16475_ }), .Y(_16411_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29872_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16240_, _16272_ }), .Y(_16208_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29873_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16442_, _16474_ }), .Y(_16410_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29874_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16239_, _16271_ }), .Y(_16207_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29875_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16054_, _16086_ }), .Y(_16022_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29876_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16441_, _16473_ }), .Y(_16409_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29877_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16238_, _16270_ }), .Y(_16206_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29878_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16440_, _16472_ }), .Y(_16408_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29879_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16237_, _16269_ }), .Y(_16205_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29880_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16438_, _16470_ }), .Y(_16406_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29881_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16267_, _16299_ }), .Y(_16235_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29882_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16437_, _16469_ }), .Y(_16405_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29883_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16266_, _16298_ }), .Y(_16234_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29884_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16053_, _16085_ }), .Y(_16021_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29885_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16436_, _16468_ }), .Y(_16404_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29886_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16265_, _16297_ }), .Y(_16233_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29887_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16052_, _16084_ }), .Y(_16020_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29888_ ( .A({ _17798_, _07122_, _17636_, _05102_ }), .Y(_17830_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29889_ ( .A({ _17796_, _07122_, _17634_, _05102_ }), .Y(_17828_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29890_ ( .A({ _17794_, _07122_, _17632_, _05102_ }), .Y(_17826_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29891_ ( .A({ _17793_, _07122_, _17631_, _05102_ }), .Y(_17825_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29892_ ( .A({ _17792_, _07122_, _17630_, _05102_ }), .Y(_17824_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29893_ ( .A({ _17791_, _07122_, _17629_, _05102_ }), .Y(_17823_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29894_ ( .A({ _17790_, _07122_, _17628_, _05102_ }), .Y(_17822_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29895_ ( .A({ _17788_, _07122_, _17626_, _05102_ }), .Y(_17820_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29896_ ( .A({ _17787_, _07122_, _17625_, _05102_ }), .Y(_17819_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29897_ ( .A({ _17785_, _07122_, _17623_, _05102_ }), .Y(_17817_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29898_ ( .A({ _17784_, _07122_, _17622_, _05102_ }), .Y(_17816_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29899_ ( .A({ _17783_, _07122_, _17621_, _05102_ }), .Y(_17815_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29900_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17220_, _17252_ }), .Y(_17188_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29901_ ( .A({ _17781_, _07122_, _17619_, _05102_ }), .Y(_17813_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29902_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17217_, _17249_ }), .Y(_17185_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29903_ ( .A({ _17779_, _07122_, _17617_, _05102_ }), .Y(_17811_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29904_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17216_, _17248_ }), .Y(_17184_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29905_ ( .A({ _17778_, _07122_, _17616_, _05102_ }), .Y(_17810_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29906_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17215_, _17247_ }), .Y(_17183_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29907_ ( .A({ _17777_, _07122_, _17615_, _05102_ }), .Y(_17809_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29908_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17214_, _17246_ }), .Y(_17182_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29909_ ( .A({ _17805_, _07122_, _17643_, _05102_ }), .Y(_17837_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29910_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17212_, _17244_ }), .Y(_17180_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29911_ ( .A({ _17804_, _07122_, _17642_, _05102_ }), .Y(_17836_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29912_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17211_, _17243_ }), .Y(_17179_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29913_ ( .A({ _17802_, _07122_, _17640_, _05102_ }), .Y(_17834_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29914_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17210_, _17242_ }), .Y(_17178_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29915_ ( .A({ _17801_, _07122_, _17639_, _05102_ }), .Y(_17833_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29916_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17209_, _17241_ }), .Y(_17177_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29917_ ( .A({ _17797_, _07122_, _17635_, _05102_ }), .Y(_17829_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29918_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17208_, _17240_ }), .Y(_17176_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29919_ ( .A({ _17786_, _07122_, _17624_, _05102_ }), .Y(_17818_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29920_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17205_, _17237_ }), .Y(_17173_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29921_ ( .A({ _17775_, _07122_, _17613_, _05102_ }), .Y(_17807_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29922_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17204_, _17236_ }), .Y(_17172_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29923_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17203_, _17235_ }), .Y(_17171_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29924_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16458_, _16490_ }), .Y(_16426_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29925_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16258_, _16290_ }), .Y(_16226_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29926_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17201_, _17233_ }), .Y(_17169_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29927_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16456_, _16488_ }), .Y(_16424_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29928_ ( .A({ _07441_, _stream_conv2d_8_source_28_source_pat_fsm_11[0], _16247_, _16279_ }), .Y(_16215_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29929_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17200_, _17232_ }), .Y(_17168_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29930_ ( .A({ _06555_, _stream_conv2d_8_source_26_source_pat_fsm_9[0], _16453_, _16485_ }), .Y(_16421_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29931_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17199_, _17231_ }), .Y(_17167_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29932_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17197_, _17229_ }), .Y(_17165_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29933_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17227_, _17259_ }), .Y(_17195_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29934_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17226_, _17258_ }), .Y(_17194_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29935_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17224_, _17256_ }), .Y(_17192_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29936_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17223_, _17255_ }), .Y(_17191_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29937_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17222_, _17254_ }), .Y(_17190_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29938_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17221_, _17253_ }), .Y(_17189_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29939_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17218_, _17250_ }), .Y(_17186_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29940_ ( .A({ _07761_, _stream_conv2d_8_source_8_source_pat_fsm_1[0], _17196_, _17228_ }), .Y(_17164_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29941_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16048_, _16080_ }), .Y(_16016_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29942_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16046_, _16078_ }), .Y(_16014_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29943_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16045_, _16077_ }), .Y(_16013_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29944_ ( .A({ _05096_, _07761_ }), .Y(_21919_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29945_ ( .A({ _stream_conv2d_8_source_8_source_pat_fsm_1[1], _07762_, _07770_, _stream_conv2d_8_source_8_source_pat_fsm_1[0] }), .Y(_05096_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29946_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16075_, _16107_ }), .Y(_16043_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29947_ ( .A({ _15983_, _07334_, _15951_, _05071_ }), .Y(_15919_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29948_ ( .A({ _15994_, _07334_, _15962_, _05071_ }), .Y(_15930_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29949_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16074_, _16106_ }), .Y(_16042_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29950_ ( .A({ _15982_, _07334_, _15950_, _05071_ }), .Y(_15918_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29951_ ( .A({ _15993_, _07334_, _15961_, _05071_ }), .Y(_15929_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29952_ ( .A({ _16004_, _07334_, _15972_, _05071_ }), .Y(_15940_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29953_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16073_, _16105_ }), .Y(_16041_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29954_ ( .A({ _15981_, _07334_, _15949_, _05071_ }), .Y(_15917_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29955_ ( .A({ _15992_, _07334_, _15960_, _05071_ }), .Y(_15928_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29956_ ( .A({ _16003_, _07334_, _15971_, _05071_ }), .Y(_15939_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29957_ ( .A({ _07032_, _stream_conv2d_8_source_30_source_pat_fsm_13[0], _16072_, _16104_ }), .Y(_16040_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29958_ ( .A({ _16011_, _07334_, _15979_, _05071_ }), .Y(_15947_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29959_ ( .A({ _15990_, _07334_, _15958_, _05071_ }), .Y(_15926_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29960_ ( .A({ _16001_, _07334_, _15969_, _05071_ }), .Y(_15937_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29961_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17123_, _17155_ }), .Y(_17091_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29962_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17121_, _17153_ }), .Y(_17089_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29963_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17120_, _17152_ }), .Y(_17088_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29964_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17119_, _17151_ }), .Y(_17087_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29965_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17118_, _17150_ }), .Y(_17086_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29966_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17117_, _17149_ }), .Y(_17085_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29967_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17116_, _17148_ }), .Y(_17084_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29968_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17115_, _17147_ }), .Y(_17083_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29969_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17114_, _17146_ }), .Y(_17082_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29970_ ( .A({ _05064_, _07772_ }), .Y(_21902_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29971_ ( .A({ _07773_, _07778_, _stream_conv2d_8_source_35_source_pat_fsm_18[0] }), .Y(_07772_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29972_ ( .A({ _07777_, _07776_, _07774_ }), .Y(_07773_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29973_ ( .A({ _07775_, _stream_conv2d_8_source_35_source_pat_fsm_18[3:2] }), .Y(_07774_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29974_ ( .A(_stream_conv2d_8_source_35_source_pat_fsm_18[7:4]), .Y(_07775_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29975_ ( .A(_stream_conv2d_8_source_35_source_pat_fsm_18[15:12]), .Y(_07776_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29976_ ( .A(_stream_conv2d_8_source_35_source_pat_fsm_18[11:8]), .Y(_07777_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29977_ ( .A({ _07782_, _07781_, _07780_, _07779_ }), .Y(_07778_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29978_ ( .A(_stream_conv2d_8_source_35_source_pat_fsm_18[23:20]), .Y(_07779_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29979_ ( .A(_stream_conv2d_8_source_35_source_pat_fsm_18[19:16]), .Y(_07780_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29980_ ( .A(_stream_conv2d_8_source_35_source_pat_fsm_18[31:28]), .Y(_07781_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29981_ ( .A(_stream_conv2d_8_source_35_source_pat_fsm_18[27:24]), .Y(_07782_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29982_ ( .A({ _07773_, _stream_conv2d_8_source_35_source_pat_fsm_18[0], _07778_, _stream_conv2d_8_source_35_source_pat_fsm_18[1] }), .Y(_05064_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29983_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17113_, _17145_ }), .Y(_17081_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29984_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17112_, _17144_ }), .Y(_17080_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29985_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17110_, _17142_ }), .Y(_17078_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29986_ ( .A({ _07056_, _stream_conv2d_8_source_19_source_pat_fsm_2[0], _17109_, _17141_ }), .Y(_17077_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29987_ ( .A({ _15596_, _07783_, _15564_, _05064_ }), .Y(_15532_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29988_ ( .A({ _07772_, _stream_conv2d_8_source_35_source_pat_fsm_18[1] }), .Y(_07783_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29989_ ( .A({ _15607_, _07783_, _15575_, _05064_ }), .Y(_15543_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29990_ ( .A({ _15618_, _07783_, _15586_, _05064_ }), .Y(_15554_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29991_ ( .A({ _15621_, _07783_, _15589_, _05064_ }), .Y(_15557_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29992_ ( .A({ _15622_, _07783_, _15590_, _05064_ }), .Y(_15558_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29993_ ( .A({ _15623_, _07783_, _15591_, _05064_ }), .Y(_15559_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29994_ ( .A({ _15624_, _07783_, _15592_, _05064_ }), .Y(_15560_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29995_ ( .A({ _15625_, _07783_, _15593_, _05064_ }), .Y(_15561_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29996_ ( .A({ _15626_, _07783_, _15594_, _05064_ }), .Y(_15562_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29997_ ( .A({ _15627_, _07783_, _15595_, _05064_ }), .Y(_15563_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29998_ ( .A({ _15597_, _07783_, _15565_, _05064_ }), .Y(_15533_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29999_ ( .A({ _15598_, _07783_, _15566_, _05064_ }), .Y(_15534_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30000_ ( .A({ _15599_, _07783_, _15567_, _05064_ }), .Y(_15535_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30001_ ( .A({ _15600_, _07783_, _15568_, _05064_ }), .Y(_15536_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30002_ ( .A({ _15601_, _07783_, _15569_, _05064_ }), .Y(_15537_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30003_ ( .A({ _15602_, _07783_, _15570_, _05064_ }), .Y(_15538_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30004_ ( .A({ _15603_, _07783_, _15571_, _05064_ }), .Y(_15539_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30005_ ( .A({ _15604_, _07783_, _15572_, _05064_ }), .Y(_15540_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30006_ ( .A({ _15605_, _07783_, _15573_, _05064_ }), .Y(_15541_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30007_ ( .A({ _15606_, _07783_, _15574_, _05064_ }), .Y(_15542_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30008_ ( .A({ _15608_, _07783_, _15576_, _05064_ }), .Y(_15544_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30009_ ( .A({ _15609_, _07783_, _15577_, _05064_ }), .Y(_15545_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30010_ ( .A({ _15610_, _07783_, _15578_, _05064_ }), .Y(_15546_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30011_ ( .A({ _15611_, _07783_, _15579_, _05064_ }), .Y(_15547_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30012_ ( .A({ _15612_, _07783_, _15580_, _05064_ }), .Y(_15548_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30013_ ( .A({ _18251_, _05107_, _18317_, _07019_ }), .Y(_18284_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30014_ ( .A({ _15613_, _07783_, _15581_, _05064_ }), .Y(_15549_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30015_ ( .A({ _18250_, _05107_, _18316_, _07019_ }), .Y(_18283_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30016_ ( .A({ _18248_, _05107_, _18314_, _07019_ }), .Y(_18281_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30017_ ( .A({ _18246_, _05107_, _18312_, _07019_ }), .Y(_18279_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30018_ ( .A({ _15614_, _07783_, _15582_, _05064_ }), .Y(_15550_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30019_ ( .A({ _18245_, _05107_, _18311_, _07019_ }), .Y(_18278_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30020_ ( .A({ _18244_, _05107_, _18310_, _07019_ }), .Y(_18277_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30021_ ( .A({ _18242_, _05107_, _18308_, _07019_ }), .Y(_18275_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30022_ ( .A({ _15615_, _07783_, _15583_, _05064_ }), .Y(_15551_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30023_ ( .A({ _18241_, _05107_, _18307_, _07019_ }), .Y(_18274_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30024_ ( .A({ _18240_, _05107_, _18306_, _07019_ }), .Y(_18273_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30025_ ( .A({ _18239_, _05107_, _18305_, _07019_ }), .Y(_18272_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30026_ ( .A({ _15616_, _07783_, _15584_, _05064_ }), .Y(_15552_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30027_ ( .A({ _18237_, _05107_, _18303_, _07019_ }), .Y(_18270_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30028_ ( .A({ _15617_, _07783_, _15585_, _05064_ }), .Y(_15553_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30029_ ( .A({ _18236_, _05107_, _18302_, _07019_ }), .Y(_18269_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30030_ ( .A({ _18235_, _05107_, _18301_, _07019_ }), .Y(_18268_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30031_ ( .A({ _15619_, _07783_, _15587_, _05064_ }), .Y(_15555_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30032_ ( .A({ _18234_, _05107_, _18300_, _07019_ }), .Y(_18267_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30033_ ( .A({ _18233_, _05107_, _18299_, _07019_ }), .Y(_18266_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30034_ ( .A({ _18231_, _05107_, _18297_, _07019_ }), .Y(_18264_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30035_ ( .A({ _18230_, _05107_, _18296_, _07019_ }), .Y(_18263_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30036_ ( .A({ _15620_, _07783_, _15588_, _05064_ }), .Y(_15556_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30037_ ( .A({ _18229_, _05107_, _18295_, _07019_ }), .Y(_18262_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30038_ ( .A({ _18228_, _05107_, _18294_, _07019_ }), .Y(_18261_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30039_ ( .A({ _18256_, _05107_, _18322_, _07019_ }), .Y(_18289_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30040_ ( .A({ _18255_, _05107_, _18321_, _07019_ }), .Y(_18288_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30041_ ( .A({ _18254_, _05107_, _18320_, _07019_ }), .Y(_18287_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30042_ ( .A({ _18253_, _05107_, _18319_, _07019_ }), .Y(_18286_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30043_ ( .A({ _18252_, _05107_, _18318_, _07019_ }), .Y(_18285_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30044_ ( .A({ _18247_, _05107_, _18313_, _07019_ }), .Y(_18280_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30045_ ( .A({ _18243_, _05107_, _18309_, _07019_ }), .Y(_18276_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30046_ ( .A({ _18259_, _05107_, _18325_, _07019_ }), .Y(_18292_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30047_ ( .A({ _18249_, _05107_, _18315_, _07019_ }), .Y(_18282_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30048_ ( .A({ _18238_, _05107_, _18304_, _07019_ }), .Y(_18271_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30049_ ( .A({ _18257_, _05107_, _18323_, _07019_ }), .Y(_18290_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30050_ ( .A({ _18258_, _05107_, _18324_, _07019_ }), .Y(_18291_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30051_ ( .A({ _18232_, _05107_, _18298_, _07019_ }), .Y(_18265_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30052_ ( .A({ _05061_, _07784_ }), .Y(_21901_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30053_ ( .A({ _07785_, _07790_, _stream_conv2d_8_source_36_source_pat_fsm_19[0] }), .Y(_07784_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30054_ ( .A({ _07789_, _07788_, _07786_ }), .Y(_07785_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30055_ ( .A({ _07787_, _stream_conv2d_8_source_36_source_pat_fsm_19[3:2] }), .Y(_07786_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30056_ ( .A(_stream_conv2d_8_source_36_source_pat_fsm_19[7:4]), .Y(_07787_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30057_ ( .A(_stream_conv2d_8_source_36_source_pat_fsm_19[15:12]), .Y(_07788_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30058_ ( .A(_stream_conv2d_8_source_36_source_pat_fsm_19[11:8]), .Y(_07789_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30059_ ( .A({ _07794_, _07793_, _07792_, _07791_ }), .Y(_07790_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30060_ ( .A(_stream_conv2d_8_source_36_source_pat_fsm_19[23:20]), .Y(_07791_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30061_ ( .A(_stream_conv2d_8_source_36_source_pat_fsm_19[19:16]), .Y(_07792_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30062_ ( .A(_stream_conv2d_8_source_36_source_pat_fsm_19[31:28]), .Y(_07793_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30063_ ( .A(_stream_conv2d_8_source_36_source_pat_fsm_19[27:24]), .Y(_07794_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _30064_ ( .A({ _07785_, _stream_conv2d_8_source_36_source_pat_fsm_19[0], _07790_, _stream_conv2d_8_source_36_source_pat_fsm_19[1] }), .Y(_05061_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30065_ ( .A({ _15500_, _07795_, _15468_, _05061_ }), .Y(_15436_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30066_ ( .A({ _07784_, _stream_conv2d_8_source_36_source_pat_fsm_19[1] }), .Y(_07795_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30067_ ( .A({ _15511_, _07795_, _15479_, _05061_ }), .Y(_15447_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30068_ ( .A({ _15522_, _07795_, _15490_, _05061_ }), .Y(_15458_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30069_ ( .A({ _15525_, _07795_, _15493_, _05061_ }), .Y(_15461_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30070_ ( .A({ _17803_, _07122_, _17641_, _05102_ }), .Y(_17835_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30071_ ( .A({ _15526_, _07795_, _15494_, _05061_ }), .Y(_15462_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30072_ ( .A({ _15527_, _07795_, _15495_, _05061_ }), .Y(_15463_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30073_ ( .A({ _17780_, _07122_, _17618_, _05102_ }), .Y(_17812_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30074_ ( .A({ _15528_, _07795_, _15496_, _05061_ }), .Y(_15464_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30075_ ( .A({ _15529_, _07795_, _15497_, _05061_ }), .Y(_15465_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30076_ ( .A({ _15530_, _07795_, _15498_, _05061_ }), .Y(_15466_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30077_ ( .A({ _15531_, _07795_, _15499_, _05061_ }), .Y(_15467_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30078_ ( .A({ _15501_, _07795_, _15469_, _05061_ }), .Y(_15437_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30079_ ( .A({ _15502_, _07795_, _15470_, _05061_ }), .Y(_15438_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30080_ ( .A({ _15503_, _07795_, _15471_, _05061_ }), .Y(_15439_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30081_ ( .A({ _15504_, _07795_, _15472_, _05061_ }), .Y(_15440_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30082_ ( .A({ _15505_, _07795_, _15473_, _05061_ }), .Y(_15441_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30083_ ( .A({ _18160_, _07122_, cparam_conv2d_8_col_select_initval[1], _05102_ }), .Y(_18162_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30084_ ( .A({ _15506_, _07795_, _15474_, _05061_ }), .Y(_15442_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _30085_ ( .A({ _15507_, _07795_, _15475_, _05061_ }), .Y(_15443_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30086_ ( .A({ _03762_, _07796_, _07809_, _saxi_register_10[31] }), .Y(_20962_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30087_ ( .A({ _07807_, _07797_ }), .Y(_07796_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30088_ ( .A({ _07798_, _07802_, main_fsm[4] }), .Y(_07797_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30089_ ( .A({ main_fsm[5], _07801_, _07800_, _07799_ }), .Y(_07798_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30090_ ( .A(main_fsm[15:12]), .Y(_07799_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _30091_ ( .A(main_fsm[7:6]), .Y(_07800_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30092_ ( .A(main_fsm[11:8]), .Y(_07801_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30093_ ( .A({ _07806_, _07805_, _07804_, _07803_ }), .Y(_07802_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30094_ ( .A(main_fsm[23:20]), .Y(_07803_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30095_ ( .A(main_fsm[19:16]), .Y(_07804_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30096_ ( .A(main_fsm[31:28]), .Y(_07805_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30097_ ( .A(main_fsm[27:24]), .Y(_07806_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30098_ ( .A({ main_fsm[0], _07808_, main_fsm[1] }), .Y(_07807_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _30099_ ( .A({ main_fsm[2], main_fsm[3] }), .Y(_07808_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30100_ ( .A({ _07812_, _07810_ }), .Y(_07809_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30101_ ( .A({ main_fsm[4], _07811_, _07802_ }), .Y(_07810_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30102_ ( .A({ _07799_, _07801_, _07800_, main_fsm[5] }), .Y(_07811_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30103_ ( .A({ _07808_, main_fsm[0], main_fsm[1] }), .Y(_07812_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30104_ ( .A({ _03761_, _07796_, _07809_, _saxi_register_10[30] }), .Y(_20961_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30105_ ( .A({ _03759_, _07796_, _07809_, _saxi_register_10[29] }), .Y(_20959_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30106_ ( .A({ _03758_, _07796_, _07809_, _saxi_register_10[28] }), .Y(_20958_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30107_ ( .A({ _03757_, _07796_, _07809_, _saxi_register_10[27] }), .Y(_20957_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30108_ ( .A({ _03756_, _07796_, _07809_, _saxi_register_10[26] }), .Y(_20956_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30109_ ( .A({ _03755_, _07796_, _07809_, _saxi_register_10[25] }), .Y(_20955_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30110_ ( .A({ _03754_, _07796_, _07809_, _saxi_register_10[24] }), .Y(_20954_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30111_ ( .A({ _03753_, _07796_, _07809_, _saxi_register_10[23] }), .Y(_20953_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30112_ ( .A({ _03752_, _07796_, _07809_, _saxi_register_10[22] }), .Y(_20952_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30113_ ( .A({ _03751_, _07796_, _07809_, _saxi_register_10[21] }), .Y(_20951_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30114_ ( .A({ _03750_, _07796_, _07809_, _saxi_register_10[20] }), .Y(_20950_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30115_ ( .A({ _03748_, _07796_, _07809_, _saxi_register_10[19] }), .Y(_20948_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30116_ ( .A({ _03747_, _07796_, _07809_, _saxi_register_10[18] }), .Y(_20947_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30117_ ( .A({ _03746_, _07796_, _07809_, _saxi_register_10[17] }), .Y(_20946_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30118_ ( .A({ _03745_, _07796_, _07809_, _saxi_register_10[16] }), .Y(_20945_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30119_ ( .A({ _03744_, _07796_, _07809_, _saxi_register_10[15] }), .Y(_20944_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30120_ ( .A({ _03743_, _07796_, _07809_, _saxi_register_10[14] }), .Y(_20943_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30121_ ( .A({ _03742_, _07796_, _07809_, _saxi_register_10[13] }), .Y(_20942_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30122_ ( .A({ _03741_, _07796_, _07809_, _saxi_register_10[12] }), .Y(_20941_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30123_ ( .A({ _03740_, _07796_, _07809_, _saxi_register_10[11] }), .Y(_20940_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30124_ ( .A({ _03739_, _07796_, _07809_, _saxi_register_10[10] }), .Y(_20939_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30125_ ( .A({ _03769_, _07796_, _07809_, _saxi_register_10[9] }), .Y(_20969_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30126_ ( .A({ _03768_, _07796_, _07809_, _saxi_register_10[8] }), .Y(_20968_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30127_ ( .A({ _03767_, _07796_, _07809_, _saxi_register_10[7] }), .Y(_20967_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30128_ ( .A({ _03766_, _07796_, _07809_, _saxi_register_10[6] }), .Y(_20966_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30129_ ( .A({ _03765_, _07796_, _07809_, _saxi_register_10[5] }), .Y(_20965_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30130_ ( .A({ _03764_, _07796_, _07809_, _saxi_register_10[4] }), .Y(_20964_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30131_ ( .A({ _03763_, _07796_, _07809_, _saxi_register_10[3] }), .Y(_20963_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30132_ ( .A({ _03760_, _07796_, _07809_, _saxi_register_10[2] }), .Y(_20960_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30133_ ( .A({ _03749_, _07796_, _07809_, _saxi_register_10[1] }), .Y(_20949_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30134_ ( .A({ _03738_, _07796_, _07809_, _saxi_register_10[0] }), .Y(_20938_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _30135_ ( .A({ _07809_, _07796_ }), .Y(_21928_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30136_ ( .A({ _03890_, _07813_, _07814_, _03730_ }), .Y(_20994_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30137_ ( .A({ _07812_, _07797_ }), .Y(_07813_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30138_ ( .A({ _07816_, _07815_ }), .Y(_07814_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30139_ ( .A({ _07802_, _07811_, main_fsm[4] }), .Y(_07815_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30140_ ( .A({ main_fsm[0], main_fsm[1], _07817_ }), .Y(_07816_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30141_ ( .A({ main_fsm[2], main_fsm[3] }), .Y(_07817_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30142_ ( .A({ _03889_, _07813_, _07814_, _03729_ }), .Y(_20993_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30143_ ( .A({ _03887_, _07813_, _07814_, _03727_ }), .Y(_20991_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30144_ ( .A({ _03886_, _07813_, _07814_, _03726_ }), .Y(_20990_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30145_ ( .A({ _03885_, _07813_, _07814_, _03725_ }), .Y(_20989_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30146_ ( .A({ _03884_, _07813_, _07814_, _03724_ }), .Y(_20988_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30147_ ( .A({ _03883_, _07813_, _07814_, _03723_ }), .Y(_20987_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30148_ ( .A({ _03882_, _07813_, _07814_, _03722_ }), .Y(_20986_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30149_ ( .A({ _03881_, _07813_, _07814_, _03721_ }), .Y(_20985_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30150_ ( .A({ _03880_, _07813_, _07814_, _03720_ }), .Y(_20984_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30151_ ( .A({ _03879_, _07813_, _07814_, _03719_ }), .Y(_20983_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30152_ ( .A({ _03878_, _07813_, _07814_, _03718_ }), .Y(_20982_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30153_ ( .A({ _03876_, _07813_, _07814_, _03716_ }), .Y(_20980_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30154_ ( .A({ _03875_, _07813_, _07814_, _03715_ }), .Y(_20979_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30155_ ( .A({ _03874_, _07813_, _07814_, _03714_ }), .Y(_20978_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30156_ ( .A({ _03873_, _07813_, _07814_, _03713_ }), .Y(_20977_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30157_ ( .A({ _03872_, _07813_, _07814_, _03712_ }), .Y(_20976_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30158_ ( .A({ _03871_, _07813_, _07814_, _03711_ }), .Y(_20975_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30159_ ( .A({ _03870_, _07813_, _07814_, _03710_ }), .Y(_20974_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30160_ ( .A({ _03869_, _07813_, _07814_, _03709_ }), .Y(_20973_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30161_ ( .A({ _03868_, _07813_, _07814_, _03708_ }), .Y(_20972_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30162_ ( .A({ _03867_, _07813_, _07814_, _03707_ }), .Y(_20971_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30163_ ( .A({ _03897_, _07813_, _07814_, _03737_ }), .Y(_21001_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30164_ ( .A({ _03896_, _07813_, _07814_, _03736_ }), .Y(_21000_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30165_ ( .A({ _03895_, _07813_, _07814_, _03735_ }), .Y(_20999_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30166_ ( .A({ _03894_, _07813_, _07814_, _03734_ }), .Y(_20998_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30167_ ( .A({ _03893_, _07813_, _07814_, _03733_ }), .Y(_20997_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30168_ ( .A({ _03892_, _07813_, _07814_, _03732_ }), .Y(_20996_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30169_ ( .A({ _03891_, _07813_, _07814_, _03731_ }), .Y(_20995_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30170_ ( .A({ _03888_, _07813_, _07814_, _03728_ }), .Y(_20992_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30171_ ( .A({ _03877_, _07813_, _07814_, _03717_ }), .Y(_20981_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30172_ ( .A({ _03866_, _07813_, _07814_, _03706_ }), .Y(_20970_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _30173_ ( .A({ _07814_, _07813_ }), .Y(_21929_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30174_ ( .A({ _03858_, _07818_, _07821_, _03698_ }), .Y(_21026_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30175_ ( .A({ _07819_, _07810_ }), .Y(_07818_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30176_ ( .A({ _07820_, main_fsm[1:0] }), .Y(_07819_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30177_ ( .A(main_fsm[3:2]), .Y(_07820_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30178_ ( .A({ _07822_, _07815_ }), .Y(_07821_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30179_ ( .A({ main_fsm[0], _07820_, main_fsm[1] }), .Y(_07822_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30180_ ( .A({ _03857_, _07818_, _07821_, _03697_ }), .Y(_21025_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30181_ ( .A({ _03855_, _07818_, _07821_, _03695_ }), .Y(_21023_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30182_ ( .A({ _03854_, _07818_, _07821_, _03694_ }), .Y(_21022_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30183_ ( .A({ _03853_, _07818_, _07821_, _03693_ }), .Y(_21021_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30184_ ( .A({ _03852_, _07818_, _07821_, _03692_ }), .Y(_21020_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30185_ ( .A({ _03851_, _07818_, _07821_, _03691_ }), .Y(_21019_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30186_ ( .A({ _03850_, _07818_, _07821_, _03690_ }), .Y(_21018_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30187_ ( .A({ _03849_, _07818_, _07821_, _03689_ }), .Y(_21017_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30188_ ( .A({ _03848_, _07818_, _07821_, _03688_ }), .Y(_21016_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30189_ ( .A({ _03847_, _07818_, _07821_, _03687_ }), .Y(_21015_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30190_ ( .A({ _03846_, _07818_, _07821_, _03686_ }), .Y(_21014_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30191_ ( .A({ _03844_, _07818_, _07821_, _03684_ }), .Y(_21012_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30192_ ( .A({ _03843_, _07818_, _07821_, _03683_ }), .Y(_21011_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30193_ ( .A({ _03842_, _07818_, _07821_, _03682_ }), .Y(_21010_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30194_ ( .A({ _03841_, _07818_, _07821_, _03681_ }), .Y(_21009_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30195_ ( .A({ _03840_, _07818_, _07821_, _03680_ }), .Y(_21008_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30196_ ( .A({ _03839_, _07818_, _07821_, _03679_ }), .Y(_21007_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30197_ ( .A({ _03838_, _07818_, _07821_, _03678_ }), .Y(_21006_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30198_ ( .A({ _03837_, _07818_, _07821_, _03677_ }), .Y(_21005_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30199_ ( .A({ _03836_, _07818_, _07821_, _03676_ }), .Y(_21004_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30200_ ( .A({ _03835_, _07818_, _07821_, _03675_ }), .Y(_21003_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30201_ ( .A({ _03865_, _07818_, _07821_, _03705_ }), .Y(_21033_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30202_ ( .A({ _03864_, _07818_, _07821_, _03704_ }), .Y(_21032_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30203_ ( .A({ _03863_, _07818_, _07821_, _03703_ }), .Y(_21031_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30204_ ( .A({ _03862_, _07818_, _07821_, _03702_ }), .Y(_21030_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30205_ ( .A({ _03861_, _07818_, _07821_, _03701_ }), .Y(_21029_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30206_ ( .A({ _03860_, _07818_, _07821_, _03700_ }), .Y(_21028_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30207_ ( .A({ _03859_, _07818_, _07821_, _03699_ }), .Y(_21027_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30208_ ( .A({ _03856_, _07818_, _07821_, _03696_ }), .Y(_21024_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30209_ ( .A({ _03845_, _07818_, _07821_, _03685_ }), .Y(_21013_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30210_ ( .A({ _03834_, _07818_, _07821_, _03674_ }), .Y(_21002_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _30211_ ( .A({ _07821_, _07818_ }), .Y(_21930_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30212_ ( .A({ _03826_, _07823_, _07824_, _03666_ }), .Y(_21058_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30213_ ( .A({ _07822_, _07810_ }), .Y(_07823_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30214_ ( .A({ _07825_, _07815_ }), .Y(_07824_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30215_ ( .A({ _07820_, main_fsm[0], main_fsm[1] }), .Y(_07825_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30216_ ( .A({ _03825_, _07823_, _07824_, _03665_ }), .Y(_21057_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30217_ ( .A({ _03823_, _07823_, _07824_, _03663_ }), .Y(_21055_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30218_ ( .A({ _03822_, _07823_, _07824_, _03662_ }), .Y(_21054_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30219_ ( .A({ _03821_, _07823_, _07824_, _03661_ }), .Y(_21053_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30220_ ( .A({ _03820_, _07823_, _07824_, _03660_ }), .Y(_21052_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30221_ ( .A({ _03819_, _07823_, _07824_, _03659_ }), .Y(_21051_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30222_ ( .A({ _03818_, _07823_, _07824_, _03658_ }), .Y(_21050_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30223_ ( .A({ _03817_, _07823_, _07824_, _03657_ }), .Y(_21049_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30224_ ( .A({ _03816_, _07823_, _07824_, _03656_ }), .Y(_21048_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30225_ ( .A({ _03815_, _07823_, _07824_, _03655_ }), .Y(_21047_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30226_ ( .A({ _03814_, _07823_, _07824_, _03654_ }), .Y(_21046_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30227_ ( .A({ _03812_, _07823_, _07824_, _03652_ }), .Y(_21044_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30228_ ( .A({ _03811_, _07823_, _07824_, _03651_ }), .Y(_21043_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30229_ ( .A({ _03810_, _07823_, _07824_, _03650_ }), .Y(_21042_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30230_ ( .A({ _03809_, _07823_, _07824_, _03649_ }), .Y(_21041_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30231_ ( .A({ _03808_, _07823_, _07824_, _03648_ }), .Y(_21040_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30232_ ( .A({ _03807_, _07823_, _07824_, _03647_ }), .Y(_21039_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30233_ ( .A({ _03806_, _07823_, _07824_, _03646_ }), .Y(_21038_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30234_ ( .A({ _03805_, _07823_, _07824_, _03645_ }), .Y(_21037_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30235_ ( .A({ _03804_, _07823_, _07824_, _03644_ }), .Y(_21036_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30236_ ( .A({ _03803_, _07823_, _07824_, _03643_ }), .Y(_21035_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30237_ ( .A({ _03833_, _07823_, _07824_, _03673_ }), .Y(_21065_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30238_ ( .A({ _03832_, _07823_, _07824_, _03672_ }), .Y(_21064_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30239_ ( .A({ _03831_, _07823_, _07824_, _03671_ }), .Y(_21063_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30240_ ( .A({ _03830_, _07823_, _07824_, _03670_ }), .Y(_21062_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30241_ ( .A({ _03829_, _07823_, _07824_, _03669_ }), .Y(_21061_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30242_ ( .A({ _03828_, _07823_, _07824_, _03668_ }), .Y(_21060_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30243_ ( .A({ _03827_, _07823_, _07824_, _03667_ }), .Y(_21059_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30244_ ( .A({ _03824_, _07823_, _07824_, _03664_ }), .Y(_21056_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30245_ ( .A({ _03813_, _07823_, _07824_, _03653_ }), .Y(_21045_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30246_ ( .A({ _03802_, _07823_, _07824_, _03642_ }), .Y(_21034_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _30247_ ( .A({ _07824_, _07823_ }), .Y(_21931_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30248_ ( .A({ _03794_, _07826_, _07827_, _saxi_register_13[31] }), .Y(_21090_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30249_ ( .A({ _07825_, _07810_ }), .Y(_07826_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30250_ ( .A({ _07828_, _07815_ }), .Y(_07827_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30251_ ( .A({ main_fsm[0], main_fsm[1], _07829_ }), .Y(_07828_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30252_ ( .A({ main_fsm[2], main_fsm[3] }), .Y(_07829_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30253_ ( .A({ _03793_, _07826_, _07827_, _saxi_register_13[30] }), .Y(_21089_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30254_ ( .A({ _03791_, _07826_, _07827_, _saxi_register_13[29] }), .Y(_21087_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30255_ ( .A({ _03790_, _07826_, _07827_, _saxi_register_13[28] }), .Y(_21086_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30256_ ( .A({ _03789_, _07826_, _07827_, _saxi_register_13[27] }), .Y(_21085_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30257_ ( .A({ _03788_, _07826_, _07827_, _saxi_register_13[26] }), .Y(_21084_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30258_ ( .A({ _03787_, _07826_, _07827_, _saxi_register_13[25] }), .Y(_21083_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30259_ ( .A({ _03786_, _07826_, _07827_, _saxi_register_13[24] }), .Y(_21082_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30260_ ( .A({ _03785_, _07826_, _07827_, _saxi_register_13[23] }), .Y(_21081_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30261_ ( .A({ _03784_, _07826_, _07827_, _saxi_register_13[22] }), .Y(_21080_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30262_ ( .A({ _03783_, _07826_, _07827_, _saxi_register_13[21] }), .Y(_21079_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30263_ ( .A({ _03782_, _07826_, _07827_, _saxi_register_13[20] }), .Y(_21078_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30264_ ( .A({ _03780_, _07826_, _07827_, _saxi_register_13[19] }), .Y(_21076_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30265_ ( .A({ _03779_, _07826_, _07827_, _saxi_register_13[18] }), .Y(_21075_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30266_ ( .A({ _03778_, _07826_, _07827_, _saxi_register_13[17] }), .Y(_21074_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30267_ ( .A({ _03777_, _07826_, _07827_, _saxi_register_13[16] }), .Y(_21073_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30268_ ( .A({ _03776_, _07826_, _07827_, _saxi_register_13[15] }), .Y(_21072_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30269_ ( .A({ _03775_, _07826_, _07827_, _saxi_register_13[14] }), .Y(_21071_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30270_ ( .A({ _03774_, _07826_, _07827_, _saxi_register_13[13] }), .Y(_21070_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30271_ ( .A({ _03773_, _07826_, _07827_, _saxi_register_13[12] }), .Y(_21069_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30272_ ( .A({ _03772_, _07826_, _07827_, _saxi_register_13[11] }), .Y(_21068_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30273_ ( .A({ _03771_, _07826_, _07827_, _saxi_register_13[10] }), .Y(_21067_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30274_ ( .A({ _03801_, _07826_, _07827_, _saxi_register_13[9] }), .Y(_21097_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30275_ ( .A({ _03800_, _07826_, _07827_, _saxi_register_13[8] }), .Y(_21096_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30276_ ( .A({ _03799_, _07826_, _07827_, _saxi_register_13[7] }), .Y(_21095_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30277_ ( .A({ _03798_, _07826_, _07827_, _saxi_register_13[6] }), .Y(_21094_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30278_ ( .A({ _03797_, _07826_, _07827_, _saxi_register_13[5] }), .Y(_21093_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30279_ ( .A({ _03796_, _07826_, _07827_, _saxi_register_13[4] }), .Y(_21092_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30280_ ( .A({ _03795_, _07826_, _07827_, _saxi_register_13[3] }), .Y(_21091_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30281_ ( .A({ _03792_, _07826_, _07827_, _saxi_register_13[2] }), .Y(_21088_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30282_ ( .A({ _03781_, _07826_, _07827_, _saxi_register_13[1] }), .Y(_21077_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30283_ ( .A({ _03770_, _07826_, _07827_, _saxi_register_13[0] }), .Y(_21066_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _30284_ ( .A({ _07827_, _07826_ }), .Y(_21932_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30285_ ( .A({ _03730_, _07830_, _saxi_register_12[31], _07831_ }), .Y(_21122_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30286_ ( .A({ _07828_, _07810_ }), .Y(_07830_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30287_ ( .A({ _07832_, _07815_ }), .Y(_07831_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30288_ ( .A({ _07829_, main_fsm[1:0] }), .Y(_07832_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30289_ ( .A({ _03729_, _07830_, _saxi_register_12[30], _07831_ }), .Y(_21121_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30290_ ( .A({ _03727_, _07830_, _saxi_register_12[29], _07831_ }), .Y(_21119_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30291_ ( .A({ _03726_, _07830_, _saxi_register_12[28], _07831_ }), .Y(_21118_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30292_ ( .A({ _03725_, _07830_, _saxi_register_12[27], _07831_ }), .Y(_21117_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30293_ ( .A({ _03724_, _07830_, _saxi_register_12[26], _07831_ }), .Y(_21116_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30294_ ( .A({ _03723_, _07830_, _saxi_register_12[25], _07831_ }), .Y(_21115_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30295_ ( .A({ _03722_, _07830_, _saxi_register_12[24], _07831_ }), .Y(_21114_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30296_ ( .A({ _03721_, _07830_, _saxi_register_12[23], _07831_ }), .Y(_21113_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30297_ ( .A({ _03720_, _07830_, _saxi_register_12[22], _07831_ }), .Y(_21112_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30298_ ( .A({ _03719_, _07830_, _saxi_register_12[21], _07831_ }), .Y(_21111_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30299_ ( .A({ _03718_, _07830_, _saxi_register_12[20], _07831_ }), .Y(_21110_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30300_ ( .A({ _03716_, _07830_, _saxi_register_12[19], _07831_ }), .Y(_21108_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30301_ ( .A({ _03715_, _07830_, _saxi_register_12[18], _07831_ }), .Y(_21107_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30302_ ( .A({ _03714_, _07830_, _saxi_register_12[17], _07831_ }), .Y(_21106_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30303_ ( .A({ _03713_, _07830_, _saxi_register_12[16], _07831_ }), .Y(_21105_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30304_ ( .A({ _03712_, _07830_, _saxi_register_12[15], _07831_ }), .Y(_21104_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30305_ ( .A({ _03711_, _07830_, _saxi_register_12[14], _07831_ }), .Y(_21103_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30306_ ( .A({ _03710_, _07830_, _saxi_register_12[13], _07831_ }), .Y(_21102_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30307_ ( .A({ _03709_, _07830_, _saxi_register_12[12], _07831_ }), .Y(_21101_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30308_ ( .A({ _03708_, _07830_, _saxi_register_12[11], _07831_ }), .Y(_21100_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30309_ ( .A({ _03707_, _07830_, _saxi_register_12[10], _07831_ }), .Y(_21099_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30310_ ( .A({ _03737_, _07830_, _saxi_register_12[9], _07831_ }), .Y(_21129_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30311_ ( .A({ _03736_, _07830_, _saxi_register_12[8], _07831_ }), .Y(_21128_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30312_ ( .A({ _03735_, _07830_, _saxi_register_12[7], _07831_ }), .Y(_21127_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30313_ ( .A({ _03734_, _07830_, _saxi_register_12[6], _07831_ }), .Y(_21126_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30314_ ( .A({ _03733_, _07830_, _saxi_register_12[5], _07831_ }), .Y(_21125_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30315_ ( .A({ _03732_, _07830_, _saxi_register_12[4], _07831_ }), .Y(_21124_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30316_ ( .A({ _03731_, _07830_, _saxi_register_12[3], _07831_ }), .Y(_21123_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30317_ ( .A({ _03728_, _07830_, _saxi_register_12[2], _07831_ }), .Y(_21120_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30318_ ( .A({ _03717_, _07830_, _saxi_register_12[1], _07831_ }), .Y(_21109_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30319_ ( .A({ _03706_, _07830_, _saxi_register_12[0], _07831_ }), .Y(_21098_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _30320_ ( .A({ _07831_, _07830_ }), .Y(_21933_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30321_ ( .A({ _03762_, _07833_, _07834_, _saxi_register_10[31] }), .Y(_21154_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30322_ ( .A({ _07832_, _07810_ }), .Y(_07833_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30323_ ( .A({ _07835_, _07815_ }), .Y(_07834_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30324_ ( .A({ main_fsm[0], _07829_, main_fsm[1] }), .Y(_07835_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30325_ ( .A({ _03761_, _07833_, _07834_, _saxi_register_10[30] }), .Y(_21153_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30326_ ( .A({ _03759_, _07833_, _07834_, _saxi_register_10[29] }), .Y(_21151_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30327_ ( .A({ _03758_, _07833_, _07834_, _saxi_register_10[28] }), .Y(_21150_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30328_ ( .A({ _03757_, _07833_, _07834_, _saxi_register_10[27] }), .Y(_21149_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30329_ ( .A({ _03756_, _07833_, _07834_, _saxi_register_10[26] }), .Y(_21148_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30330_ ( .A({ _03755_, _07833_, _07834_, _saxi_register_10[25] }), .Y(_21147_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30331_ ( .A({ _03754_, _07833_, _07834_, _saxi_register_10[24] }), .Y(_21146_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30332_ ( .A({ _03753_, _07833_, _07834_, _saxi_register_10[23] }), .Y(_21145_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30333_ ( .A({ _03752_, _07833_, _07834_, _saxi_register_10[22] }), .Y(_21144_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30334_ ( .A({ _03751_, _07833_, _07834_, _saxi_register_10[21] }), .Y(_21143_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30335_ ( .A({ _03750_, _07833_, _07834_, _saxi_register_10[20] }), .Y(_21142_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30336_ ( .A({ _03748_, _07833_, _07834_, _saxi_register_10[19] }), .Y(_21140_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30337_ ( .A({ _03747_, _07833_, _07834_, _saxi_register_10[18] }), .Y(_21139_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30338_ ( .A({ _03746_, _07833_, _07834_, _saxi_register_10[17] }), .Y(_21138_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30339_ ( .A({ _03745_, _07833_, _07834_, _saxi_register_10[16] }), .Y(_21137_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30340_ ( .A({ _03744_, _07833_, _07834_, _saxi_register_10[15] }), .Y(_21136_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30341_ ( .A({ _03743_, _07833_, _07834_, _saxi_register_10[14] }), .Y(_21135_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30342_ ( .A({ _03742_, _07833_, _07834_, _saxi_register_10[13] }), .Y(_21134_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30343_ ( .A({ _03741_, _07833_, _07834_, _saxi_register_10[12] }), .Y(_21133_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30344_ ( .A({ _03740_, _07833_, _07834_, _saxi_register_10[11] }), .Y(_21132_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30345_ ( .A({ _03739_, _07833_, _07834_, _saxi_register_10[10] }), .Y(_21131_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30346_ ( .A({ _03769_, _07833_, _07834_, _saxi_register_10[9] }), .Y(_21161_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30347_ ( .A({ _03768_, _07833_, _07834_, _saxi_register_10[8] }), .Y(_21160_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30348_ ( .A({ _03767_, _07833_, _07834_, _saxi_register_10[7] }), .Y(_21159_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30349_ ( .A({ _03766_, _07833_, _07834_, _saxi_register_10[6] }), .Y(_21158_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30350_ ( .A({ _03765_, _07833_, _07834_, _saxi_register_10[5] }), .Y(_21157_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30351_ ( .A({ _03764_, _07833_, _07834_, _saxi_register_10[4] }), .Y(_21156_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30352_ ( .A({ _03763_, _07833_, _07834_, _saxi_register_10[3] }), .Y(_21155_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30353_ ( .A({ _03760_, _07833_, _07834_, _saxi_register_10[2] }), .Y(_21152_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30354_ ( .A({ _03749_, _07833_, _07834_, _saxi_register_10[1] }), .Y(_21141_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30355_ ( .A({ _03738_, _07833_, _07834_, _saxi_register_10[0] }), .Y(_21130_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _30356_ ( .A({ _07834_, _07833_ }), .Y(_21934_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30357_ ( .A({ _07844_, _07841_, _07836_ }), .Y(_21187_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30358_ ( .A({ _21315_, _07837_, _21283_, _07839_ }), .Y(_07836_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30359_ ( .A({ _07838_, _07810_ }), .Y(_07837_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30360_ ( .A({ _07829_, main_fsm[0], main_fsm[1] }), .Y(_07838_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30361_ ( .A({ _07840_, _07810_ }), .Y(_07839_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30362_ ( .A({ _07817_, main_fsm[1:0] }), .Y(_07840_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30363_ ( .A({ _21347_, _07842_, _21379_, _04900_ }), .Y(_07841_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30364_ ( .A({ _07802_, _07843_, _07811_, main_fsm[4] }), .Y(_07842_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30365_ ( .A({ main_fsm[0], _07817_, main_fsm[1] }), .Y(_07843_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _30366_ ( .A({ _07802_, _07811_, _07812_, main_fsm[4] }), .Y(_04900_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30367_ ( .A({ _21251_, _07845_, _21219_, _07846_ }), .Y(_07844_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30368_ ( .A({ _07798_, _07835_, _07802_, main_fsm[4] }), .Y(_07845_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30369_ ( .A({ main_fsm[4], _07812_, _07802_, _07798_ }), .Y(_07846_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30370_ ( .A({ _07849_, _07848_, _07847_ }), .Y(_21186_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30371_ ( .A({ _21314_, _07837_, _21282_, _07839_ }), .Y(_07847_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30372_ ( .A({ _21346_, _07842_, _21378_, _04900_ }), .Y(_07848_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30373_ ( .A({ _21250_, _07845_, _21218_, _07846_ }), .Y(_07849_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30374_ ( .A({ _07852_, _07851_, _07850_ }), .Y(_21184_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30375_ ( .A({ _21312_, _07837_, _21280_, _07839_ }), .Y(_07850_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30376_ ( .A({ _21344_, _07842_, _21376_, _04900_ }), .Y(_07851_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30377_ ( .A({ _21248_, _07845_, _21216_, _07846_ }), .Y(_07852_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30378_ ( .A({ _07855_, _07854_, _07853_ }), .Y(_21183_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30379_ ( .A({ _21311_, _07837_, _21279_, _07839_ }), .Y(_07853_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30380_ ( .A({ _21343_, _07842_, _21375_, _04900_ }), .Y(_07854_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30381_ ( .A({ _21247_, _07845_, _21215_, _07846_ }), .Y(_07855_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30382_ ( .A({ _07858_, _07857_, _07856_ }), .Y(_21182_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30383_ ( .A({ _21310_, _07837_, _21278_, _07839_ }), .Y(_07856_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30384_ ( .A({ _21342_, _07842_, _21374_, _04900_ }), .Y(_07857_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30385_ ( .A({ _21246_, _07845_, _21214_, _07846_ }), .Y(_07858_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30386_ ( .A({ _07861_, _07860_, _07859_ }), .Y(_21181_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30387_ ( .A({ _21309_, _07837_, _21277_, _07839_ }), .Y(_07859_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30388_ ( .A({ _21341_, _07842_, _21373_, _04900_ }), .Y(_07860_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30389_ ( .A({ _21245_, _07845_, _21213_, _07846_ }), .Y(_07861_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30390_ ( .A({ _07864_, _07863_, _07862_ }), .Y(_21180_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30391_ ( .A({ _21308_, _07837_, _21276_, _07839_ }), .Y(_07862_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30392_ ( .A({ _21340_, _07842_, _21372_, _04900_ }), .Y(_07863_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30393_ ( .A({ _21244_, _07845_, _21212_, _07846_ }), .Y(_07864_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30394_ ( .A({ _07867_, _07866_, _07865_ }), .Y(_21179_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30395_ ( .A({ _21307_, _07837_, _21275_, _07839_ }), .Y(_07865_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30396_ ( .A({ _21339_, _07842_, _21371_, _04900_ }), .Y(_07866_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30397_ ( .A({ _21243_, _07845_, _21211_, _07846_ }), .Y(_07867_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30398_ ( .A({ _07870_, _07869_, _07868_ }), .Y(_21178_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30399_ ( .A({ _21306_, _07837_, _21274_, _07839_ }), .Y(_07868_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30400_ ( .A({ _21338_, _07842_, _21370_, _04900_ }), .Y(_07869_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30401_ ( .A({ _21242_, _07845_, _21210_, _07846_ }), .Y(_07870_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30402_ ( .A({ _07873_, _07872_, _07871_ }), .Y(_21177_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30403_ ( .A({ _21305_, _07837_, _21273_, _07839_ }), .Y(_07871_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30404_ ( .A({ _21337_, _07842_, _21369_, _04900_ }), .Y(_07872_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30405_ ( .A({ _21241_, _07845_, _21209_, _07846_ }), .Y(_07873_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30406_ ( .A({ _07876_, _07875_, _07874_ }), .Y(_21176_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30407_ ( .A({ _21304_, _07837_, _21272_, _07839_ }), .Y(_07874_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30408_ ( .A({ _21336_, _07842_, _21368_, _04900_ }), .Y(_07875_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30409_ ( .A({ _21240_, _07845_, _21208_, _07846_ }), .Y(_07876_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30410_ ( .A({ _07879_, _07878_, _07877_ }), .Y(_21175_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30411_ ( .A({ _21303_, _07837_, _21271_, _07839_ }), .Y(_07877_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30412_ ( .A({ _21335_, _07842_, _21367_, _04900_ }), .Y(_07878_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30413_ ( .A({ _21239_, _07845_, _21207_, _07846_ }), .Y(_07879_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30414_ ( .A({ _07882_, _07881_, _07880_ }), .Y(_21173_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30415_ ( .A({ _21301_, _07837_, _21269_, _07839_ }), .Y(_07880_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30416_ ( .A({ _21333_, _07842_, _21365_, _04900_ }), .Y(_07881_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30417_ ( .A({ _21237_, _07845_, _21205_, _07846_ }), .Y(_07882_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30418_ ( .A({ _07885_, _07884_, _07883_ }), .Y(_21172_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30419_ ( .A({ _21300_, _07837_, _21268_, _07839_ }), .Y(_07883_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30420_ ( .A({ _21332_, _07842_, _21364_, _04900_ }), .Y(_07884_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30421_ ( .A({ _21236_, _07845_, _21204_, _07846_ }), .Y(_07885_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30422_ ( .A({ _07888_, _07887_, _07886_ }), .Y(_21171_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30423_ ( .A({ _21299_, _07837_, _21267_, _07839_ }), .Y(_07886_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30424_ ( .A({ _21331_, _07842_, _21363_, _04900_ }), .Y(_07887_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30425_ ( .A({ _21235_, _07845_, _21203_, _07846_ }), .Y(_07888_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30426_ ( .A({ _07891_, _07890_, _07889_ }), .Y(_21170_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30427_ ( .A({ _21298_, _07837_, _21266_, _07839_ }), .Y(_07889_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30428_ ( .A({ _21330_, _07842_, _21362_, _04900_ }), .Y(_07890_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30429_ ( .A({ _21234_, _07845_, _21202_, _07846_ }), .Y(_07891_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30430_ ( .A({ _07894_, _07893_, _07892_ }), .Y(_21169_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30431_ ( .A({ _21297_, _07837_, _21265_, _07839_ }), .Y(_07892_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30432_ ( .A({ _21329_, _07842_, _21361_, _04900_ }), .Y(_07893_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30433_ ( .A({ _21233_, _07845_, _21201_, _07846_ }), .Y(_07894_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30434_ ( .A({ _07897_, _07896_, _07895_ }), .Y(_21168_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30435_ ( .A({ _21296_, _07837_, _21264_, _07839_ }), .Y(_07895_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30436_ ( .A({ _21328_, _07842_, _21360_, _04900_ }), .Y(_07896_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30437_ ( .A({ _21232_, _07845_, _21200_, _07846_ }), .Y(_07897_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30438_ ( .A({ _07900_, _07899_, _07898_ }), .Y(_21167_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30439_ ( .A({ _21295_, _07837_, _21263_, _07839_ }), .Y(_07898_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30440_ ( .A({ _21327_, _07842_, _21359_, _04900_ }), .Y(_07899_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30441_ ( .A({ _21231_, _07845_, _21199_, _07846_ }), .Y(_07900_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30442_ ( .A({ _07903_, _07902_, _07901_ }), .Y(_21166_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30443_ ( .A({ _21294_, _07837_, _21262_, _07839_ }), .Y(_07901_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30444_ ( .A({ _21326_, _07842_, _21358_, _04900_ }), .Y(_07902_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30445_ ( .A({ _21230_, _07845_, _21198_, _07846_ }), .Y(_07903_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30446_ ( .A({ _07906_, _07905_, _07904_ }), .Y(_21165_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30447_ ( .A({ _21293_, _07837_, _21261_, _07839_ }), .Y(_07904_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30448_ ( .A({ _21325_, _07842_, _21357_, _04900_ }), .Y(_07905_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30449_ ( .A({ _21229_, _07845_, _21197_, _07846_ }), .Y(_07906_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30450_ ( .A({ _07909_, _07908_, _07907_ }), .Y(_21164_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30451_ ( .A({ _21292_, _07837_, _21260_, _07839_ }), .Y(_07907_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30452_ ( .A({ _21324_, _07842_, _21356_, _04900_ }), .Y(_07908_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30453_ ( .A({ _21228_, _07845_, _21196_, _07846_ }), .Y(_07909_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30454_ ( .A({ _07912_, _07911_, _07910_ }), .Y(_21194_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30455_ ( .A({ _21322_, _07837_, _21290_, _07839_ }), .Y(_07910_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30456_ ( .A({ _21354_, _07842_, _21386_, _04900_ }), .Y(_07911_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30457_ ( .A({ _21258_, _07845_, _21226_, _07846_ }), .Y(_07912_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30458_ ( .A({ _07915_, _07914_, _07913_ }), .Y(_21193_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30459_ ( .A({ _21321_, _07837_, _21289_, _07839_ }), .Y(_07913_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30460_ ( .A({ _21353_, _07842_, _21385_, _04900_ }), .Y(_07914_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30461_ ( .A({ _21257_, _07845_, _21225_, _07846_ }), .Y(_07915_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30462_ ( .A({ _07918_, _07917_, _07916_ }), .Y(_21192_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30463_ ( .A({ _21320_, _07837_, _21288_, _07839_ }), .Y(_07916_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30464_ ( .A({ _21352_, _07842_, _21384_, _04900_ }), .Y(_07917_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30465_ ( .A({ _21256_, _07845_, _21224_, _07846_ }), .Y(_07918_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30466_ ( .A({ _07921_, _07920_, _07919_ }), .Y(_21191_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30467_ ( .A({ _21319_, _07837_, _21287_, _07839_ }), .Y(_07919_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30468_ ( .A({ _21351_, _07842_, _21383_, _04900_ }), .Y(_07920_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30469_ ( .A({ _21255_, _07845_, _21223_, _07846_ }), .Y(_07921_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30470_ ( .A({ _07922_, _07797_ }), .Y(_04831_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30471_ ( .A({ _07808_, main_fsm[1:0] }), .Y(_07922_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30472_ ( .A({ _07940_, _07923_ }), .Y(_21190_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30473_ ( .A({ _07935_, _05141_, _07931_, _07924_ }), .Y(_07923_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30474_ ( .A({ _07930_, _07929_, _07927_, _07925_ }), .Y(_07924_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30475_ ( .A({ _07797_, _07926_, _07840_ }), .Y(_07925_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30476_ ( .A({ _07817_, main_fsm[0], main_fsm[1] }), .Y(_07926_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30477_ ( .A({ _07797_, _07928_, _07843_ }), .Y(_07927_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30478_ ( .A({ main_fsm[0], main_fsm[1], _07820_ }), .Y(_07928_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30479_ ( .A({ _07797_, _07822_, _07819_ }), .Y(_07929_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30480_ ( .A({ _07797_, _07828_, _07825_ }), .Y(_07930_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30481_ ( .A({ _07932_, _04831_, _07796_ }), .Y(_07931_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30482_ ( .A({ _07933_, _07922_, _07807_ }), .Y(_07932_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30483_ ( .A({ main_fsm[4], _07802_, _07798_ }), .Y(_07933_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30484_ ( .A({ main_fsm[1], _07934_ }), .Y(_05141_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30485_ ( .A({ _07797_, _07829_, main_fsm[0] }), .Y(_07934_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30486_ ( .A({ _05143_, _07937_, _07936_, _07813_ }), .Y(_07935_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30487_ ( .A({ _07816_, _07797_ }), .Y(_07936_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30488_ ( .A({ _07816_, _07810_ }), .Y(_05143_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30489_ ( .A({ _07933_, _07938_ }), .Y(_07937_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _30490_ ( .A({ _07939_, _07838_, _07835_ }), .Y(_07938_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30491_ ( .A({ main_fsm[0], main_fsm[1], _07808_ }), .Y(_07939_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30492_ ( .A({ _07942_, _07941_, _07839_, _21286_ }), .Y(_07940_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30493_ ( .A({ _21318_, _07837_, _07842_, _21350_ }), .Y(_07941_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _30494_ ( .A({ _07944_, _07943_, _04900_, _21382_ }), .Y(_07942_) );
  \$lut  #( .LUT(8'he0), .WIDTH(3) ) _30495_ ( .A({ _07797_, _07838_, _07939_ }), .Y(_07943_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30496_ ( .A({ _21254_, _07845_, _21222_, _07846_ }), .Y(_07944_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30497_ ( .A({ _21381_, _04900_, _21253_, _07845_ }), .Y(_07945_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30498_ ( .A({ _05144_, _21162_ }), .Y(_07946_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30499_ ( .A({ _07926_, _07810_ }), .Y(_05144_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30500_ ( .A({ _07928_, _07810_ }), .Y(_21162_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30501_ ( .A({ _05145_, _07833_ }), .Y(_07947_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30502_ ( .A({ _07948_, main_fsm[5] }), .Y(_05145_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30503_ ( .A({ main_fsm[4], _07835_, _07802_, _07949_ }), .Y(_07948_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30504_ ( .A({ _07801_, _07800_, _07799_ }), .Y(_07949_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30505_ ( .A({ _07952_, _07951_, _07814_, _07809_ }), .Y(_07950_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30506_ ( .A({ _07830_, _07826_, _07823_, _07818_ }), .Y(_07951_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30507_ ( .A({ _07810_, _07922_, _07807_ }), .Y(_07952_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _30508_ ( .A({ _07954_, _07839_, _21285_ }), .Y(_07953_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _30509_ ( .A({ _07955_, _07937_, _07846_, _21221_ }), .Y(_07954_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30510_ ( .A({ _07939_, _07810_ }), .Y(_07955_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30511_ ( .A({ _07924_, _07960_, _07956_ }), .Y(_21188_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30512_ ( .A({ _07959_, _07957_, _07951_, _07946_ }), .Y(_07956_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30513_ ( .A({ _07958_, _07827_, _07824_ }), .Y(_07957_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30514_ ( .A({ _07815_, _07822_, _07819_ }), .Y(_07958_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30515_ ( .A({ _07843_, _07810_, _07815_, _07840_ }), .Y(_07959_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30516_ ( .A({ _07964_, _07963_, _07962_, _07961_ }), .Y(_07960_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30517_ ( .A({ _21316_, _07837_, _21220_, _07846_ }), .Y(_07961_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30518_ ( .A({ _21284_, _07839_, _21380_, _04900_ }), .Y(_07962_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30519_ ( .A({ _07815_, _07928_, _07926_ }), .Y(_07963_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30520_ ( .A({ _21348_, _07842_, _21252_, _07845_ }), .Y(_07964_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30521_ ( .A({ _07970_, _07968_, _07967_, _07965_ }), .Y(_21185_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30522_ ( .A({ _05142_, _07947_, _07966_, _07934_ }), .Y(_07965_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30523_ ( .A({ _07963_, _07955_, _07937_ }), .Y(_07966_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30524_ ( .A({ _07939_, _07797_ }), .Y(_05142_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30525_ ( .A({ _07959_, _07927_, _07925_, _07946_ }), .Y(_07967_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _30526_ ( .A({ _07969_, _07845_, _21249_ }), .Y(_07968_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30527_ ( .A({ _21281_, _07839_, _07842_, _21345_ }), .Y(_07969_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30528_ ( .A({ _07972_, _07971_, _07846_, _21217_ }), .Y(_07970_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30529_ ( .A({ _21313_, _07837_, _21377_, _04900_ }), .Y(_07971_) );
  \$lut  #( .LUT(8'h4f), .WIDTH(3) ) _30530_ ( .A({ _07815_, _07938_, _07832_ }), .Y(_07972_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30531_ ( .A({ _07982_, _07979_, _07976_, _07973_ }), .Y(_21174_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30532_ ( .A({ _07974_, _05141_, _07931_, _21934_ }), .Y(_07973_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30533_ ( .A({ _07975_, _07948_, _07831_ }), .Y(_07974_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30534_ ( .A({ _07797_, _07843_, _07840_ }), .Y(_07975_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30535_ ( .A({ _07978_, _07977_ }), .Y(_07976_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30536_ ( .A({ _21270_, _07839_, _07842_, _21334_ }), .Y(_07977_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30537_ ( .A({ _21238_, _07845_, _21206_, _07846_ }), .Y(_07978_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _30538_ ( .A({ _07958_, _07980_, _04900_, _21366_ }), .Y(_07979_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _30539_ ( .A({ _07981_, _07837_, _21302_ }), .Y(_07980_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30540_ ( .A({ _07815_, _07922_, _07807_ }), .Y(_07981_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30541_ ( .A({ _07952_, _07929_, _07983_ }), .Y(_07982_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30542_ ( .A({ _07959_, _07823_, _07818_ }), .Y(_07983_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _30543_ ( .A({ _07985_, _07815_, _07926_, _07922_ }), .Y(_07984_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30544_ ( .A({ _07815_, _07840_, _07819_ }), .Y(_07985_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30545_ ( .A({ _07987_, _05146_, _05144_ }), .Y(_07986_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30546_ ( .A({ _07922_, _07810_ }), .Y(_05146_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30547_ ( .A({ _07797_, _07825_, _07819_ }), .Y(_07987_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _30548_ ( .A({ _07989_, _04900_, _21355_ }), .Y(_07988_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30549_ ( .A({ _21291_, _07837_, _07842_, _21323_ }), .Y(_07989_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _30550_ ( .A({ _07991_, _07992_, _07846_, _21195_ }), .Y(_07990_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30551_ ( .A({ _21259_, _07839_, _21227_, _07845_ }), .Y(_07991_) );
  \$lut  #( .LUT(8'he0), .WIDTH(3) ) _30552_ ( .A({ _07838_, _07815_, _07933_ }), .Y(_07992_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30553_ ( .A({ _07925_, _07994_, _07813_, _07809_ }), .Y(_07993_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30554_ ( .A({ _07831_, _07826_, _07824_, _07818_ }), .Y(_07994_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30555_ ( .A({ _07997_, _07995_, _07950_, _07923_ }), .Y(_21935_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30556_ ( .A({ _07996_, _07957_, _07947_, _07946_ }), .Y(_07995_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _30557_ ( .A({ _07955_, _07943_, _07933_, _07832_ }), .Y(_07996_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30558_ ( .A({ _07981_, _07972_, _07963_, _07998_ }), .Y(_07997_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30559_ ( .A({ _07999_, _07959_, _07839_, _07837_ }), .Y(_07998_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30560_ ( .A({ _04900_, _07846_, _07845_, _07842_ }), .Y(_07999_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _30561_ ( .A({ _04831_, _07807_, _07810_ }), .Y(_21936_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _30562_ ( .A({ _21162_, _07819_, _07815_ }), .Y(_21937_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30563_ ( .A({ _08005_, _08000_ }), .Y(_tmp_1091) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30564_ ( .A({ _stream_matmul_15_fsm[1], _08004_, _08001_ }), .Y(_08000_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30565_ ( .A({ _08003_, _08002_, _stream_matmul_15_fsm[3:2] }), .Y(_08001_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30566_ ( .A(_stream_matmul_15_fsm[15:12]), .Y(_08002_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30567_ ( .A(_stream_matmul_15_fsm[11:8]), .Y(_08003_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30568_ ( .A(_stream_matmul_15_fsm[7:4]), .Y(_08004_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30569_ ( .A({ _stream_matmul_15_fsm[0], _08006_ }), .Y(_08005_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30570_ ( .A({ _08010_, _08009_, _08008_, _08007_ }), .Y(_08006_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30571_ ( .A(_stream_matmul_15_fsm[23:20]), .Y(_08007_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30572_ ( .A(_stream_matmul_15_fsm[19:16]), .Y(_08008_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30573_ ( .A(_stream_matmul_15_fsm[31:28]), .Y(_08009_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30574_ ( .A(_stream_matmul_15_fsm[27:24]), .Y(_08010_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30575_ ( .A({ _04901_, _tmp_1091 }), .Y(_21938_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30576_ ( .A({ _08012_, _08011_ }), .Y(_04901_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30577_ ( .A({ _08006_, _stream_matmul_15_fsm[0] }), .Y(_08011_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30578_ ( .A({ _08001_, _08004_, _stream_matmul_15_fsm[1] }), .Y(_08012_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30579_ ( .A({ _21477_, _04901_, _21445_, _08013_ }), .Y(_21413_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30580_ ( .A({ _08011_, _08000_ }), .Y(_08013_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30581_ ( .A({ _21476_, _04901_, _21444_, _08013_ }), .Y(_21412_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30582_ ( .A({ _21474_, _04901_, _21442_, _08013_ }), .Y(_21410_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30583_ ( .A({ _21473_, _04901_, _21441_, _08013_ }), .Y(_21409_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30584_ ( .A({ _21472_, _04901_, _21440_, _08013_ }), .Y(_21408_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30585_ ( .A({ _21471_, _04901_, _21439_, _08013_ }), .Y(_21407_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30586_ ( .A({ _21470_, _04901_, _21438_, _08013_ }), .Y(_21406_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30587_ ( .A({ _21469_, _04901_, _21437_, _08013_ }), .Y(_21405_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30588_ ( .A({ _21468_, _04901_, _21436_, _08013_ }), .Y(_21404_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30589_ ( .A({ _21467_, _04901_, _21435_, _08013_ }), .Y(_21403_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30590_ ( .A({ _21466_, _04901_, _21434_, _08013_ }), .Y(_21402_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30591_ ( .A({ _21465_, _04901_, _21433_, _08013_ }), .Y(_21401_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30592_ ( .A({ _21463_, _04901_, _21431_, _08013_ }), .Y(_21399_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30593_ ( .A({ _21462_, _04901_, _21430_, _08013_ }), .Y(_21398_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30594_ ( .A({ _21461_, _04901_, _21429_, _08013_ }), .Y(_21397_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30595_ ( .A({ _21460_, _04901_, _21428_, _08013_ }), .Y(_21396_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30596_ ( .A({ _21459_, _04901_, _21427_, _08013_ }), .Y(_21395_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30597_ ( .A({ _21458_, _04901_, _21426_, _08013_ }), .Y(_21394_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30598_ ( .A({ _21457_, _04901_, _21425_, _08013_ }), .Y(_21393_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30599_ ( .A({ _21456_, _04901_, _21424_, _08013_ }), .Y(_21392_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30600_ ( .A({ _21455_, _04901_, _21423_, _08013_ }), .Y(_21391_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30601_ ( .A({ _21454_, _04901_, _21422_, _08013_ }), .Y(_21390_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30602_ ( .A({ _21484_, _04901_, _21452_, _08013_ }), .Y(_21420_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30603_ ( .A({ _21483_, _04901_, _21451_, _08013_ }), .Y(_21419_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30604_ ( .A({ _21482_, _04901_, _21450_, _08013_ }), .Y(_21418_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30605_ ( .A({ _21481_, _04901_, _21449_, _08013_ }), .Y(_21417_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30606_ ( .A({ _21480_, _04901_, _21448_, _08013_ }), .Y(_21416_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30607_ ( .A({ _21479_, _04901_, _21447_, _08013_ }), .Y(_21415_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30608_ ( .A({ _21478_, _04901_, _21446_, _08013_ }), .Y(_21414_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30609_ ( .A({ _21475_, _04901_, _21443_, _08013_ }), .Y(_21411_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30610_ ( .A({ _08014_, _21432_, _08013_ }), .Y(_21400_) );
  \$lut  #( .LUT(16'h07ff), .WIDTH(4) ) _30611_ ( .A({ _08012_, _08005_, _21464_, _08011_ }), .Y(_08014_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30612_ ( .A({ _21453_, _04901_, _21421_, _08013_ }), .Y(_21389_) );
  \$lut  #( .LUT(8'he0), .WIDTH(3) ) _30613_ ( .A({ _08006_, _08000_, _08012_ }), .Y(_21939_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30614_ ( .A({ _08020_, _08015_ }), .Y(_tmp_894) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30615_ ( .A({ _stream_max_pool_serial_9_fsm[1], _08019_, _08016_ }), .Y(_08015_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30616_ ( .A({ _08018_, _08017_, _stream_max_pool_serial_9_fsm[3:2] }), .Y(_08016_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30617_ ( .A(_stream_max_pool_serial_9_fsm[15:12]), .Y(_08017_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30618_ ( .A(_stream_max_pool_serial_9_fsm[11:8]), .Y(_08018_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30619_ ( .A(_stream_max_pool_serial_9_fsm[7:4]), .Y(_08019_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30620_ ( .A({ _stream_max_pool_serial_9_fsm[0], _08021_ }), .Y(_08020_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30621_ ( .A({ _08025_, _08024_, _08023_, _08022_ }), .Y(_08021_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30622_ ( .A(_stream_max_pool_serial_9_fsm[23:20]), .Y(_08022_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30623_ ( .A(_stream_max_pool_serial_9_fsm[19:16]), .Y(_08023_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30624_ ( .A(_stream_max_pool_serial_9_fsm[31:28]), .Y(_08024_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30625_ ( .A(_stream_max_pool_serial_9_fsm[27:24]), .Y(_08025_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30626_ ( .A({ _04902_, _tmp_894 }), .Y(_21940_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30627_ ( .A({ _08027_, _08026_ }), .Y(_04902_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30628_ ( .A({ _08021_, _stream_max_pool_serial_9_fsm[0] }), .Y(_08026_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30629_ ( .A({ _08016_, _08019_, _stream_max_pool_serial_9_fsm[1] }), .Y(_08027_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30630_ ( .A({ _21575_, _04902_, _21543_, _08028_ }), .Y(_21511_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30631_ ( .A({ _08026_, _08015_ }), .Y(_08028_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30632_ ( .A({ _21574_, _04902_, _21542_, _08028_ }), .Y(_21510_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30633_ ( .A({ _21572_, _04902_, _21540_, _08028_ }), .Y(_21508_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30634_ ( .A({ _21571_, _04902_, _21539_, _08028_ }), .Y(_21507_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30635_ ( .A({ _21570_, _04902_, _21538_, _08028_ }), .Y(_21506_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30636_ ( .A({ _21569_, _04902_, _21537_, _08028_ }), .Y(_21505_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30637_ ( .A({ _21568_, _04902_, _21536_, _08028_ }), .Y(_21504_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30638_ ( .A({ _21567_, _04902_, _21535_, _08028_ }), .Y(_21503_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30639_ ( .A({ _21566_, _04902_, _21534_, _08028_ }), .Y(_21502_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30640_ ( .A({ _21565_, _04902_, _21533_, _08028_ }), .Y(_21501_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30641_ ( .A({ _21564_, _04902_, _21532_, _08028_ }), .Y(_21500_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30642_ ( .A({ _21563_, _04902_, _21531_, _08028_ }), .Y(_21499_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30643_ ( .A({ _21561_, _04902_, _21529_, _08028_ }), .Y(_21497_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30644_ ( .A({ _21560_, _04902_, _21528_, _08028_ }), .Y(_21496_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30645_ ( .A({ _21559_, _04902_, _21527_, _08028_ }), .Y(_21495_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30646_ ( .A({ _21558_, _04902_, _21526_, _08028_ }), .Y(_21494_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30647_ ( .A({ _21557_, _04902_, _21525_, _08028_ }), .Y(_21493_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30648_ ( .A({ _21556_, _04902_, _21524_, _08028_ }), .Y(_21492_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30649_ ( .A({ _21555_, _04902_, _21523_, _08028_ }), .Y(_21491_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30650_ ( .A({ _21554_, _04902_, _21522_, _08028_ }), .Y(_21490_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30651_ ( .A({ _21553_, _04902_, _21521_, _08028_ }), .Y(_21489_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30652_ ( .A({ _21552_, _04902_, _21520_, _08028_ }), .Y(_21488_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30653_ ( .A({ _21582_, _04902_, _21550_, _08028_ }), .Y(_21518_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30654_ ( .A({ _21581_, _04902_, _21549_, _08028_ }), .Y(_21517_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30655_ ( .A({ _21580_, _04902_, _21548_, _08028_ }), .Y(_21516_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30656_ ( .A({ _21579_, _04902_, _21547_, _08028_ }), .Y(_21515_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30657_ ( .A({ _21578_, _04902_, _21546_, _08028_ }), .Y(_21514_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30658_ ( .A({ _21577_, _04902_, _21545_, _08028_ }), .Y(_21513_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30659_ ( .A({ _21576_, _04902_, _21544_, _08028_ }), .Y(_21512_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30660_ ( .A({ _21573_, _04902_, _21541_, _08028_ }), .Y(_21509_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30661_ ( .A({ _08029_, _21530_, _08028_ }), .Y(_21498_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _30662_ ( .A({ _08030_, _04902_, _21562_ }), .Y(_08029_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30663_ ( .A({ _08027_, _08020_ }), .Y(_08030_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30664_ ( .A({ _21551_, _04902_, _21519_, _08028_ }), .Y(_21487_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _30665_ ( .A({ _08030_, _08028_, _21940_ }), .Y(_21941_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30666_ ( .A({ _08036_, _08031_ }), .Y(_tmp_771) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30667_ ( .A({ _stream_conv2d_8_fsm[1], _08035_, _08032_ }), .Y(_08031_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30668_ ( .A({ _08034_, _08033_, _stream_conv2d_8_fsm[3:2] }), .Y(_08032_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30669_ ( .A(_stream_conv2d_8_fsm[15:12]), .Y(_08033_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30670_ ( .A(_stream_conv2d_8_fsm[11:8]), .Y(_08034_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30671_ ( .A(_stream_conv2d_8_fsm[7:4]), .Y(_08035_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30672_ ( .A({ _stream_conv2d_8_fsm[0], _08037_ }), .Y(_08036_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30673_ ( .A({ _08041_, _08040_, _08039_, _08038_ }), .Y(_08037_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30674_ ( .A(_stream_conv2d_8_fsm[23:20]), .Y(_08038_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30675_ ( .A(_stream_conv2d_8_fsm[19:16]), .Y(_08039_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30676_ ( .A(_stream_conv2d_8_fsm[31:28]), .Y(_08040_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30677_ ( .A(_stream_conv2d_8_fsm[27:24]), .Y(_08041_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30678_ ( .A({ _04903_, _tmp_771 }), .Y(_21942_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30679_ ( .A({ _08043_, _08042_ }), .Y(_04903_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30680_ ( .A({ _08037_, _stream_conv2d_8_fsm[0] }), .Y(_08042_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30681_ ( .A({ _08032_, _08035_, _stream_conv2d_8_fsm[1] }), .Y(_08043_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30682_ ( .A({ _21673_, _04903_, _21641_, _08044_ }), .Y(_21609_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30683_ ( .A({ _08042_, _08031_ }), .Y(_08044_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30684_ ( .A({ _21672_, _04903_, _21640_, _08044_ }), .Y(_21608_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30685_ ( .A({ _21670_, _04903_, _21638_, _08044_ }), .Y(_21606_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30686_ ( .A({ _21669_, _04903_, _21637_, _08044_ }), .Y(_21605_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30687_ ( .A({ _21668_, _04903_, _21636_, _08044_ }), .Y(_21604_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30688_ ( .A({ _21667_, _04903_, _21635_, _08044_ }), .Y(_21603_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30689_ ( .A({ _21666_, _04903_, _21634_, _08044_ }), .Y(_21602_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30690_ ( .A({ _21665_, _04903_, _21633_, _08044_ }), .Y(_21601_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30691_ ( .A({ _21664_, _04903_, _21632_, _08044_ }), .Y(_21600_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30692_ ( .A({ _21663_, _04903_, _21631_, _08044_ }), .Y(_21599_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30693_ ( .A({ _21662_, _04903_, _21630_, _08044_ }), .Y(_21598_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30694_ ( .A({ _21661_, _04903_, _21629_, _08044_ }), .Y(_21597_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30695_ ( .A({ _21659_, _04903_, _21627_, _08044_ }), .Y(_21595_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30696_ ( .A({ _21658_, _04903_, _21626_, _08044_ }), .Y(_21594_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30697_ ( .A({ _21657_, _04903_, _21625_, _08044_ }), .Y(_21593_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30698_ ( .A({ _21656_, _04903_, _21624_, _08044_ }), .Y(_21592_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30699_ ( .A({ _21655_, _04903_, _21623_, _08044_ }), .Y(_21591_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30700_ ( .A({ _21654_, _04903_, _21622_, _08044_ }), .Y(_21590_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30701_ ( .A({ _21653_, _04903_, _21621_, _08044_ }), .Y(_21589_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30702_ ( .A({ _21652_, _04903_, _21620_, _08044_ }), .Y(_21588_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30703_ ( .A({ _21651_, _04903_, _21619_, _08044_ }), .Y(_21587_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30704_ ( .A({ _21650_, _04903_, _21618_, _08044_ }), .Y(_21586_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30705_ ( .A({ _21680_, _04903_, _21648_, _08044_ }), .Y(_21616_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30706_ ( .A({ _21679_, _04903_, _21647_, _08044_ }), .Y(_21615_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30707_ ( .A({ _21678_, _04903_, _21646_, _08044_ }), .Y(_21614_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30708_ ( .A({ _21677_, _04903_, _21645_, _08044_ }), .Y(_21613_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30709_ ( .A({ _21676_, _04903_, _21644_, _08044_ }), .Y(_21612_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30710_ ( .A({ _21675_, _04903_, _21643_, _08044_ }), .Y(_21611_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30711_ ( .A({ _21674_, _04903_, _21642_, _08044_ }), .Y(_21610_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30712_ ( .A({ _21671_, _04903_, _21639_, _08044_ }), .Y(_21607_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30713_ ( .A({ _08045_, _21628_, _08044_ }), .Y(_21596_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _30714_ ( .A({ _08046_, _04903_, _21660_ }), .Y(_08045_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30715_ ( .A({ _08043_, _08036_ }), .Y(_08046_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30716_ ( .A({ _21649_, _04903_, _21617_, _08044_ }), .Y(_21585_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _30717_ ( .A({ _08046_, _08044_, _21942_ }), .Y(_21943_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30718_ ( .A({ _08047_, _saxi_register_fsm[0], _21737_, _21769_ }), .Y(_21705_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30719_ ( .A({ _08048_, _08056_, _saxi_register_fsm[1] }), .Y(_08047_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30720_ ( .A({ _08055_, _08054_, _08049_ }), .Y(_08048_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30721_ ( .A({ _08053_, _08052_, _08051_, _08050_ }), .Y(_08049_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30722_ ( .A(_saxi_register_fsm[23:20]), .Y(_08050_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30723_ ( .A(_saxi_register_fsm[19:16]), .Y(_08051_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30724_ ( .A(_saxi_register_fsm[31:28]), .Y(_08052_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30725_ ( .A(_saxi_register_fsm[27:24]), .Y(_08053_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30726_ ( .A(_saxi_register_fsm[15:12]), .Y(_08054_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30727_ ( .A(_saxi_register_fsm[11:8]), .Y(_08055_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30728_ ( .A({ _08057_, _saxi_register_fsm[3:2] }), .Y(_08056_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30729_ ( .A(_saxi_register_fsm[7:4]), .Y(_08057_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30730_ ( .A({ _08047_, _saxi_register_fsm[0], _21736_, _21768_ }), .Y(_21704_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30731_ ( .A({ _08047_, _saxi_register_fsm[0], _21734_, _21766_ }), .Y(_21702_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30732_ ( .A({ _08047_, _saxi_register_fsm[0], _21733_, _21765_ }), .Y(_21701_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30733_ ( .A({ _08047_, _saxi_register_fsm[0], _21732_, _21764_ }), .Y(_21700_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30734_ ( .A({ _08047_, _saxi_register_fsm[0], _21731_, _21763_ }), .Y(_21699_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30735_ ( .A({ _08047_, _saxi_register_fsm[0], _21730_, _21762_ }), .Y(_21698_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30736_ ( .A({ _08047_, _saxi_register_fsm[0], _21729_, _21761_ }), .Y(_21697_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30737_ ( .A({ _08047_, _saxi_register_fsm[0], _21728_, _21760_ }), .Y(_21696_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30738_ ( .A({ _08047_, _saxi_register_fsm[0], _21727_, _21759_ }), .Y(_21695_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30739_ ( .A({ _08047_, _saxi_register_fsm[0], _21726_, _21758_ }), .Y(_21694_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30740_ ( .A({ _08047_, _saxi_register_fsm[0], _21725_, _21757_ }), .Y(_21693_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30741_ ( .A({ _08047_, _saxi_register_fsm[0], _21723_, _21755_ }), .Y(_21691_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30742_ ( .A({ _08047_, _saxi_register_fsm[0], _21722_, _21754_ }), .Y(_21690_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30743_ ( .A({ _08047_, _saxi_register_fsm[0], _21721_, _21753_ }), .Y(_21689_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30744_ ( .A({ _08047_, _saxi_register_fsm[0], _21720_, _21752_ }), .Y(_21688_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30745_ ( .A({ _08047_, _saxi_register_fsm[0], _21719_, _21751_ }), .Y(_21687_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30746_ ( .A({ _08047_, _saxi_register_fsm[0], _21718_, _21750_ }), .Y(_21686_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30747_ ( .A({ _08047_, _saxi_register_fsm[0], _21717_, _21749_ }), .Y(_21685_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30748_ ( .A({ _08047_, _saxi_register_fsm[0], _21716_, _21748_ }), .Y(_21684_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30749_ ( .A({ _08047_, _saxi_register_fsm[0], _21715_, _21747_ }), .Y(_21683_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30750_ ( .A({ _08047_, _saxi_register_fsm[0], _21714_, _21746_ }), .Y(_21682_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30751_ ( .A({ _08047_, _saxi_register_fsm[0], _21744_, _21776_ }), .Y(_21712_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30752_ ( .A({ _08047_, _saxi_register_fsm[0], _21743_, _21775_ }), .Y(_21711_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30753_ ( .A({ _08047_, _saxi_register_fsm[0], _21742_, _21774_ }), .Y(_21710_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30754_ ( .A({ _08047_, _saxi_register_fsm[0], _21741_, _21773_ }), .Y(_21709_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30755_ ( .A({ _08047_, _saxi_register_fsm[0], _21740_, _21772_ }), .Y(_21708_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30756_ ( .A({ _08047_, _saxi_register_fsm[0], _21739_, _21771_ }), .Y(_21707_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30757_ ( .A({ _08047_, _saxi_register_fsm[0], _21738_, _21770_ }), .Y(_21706_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30758_ ( .A({ _08047_, _saxi_register_fsm[0], _21735_, _21767_ }), .Y(_21703_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30759_ ( .A({ _08047_, _saxi_register_fsm[0], _21724_, _21756_ }), .Y(_21692_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30760_ ( .A({ _08047_, _saxi_register_fsm[0], _21713_, _21745_ }), .Y(_21681_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30761_ ( .A({ _08048_, _saxi_register_fsm[1], _08056_, _saxi_register_fsm[0] }), .Y(saxi_wready) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _30762_ ( .A({ saxi_wready, _08047_ }), .Y(_21944_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30763_ ( .A({ conv2d_8_prev_row_select[0], conv2d_8_prev_row_select[1] }), .Y(_04905_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30764_ ( .A(conv2d_8_prev_row_select), .Y(_04906_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30765_ ( .A({ __tmp_339_2[0], __tmp_339_2[1] }), .Y(_04907_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30766_ ( .A(__tmp_339_2), .Y(_04908_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30767_ ( .A({ __tmp_339_2[0], __tmp_339_2[1] }), .Y(_04909_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30768_ ( .A({ __tmp_359_2[0], __tmp_359_2[1] }), .Y(_04910_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30769_ ( .A(__tmp_359_2), .Y(_04911_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30770_ ( .A({ __tmp_359_2[0], __tmp_359_2[1] }), .Y(_04912_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30771_ ( .A({ __tmp_369_2[0], __tmp_369_2[1] }), .Y(_04913_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30772_ ( .A(__tmp_369_2), .Y(_04914_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30773_ ( .A({ __tmp_369_2[0], __tmp_369_2[1] }), .Y(_04915_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30774_ ( .A({ __tmp_379_2[0], __tmp_379_2[1] }), .Y(_04916_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30775_ ( .A(__tmp_379_2), .Y(_04917_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30776_ ( .A({ __tmp_379_2[0], __tmp_379_2[1] }), .Y(_04918_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30777_ ( .A({ __tmp_389_2[0], __tmp_389_2[1] }), .Y(_04919_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30778_ ( .A(__tmp_389_2), .Y(_04920_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30779_ ( .A({ __tmp_389_2[0], __tmp_389_2[1] }), .Y(_04921_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30780_ ( .A({ __tmp_399_2[0], __tmp_399_2[1] }), .Y(_04922_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30781_ ( .A(__tmp_399_2), .Y(_04923_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30782_ ( .A({ __tmp_399_2[0], __tmp_399_2[1] }), .Y(_04924_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30783_ ( .A({ __tmp_409_2[0], __tmp_409_2[1] }), .Y(_04925_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30784_ ( .A(__tmp_409_2), .Y(_04926_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30785_ ( .A({ __tmp_409_2[0], __tmp_409_2[1] }), .Y(_04927_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30786_ ( .A({ __tmp_419_2[0], __tmp_419_2[1] }), .Y(_04928_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30787_ ( .A(__tmp_419_2), .Y(_04929_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30788_ ( .A({ __tmp_419_2[0], __tmp_419_2[1] }), .Y(_04930_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30789_ ( .A({ __tmp_429_2[0], __tmp_429_2[1] }), .Y(_04931_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30790_ ( .A(__tmp_429_2), .Y(_04932_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30791_ ( .A({ __tmp_429_2[0], __tmp_429_2[1] }), .Y(_04933_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30792_ ( .A({ __tmp_439_2[0], __tmp_439_2[1] }), .Y(_04934_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30793_ ( .A(__tmp_439_2), .Y(_04935_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30794_ ( .A({ __tmp_439_2[0], __tmp_439_2[1] }), .Y(_04936_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30795_ ( .A({ __tmp_449_2[0], __tmp_449_2[1] }), .Y(_04937_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30796_ ( .A(__tmp_449_2), .Y(_04938_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30797_ ( .A({ __tmp_449_2[0], __tmp_449_2[1] }), .Y(_04939_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30798_ ( .A({ __tmp_459_2[0], __tmp_459_2[1] }), .Y(_04940_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30799_ ( .A(__tmp_459_2), .Y(_04941_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30800_ ( .A({ __tmp_459_2[0], __tmp_459_2[1] }), .Y(_04942_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30801_ ( .A({ __tmp_469_2[0], __tmp_469_2[1] }), .Y(_04943_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30802_ ( .A(__tmp_469_2), .Y(_04944_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30803_ ( .A({ __tmp_469_2[0], __tmp_469_2[1] }), .Y(_04945_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30804_ ( .A({ __tmp_479_2[0], __tmp_479_2[1] }), .Y(_04946_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30805_ ( .A(__tmp_479_2), .Y(_04947_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30806_ ( .A({ __tmp_479_2[0], __tmp_479_2[1] }), .Y(_04948_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30807_ ( .A({ __tmp_489_2[0], __tmp_489_2[1] }), .Y(_04949_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30808_ ( .A(__tmp_489_2), .Y(_04950_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30809_ ( .A({ __tmp_489_2[0], __tmp_489_2[1] }), .Y(_04951_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30810_ ( .A({ __tmp_499_2[0], __tmp_499_2[1] }), .Y(_04952_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30811_ ( .A(__tmp_499_2), .Y(_04953_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30812_ ( .A({ __tmp_499_2[0], __tmp_499_2[1] }), .Y(_04954_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30813_ ( .A({ __tmp_509_2[0], __tmp_509_2[1] }), .Y(_04955_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30814_ ( .A(__tmp_509_2), .Y(_04956_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30815_ ( .A({ __tmp_509_2[0], __tmp_509_2[1] }), .Y(_04957_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30816_ ( .A({ __tmp_519_2[0], __tmp_519_2[1] }), .Y(_04958_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30817_ ( .A(__tmp_519_2), .Y(_04959_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30818_ ( .A({ __tmp_519_2[0], __tmp_519_2[1] }), .Y(_04960_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30819_ ( .A({ __tmp_529_2[0], __tmp_529_2[1] }), .Y(_04961_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30820_ ( .A(__tmp_529_2), .Y(_04962_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30821_ ( .A({ __tmp_529_2[0], __tmp_529_2[1] }), .Y(_04963_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30822_ ( .A({ conv2d_8_row_select[0], conv2d_8_row_select[1] }), .Y(_04964_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30823_ ( .A(conv2d_8_row_select), .Y(_04965_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30824_ ( .A({ __tmp_865_2[0], __tmp_865_2[1] }), .Y(_04966_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30825_ ( .A(__tmp_865_2), .Y(_04967_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30826_ ( .A({ __tmp_865_2[0], __tmp_865_2[1] }), .Y(_04968_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30827_ ( .A({ __tmp_995_2[0], __tmp_995_2[1] }), .Y(_04969_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30828_ ( .A(__tmp_995_2), .Y(_04970_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30829_ ( .A({ __tmp_995_2[0], __tmp_995_2[1] }), .Y(_04971_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30830_ ( .A({ __tmp_1015_2[0], __tmp_1015_2[1] }), .Y(_04972_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30831_ ( .A(__tmp_1015_2), .Y(_04973_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30832_ ( .A({ __tmp_1015_2[0], __tmp_1015_2[1] }), .Y(_04974_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30833_ ( .A({ __tmp_1025_2[0], __tmp_1025_2[1] }), .Y(_04975_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30834_ ( .A(__tmp_1025_2), .Y(_04976_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30835_ ( .A({ __tmp_1025_2[0], __tmp_1025_2[1] }), .Y(_04977_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _30836_ ( .A({ _08058_, _tmp_5[0], _tmp_5[1] }), .Y(_04978_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _30837_ ( .A(_tmp_5[3:2]), .Y(_08058_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _30838_ ( .A({ _tmp_5[1], _08058_, _tmp_5[0] }), .Y(_04979_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30839_ ( .A({ _tmp_5[1:0], _08058_ }), .Y(_04980_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _30840_ ( .A({ _08059_, _tmp_5[1:0] }), .Y(_04981_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30841_ ( .A({ _tmp_5[2], _tmp_5[3] }), .Y(_08059_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _30842_ ( .A({ _08059_, _tmp_5[0], _tmp_5[1] }), .Y(_04982_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _30843_ ( .A({ _tmp_5[1], _08059_, _tmp_5[0] }), .Y(_04983_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30844_ ( .A({ _tmp_5[1:0], _08059_ }), .Y(_04984_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _30845_ ( .A({ _08060_, _tmp_5[1:0] }), .Y(_04985_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30846_ ( .A(_tmp_5[3:2]), .Y(_08060_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _30847_ ( .A({ _08060_, _tmp_5[0], _tmp_5[1] }), .Y(_04986_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _30848_ ( .A({ _tmp_5[1], _08060_, _tmp_5[0] }), .Y(_04987_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30849_ ( .A({ _tmp_5[1:0], _08060_ }), .Y(_04988_) );
  \$lut  #( .LUT(16'hefff), .WIDTH(4) ) _30850_ ( .A(_tmp_5), .Y(_04989_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _30851_ ( .A({ _tmp_5[2], _tmp_5[0], _tmp_5[3], _tmp_5[1] }), .Y(_04990_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30852_ ( .A({ _08062_, _08061_ }), .Y(_04991_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30853_ ( .A({ _stream_matmul_15_source_20_source_ram_sel[2], _stream_matmul_15_source_20_source_ram_sel[7:5] }), .Y(_08061_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30854_ ( .A({ _stream_matmul_15_source_20_source_ram_sel[4:3], _stream_matmul_15_source_20_source_ram_sel[1:0] }), .Y(_08062_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30855_ ( .A({ _08064_, _08063_ }), .Y(_04992_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30856_ ( .A({ _stream_conv2d_8_source_8_source_ram_sel[1], _stream_conv2d_8_source_8_source_ram_sel[7:5] }), .Y(_08063_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30857_ ( .A({ _stream_conv2d_8_source_8_source_ram_sel[4:2], _stream_conv2d_8_source_8_source_ram_sel[0] }), .Y(_08064_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30858_ ( .A({ _08066_, _08065_ }), .Y(_04993_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30859_ ( .A({ _stream_matmul_15_source_8_source_ram_sel[1], _stream_matmul_15_source_8_source_ram_sel[7:5] }), .Y(_08065_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30860_ ( .A({ _stream_matmul_15_source_8_source_ram_sel[4:2], _stream_matmul_15_source_8_source_ram_sel[0] }), .Y(_08066_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30861_ ( .A({ _08068_, _08067_ }), .Y(_04994_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30862_ ( .A({ _stream_conv2d_8_source_28_source_ram_sel[3:2], _stream_conv2d_8_source_28_source_ram_sel[7:6] }), .Y(_08067_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30863_ ( .A({ _stream_conv2d_8_source_28_source_ram_sel[5:4], _stream_conv2d_8_source_28_source_ram_sel[1:0] }), .Y(_08068_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30864_ ( .A({ _08070_, _08069_ }), .Y(_04995_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30865_ ( .A({ _stream_max_pool_serial_9_source_1_source_ram_sel[0], _stream_max_pool_serial_9_source_1_source_ram_sel[7:5] }), .Y(_08069_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30866_ ( .A(_stream_max_pool_serial_9_source_1_source_ram_sel[4:1]), .Y(_08070_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30867_ ( .A({ _08072_, _08071_ }), .Y(_04996_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30868_ ( .A({ _stream_conv2d_8_source_29_source_ram_sel[3:2], _stream_conv2d_8_source_29_source_ram_sel[0], _stream_conv2d_8_source_29_source_ram_sel[7] }), .Y(_08071_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30869_ ( .A({ _stream_conv2d_8_source_29_source_ram_sel[6:4], _stream_conv2d_8_source_29_source_ram_sel[1] }), .Y(_08072_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30870_ ( .A({ _08074_, _08073_ }), .Y(_04997_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30871_ ( .A({ _stream_matmul_15_source_19_source_ram_sel[1:0], _stream_matmul_15_source_19_source_ram_sel[7:6] }), .Y(_08073_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30872_ ( .A(_stream_matmul_15_source_19_source_ram_sel[5:2]), .Y(_08074_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30873_ ( .A({ _08076_, _08075_ }), .Y(_04998_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30874_ ( .A({ _stream_conv2d_8_source_30_source_ram_sel[3:1], _stream_conv2d_8_source_30_source_ram_sel[7] }), .Y(_08075_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30875_ ( .A({ _stream_conv2d_8_source_30_source_ram_sel[6:4], _stream_conv2d_8_source_30_source_ram_sel[0] }), .Y(_08076_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30876_ ( .A({ _08078_, _08077_ }), .Y(_04999_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30877_ ( .A(_stream_conv2d_8_source_31_source_ram_sel[3:0]), .Y(_08077_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30878_ ( .A(_stream_conv2d_8_source_31_source_ram_sel[7:4]), .Y(_08078_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30879_ ( .A({ _08080_, _08079_ }), .Y(_05000_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30880_ ( .A({ _stream_conv2d_8_source_32_source_ram_sel[4], _stream_conv2d_8_source_32_source_ram_sel[7:5] }), .Y(_08079_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30881_ ( .A(_stream_conv2d_8_source_32_source_ram_sel[3:0]), .Y(_08080_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30882_ ( .A({ _08082_, _08081_ }), .Y(_05001_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30883_ ( .A({ _stream_conv2d_8_source_33_source_ram_sel[4], _stream_conv2d_8_source_33_source_ram_sel[0], _stream_conv2d_8_source_33_source_ram_sel[7:6] }), .Y(_08081_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30884_ ( .A({ _stream_conv2d_8_source_33_source_ram_sel[5], _stream_conv2d_8_source_33_source_ram_sel[3:1] }), .Y(_08082_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30885_ ( .A({ _08084_, _08083_ }), .Y(_05002_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30886_ ( .A({ _stream_conv2d_8_source_34_source_ram_sel[4], _stream_conv2d_8_source_34_source_ram_sel[1], _stream_conv2d_8_source_34_source_ram_sel[7:6] }), .Y(_08083_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30887_ ( .A({ _stream_conv2d_8_source_34_source_ram_sel[5], _stream_conv2d_8_source_34_source_ram_sel[3:2], _stream_conv2d_8_source_34_source_ram_sel[0] }), .Y(_08084_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30888_ ( .A({ _08086_, _08085_ }), .Y(_05003_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30889_ ( .A({ _stream_conv2d_8_source_35_source_ram_sel[4], _stream_conv2d_8_source_35_source_ram_sel[1:0], _stream_conv2d_8_source_35_source_ram_sel[7] }), .Y(_08085_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30890_ ( .A({ _stream_conv2d_8_source_35_source_ram_sel[6:5], _stream_conv2d_8_source_35_source_ram_sel[3:2] }), .Y(_08086_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30891_ ( .A({ _08088_, _08087_ }), .Y(_05004_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30892_ ( .A({ _stream_conv2d_8_source_36_source_ram_sel[4], _stream_conv2d_8_source_36_source_ram_sel[2], _stream_conv2d_8_source_36_source_ram_sel[7:6] }), .Y(_08087_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30893_ ( .A({ _stream_conv2d_8_source_36_source_ram_sel[5], _stream_conv2d_8_source_36_source_ram_sel[3], _stream_conv2d_8_source_36_source_ram_sel[1:0] }), .Y(_08088_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30894_ ( .A({ _08090_, _08089_ }), .Y(_05005_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30895_ ( .A({ _stream_conv2d_8_source_19_source_ram_sel[1:0], _stream_conv2d_8_source_19_source_ram_sel[7:6] }), .Y(_08089_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30896_ ( .A(_stream_conv2d_8_source_19_source_ram_sel[5:2]), .Y(_08090_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30897_ ( .A({ _08092_, _08091_ }), .Y(_05006_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30898_ ( .A({ _stream_conv2d_8_source_20_source_ram_sel[2], _stream_conv2d_8_source_20_source_ram_sel[7:5] }), .Y(_08091_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30899_ ( .A({ _stream_conv2d_8_source_20_source_ram_sel[4:3], _stream_conv2d_8_source_20_source_ram_sel[1:0] }), .Y(_08092_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30900_ ( .A({ _08094_, _08093_ }), .Y(_05007_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30901_ ( .A({ _stream_conv2d_8_source_21_source_ram_sel[2], _stream_conv2d_8_source_21_source_ram_sel[0], _stream_conv2d_8_source_21_source_ram_sel[7:6] }), .Y(_08093_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30902_ ( .A({ _stream_conv2d_8_source_21_source_ram_sel[5:3], _stream_conv2d_8_source_21_source_ram_sel[1] }), .Y(_08094_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30903_ ( .A({ _08096_, _08095_ }), .Y(_05008_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30904_ ( .A({ _stream_conv2d_8_source_22_source_ram_sel[2:1], _stream_conv2d_8_source_22_source_ram_sel[7:6] }), .Y(_08095_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30905_ ( .A({ _stream_conv2d_8_source_22_source_ram_sel[5:3], _stream_conv2d_8_source_22_source_ram_sel[0] }), .Y(_08096_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30906_ ( .A({ _08098_, _08097_ }), .Y(_05009_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30907_ ( .A({ _stream_conv2d_8_source_23_source_ram_sel[2:0], _stream_conv2d_8_source_23_source_ram_sel[7] }), .Y(_08097_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30908_ ( .A(_stream_conv2d_8_source_23_source_ram_sel[6:3]), .Y(_08098_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30909_ ( .A({ _08100_, _08099_ }), .Y(_05010_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30910_ ( .A({ _stream_conv2d_8_source_24_source_ram_sel[3], _stream_conv2d_8_source_24_source_ram_sel[7:5] }), .Y(_08099_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30911_ ( .A({ _stream_conv2d_8_source_24_source_ram_sel[4], _stream_conv2d_8_source_24_source_ram_sel[2:0] }), .Y(_08100_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30912_ ( .A({ _08102_, _08101_ }), .Y(_05011_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30913_ ( .A({ _stream_conv2d_8_source_25_source_ram_sel[3], _stream_conv2d_8_source_25_source_ram_sel[0], _stream_conv2d_8_source_25_source_ram_sel[7:6] }), .Y(_08101_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30914_ ( .A({ _stream_conv2d_8_source_25_source_ram_sel[5:4], _stream_conv2d_8_source_25_source_ram_sel[2:1] }), .Y(_08102_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30915_ ( .A({ _08104_, _08103_ }), .Y(_05012_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30916_ ( .A({ _stream_conv2d_8_source_26_source_ram_sel[3], _stream_conv2d_8_source_26_source_ram_sel[1], _stream_conv2d_8_source_26_source_ram_sel[7:6] }), .Y(_08103_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30917_ ( .A({ _stream_conv2d_8_source_26_source_ram_sel[5:4], _stream_conv2d_8_source_26_source_ram_sel[2], _stream_conv2d_8_source_26_source_ram_sel[0] }), .Y(_08104_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30918_ ( .A({ _08106_, _08105_ }), .Y(_05013_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30919_ ( .A({ _stream_conv2d_8_source_27_source_ram_sel[3], _stream_conv2d_8_source_27_source_ram_sel[1:0], _stream_conv2d_8_source_27_source_ram_sel[7] }), .Y(_08105_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30920_ ( .A({ _stream_conv2d_8_source_27_source_ram_sel[6:4], _stream_conv2d_8_source_27_source_ram_sel[2] }), .Y(_08106_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30921_ ( .A({ _08108_, _08107_ }), .Y(_05014_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30922_ ( .A({ _stream_conv2d_8_source_6_source_ram_sel[0], _stream_conv2d_8_source_6_source_ram_sel[7:5] }), .Y(_08107_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30923_ ( .A(_stream_conv2d_8_source_6_source_ram_sel[4:1]), .Y(_08108_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30924_ ( .A({ _08110_, _08109_ }), .Y(_05015_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30925_ ( .A({ _stream_matmul_15_source_6_source_ram_sel[0], _stream_matmul_15_source_6_source_ram_sel[7:5] }), .Y(_08109_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30926_ ( .A(_stream_matmul_15_source_6_source_ram_sel[4:1]), .Y(_08110_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _30927_ ( .A({ _08111_, cparam_conv2d_8_bias_num[2:1] }), .Y(_05016_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30928_ ( .A({ cparam_conv2d_8_bias_num[0], cparam_conv2d_8_bias_num[4:3] }), .Y(_08111_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30929_ ( .A({ _08117_, _08112_ }), .Y(_05873_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30930_ ( .A({ _08116_, _08115_, _08114_, _08113_ }), .Y(_08112_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30931_ ( .A(_saxi_register_4[23:20]), .Y(_08113_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30932_ ( .A(_saxi_register_4[19:16]), .Y(_08114_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30933_ ( .A(_saxi_register_4[31:28]), .Y(_08115_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30934_ ( .A(_saxi_register_4[27:24]), .Y(_08116_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30935_ ( .A({ _08121_, _08120_, _08119_, _08118_ }), .Y(_08117_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30936_ ( .A(_saxi_register_4[7:4]), .Y(_08118_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30937_ ( .A(_saxi_register_4[3:0]), .Y(_08119_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30938_ ( .A(_saxi_register_4[15:12]), .Y(_08120_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30939_ ( .A(_saxi_register_4[11:8]), .Y(_08121_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30940_ ( .A({ _08127_, _08122_ }), .Y(_17710_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30941_ ( .A({ _08126_, _08125_, _08124_, _08123_ }), .Y(_08122_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30942_ ( .A({ _21960_, _21959_, _21958_, _21957_ }), .Y(_08123_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30943_ ( .A({ _21955_, _21954_, _21953_, _21952_ }), .Y(_08124_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30944_ ( .A({ _21969_, _21968_, _21966_, _21965_ }), .Y(_08125_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30945_ ( .A({ _21964_, _21963_, _21962_, _21961_ }), .Y(_08126_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30946_ ( .A({ _08131_, _08130_, _08129_, _08128_ }), .Y(_08127_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30947_ ( .A({ _21974_, _21973_, _21972_, _21971_ }), .Y(_08128_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30948_ ( .A({ _21970_, _21967_, _21956_, _21945_ }), .Y(_08129_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30949_ ( .A({ _21951_, _21950_, _21949_, _21948_ }), .Y(_08130_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30950_ ( .A({ _21947_, _21946_, _21976_, _21975_ }), .Y(_08131_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30951_ ( .A({ _08137_, _08132_ }), .Y(_17645_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30952_ ( .A({ _08136_, _08135_, _08134_, _08133_ }), .Y(_08132_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30953_ ( .A({ _21992_, _21991_, _21990_, _21989_ }), .Y(_08133_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30954_ ( .A({ _21987_, _21986_, _21985_, _21984_ }), .Y(_08134_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30955_ ( .A({ _22001_, _22000_, _21998_, _21997_ }), .Y(_08135_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30956_ ( .A({ _21996_, _21995_, _21994_, _21993_ }), .Y(_08136_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30957_ ( .A({ _08141_, _08140_, _08139_, _08138_ }), .Y(_08137_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30958_ ( .A({ _22006_, _22005_, _22004_, _22003_ }), .Y(_08138_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30959_ ( .A({ _22002_, _21999_, _21988_, _21977_ }), .Y(_08139_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30960_ ( .A({ _21983_, _21982_, _21981_, _21980_ }), .Y(_08140_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30961_ ( .A({ _21979_, _21978_, _22008_, _22007_ }), .Y(_08141_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30962_ ( .A({ conv2d_8_col_select[0], conv2d_8_col_select[1] }), .Y(_05017_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30963_ ( .A(conv2d_8_col_select), .Y(_05018_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30964_ ( .A({ _08147_, _08142_ }), .Y(_17548_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30965_ ( .A({ _08146_, _08145_, _08144_, _08143_ }), .Y(_08142_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30966_ ( .A({ _22024_, _22023_, _22022_, _22021_ }), .Y(_08143_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30967_ ( .A({ _22019_, _22018_, _22017_, _22016_ }), .Y(_08144_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30968_ ( .A({ _22033_, _22032_, _22030_, _22029_ }), .Y(_08145_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30969_ ( .A({ _22028_, _22027_, _22026_, _22025_ }), .Y(_08146_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30970_ ( .A({ _08151_, _08150_, _08149_, _08148_ }), .Y(_08147_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30971_ ( .A({ _22038_, _22037_, _22036_, _22035_ }), .Y(_08148_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30972_ ( .A({ _22034_, _22031_, _22020_, _22009_ }), .Y(_08149_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30973_ ( .A({ _22015_, _22014_, _22013_, _22012_ }), .Y(_08150_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30974_ ( .A({ _22011_, _22010_, _22040_, _22039_ }), .Y(_08151_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30975_ ( .A({ _stream_matmul_15_source_20_source_pat_fsm_3[1], _07089_ }), .Y(_05019_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30976_ ( .A({ _stream_matmul_15_source_19_source_pat_fsm_2[1], _07043_ }), .Y(_05022_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30977_ ( .A({ _stream_matmul_15_source_8_source_pat_fsm_1[1], _07020_ }), .Y(_05024_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30978_ ( .A({ _stream_matmul_15_source_6_source_pat_fsm_0[1], _06995_ }), .Y(_05026_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30979_ ( .A({ _08161_, _08160_, _08157_, _08152_ }), .Y(_05029_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30980_ ( .A({ _08156_, _08155_, _08154_, _08153_ }), .Y(_08152_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30981_ ( .A(_d1_control_matmul_15[23:20]), .Y(_08153_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30982_ ( .A(_d1_control_matmul_15[19:16]), .Y(_08154_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30983_ ( .A(_d1_control_matmul_15[31:28]), .Y(_08155_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30984_ ( .A(_d1_control_matmul_15[27:24]), .Y(_08156_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30985_ ( .A({ _08159_, _08158_ }), .Y(_08157_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30986_ ( .A(_d1_control_matmul_15[15:12]), .Y(_08158_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30987_ ( .A(_d1_control_matmul_15[11:8]), .Y(_08159_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30988_ ( .A({ _d1_control_matmul_15[5], _d1_control_matmul_15[1:0], _d1_control_matmul_15[4] }), .Y(_08160_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30989_ ( .A({ _d1_control_matmul_15[7:6], _d1_control_matmul_15[2], _d1_control_matmul_15[3] }), .Y(_08161_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30990_ ( .A({ _08163_, _08152_, _08162_ }), .Y(_05031_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30991_ ( .A({ _d1_control_matmul_15[2:1], _08157_, _d1_control_matmul_15[0] }), .Y(_08162_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30992_ ( .A({ _08164_, _d1_control_matmul_15[4:3] }), .Y(_08163_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _30993_ ( .A(_d1_control_matmul_15[7:5]), .Y(_08164_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30994_ ( .A({ _08165_, _08162_ }), .Y(_05032_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30995_ ( .A({ _d1_control_matmul_15[3], _08166_, _08152_ }), .Y(_08165_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30996_ ( .A({ _08164_, _d1_control_matmul_15[4] }), .Y(_08166_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30997_ ( .A({ _08167_, _08165_ }), .Y(_05033_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30998_ ( .A({ _08157_, _d1_control_matmul_15[2:0] }), .Y(_08167_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30999_ ( .A({ _08168_, _08166_, _08157_, _08152_ }), .Y(_05034_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31000_ ( .A({ _d1_control_matmul_15[0], _d1_control_matmul_15[1], _d1_control_matmul_15[2], _d1_control_matmul_15[3] }), .Y(_08168_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31001_ ( .A({ _06586_, _06601_ }), .Y(_05036_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31002_ ( .A({ _06582_, _06584_ }), .Y(_05037_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31003_ ( .A({ _stream_max_pool_serial_9_source_1_source_pat_fsm_0[1], _06533_ }), .Y(_05044_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31004_ ( .A({ _06497_, _06490_ }), .Y(_05047_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _31005_ ( .A({ _08178_, _08173_, _08169_ }), .Y(_05049_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31006_ ( .A({ _d1_control_max_pool_serial_9[0], _d1_control_max_pool_serial_9[1], _08170_, _d1_control_max_pool_serial_9[2] }), .Y(_08169_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31007_ ( .A({ _08172_, _08171_ }), .Y(_08170_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31008_ ( .A(_d1_control_max_pool_serial_9[15:12]), .Y(_08171_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31009_ ( .A(_d1_control_max_pool_serial_9[11:8]), .Y(_08172_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31010_ ( .A({ _08177_, _08176_, _08175_, _08174_ }), .Y(_08173_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31011_ ( .A(_d1_control_max_pool_serial_9[23:20]), .Y(_08174_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31012_ ( .A(_d1_control_max_pool_serial_9[19:16]), .Y(_08175_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31013_ ( .A(_d1_control_max_pool_serial_9[31:28]), .Y(_08176_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31014_ ( .A(_d1_control_max_pool_serial_9[27:24]), .Y(_08177_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _31015_ ( .A({ _08179_, _d1_control_max_pool_serial_9[7:6] }), .Y(_08178_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _31016_ ( .A({ _d1_control_max_pool_serial_9[4], _d1_control_max_pool_serial_9[5], _d1_control_max_pool_serial_9[3] }), .Y(_08179_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31017_ ( .A({ _d1_control_max_pool_serial_9[3], _08180_, _08173_, _08169_ }), .Y(_05050_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31018_ ( .A({ _d1_control_max_pool_serial_9[7:6], _d1_control_max_pool_serial_9[4], _d1_control_max_pool_serial_9[5] }), .Y(_08180_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31019_ ( .A({ _08181_, _08180_, _08170_, _08173_ }), .Y(_05051_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31020_ ( .A({ _d1_control_max_pool_serial_9[0], _d1_control_max_pool_serial_9[2:1], _d1_control_max_pool_serial_9[3] }), .Y(_08181_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _31021_ ( .A({ _08183_, _08182_, _05875_ }), .Y(_05052_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31022_ ( .A(control_max_pool_serial_9[3:2]), .Y(_08182_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31023_ ( .A({ control_max_pool_serial_9[0], control_max_pool_serial_9[1] }), .Y(_08183_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31024_ ( .A({ control_max_pool_serial_9[1:0], _05887_, _05875_ }), .Y(_05053_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31025_ ( .A({ control_max_pool_serial_9[1:0], _08182_, _05886_ }), .Y(_05054_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _31026_ ( .A({ _08183_, _05885_, _05886_ }), .Y(_05056_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31027_ ( .A({ _08189_, _08184_ }), .Y(_05057_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31028_ ( .A({ _08188_, _08187_, _08186_, _08185_ }), .Y(_08184_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31029_ ( .A(_d1__maxi_write_fsm[24:21]), .Y(_08185_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31030_ ( .A(_d1__maxi_write_fsm[20:17]), .Y(_08186_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31031_ ( .A({ _d1__maxi_write_fsm[2], _d1__maxi_write_fsm[31:29] }), .Y(_08187_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31032_ ( .A(_d1__maxi_write_fsm[28:25]), .Y(_08188_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31033_ ( .A({ _08193_, _08192_, _08191_, _08190_ }), .Y(_08189_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31034_ ( .A(_d1__maxi_write_fsm[8:5]), .Y(_08190_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31035_ ( .A({ _d1__maxi_write_fsm[4:3], _d1__maxi_write_fsm[1:0] }), .Y(_08191_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31036_ ( .A(_d1__maxi_write_fsm[16:13]), .Y(_08192_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31037_ ( .A(_d1__maxi_write_fsm[12:9]), .Y(_08193_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _31038_ ( .A({ _maxi_write_fsm[2], _08194_, _maxi_write_fsm[3] }), .Y(_05058_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31039_ ( .A({ _08202_, _08195_, _maxi_write_fsm[1:0] }), .Y(_08194_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31040_ ( .A({ _08201_, _08196_ }), .Y(_08195_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31041_ ( .A({ _08200_, _08199_, _08198_, _08197_ }), .Y(_08196_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31042_ ( .A(_maxi_write_fsm[23:20]), .Y(_08197_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31043_ ( .A(_maxi_write_fsm[19:16]), .Y(_08198_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31044_ ( .A(_maxi_write_fsm[31:28]), .Y(_08199_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31045_ ( .A(_maxi_write_fsm[27:24]), .Y(_08200_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31046_ ( .A(_maxi_write_fsm[7:4]), .Y(_08201_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31047_ ( .A({ _08204_, _08203_ }), .Y(_08202_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31048_ ( .A(_maxi_write_fsm[15:12]), .Y(_08203_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31049_ ( .A(_maxi_write_fsm[11:8]), .Y(_08204_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _31050_ ( .A({ _08205_, _maxi_write_fsm[2], _maxi_write_fsm[3] }), .Y(_05059_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31051_ ( .A({ _08195_, _maxi_write_fsm[0], _08202_, _maxi_write_fsm[1] }), .Y(_08205_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31052_ ( .A({ _stream_conv2d_8_source_36_source_pat_fsm_19[1], _07784_ }), .Y(_05060_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31053_ ( .A({ _stream_conv2d_8_source_35_source_pat_fsm_18[1], _07772_ }), .Y(_05062_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31054_ ( .A({ _stream_conv2d_8_source_34_source_pat_fsm_17[1], _07688_ }), .Y(_05063_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31055_ ( .A({ _stream_conv2d_8_source_33_source_pat_fsm_16[1], _07676_ }), .Y(_05065_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31056_ ( .A({ _08215_, _08214_, _08211_, _08206_ }), .Y(_05068_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31057_ ( .A({ _08210_, _08209_, _08208_, _08207_ }), .Y(_08206_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31058_ ( .A(_stream_conv2d_8_source_32_source_pat_fsm_15[23:20]), .Y(_08207_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31059_ ( .A(_stream_conv2d_8_source_32_source_pat_fsm_15[19:16]), .Y(_08208_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31060_ ( .A(_stream_conv2d_8_source_32_source_pat_fsm_15[31:28]), .Y(_08209_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31061_ ( .A(_stream_conv2d_8_source_32_source_pat_fsm_15[27:24]), .Y(_08210_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31062_ ( .A({ _08213_, _08212_ }), .Y(_08211_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31063_ ( .A(_stream_conv2d_8_source_32_source_pat_fsm_15[15:12]), .Y(_08212_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31064_ ( .A(_stream_conv2d_8_source_32_source_pat_fsm_15[11:8]), .Y(_08213_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31065_ ( .A(_stream_conv2d_8_source_32_source_pat_fsm_15[7:4]), .Y(_08214_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31066_ ( .A({ _stream_conv2d_8_source_32_source_pat_fsm_15[1], _stream_conv2d_8_source_32_source_pat_fsm_15[3:2], _stream_conv2d_8_source_32_source_pat_fsm_15[0] }), .Y(_08215_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31067_ ( .A({ _stream_conv2d_8_source_32_source_pat_fsm_15[0], _08216_ }), .Y(_05069_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31068_ ( .A({ _08217_, _08211_, _08206_ }), .Y(_08216_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31069_ ( .A({ _08214_, _stream_conv2d_8_source_32_source_pat_fsm_15[3:1] }), .Y(_08217_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31070_ ( .A({ _stream_conv2d_8_source_31_source_pat_fsm_14[1], _07067_ }), .Y(_05070_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31071_ ( .A({ _stream_conv2d_8_source_30_source_pat_fsm_13[0], _07032_ }), .Y(_05073_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31072_ ( .A({ _stream_conv2d_8_source_29_source_pat_fsm_12[0], _07148_ }), .Y(_05075_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31073_ ( .A({ _stream_conv2d_8_source_28_source_pat_fsm_11[0], _07441_ }), .Y(_05077_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31074_ ( .A({ _stream_conv2d_8_source_27_source_pat_fsm_10[0], _07127_ }), .Y(_05079_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31075_ ( .A({ _stream_conv2d_8_source_26_source_pat_fsm_9[0], _06555_ }), .Y(_05081_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31076_ ( .A({ _stream_conv2d_8_source_25_source_pat_fsm_8[0], _07078_ }), .Y(_05083_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31077_ ( .A({ _stream_conv2d_8_source_24_source_pat_fsm_7[0], _07358_ }), .Y(_05085_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31078_ ( .A({ _stream_conv2d_8_source_23_source_pat_fsm_6[0], _07402_ }), .Y(_05087_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31079_ ( .A({ _stream_conv2d_8_source_22_source_pat_fsm_5[0], _07369_ }), .Y(_05089_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31080_ ( .A({ _stream_conv2d_8_source_21_source_pat_fsm_4[0], _07347_ }), .Y(_05091_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31081_ ( .A({ _stream_conv2d_8_source_20_source_pat_fsm_3[0], _07335_ }), .Y(_05093_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31082_ ( .A({ _stream_conv2d_8_source_19_source_pat_fsm_2[0], _07056_ }), .Y(_05095_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31083_ ( .A({ _stream_conv2d_8_source_8_source_pat_fsm_1[0], _07761_ }), .Y(_05097_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31084_ ( .A({ _stream_conv2d_8_source_6_source_pat_fsm_0[0], _07750_ }), .Y(_05099_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31085_ ( .A({ _08226_, _08218_ }), .Y(_05103_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31086_ ( .A({ _08219_, _08225_, _08224_, _d1__maxi_read_fsm[3] }), .Y(_08218_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31087_ ( .A({ _08223_, _08222_, _08221_, _08220_ }), .Y(_08219_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31088_ ( .A({ _d1__maxi_read_fsm[22:21], _d1__maxi_read_fsm[19], _d1__maxi_read_fsm[16] }), .Y(_08220_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31089_ ( .A({ _d1__maxi_read_fsm[31], _d1__maxi_read_fsm[28], _d1__maxi_read_fsm[26:25] }), .Y(_08221_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31090_ ( .A({ _d1__maxi_read_fsm[23], _d1__maxi_read_fsm[20], _d1__maxi_read_fsm[18:17] }), .Y(_08222_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31091_ ( .A({ _d1__maxi_read_fsm[30:29], _d1__maxi_read_fsm[27], _d1__maxi_read_fsm[24] }), .Y(_08223_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31092_ ( .A({ _d1__maxi_read_fsm[15], _d1__maxi_read_fsm[13], _d1__maxi_read_fsm[11], _d1__maxi_read_fsm[9] }), .Y(_08224_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31093_ ( .A({ _d1__maxi_read_fsm[14], _d1__maxi_read_fsm[12], _d1__maxi_read_fsm[10], _d1__maxi_read_fsm[8] }), .Y(_08225_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31094_ ( .A({ _d1__maxi_read_fsm[2], _08227_, _d1__maxi_read_fsm[1:0] }), .Y(_08226_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31095_ ( .A(_d1__maxi_read_fsm[7:4]), .Y(_08227_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31096_ ( .A({ _08228_, _08218_ }), .Y(_05104_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31097_ ( .A({ _08227_, _d1__maxi_read_fsm[1:0], _d1__maxi_read_fsm[2] }), .Y(_08228_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _31098_ ( .A({ _d1_control_conv2d_8[5], _08238_, _08229_ }), .Y(_05108_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31099_ ( .A({ _d1_control_conv2d_8[4], _08235_, _08230_ }), .Y(_08229_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31100_ ( .A({ _08234_, _08233_, _08232_, _08231_ }), .Y(_08230_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31101_ ( .A(_d1_control_conv2d_8[23:20]), .Y(_08231_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31102_ ( .A(_d1_control_conv2d_8[19:16]), .Y(_08232_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31103_ ( .A(_d1_control_conv2d_8[31:28]), .Y(_08233_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31104_ ( .A(_d1_control_conv2d_8[27:24]), .Y(_08234_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31105_ ( .A({ _08237_, _08236_, _d1_control_conv2d_8[7:6] }), .Y(_08235_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31106_ ( .A(_d1_control_conv2d_8[15:12]), .Y(_08236_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31107_ ( .A(_d1_control_conv2d_8[11:8]), .Y(_08237_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _31108_ ( .A({ _08239_, _d1_control_conv2d_8[2], _d1_control_conv2d_8[3] }), .Y(_08238_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31109_ ( .A({ _d1_control_conv2d_8[0], _d1_control_conv2d_8[1] }), .Y(_08239_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _31110_ ( .A({ _08240_, _d1_control_conv2d_8[1:0] }), .Y(_05109_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31111_ ( .A({ _08242_, _08241_ }), .Y(_08240_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31112_ ( .A({ _08235_, _d1_control_conv2d_8[4] }), .Y(_08241_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31113_ ( .A({ _d1_control_conv2d_8[2], _d1_control_conv2d_8[5], _08230_, _d1_control_conv2d_8[3] }), .Y(_08242_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _31114_ ( .A({ _d1_control_conv2d_8[0], _08240_, _d1_control_conv2d_8[1] }), .Y(_05110_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31115_ ( .A({ _d1_control_conv2d_8[2], _d1_control_conv2d_8[3], _08244_, _08243_ }), .Y(_05111_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31116_ ( .A({ _08229_, _d1_control_conv2d_8[5] }), .Y(_08243_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31117_ ( .A({ _d1_control_conv2d_8[0], _d1_control_conv2d_8[1] }), .Y(_08244_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31118_ ( .A({ _08245_, _08243_ }), .Y(_05112_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31119_ ( .A({ _d1_control_conv2d_8[2:1], _d1_control_conv2d_8[3], _d1_control_conv2d_8[0] }), .Y(_08245_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _31120_ ( .A({ _08243_, _d1_control_conv2d_8[3], _08239_, _d1_control_conv2d_8[2] }), .Y(_05113_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _31121_ ( .A({ _d1_control_conv2d_8[2], _08243_, _08244_, _d1_control_conv2d_8[3] }), .Y(_05114_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31122_ ( .A({ _d1_control_conv2d_8[2], _d1_control_conv2d_8[3], _08244_, _08246_ }), .Y(_05115_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31123_ ( .A({ _08241_, _08230_, _d1_control_conv2d_8[5] }), .Y(_08246_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31124_ ( .A({ _08245_, _08246_ }), .Y(_05116_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _31125_ ( .A({ _08246_, _d1_control_conv2d_8[3], _08239_, _d1_control_conv2d_8[2] }), .Y(_05117_) );
  \$lut  #( .LUT(16'hefff), .WIDTH(4) ) _31126_ ( .A({ _08244_, _08246_, _d1_control_conv2d_8[2], _d1_control_conv2d_8[3] }), .Y(_05118_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31127_ ( .A({ _05907_, _06348_ }), .Y(_05120_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31128_ ( .A({ _05926_, _06342_ }), .Y(_05123_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31129_ ( .A({ _05915_, _06391_ }), .Y(_05128_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31130_ ( .A({ _05904_, _06391_ }), .Y(_05129_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31131_ ( .A({ _05949_, _06391_ }), .Y(_05131_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31132_ ( .A({ _07939_, _07933_ }), .Y(_05133_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31133_ ( .A({ _07807_, _07933_ }), .Y(_05134_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31134_ ( .A({ _07840_, _07797_ }), .Y(_05135_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31135_ ( .A({ _07843_, _07797_ }), .Y(_05136_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31136_ ( .A({ _07926_, _07797_ }), .Y(_05137_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31137_ ( .A({ _07928_, _07797_ }), .Y(_05138_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31138_ ( .A({ _07819_, _07797_ }), .Y(_05139_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31139_ ( .A({ _07822_, _07797_ }), .Y(_05140_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31140_ ( .A({ _07840_, _07815_ }), .Y(_05147_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31141_ ( .A({ _07928_, _07815_ }), .Y(_05148_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31142_ ( .A({ _07922_, _07815_ }), .Y(_05149_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31143_ ( .A({ _07807_, _07815_ }), .Y(_05150_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _31144_ ( .A({ _05132_, _05909_ }), .Y(_04700_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31145_ ( .A({ _15508_, _07795_, _15476_, _05061_ }), .Y(_15444_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31146_ ( .A({ _15509_, _07795_, _15477_, _05061_ }), .Y(_15445_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31147_ ( .A({ _15510_, _07795_, _15478_, _05061_ }), .Y(_15446_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31148_ ( .A({ _15512_, _07795_, _15480_, _05061_ }), .Y(_15448_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31149_ ( .A({ _15513_, _07795_, _15481_, _05061_ }), .Y(_15449_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31150_ ( .A({ _15514_, _07795_, _15482_, _05061_ }), .Y(_15450_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31151_ ( .A({ _15515_, _07795_, _15483_, _05061_ }), .Y(_15451_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31152_ ( .A({ _15516_, _07795_, _15484_, _05061_ }), .Y(_15452_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31153_ ( .A({ _15517_, _07795_, _15485_, _05061_ }), .Y(_15453_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31154_ ( .A({ _15518_, _07795_, _15486_, _05061_ }), .Y(_15454_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31155_ ( .A({ _15519_, _07795_, _15487_, _05061_ }), .Y(_15455_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31156_ ( .A({ _15520_, _07795_, _15488_, _05061_ }), .Y(_15456_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31157_ ( .A({ _15521_, _07795_, _15489_, _05061_ }), .Y(_15457_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31158_ ( .A({ _15523_, _07795_, _15491_, _05061_ }), .Y(_15459_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _31159_ ( .A({ _15524_, _07795_, _15492_, _05061_ }), .Y(_15460_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31160_ ( .A({ _08255_, _08254_, _08249_, _08247_ }), .Y(_21900_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31161_ ( .A({ _08248_, _stream_conv2d_8_sink_37_sink_fsm_20[31:29] }), .Y(_08247_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31162_ ( .A(_stream_conv2d_8_sink_37_sink_fsm_20[28:25]), .Y(_08248_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31163_ ( .A({ _08253_, _08252_, _08251_, _08250_ }), .Y(_08249_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31164_ ( .A(_stream_conv2d_8_sink_37_sink_fsm_20[8:5]), .Y(_08250_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31165_ ( .A(_stream_conv2d_8_sink_37_sink_fsm_20[4:1]), .Y(_08251_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31166_ ( .A(_stream_conv2d_8_sink_37_sink_fsm_20[16:13]), .Y(_08252_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31167_ ( .A(_stream_conv2d_8_sink_37_sink_fsm_20[12:9]), .Y(_08253_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31168_ ( .A(_stream_conv2d_8_sink_37_sink_fsm_20[24:21]), .Y(_08254_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31169_ ( .A(_stream_conv2d_8_sink_37_sink_fsm_20[20:17]), .Y(_08255_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31170_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15340_, _15404_ }), .Y(_15372_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31171_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15351_, _15415_ }), .Y(_15383_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31172_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15362_, _15426_ }), .Y(_15394_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31173_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15365_, _15429_ }), .Y(_15397_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31174_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15366_, _15430_ }), .Y(_15398_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31175_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15367_, _15431_ }), .Y(_15399_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31176_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15368_, _15432_ }), .Y(_15400_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31177_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15369_, _15433_ }), .Y(_15401_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31178_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15370_, _15434_ }), .Y(_15402_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31179_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15371_, _15435_ }), .Y(_15403_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31180_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15341_, _15405_ }), .Y(_15373_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31181_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15342_, _15406_ }), .Y(_15374_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31182_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15343_, _15407_ }), .Y(_15375_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31183_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15344_, _15408_ }), .Y(_15376_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31184_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15345_, _15409_ }), .Y(_15377_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31185_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15346_, _15410_ }), .Y(_15378_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31186_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15347_, _15411_ }), .Y(_15379_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31187_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15348_, _15412_ }), .Y(_15380_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31188_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15349_, _15413_ }), .Y(_15381_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31189_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15350_, _15414_ }), .Y(_15382_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31190_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15352_, _15416_ }), .Y(_15384_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31191_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15353_, _15417_ }), .Y(_15385_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31192_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15354_, _15418_ }), .Y(_15386_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31193_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15355_, _15419_ }), .Y(_15387_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31194_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15356_, _15420_ }), .Y(_15388_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31195_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15357_, _15421_ }), .Y(_15389_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31196_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15358_, _15422_ }), .Y(_15390_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31197_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15359_, _15423_ }), .Y(_15391_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31198_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15360_, _15424_ }), .Y(_15392_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31199_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15361_, _15425_ }), .Y(_15393_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31200_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15363_, _15427_ }), .Y(_15395_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31201_ ( .A({ _21900_, _stream_conv2d_8_sink_37_sink_fsm_20[0], _15364_, _15428_ }), .Y(_15396_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31202_ ( .A({ _08257_, _08256_ }), .Y(_21898_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _31203_ ( .A({ _08194_, _maxi_write_fsm[2], _maxi_write_fsm[3] }), .Y(_08256_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31204_ ( .A({ _maxi_write_fsm[0], _08196_, _08258_ }), .Y(_08257_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31205_ ( .A({ _08259_, _08202_ }), .Y(_08258_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31206_ ( .A({ _08201_, _maxi_write_fsm[1], _maxi_write_fsm[2], _maxi_write_fsm[3] }), .Y(_08259_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31207_ ( .A({ _15180_, _08256_, _08257_, _15116_ }), .Y(_15148_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31208_ ( .A({ _15191_, _08256_, _08257_, _15127_ }), .Y(_15159_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31209_ ( .A({ _15202_, _08256_, _08257_, _15138_ }), .Y(_15170_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31210_ ( .A({ _15205_, _08256_, _08257_, _15141_ }), .Y(_15173_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31211_ ( .A({ _15206_, _08256_, _08257_, _15142_ }), .Y(_15174_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31212_ ( .A({ _15207_, _08256_, _08257_, _15143_ }), .Y(_15175_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31213_ ( .A({ _15208_, _08256_, _08257_, _15144_ }), .Y(_15176_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31214_ ( .A({ _15209_, _08256_, _08257_, _15145_ }), .Y(_15177_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31215_ ( .A({ _15210_, _08256_, _08257_, _15146_ }), .Y(_15178_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31216_ ( .A({ _15211_, _08256_, _08257_, _15147_ }), .Y(_15179_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31217_ ( .A({ _15181_, _08256_, _08257_, _15117_ }), .Y(_15149_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31218_ ( .A({ _15182_, _08256_, _08257_, _15118_ }), .Y(_15150_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31219_ ( .A({ _15183_, _08256_, _08257_, _15119_ }), .Y(_15151_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31220_ ( .A({ _15184_, _08256_, _08257_, _15120_ }), .Y(_15152_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31221_ ( .A({ _15185_, _08256_, _08257_, _15121_ }), .Y(_15153_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31222_ ( .A({ _15186_, _08256_, _08257_, _15122_ }), .Y(_15154_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31223_ ( .A({ _15187_, _08256_, _08257_, _15123_ }), .Y(_15155_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31224_ ( .A({ _15188_, _08256_, _08257_, _15124_ }), .Y(_15156_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31225_ ( .A({ _15189_, _08256_, _08257_, _15125_ }), .Y(_15157_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31226_ ( .A({ _15190_, _08256_, _08257_, _15126_ }), .Y(_15158_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31227_ ( .A({ _15192_, _08256_, _08257_, _15128_ }), .Y(_15160_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31228_ ( .A({ _15193_, _08256_, _08257_, _15129_ }), .Y(_15161_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31229_ ( .A({ _15194_, _08256_, _08257_, _15130_ }), .Y(_15162_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31230_ ( .A({ _15195_, _08256_, _08257_, _15131_ }), .Y(_15163_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31231_ ( .A({ _15196_, _08256_, _08257_, _15132_ }), .Y(_15164_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31232_ ( .A({ _15197_, _08256_, _08257_, _15133_ }), .Y(_15165_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31233_ ( .A({ _15198_, _08256_, _08257_, _15134_ }), .Y(_15166_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31234_ ( .A({ _15199_, _08256_, _08257_, _15135_ }), .Y(_15167_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31235_ ( .A({ _15200_, _08256_, _08257_, _15136_ }), .Y(_15168_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31236_ ( .A({ _15201_, _08256_, _08257_, _15137_ }), .Y(_15169_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31237_ ( .A({ _15203_, _08256_, _08257_, _15139_ }), .Y(_15171_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31238_ ( .A({ _15204_, _08256_, _08257_, _15140_ }), .Y(_15172_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _31239_ ( .A({ _05059_, _08256_ }), .Y(_04832_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31240_ ( .A({ _08258_, _08196_, _maxi_write_fsm[0] }), .Y(_08260_) );
  \$lut  #( .LUT(16'hf8ff), .WIDTH(4) ) _31241_ ( .A({ _08261_, _08262_, _08256_, _15308_ }), .Y(_15212_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31242_ ( .A({ _05058_, _08257_, _15244_ }), .Y(_08261_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31243_ ( .A({ _15276_, _08260_ }), .Y(_08262_) );
  \$lut  #( .LUT(16'hf8ff), .WIDTH(4) ) _31244_ ( .A({ _08263_, _08264_, _08256_, _15319_ }), .Y(_15223_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31245_ ( .A({ _05059_, _08260_, _15287_ }), .Y(_08263_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31246_ ( .A({ _15255_, _08257_ }), .Y(_08264_) );
  \$lut  #( .LUT(16'hf8ff), .WIDTH(4) ) _31247_ ( .A({ _08265_, _08266_, _08256_, _15330_ }), .Y(_15234_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31248_ ( .A({ _05058_, _08257_, _15266_ }), .Y(_08265_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31249_ ( .A({ _15298_, _08260_ }), .Y(_08266_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31250_ ( .A({ _08267_, _15333_, _08256_ }), .Y(_15237_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31251_ ( .A({ _15269_, _08257_, _15301_, _08260_ }), .Y(_08267_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31252_ ( .A({ _08268_, _15334_, _08256_ }), .Y(_15238_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31253_ ( .A({ _15270_, _08257_, _15302_, _08260_ }), .Y(_08268_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31254_ ( .A({ _08269_, _15335_, _08256_ }), .Y(_15239_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31255_ ( .A({ _15271_, _08257_, _15303_, _08260_ }), .Y(_08269_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31256_ ( .A({ _08270_, _15336_, _08256_ }), .Y(_15240_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31257_ ( .A({ _15272_, _08257_, _15304_, _08260_ }), .Y(_08270_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31258_ ( .A({ _08271_, _15337_, _08256_ }), .Y(_15241_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31259_ ( .A({ _15273_, _08257_, _15305_, _08260_ }), .Y(_08271_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31260_ ( .A({ _08272_, _15338_, _08256_ }), .Y(_15242_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31261_ ( .A({ _15274_, _08257_, _15306_, _08260_ }), .Y(_08272_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31262_ ( .A({ _08273_, _15339_, _08256_ }), .Y(_15243_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31263_ ( .A({ _15275_, _08257_, _15307_, _08260_ }), .Y(_08273_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31264_ ( .A({ _08274_, _15309_, _08256_ }), .Y(_15213_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31265_ ( .A({ _15245_, _08257_, _15277_, _08260_ }), .Y(_08274_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31266_ ( .A({ _08275_, _15310_, _08256_ }), .Y(_15214_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31267_ ( .A({ _15246_, _08257_, _15278_, _08260_ }), .Y(_08275_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31268_ ( .A({ _08276_, _15311_, _08256_ }), .Y(_15215_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31269_ ( .A({ _15247_, _08257_, _15279_, _08260_ }), .Y(_08276_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31270_ ( .A({ _08277_, _15312_, _08256_ }), .Y(_15216_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31271_ ( .A({ _15248_, _08257_, _15280_, _08260_ }), .Y(_08277_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31272_ ( .A({ _08278_, _15313_, _08256_ }), .Y(_15217_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31273_ ( .A({ _15249_, _08257_, _15281_, _08260_ }), .Y(_08278_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31274_ ( .A({ _08279_, _15314_, _08256_ }), .Y(_15218_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31275_ ( .A({ _15250_, _08257_, _15282_, _08260_ }), .Y(_08279_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31276_ ( .A({ _08280_, _15315_, _08256_ }), .Y(_15219_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31277_ ( .A({ _15251_, _08257_, _15283_, _08260_ }), .Y(_08280_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31278_ ( .A({ _08281_, _15316_, _08256_ }), .Y(_15220_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31279_ ( .A({ _15252_, _08257_, _15284_, _08260_ }), .Y(_08281_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31280_ ( .A({ _08282_, _15317_, _08256_ }), .Y(_15221_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31281_ ( .A({ _15253_, _08257_, _15285_, _08260_ }), .Y(_08282_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31282_ ( .A({ _08283_, _15318_, _08256_ }), .Y(_15222_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31283_ ( .A({ _15254_, _08257_, _15286_, _08260_ }), .Y(_08283_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31284_ ( .A({ _08284_, _15320_, _08256_ }), .Y(_15224_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31285_ ( .A({ _15256_, _08257_, _15288_, _08260_ }), .Y(_08284_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31286_ ( .A({ _08285_, _15321_, _08256_ }), .Y(_15225_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31287_ ( .A({ _15257_, _08257_, _15289_, _08260_ }), .Y(_08285_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31288_ ( .A({ _08286_, _15322_, _08256_ }), .Y(_15226_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31289_ ( .A({ _15258_, _08257_, _15290_, _08260_ }), .Y(_08286_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31290_ ( .A({ _08287_, _15323_, _08256_ }), .Y(_15227_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31291_ ( .A({ _15259_, _08257_, _15291_, _08260_ }), .Y(_08287_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31292_ ( .A({ _08288_, _15324_, _08256_ }), .Y(_15228_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31293_ ( .A({ _15260_, _08257_, _15292_, _08260_ }), .Y(_08288_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31294_ ( .A({ _08289_, _15325_, _08256_ }), .Y(_15229_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31295_ ( .A({ _15261_, _08257_, _15293_, _08260_ }), .Y(_08289_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31296_ ( .A({ _08290_, _15326_, _08256_ }), .Y(_15230_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31297_ ( .A({ _15262_, _08257_, _15294_, _08260_ }), .Y(_08290_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31298_ ( .A({ _08291_, _15327_, _08256_ }), .Y(_15231_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31299_ ( .A({ _15263_, _08257_, _15295_, _08260_ }), .Y(_08291_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31300_ ( .A({ _08292_, _15328_, _08256_ }), .Y(_15232_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31301_ ( .A({ _15264_, _08257_, _15296_, _08260_ }), .Y(_08292_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31302_ ( .A({ _08293_, _15329_, _08256_ }), .Y(_15233_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31303_ ( .A({ _15265_, _08257_, _15297_, _08260_ }), .Y(_08293_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31304_ ( .A({ _08294_, _15331_, _08256_ }), .Y(_15235_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31305_ ( .A({ _15267_, _08257_, _15299_, _08260_ }), .Y(_08294_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31306_ ( .A({ _08295_, _15332_, _08256_ }), .Y(_15236_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31307_ ( .A({ _15268_, _08257_, _15300_, _08260_ }), .Y(_08295_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31308_ ( .A({ _15017_, _05059_, _15083_, _08256_ }), .Y(_15050_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31309_ ( .A({ _15028_, _05059_, _15094_, _08256_ }), .Y(_15061_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31310_ ( .A({ _15039_, _05059_, _15105_, _08256_ }), .Y(_15072_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31311_ ( .A({ _15043_, _05059_, _15109_, _08256_ }), .Y(_15076_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31312_ ( .A({ _15044_, _05059_, _15110_, _08256_ }), .Y(_15077_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31313_ ( .A({ _15045_, _05059_, _15111_, _08256_ }), .Y(_15078_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31314_ ( .A({ _15046_, _05059_, _15112_, _08256_ }), .Y(_15079_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31315_ ( .A({ _15047_, _05059_, _15113_, _08256_ }), .Y(_15080_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31316_ ( .A({ _15048_, _05059_, _15114_, _08256_ }), .Y(_15081_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31317_ ( .A({ _15049_, _05059_, _15115_, _08256_ }), .Y(_15082_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31318_ ( .A({ _15018_, _05059_, _15084_, _08256_ }), .Y(_15051_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31319_ ( .A({ _15019_, _05059_, _15085_, _08256_ }), .Y(_15052_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31320_ ( .A({ _15020_, _05059_, _15086_, _08256_ }), .Y(_15053_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31321_ ( .A({ _15021_, _05059_, _15087_, _08256_ }), .Y(_15054_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31322_ ( .A({ _15022_, _05059_, _15088_, _08256_ }), .Y(_15055_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31323_ ( .A({ _15023_, _05059_, _15089_, _08256_ }), .Y(_15056_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31324_ ( .A({ _15024_, _05059_, _15090_, _08256_ }), .Y(_15057_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31325_ ( .A({ _15025_, _05059_, _15091_, _08256_ }), .Y(_15058_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31326_ ( .A({ _15026_, _05059_, _15092_, _08256_ }), .Y(_15059_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31327_ ( .A({ _15027_, _05059_, _15093_, _08256_ }), .Y(_15060_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31328_ ( .A({ _15029_, _05059_, _15095_, _08256_ }), .Y(_15062_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31329_ ( .A({ _15030_, _05059_, _15096_, _08256_ }), .Y(_15063_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31330_ ( .A({ _15031_, _05059_, _15097_, _08256_ }), .Y(_15064_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31331_ ( .A({ _15032_, _05059_, _15098_, _08256_ }), .Y(_15065_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31332_ ( .A({ _15033_, _05059_, _15099_, _08256_ }), .Y(_15066_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31333_ ( .A({ _15034_, _05059_, _15100_, _08256_ }), .Y(_15067_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31334_ ( .A({ _15035_, _05059_, _15101_, _08256_ }), .Y(_15068_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31335_ ( .A({ _15036_, _05059_, _15102_, _08256_ }), .Y(_15069_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31336_ ( .A({ _15037_, _05059_, _15103_, _08256_ }), .Y(_15070_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31337_ ( .A({ _15038_, _05059_, _15104_, _08256_ }), .Y(_15071_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31338_ ( .A({ _15040_, _05059_, _15106_, _08256_ }), .Y(_15073_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31339_ ( .A({ _15041_, _05059_, _15107_, _08256_ }), .Y(_15074_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _31340_ ( .A({ _15042_, _05059_, _15108_, _08256_ }), .Y(_15075_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31341_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15876_, _15908_ }), .Y(_15844_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31342_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15875_, _15907_ }), .Y(_15843_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31343_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15871_, _15903_ }), .Y(_15839_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31344_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15873_, _15905_ }), .Y(_15841_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31345_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15872_, _15904_ }), .Y(_15840_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31346_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15870_, _15902_ }), .Y(_15838_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31347_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15869_, _15901_ }), .Y(_15837_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31348_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15866_, _15898_ }), .Y(_15834_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31349_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15868_, _15900_ }), .Y(_15836_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31350_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15867_, _15899_ }), .Y(_15835_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31351_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15865_, _15897_ }), .Y(_15833_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31352_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15864_, _15896_ }), .Y(_15832_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31353_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15860_, _15892_ }), .Y(_15828_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31354_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15862_, _15894_ }), .Y(_15830_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31355_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15861_, _15893_ }), .Y(_15829_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31356_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15859_, _15891_ }), .Y(_15827_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31357_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15858_, _15890_ }), .Y(_15826_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31358_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15855_, _15887_ }), .Y(_15823_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31359_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15857_, _15889_ }), .Y(_15825_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31360_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15856_, _15888_ }), .Y(_15824_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31361_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15854_, _15886_ }), .Y(_15822_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31362_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15853_, _15885_ }), .Y(_15821_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31363_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15881_, _15913_ }), .Y(_15849_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31364_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15883_, _15915_ }), .Y(_15851_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31365_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15882_, _15914_ }), .Y(_15850_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31366_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15880_, _15912_ }), .Y(_15848_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31367_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15879_, _15911_ }), .Y(_15847_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31368_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15874_, _15906_ }), .Y(_15842_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31369_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15878_, _15910_ }), .Y(_15846_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31370_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15877_, _15909_ }), .Y(_15845_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31371_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15863_, _15895_ }), .Y(_15831_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31372_ ( .A({ _08216_, _stream_conv2d_8_source_32_source_pat_fsm_15[0], _15852_, _15884_ }), .Y(_15820_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _31373_ ( .A({ _05068_, _08216_ }), .Y(_21905_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31374_ ( .A({ _18582_, _05909_, _06338_, _18614_ }), .Y(_04833_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31375_ ( .A({ _18581_, _05909_, _06338_, _18613_ }), .Y(_04834_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31376_ ( .A({ _18579_, _05909_, _06338_, _18611_ }), .Y(_04835_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31377_ ( .A({ _18578_, _05909_, _06338_, _18610_ }), .Y(_04836_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31378_ ( .A({ _18577_, _05909_, _06338_, _18609_ }), .Y(_04837_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31379_ ( .A({ _18576_, _05909_, _06338_, _18608_ }), .Y(_04838_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31380_ ( .A({ _18575_, _05909_, _06338_, _18607_ }), .Y(_04839_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31381_ ( .A({ _18574_, _05909_, _06338_, _18606_ }), .Y(_04840_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31382_ ( .A({ _18573_, _05909_, _06338_, _18605_ }), .Y(_04841_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31383_ ( .A({ _18572_, _05909_, _06338_, _18604_ }), .Y(_04842_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31384_ ( .A({ _18571_, _05909_, _06338_, _18603_ }), .Y(_04843_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31385_ ( .A({ _18570_, _05909_, _06338_, _18602_ }), .Y(_04844_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31386_ ( .A({ _18568_, _05909_, _06338_, _18600_ }), .Y(_04845_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31387_ ( .A({ _18567_, _05909_, _06338_, _18599_ }), .Y(_04846_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31388_ ( .A({ _18566_, _05909_, _06338_, _18598_ }), .Y(_04847_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31389_ ( .A({ _18565_, _05909_, _06338_, _18597_ }), .Y(_04848_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31390_ ( .A({ _18564_, _05909_, _06338_, _18596_ }), .Y(_04849_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31391_ ( .A({ _18563_, _05909_, _06338_, _18595_ }), .Y(_04850_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31392_ ( .A({ _18562_, _05909_, _06338_, _18594_ }), .Y(_04851_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31393_ ( .A({ _18561_, _05909_, _06338_, _18593_ }), .Y(_04852_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31394_ ( .A({ _18560_, _05909_, _06338_, _18592_ }), .Y(_04853_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31395_ ( .A({ _18559_, _05909_, _06338_, _18591_ }), .Y(_04854_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31396_ ( .A({ _18589_, _05909_, _06338_, _18621_ }), .Y(_04855_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31397_ ( .A({ _18588_, _05909_, _06338_, _18620_ }), .Y(_04856_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31398_ ( .A({ _18587_, _05909_, _06338_, _18619_ }), .Y(_04857_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31399_ ( .A({ _18586_, _05909_, _06338_, _18618_ }), .Y(_04858_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31400_ ( .A({ _18585_, _05909_, _06338_, _18617_ }), .Y(_04859_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31401_ ( .A({ _18584_, _05909_, _06338_, _18616_ }), .Y(_04860_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31402_ ( .A({ _18583_, _05909_, _06338_, _18615_ }), .Y(_04861_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31403_ ( .A({ _18580_, _05909_, _06338_, _18612_ }), .Y(_04862_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31404_ ( .A({ _18569_, _05909_, _06338_, _18601_ }), .Y(_04863_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31405_ ( .A({ _18558_, _05909_, _06338_, _18590_ }), .Y(_04864_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31406_ ( .A({ _05909_, _21926_ }), .Y(_21925_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _31407_ ( .A({ _05132_, _06338_ }), .Y(_21926_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31408_ ( .A({ _05132_, _19720_, _05909_ }), .Y(_19721_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31409_ ( .A({ _08297_, _08182_, _05886_ }), .Y(_08296_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31410_ ( .A(control_max_pool_serial_9[1:0]), .Y(_08297_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31411_ ( .A({ _05884_, _08299_, _05881_, _05876_ }), .Y(_08298_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31412_ ( .A({ control_max_pool_serial_9[1], _05887_, control_max_pool_serial_9[0] }), .Y(_08299_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31413_ ( .A({ _05885_, _05875_ }), .Y(_08300_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31414_ ( .A({ control_max_pool_serial_9[1:0], _05886_ }), .Y(_08301_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31415_ ( .A({ control_max_pool_serial_9[1], _05886_, _08303_, control_max_pool_serial_9[0] }), .Y(_08302_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31416_ ( .A(control_max_pool_serial_9[3:2]), .Y(_08303_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31417_ ( .A({ control_max_pool_serial_9[1], _05886_, _08182_, control_max_pool_serial_9[0] }), .Y(_08304_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31418_ ( .A({ control_max_pool_serial_9[1], _05886_, _05885_, control_max_pool_serial_9[0] }), .Y(_08305_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31419_ ( .A({ _08183_, _05887_, _05875_ }), .Y(_08306_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31420_ ( .A({ _08297_, _05885_, _05886_ }), .Y(_08307_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31421_ ( .A({ _08297_, _05887_, _05886_ }), .Y(_08308_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31422_ ( .A({ _08310_, _05056_, _05054_ }), .Y(_08309_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _31423_ ( .A({ _05886_, _08303_, control_max_pool_serial_9[1] }), .Y(_08310_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31424_ ( .A({ _08183_, _08182_, _05886_ }), .Y(_08311_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31425_ ( .A({ _08297_, _05875_, control_max_pool_serial_9[3:2] }), .Y(_08312_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31426_ ( .A({ control_max_pool_serial_9[3], _05875_, _08297_, control_max_pool_serial_9[2] }), .Y(_08313_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31427_ ( .A({ _08315_, _08306_, _14729_ }), .Y(_08314_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31428_ ( .A({ _14569_, _05052_, _14985_, _08308_ }), .Y(_08315_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31429_ ( .A({ _08318_, _08317_ }), .Y(_08316_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31430_ ( .A({ _14889_, _08296_, _08302_, _14793_ }), .Y(_08317_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31431_ ( .A({ _14921_, _08307_, _08311_, _14857_ }), .Y(_08318_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _31432_ ( .A({ _08320_, _21895_, _08321_, _14953_ }), .Y(_08319_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31433_ ( .A({ _14665_, _06012_, _14825_, _08304_ }), .Y(_08320_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31434_ ( .A({ control_max_pool_serial_9[1:0], _05887_, _05886_ }), .Y(_08321_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31435_ ( .A({ _14658_, _08313_ }), .Y(_08322_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31436_ ( .A({ _14786_, _08312_ }), .Y(_08323_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31437_ ( .A({ _05054_, _08298_, _14722_ }), .Y(_08324_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31438_ ( .A({ _08326_, _08304_, _14850_ }), .Y(_08325_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31439_ ( .A({ _14882_, _08311_, _14978_, _08321_ }), .Y(_08326_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31440_ ( .A({ _14914_, _08296_, _08302_, _14818_ }), .Y(_08327_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _31441_ ( .A({ _08329_, _08310_, _06012_, _14690_ }), .Y(_08328_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31442_ ( .A({ _15010_, _08308_, _08306_, _14754_ }), .Y(_08329_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31443_ ( .A({ _14772_, _08312_, _08313_, _14644_ }), .Y(_08330_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31444_ ( .A({ _08332_, _08311_, _14868_ }), .Y(_08331_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31445_ ( .A({ _14900_, _08296_, _14932_, _08307_ }), .Y(_08332_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31446_ ( .A({ _08337_, _08336_, _08335_, _08334_ }), .Y(_08333_) );
  \$lut  #( .LUT(16'h4fff), .WIDTH(4) ) _31447_ ( .A({ control_max_pool_serial_9[0], _08300_, control_max_pool_serial_9[1], _14676_ }), .Y(_08334_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31448_ ( .A({ _14836_, _08304_, _08306_, _14740_ }), .Y(_08335_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31449_ ( .A({ _14996_, _08308_, _08302_, _14804_ }), .Y(_08336_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31450_ ( .A({ _14580_, _05052_, _14964_, _08321_ }), .Y(_08337_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _31451_ ( .A({ _08343_, _08341_, _08338_ }), .Y(_14623_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31452_ ( .A({ _08340_, _08339_, _08309_ }), .Y(_08338_) );
  \$lut  #( .LUT(16'h8f00), .WIDTH(4) ) _31453_ ( .A({ _05053_, _08300_, control_max_pool_serial_9[1:0] }), .Y(_08339_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31454_ ( .A({ _14783_, _08312_, _08313_, _14655_ }), .Y(_08340_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31455_ ( .A({ _08342_, _08306_, _14751_ }), .Y(_08341_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31456_ ( .A({ _14815_, _08302_, _14879_, _08311_ }), .Y(_08342_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31457_ ( .A({ _08348_, _08346_, _08345_, _08344_ }), .Y(_08343_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31458_ ( .A({ _14591_, _05052_, _14975_, _08321_ }), .Y(_08344_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31459_ ( .A({ _14687_, _06012_, _14943_, _08307_ }), .Y(_08345_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _31460_ ( .A({ _08305_, _08347_, _08296_, _14911_ }), .Y(_08346_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31461_ ( .A({ _14719_, _08298_ }), .Y(_08347_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31462_ ( .A({ _15007_, _08308_, _08304_, _14847_ }), .Y(_08348_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31463_ ( .A({ _08356_, _08353_, _08351_, _08349_ }), .Y(_14627_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _31464_ ( .A({ _08339_, _08350_, _08312_, _14787_ }), .Y(_08349_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31465_ ( .A({ _14659_, _08313_ }), .Y(_08350_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31466_ ( .A({ _08352_, _08307_, _14947_ }), .Y(_08351_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31467_ ( .A({ _14595_, _05052_, _14819_, _08302_ }), .Y(_08352_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31468_ ( .A({ _08355_, _08354_ }), .Y(_08353_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31469_ ( .A({ _14915_, _08296_, _08306_, _14755_ }), .Y(_08354_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31470_ ( .A({ _15011_, _08308_, _08321_, _14979_ }), .Y(_08355_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _31471_ ( .A({ _08358_, _08357_, _06012_, _14691_ }), .Y(_08356_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31472_ ( .A({ _08303_, _08301_, _14723_, _08298_ }), .Y(_08357_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31473_ ( .A({ _14851_, _08304_, _14883_, _08311_ }), .Y(_08358_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31474_ ( .A({ _08366_, _08365_, _08363_, _08359_ }), .Y(_14628_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31475_ ( .A({ _08362_, _08361_, _08360_ }), .Y(_08359_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31476_ ( .A({ _14756_, _08306_, _08298_, _14724_ }), .Y(_08360_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31477_ ( .A({ _14692_, _06012_, _14948_, _08307_ }), .Y(_08361_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31478_ ( .A({ _14788_, _08312_, _08313_, _14660_ }), .Y(_08362_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31479_ ( .A({ _08364_, _08321_, _14980_ }), .Y(_08363_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31480_ ( .A({ _14916_, _08296_, _08304_, _14852_ }), .Y(_08364_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31481_ ( .A({ _14596_, _05052_, _14884_, _08311_ }), .Y(_08365_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31482_ ( .A({ _15012_, _08308_, _08302_, _14820_ }), .Y(_08366_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31483_ ( .A({ _08374_, _08373_, _08371_, _08367_ }), .Y(_14631_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31484_ ( .A({ _08370_, _08369_, _08368_ }), .Y(_08367_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31485_ ( .A({ _14759_, _08306_, _08298_, _14727_ }), .Y(_08368_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31486_ ( .A({ _14695_, _06012_, _14983_, _08321_ }), .Y(_08369_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31487_ ( .A({ _14791_, _08312_, _08313_, _14663_ }), .Y(_08370_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31488_ ( .A({ _08372_, _08307_, _14951_ }), .Y(_08371_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31489_ ( .A({ _14919_, _08296_, _08304_, _14855_ }), .Y(_08372_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31490_ ( .A({ _14599_, _05052_, _14887_, _08311_ }), .Y(_08373_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31491_ ( .A({ _15015_, _08308_, _08302_, _14823_ }), .Y(_08374_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31492_ ( .A({ _08382_, _08381_, _08379_, _08375_ }), .Y(_14629_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31493_ ( .A({ _08378_, _08377_, _08376_ }), .Y(_08375_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31494_ ( .A({ _14757_, _08306_, _08298_, _14725_ }), .Y(_08376_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31495_ ( .A({ _14693_, _06012_, _14981_, _08321_ }), .Y(_08377_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31496_ ( .A({ _14789_, _08312_, _08313_, _14661_ }), .Y(_08378_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31497_ ( .A({ _08380_, _08307_, _14949_ }), .Y(_08379_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31498_ ( .A({ _14917_, _08296_, _08304_, _14853_ }), .Y(_08380_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31499_ ( .A({ _14597_, _05052_, _14885_, _08311_ }), .Y(_08381_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31500_ ( .A({ _15013_, _08308_, _08302_, _14821_ }), .Y(_08382_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31501_ ( .A({ _08390_, _08389_, _08387_, _08383_ }), .Y(_14602_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31502_ ( .A({ _08386_, _08385_, _08384_ }), .Y(_08383_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31503_ ( .A({ _14730_, _08306_, _08298_, _14698_ }), .Y(_08384_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31504_ ( .A({ _14666_, _06012_, _14954_, _08321_ }), .Y(_08385_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31505_ ( .A({ _14762_, _08312_, _08313_, _14634_ }), .Y(_08386_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31506_ ( .A({ _08388_, _08307_, _14922_ }), .Y(_08387_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31507_ ( .A({ _14890_, _08296_, _08304_, _14826_ }), .Y(_08388_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31508_ ( .A({ _14570_, _05052_, _14858_, _08311_ }), .Y(_08389_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31509_ ( .A({ _14986_, _08308_, _08302_, _14794_ }), .Y(_08390_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31510_ ( .A({ _08398_, _08397_, _08395_, _08391_ }), .Y(_14630_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31511_ ( .A({ _08394_, _08393_, _08392_ }), .Y(_08391_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31512_ ( .A({ _14758_, _08306_, _08298_, _14726_ }), .Y(_08392_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31513_ ( .A({ _14694_, _06012_, _14982_, _08321_ }), .Y(_08393_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31514_ ( .A({ _14790_, _08312_, _08313_, _14662_ }), .Y(_08394_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31515_ ( .A({ _08396_, _08307_, _14950_ }), .Y(_08395_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31516_ ( .A({ _14918_, _08296_, _08304_, _14854_ }), .Y(_08396_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31517_ ( .A({ _14598_, _05052_, _14886_, _08311_ }), .Y(_08397_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31518_ ( .A({ _15014_, _08308_, _08302_, _14822_ }), .Y(_08398_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31519_ ( .A({ _08406_, _08405_, _08403_, _08399_ }), .Y(_14632_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31520_ ( .A({ _08402_, _08401_, _08400_ }), .Y(_08399_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31521_ ( .A({ _14760_, _08306_, _08298_, _14728_ }), .Y(_08400_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31522_ ( .A({ _14696_, _06012_, _14984_, _08321_ }), .Y(_08401_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31523_ ( .A({ _14792_, _08312_, _08313_, _14664_ }), .Y(_08402_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31524_ ( .A({ _08404_, _08307_, _14952_ }), .Y(_08403_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31525_ ( .A({ _14920_, _08296_, _08304_, _14856_ }), .Y(_08404_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31526_ ( .A({ _14600_, _05052_, _14888_, _08311_ }), .Y(_08405_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31527_ ( .A({ _15016_, _08308_, _08302_, _14824_ }), .Y(_08406_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31528_ ( .A({ _08414_, _08413_, _08411_, _08407_ }), .Y(_14603_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31529_ ( .A({ _08410_, _08409_, _08408_ }), .Y(_08407_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31530_ ( .A({ _14955_, _08321_, _08298_, _14699_ }), .Y(_08408_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31531_ ( .A({ _14667_, _06012_, _14891_, _08296_ }), .Y(_08409_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31532_ ( .A({ _14763_, _08312_, _08313_, _14635_ }), .Y(_08410_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31533_ ( .A({ _08412_, _08308_, _14987_ }), .Y(_08411_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31534_ ( .A({ _14923_, _08307_, _08302_, _14795_ }), .Y(_08412_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31535_ ( .A({ _14827_, _08304_, _08306_, _14731_ }), .Y(_08413_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31536_ ( .A({ _14571_, _05052_, _14859_, _08311_ }), .Y(_08414_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31537_ ( .A({ _08422_, _08421_, _08419_, _08415_ }), .Y(_14605_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31538_ ( .A({ _08418_, _08417_, _08416_ }), .Y(_08415_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31539_ ( .A({ _14733_, _08306_, _08298_, _14701_ }), .Y(_08416_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31540_ ( .A({ _14669_, _06012_, _14925_, _08307_ }), .Y(_08417_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31541_ ( .A({ _14765_, _08312_, _08313_, _14637_ }), .Y(_08418_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31542_ ( .A({ _08420_, _08321_, _14957_ }), .Y(_08419_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31543_ ( .A({ _14893_, _08296_, _08304_, _14829_ }), .Y(_08420_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31544_ ( .A({ _14573_, _05052_, _14861_, _08311_ }), .Y(_08421_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31545_ ( .A({ _14989_, _08308_, _08302_, _14797_ }), .Y(_08422_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31546_ ( .A({ _08430_, _08429_, _08427_, _08423_ }), .Y(_14607_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31547_ ( .A({ _08426_, _08425_, _08424_ }), .Y(_08423_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31548_ ( .A({ _14735_, _08306_, _08298_, _14703_ }), .Y(_08424_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31549_ ( .A({ _14671_, _06012_, _14959_, _08321_ }), .Y(_08425_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31550_ ( .A({ _14767_, _08312_, _08313_, _14639_ }), .Y(_08426_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31551_ ( .A({ _08428_, _08307_, _14927_ }), .Y(_08427_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31552_ ( .A({ _14895_, _08296_, _08304_, _14831_ }), .Y(_08428_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31553_ ( .A({ _14575_, _05052_, _14863_, _08311_ }), .Y(_08429_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31554_ ( .A({ _14991_, _08308_, _08302_, _14799_ }), .Y(_08430_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31555_ ( .A({ _08438_, _08437_, _08435_, _08431_ }), .Y(_14604_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31556_ ( .A({ _08434_, _08433_, _08432_ }), .Y(_08431_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31557_ ( .A({ _14732_, _08306_, _08298_, _14700_ }), .Y(_08432_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31558_ ( .A({ _14668_, _06012_, _14956_, _08321_ }), .Y(_08433_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31559_ ( .A({ _14764_, _08312_, _08313_, _14636_ }), .Y(_08434_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31560_ ( .A({ _08436_, _08307_, _14924_ }), .Y(_08435_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31561_ ( .A({ _14892_, _08296_, _08304_, _14828_ }), .Y(_08436_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31562_ ( .A({ _14572_, _05052_, _14860_, _08311_ }), .Y(_08437_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31563_ ( .A({ _14988_, _08308_, _08302_, _14796_ }), .Y(_08438_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31564_ ( .A({ _08446_, _08445_, _08443_, _08439_ }), .Y(_14606_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31565_ ( .A({ _08442_, _08441_, _08440_ }), .Y(_08439_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31566_ ( .A({ _14830_, _08304_, _08298_, _14702_ }), .Y(_08440_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31567_ ( .A({ _14990_, _08308_, _08321_, _14958_ }), .Y(_08441_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31568_ ( .A({ _14766_, _08312_, _08313_, _14638_ }), .Y(_08442_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31569_ ( .A({ _08444_, _06012_, _14670_ }), .Y(_08443_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31570_ ( .A({ _14894_, _08296_, _08306_, _14734_ }), .Y(_08444_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31571_ ( .A({ _14926_, _08307_, _08311_, _14862_ }), .Y(_08445_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31572_ ( .A({ _14574_, _05052_, _14798_, _08302_ }), .Y(_08446_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31573_ ( .A({ _08454_, _08453_, _08451_, _08447_ }), .Y(_14608_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31574_ ( .A({ _08450_, _08449_, _08448_ }), .Y(_08447_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31575_ ( .A({ _14736_, _08306_, _08298_, _14704_ }), .Y(_08448_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31576_ ( .A({ _14672_, _06012_, _14928_, _08307_ }), .Y(_08449_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31577_ ( .A({ _14768_, _08312_, _08313_, _14640_ }), .Y(_08450_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31578_ ( .A({ _08452_, _08321_, _14960_ }), .Y(_08451_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31579_ ( .A({ _14896_, _08296_, _08304_, _14832_ }), .Y(_08452_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31580_ ( .A({ _14576_, _05052_, _14864_, _08311_ }), .Y(_08453_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31581_ ( .A({ _14992_, _08308_, _08302_, _14800_ }), .Y(_08454_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31582_ ( .A({ _08462_, _08461_, _08459_, _08455_ }), .Y(_14613_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31583_ ( .A({ _08458_, _08457_, _08456_ }), .Y(_08455_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31584_ ( .A({ _14741_, _08306_, _08298_, _14709_ }), .Y(_08456_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31585_ ( .A({ _14677_, _06012_, _14965_, _08321_ }), .Y(_08457_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31586_ ( .A({ _14773_, _08312_, _08313_, _14645_ }), .Y(_08458_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31587_ ( .A({ _08460_, _08307_, _14933_ }), .Y(_08459_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31588_ ( .A({ _14901_, _08296_, _08304_, _14837_ }), .Y(_08460_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31589_ ( .A({ _14581_, _05052_, _14869_, _08311_ }), .Y(_08461_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31590_ ( .A({ _14997_, _08308_, _08302_, _14805_ }), .Y(_08462_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31591_ ( .A({ _08470_, _08469_, _08467_, _08463_ }), .Y(_14609_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31592_ ( .A({ _08466_, _08465_, _08464_ }), .Y(_08463_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31593_ ( .A({ _14737_, _08306_, _08298_, _14705_ }), .Y(_08464_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31594_ ( .A({ _14673_, _06012_, _14929_, _08307_ }), .Y(_08465_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31595_ ( .A({ _14769_, _08312_, _08313_, _14641_ }), .Y(_08466_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31596_ ( .A({ _08468_, _08321_, _14961_ }), .Y(_08467_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31597_ ( .A({ _14897_, _08296_, _08304_, _14833_ }), .Y(_08468_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31598_ ( .A({ _14577_, _05052_, _14865_, _08311_ }), .Y(_08469_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31599_ ( .A({ _14993_, _08308_, _08302_, _14801_ }), .Y(_08470_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31600_ ( .A({ _08478_, _08477_, _08475_, _08471_ }), .Y(_14610_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31601_ ( .A({ _08474_, _08473_, _08472_ }), .Y(_08471_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31602_ ( .A({ _14738_, _08306_, _08298_, _14706_ }), .Y(_08472_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31603_ ( .A({ _14674_, _06012_, _14962_, _08321_ }), .Y(_08473_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31604_ ( .A({ _14770_, _08312_, _08313_, _14642_ }), .Y(_08474_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31605_ ( .A({ _08476_, _08307_, _14930_ }), .Y(_08475_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31606_ ( .A({ _14898_, _08296_, _08304_, _14834_ }), .Y(_08476_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31607_ ( .A({ _14578_, _05052_, _14866_, _08311_ }), .Y(_08477_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31608_ ( .A({ _14994_, _08308_, _08302_, _14802_ }), .Y(_08478_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31609_ ( .A({ _08486_, _08485_, _08483_, _08479_ }), .Y(_14611_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31610_ ( .A({ _08482_, _08481_, _08480_ }), .Y(_08479_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31611_ ( .A({ _14835_, _08304_, _08298_, _14707_ }), .Y(_08480_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31612_ ( .A({ _14675_, _06012_, _14995_, _08308_ }), .Y(_08481_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31613_ ( .A({ _14771_, _08312_, _08313_, _14643_ }), .Y(_08482_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _31614_ ( .A({ _08484_, _05052_, _14579_ }), .Y(_08483_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31615_ ( .A({ _14899_, _08296_, _08311_, _14867_ }), .Y(_08484_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31616_ ( .A({ _14931_, _08307_, _08302_, _14803_ }), .Y(_08485_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31617_ ( .A({ _14739_, _08306_, _14963_, _08321_ }), .Y(_08486_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31618_ ( .A({ _08494_, _08493_, _08491_, _08487_ }), .Y(_14614_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31619_ ( .A({ _08490_, _08489_, _08488_ }), .Y(_08487_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31620_ ( .A({ _14838_, _08304_, _08298_, _14710_ }), .Y(_08488_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31621_ ( .A({ _14678_, _06012_, _14998_, _08308_ }), .Y(_08489_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31622_ ( .A({ _14774_, _08312_, _08313_, _14646_ }), .Y(_08490_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _31623_ ( .A({ _08492_, _05052_, _14582_ }), .Y(_08491_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31624_ ( .A({ _14902_, _08296_, _08311_, _14870_ }), .Y(_08492_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31625_ ( .A({ _14806_, _08302_, _14966_, _08321_ }), .Y(_08493_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31626_ ( .A({ _14934_, _08307_, _08306_, _14742_ }), .Y(_08494_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31627_ ( .A({ _08502_, _08501_, _08499_, _08495_ }), .Y(_14615_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31628_ ( .A({ _08498_, _08497_, _08496_ }), .Y(_08495_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31629_ ( .A({ _14743_, _08306_, _08298_, _14711_ }), .Y(_08496_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31630_ ( .A({ _14679_, _06012_, _14967_, _08321_ }), .Y(_08497_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31631_ ( .A({ _14775_, _08312_, _08313_, _14647_ }), .Y(_08498_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31632_ ( .A({ _08500_, _08307_, _14935_ }), .Y(_08499_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31633_ ( .A({ _14903_, _08296_, _08304_, _14839_ }), .Y(_08500_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31634_ ( .A({ _14583_, _05052_, _14871_, _08311_ }), .Y(_08501_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31635_ ( .A({ _14999_, _08308_, _08302_, _14807_ }), .Y(_08502_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31636_ ( .A({ _08510_, _08509_, _08507_, _08503_ }), .Y(_14616_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31637_ ( .A({ _08506_, _08505_, _08504_ }), .Y(_08503_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31638_ ( .A({ _14840_, _08304_, _08298_, _14712_ }), .Y(_08504_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31639_ ( .A({ _15000_, _08308_, _08321_, _14968_ }), .Y(_08505_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31640_ ( .A({ _14776_, _08312_, _08313_, _14648_ }), .Y(_08506_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _31641_ ( .A({ _08508_, _05052_, _14584_ }), .Y(_08507_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31642_ ( .A({ _14904_, _08296_, _08311_, _14872_ }), .Y(_08508_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31643_ ( .A({ _14680_, _06012_, _14808_, _08302_ }), .Y(_08509_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31644_ ( .A({ _14936_, _08307_, _08306_, _14744_ }), .Y(_08510_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31645_ ( .A({ _08518_, _08517_, _08515_, _08511_ }), .Y(_14617_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31646_ ( .A({ _08514_, _08513_, _08512_ }), .Y(_08511_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31647_ ( .A({ _14745_, _08306_, _08298_, _14713_ }), .Y(_08512_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31648_ ( .A({ _14681_, _06012_, _14937_, _08307_ }), .Y(_08513_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31649_ ( .A({ _14777_, _08312_, _08313_, _14649_ }), .Y(_08514_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31650_ ( .A({ _08516_, _08321_, _14969_ }), .Y(_08515_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31651_ ( .A({ _14905_, _08296_, _08304_, _14841_ }), .Y(_08516_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31652_ ( .A({ _14585_, _05052_, _14873_, _08311_ }), .Y(_08517_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31653_ ( .A({ _15001_, _08308_, _08302_, _14809_ }), .Y(_08518_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31654_ ( .A({ _08526_, _08525_, _08523_, _08519_ }), .Y(_14618_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31655_ ( .A({ _08522_, _08521_, _08520_ }), .Y(_08519_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31656_ ( .A({ _14746_, _08306_, _08298_, _14714_ }), .Y(_08520_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31657_ ( .A({ _14682_, _06012_, _14970_, _08321_ }), .Y(_08521_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31658_ ( .A({ _14778_, _08312_, _08313_, _14650_ }), .Y(_08522_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31659_ ( .A({ _08524_, _08307_, _14938_ }), .Y(_08523_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31660_ ( .A({ _14906_, _08296_, _08304_, _14842_ }), .Y(_08524_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31661_ ( .A({ _14586_, _05052_, _14874_, _08311_ }), .Y(_08525_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31662_ ( .A({ _15002_, _08308_, _08302_, _14810_ }), .Y(_08526_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31663_ ( .A({ _08534_, _08533_, _08531_, _08527_ }), .Y(_14619_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31664_ ( .A({ _08530_, _08529_, _08528_ }), .Y(_08527_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31665_ ( .A({ _14843_, _08304_, _08298_, _14715_ }), .Y(_08528_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31666_ ( .A({ _14683_, _06012_, _15003_, _08308_ }), .Y(_08529_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31667_ ( .A({ _14779_, _08312_, _08313_, _14651_ }), .Y(_08530_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _31668_ ( .A({ _08532_, _05052_, _14587_ }), .Y(_08531_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31669_ ( .A({ _14907_, _08296_, _08311_, _14875_ }), .Y(_08532_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31670_ ( .A({ _14939_, _08307_, _08302_, _14811_ }), .Y(_08533_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31671_ ( .A({ _14747_, _08306_, _14971_, _08321_ }), .Y(_08534_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31672_ ( .A({ _08542_, _08541_, _08539_, _08535_ }), .Y(_14620_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31673_ ( .A({ _08538_, _08537_, _08536_ }), .Y(_08535_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31674_ ( .A({ _14844_, _08304_, _08298_, _14716_ }), .Y(_08536_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31675_ ( .A({ _14940_, _08307_, _15004_, _08308_ }), .Y(_08537_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31676_ ( .A({ _14780_, _08312_, _08313_, _14652_ }), .Y(_08538_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31677_ ( .A({ _08540_, _06012_, _14684_ }), .Y(_08539_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31678_ ( .A({ _14908_, _08296_, _08306_, _14748_ }), .Y(_08540_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31679_ ( .A({ _14876_, _08311_, _14972_, _08321_ }), .Y(_08541_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31680_ ( .A({ _14588_, _05052_, _14812_, _08302_ }), .Y(_08542_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31681_ ( .A({ _08550_, _08549_, _08547_, _08543_ }), .Y(_14621_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31682_ ( .A({ _08546_, _08545_, _08544_ }), .Y(_08543_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31683_ ( .A({ _14749_, _08306_, _08298_, _14717_ }), .Y(_08544_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31684_ ( .A({ _14685_, _06012_, _14973_, _08321_ }), .Y(_08545_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31685_ ( .A({ _14781_, _08312_, _08313_, _14653_ }), .Y(_08546_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31686_ ( .A({ _08548_, _08307_, _14941_ }), .Y(_08547_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31687_ ( .A({ _14909_, _08296_, _08304_, _14845_ }), .Y(_08548_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31688_ ( .A({ _14589_, _05052_, _14877_, _08311_ }), .Y(_08549_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31689_ ( .A({ _15005_, _08308_, _08302_, _14813_ }), .Y(_08550_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31690_ ( .A({ _08558_, _08557_, _08555_, _08551_ }), .Y(_14622_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31691_ ( .A({ _08554_, _08553_, _08552_ }), .Y(_08551_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31692_ ( .A({ _14750_, _08306_, _08298_, _14718_ }), .Y(_08552_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31693_ ( .A({ _14686_, _06012_, _14942_, _08307_ }), .Y(_08553_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31694_ ( .A({ _14782_, _08312_, _08313_, _14654_ }), .Y(_08554_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31695_ ( .A({ _08556_, _08321_, _14974_ }), .Y(_08555_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31696_ ( .A({ _14910_, _08296_, _08304_, _14846_ }), .Y(_08556_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31697_ ( .A({ _14590_, _05052_, _14878_, _08311_ }), .Y(_08557_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31698_ ( .A({ _15006_, _08308_, _08302_, _14814_ }), .Y(_08558_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31699_ ( .A({ _08566_, _08565_, _08563_, _08559_ }), .Y(_14624_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31700_ ( .A({ _08562_, _08561_, _08560_ }), .Y(_08559_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31701_ ( .A({ _15008_, _08308_, _08298_, _14720_ }), .Y(_08560_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31702_ ( .A({ _14912_, _08296_, _08306_, _14752_ }), .Y(_08561_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31703_ ( .A({ _14784_, _08312_, _08313_, _14656_ }), .Y(_08562_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31704_ ( .A({ _08564_, _06012_, _14688_ }), .Y(_08563_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31705_ ( .A({ _14944_, _08307_, _08302_, _14816_ }), .Y(_08564_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31706_ ( .A({ _14592_, _05052_, _14880_, _08311_ }), .Y(_08565_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31707_ ( .A({ _14848_, _08304_, _14976_, _08321_ }), .Y(_08566_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31708_ ( .A({ _08574_, _08573_, _08571_, _08567_ }), .Y(_14625_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31709_ ( .A({ _08570_, _08569_, _08568_ }), .Y(_08567_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31710_ ( .A({ _14753_, _08306_, _08298_, _14721_ }), .Y(_08568_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31711_ ( .A({ _14689_, _06012_, _14977_, _08321_ }), .Y(_08569_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31712_ ( .A({ _14785_, _08312_, _08313_, _14657_ }), .Y(_08570_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31713_ ( .A({ _08572_, _08307_, _14945_ }), .Y(_08571_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31714_ ( .A({ _14913_, _08296_, _08304_, _14849_ }), .Y(_08572_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31715_ ( .A({ _14593_, _05052_, _14881_, _08311_ }), .Y(_08573_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31716_ ( .A({ _15009_, _08308_, _08302_, _14817_ }), .Y(_08574_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31717_ ( .A({ conv2d_8_prev_row_select[0], conv2d_8_prev_row_select[1] }), .Y(_04865_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31718_ ( .A({ __tmp_339_2[0], __tmp_339_2[1] }), .Y(_04866_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31719_ ( .A({ __tmp_359_2[0], __tmp_359_2[1] }), .Y(_04867_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31720_ ( .A({ __tmp_369_2[0], __tmp_369_2[1] }), .Y(_04868_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31721_ ( .A({ __tmp_379_2[0], __tmp_379_2[1] }), .Y(_04869_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31722_ ( .A({ __tmp_389_2[0], __tmp_389_2[1] }), .Y(_04870_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31723_ ( .A({ __tmp_399_2[0], __tmp_399_2[1] }), .Y(_04871_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31724_ ( .A({ __tmp_409_2[0], __tmp_409_2[1] }), .Y(_04872_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31725_ ( .A({ __tmp_419_2[0], __tmp_419_2[1] }), .Y(_04873_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31726_ ( .A({ __tmp_429_2[0], __tmp_429_2[1] }), .Y(_04874_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31727_ ( .A({ __tmp_439_2[0], __tmp_439_2[1] }), .Y(_04875_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31728_ ( .A({ __tmp_449_2[0], __tmp_449_2[1] }), .Y(_04876_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31729_ ( .A({ __tmp_459_2[0], __tmp_459_2[1] }), .Y(_04877_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31730_ ( .A({ __tmp_469_2[0], __tmp_469_2[1] }), .Y(_04878_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31731_ ( .A({ __tmp_479_2[0], __tmp_479_2[1] }), .Y(_04879_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31732_ ( .A({ __tmp_489_2[0], __tmp_489_2[1] }), .Y(_04880_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31733_ ( .A({ __tmp_499_2[0], __tmp_499_2[1] }), .Y(_04881_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31734_ ( .A({ __tmp_509_2[0], __tmp_509_2[1] }), .Y(_04882_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31735_ ( .A({ __tmp_519_2[0], __tmp_519_2[1] }), .Y(_04883_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31736_ ( .A({ __tmp_529_2[0], __tmp_529_2[1] }), .Y(_04884_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31737_ ( .A({ conv2d_8_row_select[0], conv2d_8_row_select[1] }), .Y(_04885_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31738_ ( .A({ __tmp_865_2[0], __tmp_865_2[1] }), .Y(_04886_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31739_ ( .A({ __tmp_995_2[0], __tmp_995_2[1] }), .Y(_04887_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31740_ ( .A({ __tmp_1015_2[0], __tmp_1015_2[1] }), .Y(_04888_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31741_ ( .A({ __tmp_1025_2[0], __tmp_1025_2[1] }), .Y(_04889_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _31742_ ( .A({ _08058_, _tmp_5[1:0] }), .Y(_04890_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31743_ ( .A({ _08584_, _08583_, _08582_, _08575_ }), .Y(_04891_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31744_ ( .A({ _08581_, _08576_, _reduceadd_count_15[1:0] }), .Y(_08575_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31745_ ( .A({ _08580_, _08579_, _08578_, _08577_ }), .Y(_08576_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31746_ ( .A(_reduceadd_count_15[13:10]), .Y(_08577_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31747_ ( .A(_reduceadd_count_15[9:6]), .Y(_08578_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31748_ ( .A(_reduceadd_count_15[21:18]), .Y(_08579_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31749_ ( .A(_reduceadd_count_15[17:14]), .Y(_08580_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31750_ ( .A(_reduceadd_count_15[5:2]), .Y(_08581_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _31751_ ( .A(_reduceadd_count_15[32:30]), .Y(_08582_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31752_ ( .A(_reduceadd_count_15[29:26]), .Y(_08583_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31753_ ( .A(_reduceadd_count_15[25:22]), .Y(_08584_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _31754_ ( .A({ _08585_, _reducecustom_count_191[4:3] }), .Y(_04892_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31755_ ( .A({ _08586_, _reducecustom_count_191[8:6] }), .Y(_08585_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31756_ ( .A({ _reducecustom_count_191[5], _reducecustom_count_191[2:0] }), .Y(_08586_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _31757_ ( .A(_counter_count_762), .Y(_04893_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31758_ ( .A({ _08592_, _08587_ }), .Y(_04894_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31759_ ( .A({ _08591_, _08590_, _08589_, _08588_ }), .Y(_08587_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31760_ ( .A(conv2d_8_out_ram_select[23:20]), .Y(_08588_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31761_ ( .A(conv2d_8_out_ram_select[19:16]), .Y(_08589_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31762_ ( .A(conv2d_8_out_ram_select[31:28]), .Y(_08590_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31763_ ( .A(conv2d_8_out_ram_select[27:24]), .Y(_08591_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31764_ ( .A({ _08596_, _08595_, _08594_, _08593_ }), .Y(_08592_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31765_ ( .A(conv2d_8_out_ram_select[7:4]), .Y(_08593_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31766_ ( .A(conv2d_8_out_ram_select[3:0]), .Y(_08594_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31767_ ( .A(conv2d_8_out_ram_select[15:12]), .Y(_08595_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31768_ ( .A(conv2d_8_out_ram_select[11:8]), .Y(_08596_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31769_ ( .A({ conv2d_8_col_select[0], conv2d_8_col_select[1] }), .Y(_04895_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31770_ ( .A({ _08602_, _08597_ }), .Y(_04896_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31771_ ( .A({ _08601_, _08600_, _08599_, _08598_ }), .Y(_08597_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31772_ ( .A(matmul_15_out_ram_select[23:20]), .Y(_08598_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31773_ ( .A(matmul_15_out_ram_select[19:16]), .Y(_08599_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31774_ ( .A(matmul_15_out_ram_select[31:28]), .Y(_08600_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31775_ ( .A(matmul_15_out_ram_select[27:24]), .Y(_08601_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31776_ ( .A({ _08606_, _08605_, _08604_, _08603_ }), .Y(_08602_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31777_ ( .A(matmul_15_out_ram_select[7:4]), .Y(_08603_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31778_ ( .A(matmul_15_out_ram_select[3:0]), .Y(_08604_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31779_ ( .A(matmul_15_out_ram_select[15:12]), .Y(_08605_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31780_ ( .A(matmul_15_out_ram_select[11:8]), .Y(_08606_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _31781_ ( .A({ _08047_, _saxi_register_fsm[0] }), .Y(_04904_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31782_ ( .A({ _tmp_62[0], _tmp_62[1], _tmp_62[3:2] }), .Y(_05153_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31783_ ( .A({ _tmp_93[0], _tmp_93[1], _tmp_93[3:2] }), .Y(_05162_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31784_ ( .A({ _tmp_124[0], _tmp_124[1], _tmp_124[3:2] }), .Y(_05171_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31785_ ( .A({ _tmp_155[0], _tmp_155[1], _tmp_155[3:2] }), .Y(_05180_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31786_ ( .A({ _tmp_62[0], _tmp_62[1], _tmp_62[3:2] }), .Y(_05154_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31787_ ( .A({ _tmp_93[0], _tmp_93[1], _tmp_93[3:2] }), .Y(_05163_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31788_ ( .A({ _tmp_124[0], _tmp_124[1], _tmp_124[3:2] }), .Y(_05172_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31789_ ( .A({ _tmp_155[0], _tmp_155[1], _tmp_155[3:2] }), .Y(_05181_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31790_ ( .A({ _tmp_62[1:0], _tmp_62[3:2] }), .Y(_05155_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31791_ ( .A({ _tmp_93[1:0], _tmp_93[3:2] }), .Y(_05164_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31792_ ( .A({ _tmp_124[1:0], _tmp_124[3:2] }), .Y(_05173_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31793_ ( .A({ _tmp_155[1:0], _tmp_155[3:2] }), .Y(_05182_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31794_ ( .A({ _tmp_62[0], _tmp_62[1], _tmp_62[3:2] }), .Y(_05156_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31795_ ( .A({ _tmp_93[0], _tmp_93[1], _tmp_93[3:2] }), .Y(_05165_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31796_ ( .A({ _tmp_124[0], _tmp_124[1], _tmp_124[3:2] }), .Y(_05174_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31797_ ( .A({ _tmp_155[0], _tmp_155[1], _tmp_155[3:2] }), .Y(_05183_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31798_ ( .A({ _tmp_62[2], _tmp_62[0], _tmp_62[1], _tmp_62[3] }), .Y(_05157_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31799_ ( .A({ _tmp_93[2], _tmp_93[0], _tmp_93[1], _tmp_93[3] }), .Y(_05166_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31800_ ( .A({ _tmp_124[2], _tmp_124[0], _tmp_124[1], _tmp_124[3] }), .Y(_05175_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31801_ ( .A({ _tmp_155[2], _tmp_155[0], _tmp_155[1], _tmp_155[3] }), .Y(_05184_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31802_ ( .A({ _tmp_62[0], _tmp_62[2:1], _tmp_62[3] }), .Y(_05158_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31803_ ( .A({ _tmp_93[0], _tmp_93[2:1], _tmp_93[3] }), .Y(_05167_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31804_ ( .A({ _tmp_124[0], _tmp_124[2:1], _tmp_124[3] }), .Y(_05176_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31805_ ( .A({ _tmp_155[0], _tmp_155[2:1], _tmp_155[3] }), .Y(_05185_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31806_ ( .A({ _tmp_62[2:0], _tmp_62[3] }), .Y(_05159_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31807_ ( .A({ _tmp_93[2:0], _tmp_93[3] }), .Y(_05168_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31808_ ( .A({ _tmp_124[2:0], _tmp_124[3] }), .Y(_05177_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31809_ ( .A({ _tmp_155[2:0], _tmp_155[3] }), .Y(_05186_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31810_ ( .A({ _tmp_62[0], _tmp_62[1], _tmp_62[2], _tmp_62[3] }), .Y(_05160_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31811_ ( .A({ _tmp_93[0], _tmp_93[1], _tmp_93[2], _tmp_93[3] }), .Y(_05169_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31812_ ( .A({ _tmp_124[0], _tmp_124[1], _tmp_124[2], _tmp_124[3] }), .Y(_05178_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31813_ ( .A({ _tmp_155[0], _tmp_155[1], _tmp_155[2], _tmp_155[3] }), .Y(_05187_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31814_ ( .A({ _tmp_62[3], _tmp_62[0], _tmp_62[1], _tmp_62[2] }), .Y(_05152_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31815_ ( .A({ _tmp_93[3], _tmp_93[0], _tmp_93[1], _tmp_93[2] }), .Y(_05161_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31816_ ( .A({ _tmp_124[3], _tmp_124[0], _tmp_124[1], _tmp_124[2] }), .Y(_05170_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31817_ ( .A({ _tmp_155[3], _tmp_155[0], _tmp_155[1], _tmp_155[2] }), .Y(_05179_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31818_ ( .A({ _tmp_173[0], _tmp_173[1] }), .Y(_05189_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31819_ ( .A({ _tmp_186[0], _tmp_186[1] }), .Y(_05192_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31820_ ( .A({ _tmp_199[0], _tmp_199[1] }), .Y(_05195_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31821_ ( .A({ _tmp_212[0], _tmp_212[1] }), .Y(_05198_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31822_ ( .A({ _tmp_173[0], _tmp_173[1] }), .Y(_05190_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31823_ ( .A({ _tmp_186[0], _tmp_186[1] }), .Y(_05193_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31824_ ( .A({ _tmp_199[0], _tmp_199[1] }), .Y(_05196_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31825_ ( .A({ _tmp_212[0], _tmp_212[1] }), .Y(_05199_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31826_ ( .A(_tmp_173), .Y(_05188_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31827_ ( .A(_tmp_186), .Y(_05191_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31828_ ( .A(_tmp_199), .Y(_05194_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31829_ ( .A(_tmp_212), .Y(_05197_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31830_ ( .A({ _tmp_230[0], _tmp_230[1] }), .Y(_05201_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31831_ ( .A({ _tmp_243[0], _tmp_243[1] }), .Y(_05204_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31832_ ( .A({ _tmp_256[0], _tmp_256[1] }), .Y(_05207_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31833_ ( .A({ _tmp_269[0], _tmp_269[1] }), .Y(_05210_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31834_ ( .A({ _tmp_230[0], _tmp_230[1] }), .Y(_05202_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31835_ ( .A({ _tmp_243[0], _tmp_243[1] }), .Y(_05205_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31836_ ( .A({ _tmp_256[0], _tmp_256[1] }), .Y(_05208_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31837_ ( .A({ _tmp_269[0], _tmp_269[1] }), .Y(_05211_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31838_ ( .A(_tmp_230), .Y(_05200_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31839_ ( .A(_tmp_243), .Y(_05203_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31840_ ( .A(_tmp_256), .Y(_05206_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31841_ ( .A(_tmp_269), .Y(_05209_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31842_ ( .A({ _tmp_287[0], _tmp_287[1] }), .Y(_05213_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31843_ ( .A({ _tmp_300[0], _tmp_300[1] }), .Y(_05216_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31844_ ( .A({ _tmp_313[0], _tmp_313[1] }), .Y(_05219_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31845_ ( .A({ _tmp_326[0], _tmp_326[1] }), .Y(_05222_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31846_ ( .A({ _tmp_287[0], _tmp_287[1] }), .Y(_05214_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31847_ ( .A({ _tmp_300[0], _tmp_300[1] }), .Y(_05217_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31848_ ( .A({ _tmp_313[0], _tmp_313[1] }), .Y(_05220_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31849_ ( .A({ _tmp_326[0], _tmp_326[1] }), .Y(_05223_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31850_ ( .A(_tmp_287), .Y(_05212_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31851_ ( .A(_tmp_300), .Y(_05215_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31852_ ( .A(_tmp_313), .Y(_05218_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31853_ ( .A(_tmp_326), .Y(_05221_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31854_ ( .A({ _08616_, _08614_, _08607_ }), .Y(_05151_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31855_ ( .A({ _08613_, _08608_, _maxi_write_size[2:1] }), .Y(_08607_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31856_ ( .A({ _08612_, _08611_, _08610_, _08609_ }), .Y(_08608_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31857_ ( .A(_maxi_write_size[14:11]), .Y(_08609_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31858_ ( .A(_maxi_write_size[10:7]), .Y(_08610_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31859_ ( .A(_maxi_write_size[22:19]), .Y(_08611_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31860_ ( .A(_maxi_write_size[18:15]), .Y(_08612_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31861_ ( .A(_maxi_write_size[6:3]), .Y(_08613_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31862_ ( .A({ _maxi_write_size[0], _08615_, _maxi_write_size[32:31] }), .Y(_08614_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31863_ ( .A({ _maxi_write_size[29:28], _maxi_write_size[26], _maxi_write_size[23] }), .Y(_08615_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31864_ ( .A({ _maxi_write_size[30], _maxi_write_size[27], _maxi_write_size[25:24] }), .Y(_08616_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31865_ ( .A(__variable_wdata_195), .Y(_05224_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31866_ ( .A({ __variable_wdata_195[0], __variable_wdata_195[1] }), .Y(_05225_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31867_ ( .A(__variable_wdata_195), .Y(_05226_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31868_ ( .A(__variable_wdata_196), .Y(_05227_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31869_ ( .A({ __variable_wdata_196[0], __variable_wdata_196[1] }), .Y(_05228_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31870_ ( .A(__variable_wdata_196), .Y(_05229_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31871_ ( .A({ _tmp_3, saxi_bvalid, _05867_, _04904_ }), .Y(saxi_awready) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31872_ ( .A({ _tmp_1, _tmp_2 }), .Y(_05867_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _31873_ ( .A({ _tmp_4, _05867_, _04904_ }), .Y(saxi_arready) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _31874_ ( .A({ _08621_, _08620_, _08618_, _08619_ }), .Y(_08617_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31875_ ( .A({ conv2d_8_row_count[2], _04498_ }), .Y(_08618_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _31876_ ( .A({ _04476_, _04487_, conv2d_8_row_count[0], conv2d_8_row_count[1] }), .Y(_08619_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31877_ ( .A({ _04498_, conv2d_8_row_count[2], _04501_, conv2d_8_row_count[3] }), .Y(_08620_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31878_ ( .A({ conv2d_8_row_count[3], _04501_, conv2d_8_row_count[4], _04502_ }), .Y(_08621_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31879_ ( .A({ _04502_, conv2d_8_row_count[4] }), .Y(_08622_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31880_ ( .A({ _04505_, conv2d_8_row_count[7], _04506_, conv2d_8_row_count[8] }), .Y(_08623_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31881_ ( .A({ _04478_, conv2d_8_row_count[11], _04477_, conv2d_8_row_count[10] }), .Y(_08624_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31882_ ( .A({ conv2d_8_row_count[8], _04506_, conv2d_8_row_count[9], _04507_ }), .Y(_08625_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31883_ ( .A({ conv2d_8_row_count[6], _04504_, conv2d_8_row_count[7], _04505_ }), .Y(_08626_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _31884_ ( .A({ _08630_, _08628_, conv2d_8_row_count[13], _04480_ }), .Y(_08627_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _31885_ ( .A({ _08629_, conv2d_8_row_count[12], _04479_ }), .Y(_08628_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31886_ ( .A({ _04482_, conv2d_8_row_count[15:14], _04481_ }), .Y(_08629_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31887_ ( .A({ conv2d_8_row_count[12], _04479_, conv2d_8_row_count[13], _04480_ }), .Y(_08630_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _31888_ ( .A({ conv2d_8_row_count[10], _04477_, _04478_, conv2d_8_row_count[11] }), .Y(_08631_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31889_ ( .A({ _08638_, _08637_, _08633_ }), .Y(_08632_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _31890_ ( .A({ _08636_, _08634_, conv2d_8_row_count[28], _04496_ }), .Y(_08633_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _31891_ ( .A({ _08635_, conv2d_8_row_count[29], _04497_ }), .Y(_08634_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31892_ ( .A({ _04500_, conv2d_8_row_count[31], _04499_, conv2d_8_row_count[30] }), .Y(_08635_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31893_ ( .A({ conv2d_8_row_count[28], _04496_, conv2d_8_row_count[29], _04497_ }), .Y(_08636_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31894_ ( .A({ conv2d_8_row_count[27], _04495_, _04494_, conv2d_8_row_count[26] }), .Y(_08637_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31895_ ( .A({ _04493_, conv2d_8_row_count[25], _04492_, conv2d_8_row_count[24] }), .Y(_08638_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31896_ ( .A({ conv2d_8_row_count[16], _04483_, conv2d_8_row_count[17], _04484_ }), .Y(_08639_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _31897_ ( .A({ _08641_, _04485_, conv2d_8_row_count[18] }), .Y(_08640_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _31898_ ( .A({ _04486_, conv2d_8_row_count[19], _04484_, conv2d_8_row_count[17] }), .Y(_08641_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _31899_ ( .A({ _08629_, _08630_, conv2d_8_row_count[13], _04480_ }), .Y(_08642_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _31900_ ( .A({ conv2d_8_row_count[14], _04481_, _04482_, conv2d_8_row_count[15] }), .Y(_08643_) );
  \$lut  #( .LUT(16'h000b), .WIDTH(4) ) _31901_ ( .A({ _08648_, _08645_, _08634_, _08636_ }), .Y(_08644_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _31902_ ( .A({ _08633_, _08647_, _08637_, _08646_ }), .Y(_08645_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _31903_ ( .A({ conv2d_8_row_count[24], _04492_, _04493_, conv2d_8_row_count[25] }), .Y(_08646_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _31904_ ( .A({ conv2d_8_row_count[26], conv2d_8_row_count[27], _04494_, _04495_ }), .Y(_08647_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _31905_ ( .A({ conv2d_8_row_count[30], _04499_, _04500_, conv2d_8_row_count[31] }), .Y(_08648_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _31906_ ( .A({ _08652_, _08650_, _08640_, _08639_ }), .Y(_08649_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _31907_ ( .A({ _08651_, conv2d_8_row_count[20], _04488_ }), .Y(_08650_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _31908_ ( .A({ conv2d_8_row_count[18], _04485_, _04486_, conv2d_8_row_count[19] }), .Y(_08651_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31909_ ( .A({ _04488_, conv2d_8_row_count[20], _04489_, conv2d_8_row_count[21] }), .Y(_08652_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31910_ ( .A({ conv2d_8_row_count[21], _04489_, conv2d_8_row_count[22], _04490_ }), .Y(_08653_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31911_ ( .A({ cparam_conv2d_8_pad_col_left, _08655_, conv2d_8_row_count[4:3] }), .Y(_08654_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31912_ ( .A({ _07440_, conv2d_8_row_count[2:0] }), .Y(_08655_) );
  \$lut  #( .LUT(16'hfeff), .WIDTH(4) ) _31913_ ( .A({ _08698_, _08713_, _08710_, _08656_ }), .Y(conv2d_8_dma_pad_mask_1) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _31914_ ( .A({ _08692_, _08680_, _08690_, _08657_ }), .Y(_08656_) );
  \$lut  #( .LUT(16'hbf00), .WIDTH(4) ) _31915_ ( .A({ _08675_, _08679_, _08676_, _08658_ }), .Y(_08657_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _31916_ ( .A({ _08671_, _08668_, _08674_, _08659_ }), .Y(_08658_) );
  \$lut  #( .LUT(16'h00f4), .WIDTH(4) ) _31917_ ( .A({ _08665_, _08666_, _08667_, _08660_ }), .Y(_08659_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _31918_ ( .A({ _08664_, _08663_, _08661_, _08662_ }), .Y(_08660_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31919_ ( .A({ _04530_, _04498_ }), .Y(_08661_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _31920_ ( .A({ _04476_, _04508_, _04519_, _04487_ }), .Y(_08662_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31921_ ( .A({ _04498_, _04530_, _04501_, _04533_ }), .Y(_08663_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31922_ ( .A({ _04534_, _04502_, _04533_, _04501_ }), .Y(_08664_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31923_ ( .A({ _04504_, _04536_ }), .Y(_08665_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31924_ ( .A({ _04535_, _04503_ }), .Y(_08666_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31925_ ( .A({ _04502_, _04534_, _04503_, _04535_ }), .Y(_08667_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _31926_ ( .A({ _08670_, _08669_, _04537_, _04505_ }), .Y(_08668_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31927_ ( .A({ _04478_, _04510_, _04509_, _04477_ }), .Y(_08669_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31928_ ( .A({ _04539_, _04507_, _04538_, _04506_ }), .Y(_08670_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _31929_ ( .A({ _08672_, _08669_, _08673_ }), .Y(_08671_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _31930_ ( .A({ _04509_, _04477_, _04478_, _04510_ }), .Y(_08672_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _31931_ ( .A({ _04538_, _04539_, _04506_, _04507_ }), .Y(_08673_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31932_ ( .A({ _04536_, _04504_, _04537_, _04505_ }), .Y(_08674_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _31933_ ( .A({ _08677_, _08676_, _08678_ }), .Y(_08675_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31934_ ( .A({ _04514_, _04482_, _04513_, _04481_ }), .Y(_08676_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _31935_ ( .A({ _04513_, _04514_, _04481_, _04482_ }), .Y(_08677_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _31936_ ( .A({ _04511_, _04512_, _04479_, _04480_ }), .Y(_08678_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31937_ ( .A({ _04512_, _04480_, _04511_, _04479_ }), .Y(_08679_) );
  \$lut  #( .LUT(16'h000b), .WIDTH(4) ) _31938_ ( .A({ _08689_, _08681_, _08683_, _08685_ }), .Y(_08680_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _31939_ ( .A({ _08682_, _08687_, _08688_, _08686_ }), .Y(_08681_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _31940_ ( .A({ _08685_, _08683_, _04488_, _04520_ }), .Y(_08682_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _31941_ ( .A({ _08684_, _04522_, _04490_ }), .Y(_08683_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _31942_ ( .A({ _04523_, _04491_, _04489_, _04521_ }), .Y(_08684_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31943_ ( .A({ _04520_, _04488_, _04521_, _04489_ }), .Y(_08685_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31944_ ( .A({ _04518_, _04486_, _04517_, _04485_ }), .Y(_08686_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _31945_ ( .A({ _04517_, _04518_, _04485_, _04486_ }), .Y(_08687_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _31946_ ( .A({ _04515_, _04516_, _04483_, _04484_ }), .Y(_08688_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _31947_ ( .A({ _04522_, _04523_, _04490_, _04491_ }), .Y(_08689_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31948_ ( .A({ _08691_, _08686_, _08682_ }), .Y(_08690_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31949_ ( .A({ _04516_, _04484_, _04515_, _04483_ }), .Y(_08691_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31950_ ( .A({ _08697_, _08696_, _08693_ }), .Y(_08692_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31951_ ( .A({ _08695_, _08694_ }), .Y(_08693_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31952_ ( .A({ _04532_, _04500_, _04531_, _04499_ }), .Y(_08694_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31953_ ( .A({ _04496_, _04528_, _04529_, _04497_ }), .Y(_08695_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31954_ ( .A({ _04527_, _04495_, _04526_, _04494_ }), .Y(_08696_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31955_ ( .A({ _04525_, _04493_, _04524_, _04492_ }), .Y(_08697_) );
  \$lut  #( .LUT(16'h7f00), .WIDTH(4) ) _31956_ ( .A({ _08709_, _08707_, _08703_, _08699_ }), .Y(_08698_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31957_ ( .A({ _08702_, _08700_, _04529_, _04526_ }), .Y(_08699_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31958_ ( .A({ _08701_, _04517_, _04516_, _04537_ }), .Y(_08700_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31959_ ( .A({ cparam_conv2d_8_pad_col_left, _04520_, _04518_, _04533_ }), .Y(_08701_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31960_ ( .A({ _04510_, _04509_, _04539_, _04538_ }), .Y(_08702_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31961_ ( .A({ _08706_, _08704_, _04532_, _04525_ }), .Y(_08703_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31962_ ( .A({ _08705_, _04524_, _04522_, _04534_ }), .Y(_08704_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31963_ ( .A({ _04531_, _04523_, _04536_, _04519_ }), .Y(_08705_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31964_ ( .A({ _04515_, _04512_, _04530_, _04508_ }), .Y(_08706_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31965_ ( .A({ _08708_, _04528_, _04527_, _04521_ }), .Y(_08707_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31966_ ( .A({ _04514_, _04513_, _04511_, _04535_ }), .Y(_08708_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _31967_ ( .A({ _04531_, _04532_, _04499_, _04500_ }), .Y(_08709_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _31968_ ( .A({ _08693_, _08712_, _08711_, _08696_ }), .Y(_08710_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _31969_ ( .A({ _04524_, _04525_, _04492_, _04493_ }), .Y(_08711_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _31970_ ( .A({ _04526_, _04527_, _04494_, _04495_ }), .Y(_08712_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31971_ ( .A({ _08714_, _08694_ }), .Y(_08713_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _31972_ ( .A({ _04528_, _04529_, _04496_, _04497_ }), .Y(_08714_) );
  \$lut  #( .LUT(16'hf2ff), .WIDTH(4) ) _31973_ ( .A({ _08753_, _08766_, _08715_, _08738_ }), .Y(conv2d_8_dma_pad_mask_2) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _31974_ ( .A({ _08735_, _08732_, _08716_, _08730_ }), .Y(_08715_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _31975_ ( .A({ _08728_, _08725_, _08729_, _08717_ }), .Y(_08716_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _31976_ ( .A({ _08718_, _04568_, _04504_ }), .Y(_08717_) );
  \$lut  #( .LUT(16'hddd4), .WIDTH(4) ) _31977_ ( .A({ _08724_, _08719_, _04503_, _04567_ }), .Y(_08718_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _31978_ ( .A({ _08723_, _08722_, _08721_, _08720_ }), .Y(_08719_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31979_ ( .A({ _04487_, _04551_, _04476_, _04540_ }), .Y(_08720_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31980_ ( .A({ _04551_, _04487_, _04562_, _04498_ }), .Y(_08721_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31981_ ( .A({ _04498_, _04562_, _04501_, _04565_ }), .Y(_08722_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31982_ ( .A({ _04566_, _04502_, _04565_, _04501_ }), .Y(_08723_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31983_ ( .A({ _04502_, _04566_ }), .Y(_08724_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _31984_ ( .A({ _08727_, _08726_, _04569_, _04505_ }), .Y(_08725_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31985_ ( .A({ _04478_, _04542_, _04541_, _04477_ }), .Y(_08726_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31986_ ( .A({ _04571_, _04507_, _04570_, _04506_ }), .Y(_08727_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _31987_ ( .A({ _04541_, _04477_, _04478_, _04542_ }), .Y(_08728_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31988_ ( .A({ _04568_, _04504_, _04569_, _04505_ }), .Y(_08729_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _31989_ ( .A({ _08726_, _04571_, _04507_, _08731_ }), .Y(_08730_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31990_ ( .A({ _04570_, _04506_ }), .Y(_08731_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31991_ ( .A({ _08734_, _08733_ }), .Y(_08732_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31992_ ( .A({ _04482_, _04546_, _04545_, _04481_ }), .Y(_08733_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _31993_ ( .A({ _04544_, _04480_, _04543_, _04479_ }), .Y(_08734_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _31994_ ( .A({ _08737_, _08733_, _08736_ }), .Y(_08735_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _31995_ ( .A({ _04543_, _04544_, _04479_, _04480_ }), .Y(_08736_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _31996_ ( .A({ _04545_, _04481_, _04482_, _04546_ }), .Y(_08737_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _31997_ ( .A({ _08749_, _08739_, _04483_, _04547_ }), .Y(_08738_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31998_ ( .A({ _08748_, _08746_, _08740_ }), .Y(_08739_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31999_ ( .A({ _08745_, _08744_, _08741_ }), .Y(_08740_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32000_ ( .A({ _08743_, _08742_ }), .Y(_08741_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32001_ ( .A({ _04564_, _04500_, _04563_, _04499_ }), .Y(_08742_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32002_ ( .A({ _04496_, _04560_, _04561_, _04497_ }), .Y(_08743_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32003_ ( .A({ _04559_, _04495_, _04558_, _04494_ }), .Y(_08744_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32004_ ( .A({ _04557_, _04493_, _04556_, _04492_ }), .Y(_08745_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _32005_ ( .A({ _08747_, _04484_, _04548_ }), .Y(_08746_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32006_ ( .A({ _04550_, _04486_, _04549_, _04485_ }), .Y(_08747_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32007_ ( .A({ _04547_, _04483_, _04548_, _04484_ }), .Y(_08748_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _32008_ ( .A({ _08752_, _08750_, _04488_, _04552_ }), .Y(_08749_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _32009_ ( .A({ _08751_, _04489_, _04553_ }), .Y(_08750_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32010_ ( .A({ _04491_, _04555_, _04554_, _04490_ }), .Y(_08751_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32011_ ( .A({ _04552_, _04488_, _04553_, _04489_ }), .Y(_08752_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _32012_ ( .A({ _08763_, _08760_, _08754_ }), .Y(_08753_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32013_ ( .A({ _08740_, _08758_, _08749_, _08755_ }), .Y(_08754_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _32014_ ( .A({ _08756_, _08746_, _08748_ }), .Y(_08755_) );
  \$lut  #( .LUT(8'h71), .WIDTH(3) ) _32015_ ( .A({ _04486_, _04550_, _08757_ }), .Y(_08756_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32016_ ( .A({ _04549_, _04485_ }), .Y(_08757_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _32017_ ( .A({ _08759_, _08750_, _08752_ }), .Y(_08758_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32018_ ( .A({ _04554_, _04490_, _04491_, _04555_ }), .Y(_08759_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _32019_ ( .A({ _08741_, _08761_, _08762_, _08744_ }), .Y(_08760_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32020_ ( .A({ _04558_, _04559_, _04494_, _04495_ }), .Y(_08761_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32021_ ( .A({ _04556_, _04557_, _04492_, _04493_ }), .Y(_08762_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _32022_ ( .A({ _08765_, _08742_, _08764_ }), .Y(_08763_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32023_ ( .A({ _04560_, _04561_, _04496_, _04497_ }), .Y(_08764_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _32024_ ( .A({ _04563_, _04564_, _04499_, _04500_ }), .Y(_08765_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32025_ ( .A({ _08777_, _08776_, _08767_ }), .Y(_08766_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32026_ ( .A({ _08775_, _08774_, _08772_, _08768_ }), .Y(_08767_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32027_ ( .A({ _08771_, _08770_, _08769_ }), .Y(_08768_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _32028_ ( .A({ _04564_, _04563_, _04561_ }), .Y(_08769_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32029_ ( .A({ _04560_, _04559_, _04558_, _04557_ }), .Y(_08770_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32030_ ( .A({ _04556_, _04555_, _04554_, _04553_ }), .Y(_08771_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32031_ ( .A({ _08773_, cparam_conv2d_8_pad_col_left, _04540_ }), .Y(_08772_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32032_ ( .A({ _04566_, _04565_, _04562_, _04551_ }), .Y(_08773_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32033_ ( .A({ _04552_, _04550_, _04549_, _04548_ }), .Y(_08774_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32034_ ( .A({ _04547_, _04546_, _04545_, _04544_ }), .Y(_08775_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32035_ ( .A({ _04543_, _04542_, _04541_, _04571_ }), .Y(_08776_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32036_ ( .A({ _04570_, _04569_, _04568_, _04567_ }), .Y(_08777_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32037_ ( .A({ _08825_, _08778_ }), .Y(conv2d_8_stream_pad_mask_0_0) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32038_ ( .A({ _11253_, _08794_, _08822_, _11249_ }), .Y(_08778_) );
  \$lut  #( .LUT(16'hf100), .WIDTH(4) ) _32039_ ( .A({ _08787_, _08785_, _08786_, _08780_ }), .Y(_08779_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32040_ ( .A({ _08784_, _08783_, _08782_, _08781_ }), .Y(_08780_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32041_ ( .A({ conv2d_8_col_count[2], _04498_ }), .Y(_08781_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32042_ ( .A({ _04476_, _04487_, conv2d_8_col_count[0], conv2d_8_col_count[1] }), .Y(_08782_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32043_ ( .A({ _04498_, conv2d_8_col_count[2], _04501_, conv2d_8_col_count[3] }), .Y(_08783_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32044_ ( .A({ conv2d_8_col_count[4], _04502_, conv2d_8_col_count[3], _04501_ }), .Y(_08784_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32045_ ( .A({ conv2d_8_col_count[5], _04503_ }), .Y(_08785_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32046_ ( .A({ _04502_, conv2d_8_col_count[4] }), .Y(_08786_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32047_ ( .A({ _04503_, conv2d_8_col_count[5], _04504_, conv2d_8_col_count[6] }), .Y(_08787_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32048_ ( .A({ _04478_, conv2d_8_col_count[11], _04477_, conv2d_8_col_count[10] }), .Y(_08788_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32049_ ( .A({ _04505_, conv2d_8_col_count[7], _04506_, conv2d_8_col_count[8] }), .Y(_08789_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32050_ ( .A({ conv2d_8_col_count[7], _04505_, conv2d_8_col_count[6], _04504_ }), .Y(_08790_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32051_ ( .A({ conv2d_8_col_count[8], _04506_, conv2d_8_col_count[9], _04507_ }), .Y(_08791_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32052_ ( .A({ _04482_, conv2d_8_col_count[15:14], _04481_ }), .Y(_08792_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32053_ ( .A({ conv2d_8_col_count[10], _04477_, _04478_, conv2d_8_col_count[11] }), .Y(_08793_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32054_ ( .A({ _08808_, _08807_, _08805_, _08795_ }), .Y(_08794_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _32055_ ( .A({ _08804_, _08796_, conv2d_8_col_count[21], _04489_ }), .Y(_08795_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32056_ ( .A({ _08803_, _08802_, _08797_ }), .Y(_08796_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _32057_ ( .A({ _08801_, _08798_, _08799_, _08800_ }), .Y(_08797_) );
  \$lut  #( .LUT(4'h9), .WIDTH(2) ) _32058_ ( .A({ _04500_, conv2d_8_col_count[31] }), .Y(_08798_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _32059_ ( .A({ _04499_, conv2d_8_col_count[30], _04497_, conv2d_8_col_count[29] }), .Y(_08799_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32060_ ( .A({ _04496_, conv2d_8_col_count[28] }), .Y(_08800_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32061_ ( .A({ conv2d_8_col_count[28], _04496_, conv2d_8_col_count[29], _04497_ }), .Y(_08801_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32062_ ( .A({ conv2d_8_col_count[27], _04495_, conv2d_8_col_count[26], _04494_ }), .Y(_08802_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32063_ ( .A({ _04493_, conv2d_8_col_count[25], _04492_, conv2d_8_col_count[24] }), .Y(_08803_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32064_ ( .A({ conv2d_8_col_count[22], _04490_, _04491_, conv2d_8_col_count[23] }), .Y(_08804_) );
  \$lut  #( .LUT(8'h41), .WIDTH(3) ) _32065_ ( .A({ _04488_, conv2d_8_col_count[20], _08806_ }), .Y(_08805_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32066_ ( .A({ conv2d_8_col_count[21], _04489_ }), .Y(_08806_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32067_ ( .A({ conv2d_8_col_count[19], _04486_, conv2d_8_col_count[18], _04485_ }), .Y(_08807_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32068_ ( .A({ _04484_, conv2d_8_col_count[17], _04483_, conv2d_8_col_count[16] }), .Y(_08808_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _32069_ ( .A({ _08815_, _08810_, _07383_, _08813_ }), .Y(_08809_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _32070_ ( .A({ _08797_, _08812_, _08811_, _08802_ }), .Y(_08810_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _32071_ ( .A({ conv2d_8_col_count[24], _04492_, _04493_, conv2d_8_col_count[25] }), .Y(_08811_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32072_ ( .A({ conv2d_8_col_count[26], conv2d_8_col_count[27], _04494_, _04495_ }), .Y(_08812_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32073_ ( .A({ _08814_, cparam_conv2d_8_pad_col_left, conv2d_8_col_count[0] }), .Y(_08813_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32074_ ( .A({ conv2d_8_col_count[3:2], conv2d_8_col_count[4], conv2d_8_col_count[1] }), .Y(_08814_) );
  \$lut  #( .LUT(16'hbf00), .WIDTH(4) ) _32075_ ( .A({ _08816_, _08798_, _08799_, _08801_ }), .Y(_08815_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32076_ ( .A({ conv2d_8_col_count[30], _04499_, _04500_, conv2d_8_col_count[31] }), .Y(_08816_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32077_ ( .A({ conv2d_8_col_count[16], _04483_, _04484_, conv2d_8_col_count[17] }), .Y(_08817_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32078_ ( .A({ conv2d_8_col_count[18], conv2d_8_col_count[19], _04485_, _04486_ }), .Y(_08818_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32079_ ( .A({ conv2d_8_col_count[23], _04491_, conv2d_8_col_count[22], _04490_ }), .Y(_08819_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32080_ ( .A({ _04489_, conv2d_8_col_count[21], _04490_, conv2d_8_col_count[22] }), .Y(_08820_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _32081_ ( .A({ _08796_, conv2d_8_col_count[23], _04491_ }), .Y(_08821_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _32082_ ( .A({ _08824_, _08792_, _08823_ }), .Y(_08822_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32083_ ( .A({ conv2d_8_col_count[12], _04479_, _04480_, conv2d_8_col_count[13] }), .Y(_08823_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32084_ ( .A({ conv2d_8_col_count[14], _04481_, _04482_, conv2d_8_col_count[15] }), .Y(_08824_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _32085_ ( .A({ _08866_, _08826_, _08860_, _08846_ }), .Y(_08825_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32086_ ( .A({ _08841_, _08857_, _08854_, _11256_ }), .Y(_08826_) );
  \$lut  #( .LUT(16'hf100), .WIDTH(4) ) _32087_ ( .A({ _08835_, _08833_, _08834_, _08828_ }), .Y(_08827_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _32088_ ( .A({ _08832_, _08831_, _08829_, _08830_ }), .Y(_08828_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32089_ ( .A({ conv2d_8_row_count_buf[2], _04498_ }), .Y(_08829_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32090_ ( .A({ _04476_, conv2d_8_row_count_buf[0], conv2d_8_row_count_buf[1], _04487_ }), .Y(_08830_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32091_ ( .A({ _04498_, conv2d_8_row_count_buf[2], _04501_, conv2d_8_row_count_buf[3] }), .Y(_08831_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32092_ ( .A({ conv2d_8_row_count_buf[4], _04502_, conv2d_8_row_count_buf[3], _04501_ }), .Y(_08832_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32093_ ( .A({ conv2d_8_row_count_buf[5], _04503_ }), .Y(_08833_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32094_ ( .A({ _04502_, conv2d_8_row_count_buf[4] }), .Y(_08834_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32095_ ( .A({ _04503_, conv2d_8_row_count_buf[5], _04504_, conv2d_8_row_count_buf[6] }), .Y(_08835_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32096_ ( .A({ _04478_, conv2d_8_row_count_buf[11:10], _04477_ }), .Y(_08836_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _32097_ ( .A({ conv2d_8_row_count_buf[10], _04477_, _04478_, conv2d_8_row_count_buf[11] }), .Y(_08837_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _32098_ ( .A({ _08839_, _08836_, conv2d_8_row_count_buf[7], _04505_ }), .Y(_08838_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32099_ ( .A({ conv2d_8_row_count_buf[9], _04507_, conv2d_8_row_count_buf[8], _04506_ }), .Y(_08839_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32100_ ( .A({ conv2d_8_row_count_buf[6], _04504_, conv2d_8_row_count_buf[7], _04505_ }), .Y(_08840_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32101_ ( .A({ _08853_, _08852_, _08846_, _08842_ }), .Y(_08841_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _32102_ ( .A({ _08845_, _08843_, _04488_, conv2d_8_row_count_buf[20] }), .Y(_08842_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _32103_ ( .A({ _08844_, _04489_, conv2d_8_row_count_buf[21] }), .Y(_08843_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32104_ ( .A({ _04491_, conv2d_8_row_count_buf[23:22], _04490_ }), .Y(_08844_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32105_ ( .A({ conv2d_8_row_count_buf[20], _04488_, conv2d_8_row_count_buf[21], _04489_ }), .Y(_08845_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32106_ ( .A({ _08851_, _08850_, _08847_ }), .Y(_08846_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32107_ ( .A({ _08849_, _08848_ }), .Y(_08847_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32108_ ( .A({ conv2d_8_row_count_buf[31], _04500_, conv2d_8_row_count_buf[30], _04499_ }), .Y(_08848_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32109_ ( .A({ _04496_, conv2d_8_row_count_buf[28], conv2d_8_row_count_buf[29], _04497_ }), .Y(_08849_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32110_ ( .A({ conv2d_8_row_count_buf[27], _04495_, conv2d_8_row_count_buf[26], _04494_ }), .Y(_08850_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32111_ ( .A({ conv2d_8_row_count_buf[25], _04493_, conv2d_8_row_count_buf[24], _04492_ }), .Y(_08851_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32112_ ( .A({ conv2d_8_row_count_buf[19], _04486_, conv2d_8_row_count_buf[18], _04485_ }), .Y(_08852_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32113_ ( .A({ conv2d_8_row_count_buf[17], _04484_, conv2d_8_row_count_buf[16], _04483_ }), .Y(_08853_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _32114_ ( .A({ _08856_, _08855_, _04480_, conv2d_8_row_count_buf[13] }), .Y(_08854_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32115_ ( .A({ _04482_, conv2d_8_row_count_buf[15:14], _04481_ }), .Y(_08855_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _32116_ ( .A({ conv2d_8_row_count_buf[12], _04479_, conv2d_8_row_count_buf[13], _04480_ }), .Y(_08856_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _32117_ ( .A({ _08859_, _08855_, _08858_ }), .Y(_08857_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32118_ ( .A({ conv2d_8_row_count_buf[12], conv2d_8_row_count_buf[13], _04479_, _04480_ }), .Y(_08858_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32119_ ( .A({ conv2d_8_row_count_buf[14], _04481_, _04482_, conv2d_8_row_count_buf[15] }), .Y(_08859_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _32120_ ( .A({ _08861_, _08843_, _08845_ }), .Y(_08860_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _32121_ ( .A({ _08865_, _08842_, _08862_ }), .Y(_08861_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _32122_ ( .A({ _08864_, _08852_, _08863_ }), .Y(_08862_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32123_ ( .A({ conv2d_8_row_count_buf[16], conv2d_8_row_count_buf[17], _04483_, _04484_ }), .Y(_08863_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _32124_ ( .A({ conv2d_8_row_count_buf[18], conv2d_8_row_count_buf[19], _04485_, _04486_ }), .Y(_08864_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _32125_ ( .A({ conv2d_8_row_count_buf[22], _04490_, _04491_, conv2d_8_row_count_buf[23] }), .Y(_08865_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32126_ ( .A({ _08885_, _08867_, _08883_ }), .Y(_08866_) );
  \$lut  #( .LUT(16'h001f), .WIDTH(4) ) _32127_ ( .A({ _08868_, _08847_, _08882_, _08880_ }), .Y(_08867_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32128_ ( .A({ _08875_, _08873_, _08869_ }), .Y(_08868_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32129_ ( .A({ _08872_, _08871_, _08870_ }), .Y(_08869_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _32130_ ( .A({ conv2d_8_row_count_buf[29], conv2d_8_row_count_buf[26], conv2d_8_row_count_buf[4] }), .Y(_08870_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32131_ ( .A({ cparam_conv2d_8_pad_col_left, conv2d_8_row_count_buf[20:19], conv2d_8_row_count_buf[3] }), .Y(_08871_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32132_ ( .A({ conv2d_8_row_count_buf[31], conv2d_8_row_count_buf[25], conv2d_8_row_count_buf[6], conv2d_8_row_count_buf[1] }), .Y(_08872_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32133_ ( .A({ _08874_, conv2d_8_row_count_buf[18:17], conv2d_8_row_count_buf[7] }), .Y(_08873_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32134_ ( .A({ conv2d_8_row_count_buf[16], conv2d_8_row_count_buf[13], conv2d_8_row_count_buf[2], conv2d_8_row_count_buf[0] }), .Y(_08874_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32135_ ( .A({ _08879_, _08878_, _08877_, _08876_ }), .Y(_08875_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32136_ ( .A(conv2d_8_row_count_buf[11:8]), .Y(_08876_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _32137_ ( .A({ conv2d_8_row_count_buf[28], conv2d_8_row_count_buf[24], conv2d_8_row_count_buf[22] }), .Y(_08877_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32138_ ( .A({ conv2d_8_row_count_buf[15:14], conv2d_8_row_count_buf[12], conv2d_8_row_count_buf[5] }), .Y(_08878_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32139_ ( .A({ conv2d_8_row_count_buf[30], conv2d_8_row_count_buf[27], conv2d_8_row_count_buf[23], conv2d_8_row_count_buf[21] }), .Y(_08879_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _32140_ ( .A({ _08850_, conv2d_8_row_count_buf[25], _04493_, _08881_ }), .Y(_08880_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32141_ ( .A({ conv2d_8_row_count_buf[24], _04492_ }), .Y(_08881_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32142_ ( .A({ conv2d_8_row_count_buf[26], conv2d_8_row_count_buf[27], _04494_, _04495_ }), .Y(_08882_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _32143_ ( .A({ _08848_, conv2d_8_row_count_buf[29], _04497_, _08884_ }), .Y(_08883_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32144_ ( .A({ conv2d_8_row_count_buf[28], _04496_ }), .Y(_08884_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _32145_ ( .A({ conv2d_8_row_count_buf[30], conv2d_8_row_count_buf[31], _04499_, _04500_ }), .Y(_08885_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32146_ ( .A({ _11258_, _08825_ }), .Y(conv2d_8_stream_pad_mask_0_1) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32147_ ( .A({ _08901_, _08896_, _08903_, _08887_ }), .Y(_08886_) );
  \$lut  #( .LUT(16'hf100), .WIDTH(4) ) _32148_ ( .A({ _08895_, _08893_, _08894_, _08888_ }), .Y(_08887_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32149_ ( .A({ _08892_, _08891_, _08890_, _08889_ }), .Y(_08888_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32150_ ( .A({ _04594_, _04498_ }), .Y(_08889_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32151_ ( .A({ _04476_, _04487_, _04572_, _04583_ }), .Y(_08890_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32152_ ( .A({ _04498_, _04594_, _04501_, _04597_ }), .Y(_08891_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32153_ ( .A({ _04597_, _04501_, _04598_, _04502_ }), .Y(_08892_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32154_ ( .A({ _04599_, _04503_ }), .Y(_08893_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32155_ ( .A({ _04502_, _04598_ }), .Y(_08894_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32156_ ( .A({ _04503_, _04599_, _04504_, _04600_ }), .Y(_08895_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32157_ ( .A({ _08900_, _08897_ }), .Y(_08896_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _32158_ ( .A({ _08898_, _04603_, _04507_ }), .Y(_08897_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32159_ ( .A({ _04478_, _04574_, _04477_, _04573_ }), .Y(_08898_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32160_ ( .A({ _04602_, _04506_, _04603_, _04507_ }), .Y(_08899_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32161_ ( .A({ _04505_, _04601_, _04506_, _04602_ }), .Y(_08900_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _32162_ ( .A({ _08902_, _08897_, _08899_ }), .Y(_08901_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32163_ ( .A({ _04573_, _04477_, _04478_, _04574_ }), .Y(_08902_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32164_ ( .A({ _04600_, _04504_, _04601_, _04505_ }), .Y(_08903_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32165_ ( .A({ _08919_, _08918_, _08912_, _08905_ }), .Y(_08904_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _32166_ ( .A({ _08909_, _08906_, _04587_, _04491_ }), .Y(_08905_) );
  \$lut  #( .LUT(16'h9000), .WIDTH(4) ) _32167_ ( .A({ _08908_, _08907_, _04596_, _04500_ }), .Y(_08906_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _32168_ ( .A({ _04595_, _04499_, _04497_, _04593_ }), .Y(_08907_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _32169_ ( .A({ _04496_, _04592_, _04593_, _04497_ }), .Y(_08908_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _32170_ ( .A({ _08911_, _08910_, _04492_, _04588_ }), .Y(_08909_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32171_ ( .A({ _04591_, _04495_, _04590_, _04494_ }), .Y(_08910_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _32172_ ( .A({ _04589_, _04493_, _04588_, _04492_ }), .Y(_08911_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32173_ ( .A({ _08917_, _08916_, _08913_ }), .Y(_08912_) );
  \$lut  #( .LUT(16'h1001), .WIDTH(4) ) _32174_ ( .A({ _04484_, _04580_, _08915_, _08914_ }), .Y(_08913_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32175_ ( .A({ _04488_, _04584_ }), .Y(_08914_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32176_ ( .A({ _04585_, _04489_ }), .Y(_08915_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32177_ ( .A({ _04586_, _04490_, _04587_, _04491_ }), .Y(_08916_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32178_ ( .A({ _04489_, _04585_, _04490_, _04586_ }), .Y(_08917_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32179_ ( .A({ _04582_, _04486_, _04581_, _04485_ }), .Y(_08918_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _32180_ ( .A({ _04579_, _04483_, _04584_, _04488_ }), .Y(_08919_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32181_ ( .A({ _04482_, _04578_, _04577_, _04481_ }), .Y(_08920_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32182_ ( .A({ _04576_, _04480_, _04575_, _04479_ }), .Y(_08921_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _32183_ ( .A({ _04577_, _04481_, _04482_, _04578_ }), .Y(_08922_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32184_ ( .A({ _04575_, _04576_, _04479_, _04480_ }), .Y(_08923_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32185_ ( .A({ _08918_, _08925_ }), .Y(_08924_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32186_ ( .A({ _04579_, _04483_, _04484_, _04580_ }), .Y(_08925_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _32187_ ( .A({ _04581_, _04582_, _04485_, _04486_ }), .Y(_08926_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32188_ ( .A({ _08928_, _04588_, _04586_, _04598_ }), .Y(_08927_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32189_ ( .A({ _04595_, _04587_, _04600_, _04583_ }), .Y(_08928_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32190_ ( .A({ _08930_, _04593_, _04590_, _04589_ }), .Y(_08929_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32191_ ( .A({ _04579_, _04576_, _04594_, _04572_ }), .Y(_08930_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32192_ ( .A({ _08932_, _04592_, _04591_, _04585_ }), .Y(_08931_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32193_ ( .A({ _04578_, _04577_, _04575_, _04599_ }), .Y(_08932_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32194_ ( .A({ _08934_, _04581_, _04580_, _04601_ }), .Y(_08933_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32195_ ( .A({ cparam_conv2d_8_pad_col_left, _04584_, _04582_, _04597_ }), .Y(_08934_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32196_ ( .A({ _04574_, _04573_, _04603_, _04602_ }), .Y(_08935_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _32197_ ( .A({ _08906_, _08937_, _08938_, _08910_ }), .Y(_08936_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32198_ ( .A({ _04590_, _04591_, _04494_, _04495_ }), .Y(_08937_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32199_ ( .A({ _04588_, _04589_, _04492_, _04493_ }), .Y(_08938_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32200_ ( .A({ _04593_, _04497_, _04592_, _04496_ }), .Y(_08939_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32201_ ( .A({ _08940_, _08825_ }), .Y(conv2d_8_stream_pad_mask_0_2) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _32202_ ( .A({ _08974_, _08995_, _08941_, _11266_ }), .Y(_08940_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32203_ ( .A({ _08949_, _08942_, _04491_, _04619_ }), .Y(_08941_) );
  \$lut  #( .LUT(16'hf400), .WIDTH(4) ) _32204_ ( .A({ _08948_, _08943_, _04617_, _04489_ }), .Y(_08942_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32205_ ( .A({ _08947_, _08944_, _04616_, _04488_ }), .Y(_08943_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32206_ ( .A({ _08946_, _08945_ }), .Y(_08944_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32207_ ( .A({ _04611_, _04483_, _04484_, _04612_ }), .Y(_08945_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32208_ ( .A({ _04614_, _04486_, _04613_, _04485_ }), .Y(_08946_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _32209_ ( .A({ _04613_, _04614_, _04485_, _04486_ }), .Y(_08947_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32210_ ( .A({ _04489_, _04617_, _04490_, _04618_ }), .Y(_08948_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32211_ ( .A({ _04618_, _04490_, _04619_, _04491_ }), .Y(_08949_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32212_ ( .A({ _08963_, _08960_, _08966_, _08951_ }), .Y(_08950_) );
  \$lut  #( .LUT(16'h00f4), .WIDTH(4) ) _32213_ ( .A({ _08957_, _08958_, _08959_, _08952_ }), .Y(_08951_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32214_ ( .A({ _08956_, _08955_, _08954_, _08953_ }), .Y(_08952_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32215_ ( .A({ _04626_, _04498_ }), .Y(_08953_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32216_ ( .A({ _04476_, _04487_, _04604_, _04615_ }), .Y(_08954_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32217_ ( .A({ _04498_, _04626_, _04501_, _04629_ }), .Y(_08955_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32218_ ( .A({ _04629_, _04501_, _04630_, _04502_ }), .Y(_08956_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32219_ ( .A({ _04504_, _04632_ }), .Y(_08957_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32220_ ( .A({ _04631_, _04503_ }), .Y(_08958_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32221_ ( .A({ _04502_, _04630_, _04503_, _04631_ }), .Y(_08959_) );
  \$lut  #( .LUT(16'h9000), .WIDTH(4) ) _32222_ ( .A({ _08962_, _08961_, _04507_, _04635_ }), .Y(_08960_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32223_ ( .A({ _04478_, _04606_, _04477_, _04605_ }), .Y(_08961_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _32224_ ( .A({ _04506_, _04634_, _04505_, _04633_ }), .Y(_08962_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _32225_ ( .A({ _08965_, _08961_, _08964_ }), .Y(_08963_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32226_ ( .A({ _04634_, _04506_, _04507_, _04635_ }), .Y(_08964_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _32227_ ( .A({ _04605_, _04477_, _04478_, _04606_ }), .Y(_08965_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32228_ ( .A({ _04632_, _04504_, _04633_, _04505_ }), .Y(_08966_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32229_ ( .A({ _04488_, _04616_, _04617_, _04489_ }), .Y(_08967_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32230_ ( .A({ _08970_, _08969_ }), .Y(_08968_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32231_ ( .A({ _04482_, _04610_, _04609_, _04481_ }), .Y(_08969_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32232_ ( .A({ _04608_, _04480_, _04607_, _04479_ }), .Y(_08970_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _32233_ ( .A({ _08973_, _08969_, _08972_ }), .Y(_08971_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32234_ ( .A({ _04607_, _04608_, _04479_, _04480_ }), .Y(_08972_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _32235_ ( .A({ _04609_, _04481_, _04482_, _04610_ }), .Y(_08973_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _32236_ ( .A({ _08994_, _08975_, _08986_, _08992_ }), .Y(_08974_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32237_ ( .A({ _08985_, _08984_, _08983_, _08976_ }), .Y(_08975_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _32238_ ( .A({ _08977_, cparam_conv2d_8_pad_col_left, _08982_, _04604_ }), .Y(_08976_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32239_ ( .A({ _08981_, _08980_, _08979_, _08978_ }), .Y(_08977_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32240_ ( .A({ _04616_, _04614_, _04613_, _04612_ }), .Y(_08978_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32241_ ( .A({ _04611_, _04610_, _04609_, _04608_ }), .Y(_08979_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32242_ ( .A({ _04607_, _04606_, _04605_, _04635_ }), .Y(_08980_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32243_ ( .A({ _04634_, _04633_, _04632_, _04631_ }), .Y(_08981_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32244_ ( .A({ _04630_, _04629_, _04626_, _04615_ }), .Y(_08982_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _32245_ ( .A({ _04628_, _04627_, _04625_ }), .Y(_08983_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32246_ ( .A({ _04624_, _04623_, _04622_, _04621_ }), .Y(_08984_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32247_ ( .A({ _04620_, _04619_, _04618_, _04617_ }), .Y(_08985_) );
  \$lut  #( .LUT(16'hf400), .WIDTH(4) ) _32248_ ( .A({ _08991_, _08987_, _04496_, _04624_ }), .Y(_08986_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _32249_ ( .A({ _08989_, _08988_, _08990_ }), .Y(_08987_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32250_ ( .A({ _04623_, _04495_, _04622_, _04494_ }), .Y(_08988_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32251_ ( .A({ _04622_, _04623_, _04494_, _04495_ }), .Y(_08989_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32252_ ( .A({ _04620_, _04621_, _04492_, _04493_ }), .Y(_08990_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32253_ ( .A({ _04625_, _04497_, _04624_, _04496_ }), .Y(_08991_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _32254_ ( .A({ _08993_, _04497_, _04625_ }), .Y(_08992_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32255_ ( .A({ _04500_, _04628_, _04499_, _04627_ }), .Y(_08993_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32256_ ( .A({ _04627_, _04499_, _04500_, _04628_ }), .Y(_08994_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32257_ ( .A({ _08997_, _08988_, _08996_ }), .Y(_08995_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _32258_ ( .A({ _08991_, _08992_, _04624_, _04496_ }), .Y(_08996_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32259_ ( .A({ _04621_, _04493_, _04620_, _04492_ }), .Y(_08997_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32260_ ( .A({ _08998_, _08778_ }), .Y(conv2d_8_stream_pad_mask_1_0) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _32261_ ( .A({ _09038_, _09062_, _08999_, _09009_ }), .Y(_08998_) );
  \$lut  #( .LUT(16'h004f), .WIDTH(4) ) _32262_ ( .A({ _09006_, _09007_, _09008_, _09000_ }), .Y(_08999_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _32263_ ( .A({ _09001_, _04649_, _04489_ }), .Y(_09000_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32264_ ( .A({ _09005_, _09002_, _04648_, _04488_ }), .Y(_09001_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32265_ ( .A({ _09004_, _09003_ }), .Y(_09002_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32266_ ( .A({ _04643_, _04483_, _04484_, _04644_ }), .Y(_09003_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32267_ ( .A({ _04646_, _04486_, _04645_, _04485_ }), .Y(_09004_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _32268_ ( .A({ _04645_, _04646_, _04485_, _04486_ }), .Y(_09005_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32269_ ( .A({ _04491_, _04651_ }), .Y(_09006_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32270_ ( .A({ _04650_, _04490_, _04651_, _04491_ }), .Y(_09007_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32271_ ( .A({ _04489_, _04649_, _04490_, _04650_ }), .Y(_09008_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32272_ ( .A({ _09027_, _09035_, _09032_, _09010_ }), .Y(_09009_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32273_ ( .A({ _09023_, _09020_, _09026_, _09011_ }), .Y(_09010_) );
  \$lut  #( .LUT(16'h00f4), .WIDTH(4) ) _32274_ ( .A({ _09017_, _09018_, _09019_, _09012_ }), .Y(_09011_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _32275_ ( .A({ _09016_, _09015_, _09013_, _09014_ }), .Y(_09012_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32276_ ( .A({ _04476_, _04636_, _04647_, _04487_ }), .Y(_09013_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _32277_ ( .A({ _04498_, _04658_, _04501_, _04661_ }), .Y(_09014_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _32278_ ( .A({ _04658_, _04498_, _04661_, _04501_ }), .Y(_09015_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32279_ ( .A({ _04662_, _04502_, _04661_, _04501_ }), .Y(_09016_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32280_ ( .A({ _04504_, _04664_ }), .Y(_09017_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32281_ ( .A({ _04663_, _04503_ }), .Y(_09018_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32282_ ( .A({ _04502_, _04662_, _04503_, _04663_ }), .Y(_09019_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _32283_ ( .A({ _09022_, _09021_, _04665_, _04505_ }), .Y(_09020_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32284_ ( .A({ _04478_, _04638_, _04637_, _04477_ }), .Y(_09021_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32285_ ( .A({ _04667_, _04507_, _04666_, _04506_ }), .Y(_09022_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _32286_ ( .A({ _09024_, _09021_, _09025_ }), .Y(_09023_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _32287_ ( .A({ _04637_, _04477_, _04478_, _04638_ }), .Y(_09024_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32288_ ( .A({ _04666_, _04667_, _04506_, _04507_ }), .Y(_09025_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32289_ ( .A({ _04664_, _04504_, _04665_, _04505_ }), .Y(_09026_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32290_ ( .A({ _09031_, _09030_, _09028_ }), .Y(_09027_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32291_ ( .A({ _09004_, _09008_, _09007_, _09029_ }), .Y(_09028_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _32292_ ( .A({ _09006_, _04649_, _04489_ }), .Y(_09029_) );
  \$lut  #( .LUT(4'h9), .WIDTH(2) ) _32293_ ( .A({ _04648_, _04488_ }), .Y(_09030_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32294_ ( .A({ _04484_, _04644_, _04643_, _04483_ }), .Y(_09031_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32295_ ( .A({ _09034_, _09033_ }), .Y(_09032_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32296_ ( .A({ _04482_, _04642_, _04641_, _04481_ }), .Y(_09033_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32297_ ( .A({ _04640_, _04480_, _04639_, _04479_ }), .Y(_09034_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _32298_ ( .A({ _09036_, _09033_, _09037_ }), .Y(_09035_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _32299_ ( .A({ _04641_, _04481_, _04482_, _04642_ }), .Y(_09036_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32300_ ( .A({ _04639_, _04640_, _04479_, _04480_ }), .Y(_09037_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _32301_ ( .A({ _09039_, _09049_, _09041_, _09043_ }), .Y(_09038_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _32302_ ( .A({ _09048_, _09040_, _09044_ }), .Y(_09039_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _32303_ ( .A({ _09043_, _09041_, _04656_, _04496_ }), .Y(_09040_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _32304_ ( .A({ _09042_, _04660_, _04500_ }), .Y(_09041_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _32305_ ( .A({ _04659_, _04499_, _04497_, _04657_ }), .Y(_09042_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32306_ ( .A({ _04657_, _04497_, _04656_, _04496_ }), .Y(_09043_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _32307_ ( .A({ _09046_, _09045_, _09047_ }), .Y(_09044_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32308_ ( .A({ _04655_, _04495_, _04654_, _04494_ }), .Y(_09045_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32309_ ( .A({ _04654_, _04655_, _04494_, _04495_ }), .Y(_09046_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32310_ ( .A({ _04652_, _04653_, _04492_, _04493_ }), .Y(_09047_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _32311_ ( .A({ _04659_, _04660_, _04499_, _04500_ }), .Y(_09048_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32312_ ( .A({ _09059_, _09056_, _09054_, _09050_ }), .Y(_09049_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32313_ ( .A({ _09053_, _09052_, _09051_ }), .Y(_09050_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _32314_ ( .A({ _04660_, _04659_, _04657_ }), .Y(_09051_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32315_ ( .A({ _04656_, _04655_, _04654_, _04653_ }), .Y(_09052_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32316_ ( .A({ _04652_, _04651_, _04650_, _04649_ }), .Y(_09053_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32317_ ( .A({ _09055_, cparam_conv2d_8_pad_col_left, _04636_ }), .Y(_09054_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32318_ ( .A({ _04662_, _04661_, _04658_, _04647_ }), .Y(_09055_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32319_ ( .A({ _09058_, _09057_ }), .Y(_09056_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32320_ ( .A({ _04639_, _04638_, _04637_, _04667_ }), .Y(_09057_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32321_ ( .A({ _04666_, _04665_, _04664_, _04663_ }), .Y(_09058_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32322_ ( .A({ _09061_, _09060_ }), .Y(_09059_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32323_ ( .A({ _04648_, _04646_, _04645_, _04644_ }), .Y(_09060_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32324_ ( .A({ _04643_, _04642_, _04641_, _04640_ }), .Y(_09061_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32325_ ( .A({ _09063_, _09045_, _09040_ }), .Y(_09062_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32326_ ( .A({ _04653_, _04493_, _04652_, _04492_ }), .Y(_09063_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32327_ ( .A({ _08998_, _11258_ }), .Y(conv2d_8_stream_pad_mask_1_1) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32328_ ( .A({ _08998_, _08940_ }), .Y(conv2d_8_stream_pad_mask_1_2) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32329_ ( .A({ _09064_, _08778_ }), .Y(conv2d_8_stream_pad_mask_2_0) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32330_ ( .A({ _09083_, _11272_, _09121_, _09065_ }), .Y(_09064_) );
  \$lut  #( .LUT(16'hf400), .WIDTH(4) ) _32331_ ( .A({ _09080_, _09081_, _09082_, _11269_ }), .Y(_09065_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32332_ ( .A({ _09074_, _09073_, _09072_, _09067_ }), .Y(_09066_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32333_ ( .A({ _09071_, _09070_, _09069_, _09068_ }), .Y(_09067_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32334_ ( .A({ _04476_, _04668_, _04487_, _04679_ }), .Y(_09068_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32335_ ( .A({ _04679_, _04487_, _04690_, _04498_ }), .Y(_09069_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32336_ ( .A({ _04498_, _04690_, _04501_, _04693_ }), .Y(_09070_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32337_ ( .A({ _04693_, _04501_, _04694_, _04502_ }), .Y(_09071_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32338_ ( .A({ _04502_, _04694_, _04503_, _04695_ }), .Y(_09072_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32339_ ( .A({ _04695_, _04503_, _04696_, _04504_ }), .Y(_09073_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32340_ ( .A({ _04504_, _04696_, _04505_, _04697_ }), .Y(_09074_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32341_ ( .A({ _04478_, _04670_, _04477_, _04669_ }), .Y(_09075_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _32342_ ( .A({ _09077_, _09075_, _09078_ }), .Y(_09076_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32343_ ( .A({ _04669_, _04477_, _04478_, _04670_ }), .Y(_09077_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32344_ ( .A({ _04698_, _04506_, _04507_, _04699_ }), .Y(_09078_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32345_ ( .A({ _04697_, _04505_ }), .Y(_09079_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32346_ ( .A({ _04482_, _04674_, _04673_, _04481_ }), .Y(_09080_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32347_ ( .A({ _04671_, _04672_, _04479_, _04480_ }), .Y(_09081_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32348_ ( .A({ _04672_, _04480_, _04671_, _04479_ }), .Y(_09082_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _32349_ ( .A({ _09108_, _09095_, _09084_ }), .Y(_09083_) );
  \$lut  #( .LUT(16'h40ff), .WIDTH(4) ) _32350_ ( .A({ _09085_, _09094_, _09088_, _09090_ }), .Y(_09084_) );
  \$lut  #( .LUT(16'h0071), .WIDTH(4) ) _32351_ ( .A({ _09086_, _04500_, _04692_, _09089_ }), .Y(_09085_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _32352_ ( .A({ _09088_, _09087_, _04497_, _04689_ }), .Y(_09086_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32353_ ( .A({ _04689_, _04497_, _04688_, _04496_ }), .Y(_09087_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32354_ ( .A({ _04500_, _04692_, _04499_, _04691_ }), .Y(_09088_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32355_ ( .A({ _04691_, _04499_ }), .Y(_09089_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _32356_ ( .A({ _09092_, _09091_, _09093_ }), .Y(_09090_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32357_ ( .A({ _04687_, _04495_, _04686_, _04494_ }), .Y(_09091_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32358_ ( .A({ _04686_, _04687_, _04494_, _04495_ }), .Y(_09092_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _32359_ ( .A({ _04684_, _04685_, _04492_, _04493_ }), .Y(_09093_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32360_ ( .A({ _04496_, _04688_, _04689_, _04497_ }), .Y(_09094_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _32361_ ( .A({ _09096_, _09106_, _09107_, _09099_ }), .Y(_09095_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _32362_ ( .A({ _09097_, _04683_, _04491_ }), .Y(_09096_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32363_ ( .A({ _09098_, _09094_, _09088_, _09091_ }), .Y(_09097_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32364_ ( .A({ _04685_, _04493_, _04684_, _04492_ }), .Y(_09098_) );
  \$lut  #( .LUT(16'h00f4), .WIDTH(4) ) _32365_ ( .A({ _09105_, _09100_, _04488_, _04680_ }), .Y(_09099_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _32366_ ( .A({ _09104_, _09101_, _09102_, _09103_ }), .Y(_09100_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32367_ ( .A({ _04680_, _04488_ }), .Y(_09101_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _32368_ ( .A({ _04486_, _04678_, _04677_, _04485_ }), .Y(_09102_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _32369_ ( .A({ _04675_, _04483_, _04484_, _04676_ }), .Y(_09103_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32370_ ( .A({ _04677_, _04485_, _04486_, _04678_ }), .Y(_09104_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32371_ ( .A({ _04681_, _04489_ }), .Y(_09105_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32372_ ( .A({ _04682_, _04490_, _04683_, _04491_ }), .Y(_09106_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32373_ ( .A({ _04489_, _04681_, _04490_, _04682_ }), .Y(_09107_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32374_ ( .A({ _09119_, _09117_, _09109_ }), .Y(_09108_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32375_ ( .A({ _09116_, _09115_, _09112_, _09110_ }), .Y(_09109_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32376_ ( .A({ _09111_, cparam_conv2d_8_pad_col_left, _04668_ }), .Y(_09110_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32377_ ( .A({ _04694_, _04693_, _04690_, _04679_ }), .Y(_09111_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32378_ ( .A({ _09114_, _09113_ }), .Y(_09112_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32379_ ( .A({ _04680_, _04678_, _04677_, _04676_ }), .Y(_09113_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32380_ ( .A({ _04675_, _04674_, _04673_, _04672_ }), .Y(_09114_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32381_ ( .A({ _04671_, _04670_, _04669_, _04699_ }), .Y(_09115_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32382_ ( .A({ _04698_, _04697_, _04696_, _04695_ }), .Y(_09116_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32383_ ( .A({ _09118_, _04683_, _04682_, _04681_ }), .Y(_09117_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32384_ ( .A({ _04688_, _04687_, _04686_, _04685_ }), .Y(_09118_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32385_ ( .A({ _04692_, _04691_, _04689_, _04684_ }), .Y(_09119_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _32386_ ( .A({ _09106_, _09101_, _09105_ }), .Y(_09120_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _32387_ ( .A({ _04673_, _04481_, _04482_, _04674_ }), .Y(_09121_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32388_ ( .A({ _09064_, _11258_ }), .Y(conv2d_8_stream_pad_mask_2_1) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32389_ ( .A({ _09064_, _08940_ }), .Y(conv2d_8_stream_pad_mask_2_2) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32390_ ( .A({ _07328_, _stream_conv2d_8_source_busy }), .Y(_05863_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32391_ ( .A({ _09128_, _09127_, _09122_ }), .Y(_stream_conv2d_8_done) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32392_ ( .A({ _09126_, _09125_, _09123_ }), .Y(_09122_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32393_ ( .A({ _stream_conv2d_8_source_8_idle, _stream_conv2d_8_source_6_idle, _stream_conv2d_8_source_36_idle, _09124_ }), .Y(_09123_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32394_ ( .A({ _stream_conv2d_8_source_35_idle, _stream_conv2d_8_source_34_idle, _stream_conv2d_8_source_33_idle, _stream_conv2d_8_source_32_idle }), .Y(_09124_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32395_ ( .A({ _stream_conv2d_8_source_31_idle, _stream_conv2d_8_source_30_idle, _stream_conv2d_8_source_29_idle, _stream_conv2d_8_source_28_idle }), .Y(_09125_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32396_ ( .A({ _stream_conv2d_8_source_27_idle, _stream_conv2d_8_source_26_idle, _stream_conv2d_8_source_25_idle, _stream_conv2d_8_source_24_idle }), .Y(_09126_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32397_ ( .A({ _stream_conv2d_8_source_23_idle, _stream_conv2d_8_source_22_idle, _stream_conv2d_8_source_21_idle, _stream_conv2d_8_source_20_idle }), .Y(_09127_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32398_ ( .A({ _stream_conv2d_8_source_19_idle, _stream_conv2d_8_source_14_idle, _stream_conv2d_8_source_12_idle, _stream_conv2d_8_source_10_idle }), .Y(_09128_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32399_ ( .A({ _11277_, _11275_ }), .Y(max_pool_serial_9_stream_pad_mask_0_0) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _32400_ ( .A({ cparam_max_pool_serial_9_act_num_col[2], _09130_, _09131_, max_pool_serial_9_col_count[2] }), .Y(_09129_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _32401_ ( .A({ cparam_max_pool_serial_9_act_num_col[0], max_pool_serial_9_col_count[0], cparam_max_pool_serial_9_act_num_col[1], max_pool_serial_9_col_count[1] }), .Y(_09130_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32402_ ( .A({ max_pool_serial_9_col_count[1], cparam_max_pool_serial_9_act_num_col[1] }), .Y(_09131_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _32403_ ( .A({ cparam_max_pool_serial_9_act_num_col[3], max_pool_serial_9_row_count_buf[3], _09133_ }), .Y(_09132_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _32404_ ( .A({ cparam_max_pool_serial_9_act_num_col[2], max_pool_serial_9_row_count_buf[2], _09134_ }), .Y(_09133_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _32405_ ( .A({ cparam_max_pool_serial_9_act_num_col[0], max_pool_serial_9_row_count_buf[0], max_pool_serial_9_row_count_buf[1], cparam_max_pool_serial_9_act_num_col[1] }), .Y(_09134_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32406_ ( .A({ _09141_, _09140_, _09136_ }), .Y(_09135_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _32407_ ( .A({ _09139_, _09137_, max_pool_serial_9_row_count_buf[8], max_pool_serial_9_row_count_buf[5] }), .Y(_09136_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32408_ ( .A({ _09138_, max_pool_serial_9_row_count_buf[30], max_pool_serial_9_row_count_buf[27:26] }), .Y(_09137_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32409_ ( .A({ max_pool_serial_9_row_count_buf[23:22], max_pool_serial_9_row_count_buf[20], max_pool_serial_9_row_count_buf[17] }), .Y(_09138_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32410_ ( .A({ max_pool_serial_9_row_count_buf[15:14], max_pool_serial_9_row_count_buf[12], max_pool_serial_9_row_count_buf[9] }), .Y(_09139_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32411_ ( .A({ max_pool_serial_9_row_count_buf[24], max_pool_serial_9_row_count_buf[21], max_pool_serial_9_row_count_buf[19:18] }), .Y(_09140_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32412_ ( .A({ max_pool_serial_9_row_count_buf[31], max_pool_serial_9_row_count_buf[29:28], max_pool_serial_9_row_count_buf[25] }), .Y(_09141_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32413_ ( .A({ max_pool_serial_9_row_count_buf[16], max_pool_serial_9_row_count_buf[13], max_pool_serial_9_row_count_buf[11:10] }), .Y(_09142_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32414_ ( .A({ _11280_, _11277_ }), .Y(max_pool_serial_9_stream_pad_mask_0_1) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32415_ ( .A({ _03608_, _03607_, _03606_, _03605_ }), .Y(_09143_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32416_ ( .A({ _03585_, _03584_, _03583_, _03582_ }), .Y(_09144_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32417_ ( .A({ _03581_, _03580_, _03579_, _03609_ }), .Y(_09145_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32418_ ( .A({ _09147_, _03602_, _03601_, _03599_ }), .Y(_09146_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32419_ ( .A({ _03598_, _03597_, _03596_, _03595_ }), .Y(_09147_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32420_ ( .A({ _03594_, _03593_, _03592_, _03591_ }), .Y(_09148_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32421_ ( .A({ _03590_, _03588_, _03587_, _03586_ }), .Y(_09149_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _32422_ ( .A({ cparam_max_pool_serial_9_act_num_col[3], _03603_, _09151_ }), .Y(_09150_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _32423_ ( .A({ cparam_max_pool_serial_9_act_num_col[2], _03600_, _09152_ }), .Y(_09151_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _32424_ ( .A({ cparam_max_pool_serial_9_act_num_col[0], _03578_, _03589_, cparam_max_pool_serial_9_act_num_col[1] }), .Y(_09152_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32425_ ( .A({ _11282_, _11275_ }), .Y(max_pool_serial_9_stream_pad_mask_1_0) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _32426_ ( .A({ cparam_max_pool_serial_9_act_num_col[3], _03635_, _09154_ }), .Y(_09153_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _32427_ ( .A({ cparam_max_pool_serial_9_act_num_col[2], _03632_, _09155_ }), .Y(_09154_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _32428_ ( .A({ cparam_max_pool_serial_9_act_num_col[0], _03610_, _03621_, cparam_max_pool_serial_9_act_num_col[1] }), .Y(_09155_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32429_ ( .A({ _09162_, _09161_, _09157_ }), .Y(_09156_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _32430_ ( .A({ _09160_, _09158_, _03640_, _03637_ }), .Y(_09157_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32431_ ( .A({ _09159_, _03633_, _03629_, _03628_ }), .Y(_09158_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32432_ ( .A({ _03625_, _03624_, _03622_, _03618_ }), .Y(_09159_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32433_ ( .A({ _03616_, _03615_, _03613_, _03641_ }), .Y(_09160_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32434_ ( .A({ _03626_, _03623_, _03620_, _03619_ }), .Y(_09161_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32435_ ( .A({ _03634_, _03631_, _03630_, _03627_ }), .Y(_09162_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32436_ ( .A({ _03617_, _03614_, _03612_, _03611_ }), .Y(_09163_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32437_ ( .A({ _11282_, _11280_ }), .Y(max_pool_serial_9_stream_pad_mask_1_1) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _32438_ ( .A({ _09179_, _09174_, _09169_, _09164_ }), .Y(matmul_15_stream_pad_mask_0_0) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32439_ ( .A({ _09168_, _09167_, _09166_, _09165_ }), .Y(_09164_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32440_ ( .A(matmul_15_row_count_buf[23:20]), .Y(_09165_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32441_ ( .A(matmul_15_row_count_buf[19:16]), .Y(_09166_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32442_ ( .A(matmul_15_row_count_buf[31:28]), .Y(_09167_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32443_ ( .A(matmul_15_row_count_buf[27:24]), .Y(_09168_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32444_ ( .A({ _09173_, _09172_, _09171_, _09170_ }), .Y(_09169_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32445_ ( .A(matmul_15_row_count_buf[7:4]), .Y(_09170_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32446_ ( .A(matmul_15_row_count_buf[3:0]), .Y(_09171_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32447_ ( .A(matmul_15_row_count_buf[15:12]), .Y(_09172_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32448_ ( .A(matmul_15_row_count_buf[11:8]), .Y(_09173_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32449_ ( .A({ _09178_, _09177_, _09176_, _09175_ }), .Y(_09174_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32450_ ( .A(matmul_15_col_count[24:21]), .Y(_09175_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32451_ ( .A(matmul_15_col_count[20:17]), .Y(_09176_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32452_ ( .A({ matmul_15_col_count[0], matmul_15_col_count[31:29] }), .Y(_09177_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32453_ ( .A(matmul_15_col_count[28:25]), .Y(_09178_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32454_ ( .A({ _09183_, _09182_, _09181_, _09180_ }), .Y(_09179_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32455_ ( .A(matmul_15_col_count[8:5]), .Y(_09180_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32456_ ( .A(matmul_15_col_count[4:1]), .Y(_09181_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32457_ ( .A(matmul_15_col_count[16:13]), .Y(_09182_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32458_ ( .A(matmul_15_col_count[12:9]), .Y(_09183_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32459_ ( .A({ _06990_, _stream_matmul_15_source_busy }), .Y(_05264_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32460_ ( .A({ _stream_matmul_15_source_8_idle, _stream_matmul_15_source_6_idle, _stream_matmul_15_source_20_idle, _09184_ }), .Y(_stream_matmul_15_done) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32461_ ( .A({ _stream_matmul_15_source_19_idle, _stream_matmul_15_source_14_idle, _stream_matmul_15_source_12_idle, _stream_matmul_15_source_10_idle }), .Y(_09184_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32462_ ( .A({ _tmp_1167, maxi_wready, maxi_wvalid }), .Y(_05265_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32463_ ( .A({ _tmp_958, maxi_wready, maxi_wvalid }), .Y(_05266_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32464_ ( .A({ _tmp_848, maxi_wready, maxi_wvalid }), .Y(_05267_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32465_ ( .A({ maxi_arvalid, maxi_arready }), .Y(_05269_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32466_ ( .A({ _07638_, _09185_, _05269_ }), .Y(_05268_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _32467_ ( .A({ _09186_, _tmp_14[4:3] }), .Y(_09185_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32468_ ( .A({ _09187_, _tmp_14[8:6] }), .Y(_09186_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32469_ ( .A({ _tmp_14[5], _tmp_14[2:0] }), .Y(_09187_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32470_ ( .A({ _09188_, _09185_ }), .Y(_05270_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32471_ ( .A({ maxi_rvalid, maxi_rready }), .Y(_09188_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32472_ ( .A({ _08260_, _09189_, _05273_ }), .Y(_05271_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32473_ ( .A({ _09190_, _tmp_847[0] }), .Y(_09189_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32474_ ( .A({ _09192_, _09191_ }), .Y(_09190_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32475_ ( .A(_tmp_847[8:5]), .Y(_09191_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32476_ ( .A(_tmp_847[4:1]), .Y(_09192_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32477_ ( .A({ maxi_awvalid, maxi_awready }), .Y(_05273_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32478_ ( .A({ _09202_, _09200_, _09193_, _05271_ }), .Y(_05272_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _32479_ ( .A({ _09199_, _09194_, _maxi_write_cur_size[1:0] }), .Y(_09193_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32480_ ( .A({ _09198_, _09197_, _09196_, _09195_ }), .Y(_09194_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32481_ ( .A(_maxi_write_cur_size[13:10]), .Y(_09195_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32482_ ( .A(_maxi_write_cur_size[9:6]), .Y(_09196_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32483_ ( .A(_maxi_write_cur_size[21:18]), .Y(_09197_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32484_ ( .A(_maxi_write_cur_size[17:14]), .Y(_09198_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32485_ ( .A(_maxi_write_cur_size[5:2]), .Y(_09199_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32486_ ( .A({ _09201_, _maxi_write_cur_size[32:30] }), .Y(_09200_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32487_ ( .A({ _maxi_write_cur_size[28:27], _maxi_write_cur_size[25], _maxi_write_cur_size[22] }), .Y(_09201_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32488_ ( .A({ _maxi_write_cur_size[29], _maxi_write_cur_size[26], _maxi_write_cur_size[24:23] }), .Y(_09202_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32489_ ( .A({ _dataflow_cat_valid_74, _09204_, _09203_ }), .Y(_05274_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _32490_ ( .A({ _08257_, _05276_, _09189_ }), .Y(_09203_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32491_ ( .A({ maxi_wvalid, maxi_wready }), .Y(_05276_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _32492_ ( .A({ _maxi_write_op_sel[0], _09205_, _09206_, _maxi_write_op_sel[1] }), .Y(_09204_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32493_ ( .A(_maxi_write_op_sel[7:4]), .Y(_09205_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32494_ ( .A(_maxi_write_op_sel[3:2]), .Y(_09206_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32495_ ( .A({ _09207_, _05274_ }), .Y(_05275_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32496_ ( .A({ _tmp_847[0], _09190_ }), .Y(_09207_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32497_ ( .A({ _dataflow_cat_valid_96, _09208_, _09203_ }), .Y(_05277_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _32498_ ( .A({ _09205_, _maxi_write_op_sel[1], _09206_, _maxi_write_op_sel[0] }), .Y(_09208_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32499_ ( .A({ _09207_, _05277_ }), .Y(_05278_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32500_ ( .A({ _dataflow_cat_valid_131, _09209_, _09203_ }), .Y(_05279_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32501_ ( .A({ _maxi_write_op_sel[0], _maxi_write_op_sel[1], _09206_, _09205_ }), .Y(_09209_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32502_ ( .A({ _09207_, _05279_ }), .Y(_05280_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32503_ ( .A({ _dataflow_slice_valid_4, _09210_ }), .Y(_05281_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32504_ ( .A({ _tmp_20, _09211_ }), .Y(_09210_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32505_ ( .A({ _09212_, _tmp_19[0], _tmp_19[33:32] }), .Y(_09211_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32506_ ( .A({ _09221_, _09220_, _09218_, _09213_ }), .Y(_09212_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32507_ ( .A({ _09217_, _09216_, _09215_, _09214_ }), .Y(_09213_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32508_ ( .A({ _tmp_19[24], _tmp_19[21], _tmp_19[19:18] }), .Y(_09214_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32509_ ( .A({ _tmp_19[31], _tmp_19[29:28], _tmp_19[25] }), .Y(_09215_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32510_ ( .A({ _tmp_19[7:6], _tmp_19[4], _tmp_19[1] }), .Y(_09216_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32511_ ( .A({ _tmp_19[16], _tmp_19[13], _tmp_19[11:10] }), .Y(_09217_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32512_ ( .A({ _09219_, _tmp_19[30], _tmp_19[27:26] }), .Y(_09218_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32513_ ( .A({ _tmp_19[23:22], _tmp_19[20], _tmp_19[17] }), .Y(_09219_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32514_ ( .A({ _tmp_19[8], _tmp_19[5], _tmp_19[3:2] }), .Y(_09220_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32515_ ( .A({ _tmp_19[15:14], _tmp_19[12], _tmp_19[9] }), .Y(_09221_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32516_ ( .A({ _wvalid_18, _05281_ }), .Y(_05282_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32517_ ( .A({ _dataflow_slice_valid_7, _09222_ }), .Y(_05284_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32518_ ( .A({ _tmp_22, _09223_ }), .Y(_09222_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32519_ ( .A({ _09224_, _tmp_21[0], _tmp_21[33:32] }), .Y(_09223_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32520_ ( .A({ _09233_, _09232_, _09230_, _09225_ }), .Y(_09224_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32521_ ( .A({ _09229_, _09228_, _09227_, _09226_ }), .Y(_09225_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32522_ ( .A({ _tmp_21[24], _tmp_21[21], _tmp_21[19:18] }), .Y(_09226_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32523_ ( .A({ _tmp_21[31], _tmp_21[29:28], _tmp_21[25] }), .Y(_09227_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32524_ ( .A({ _tmp_21[7:6], _tmp_21[4], _tmp_21[1] }), .Y(_09228_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32525_ ( .A({ _tmp_21[16], _tmp_21[13], _tmp_21[11:10] }), .Y(_09229_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32526_ ( .A({ _09231_, _tmp_21[30], _tmp_21[27:26] }), .Y(_09230_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32527_ ( .A({ _tmp_21[23:22], _tmp_21[20], _tmp_21[17] }), .Y(_09231_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32528_ ( .A({ _tmp_21[8], _tmp_21[5], _tmp_21[3:2] }), .Y(_09232_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32529_ ( .A({ _tmp_21[15:14], _tmp_21[12], _tmp_21[9] }), .Y(_09233_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32530_ ( .A({ _wvalid_18, _05284_ }), .Y(_05285_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32531_ ( .A({ _dataflow_slice_valid_10, _09234_ }), .Y(_05287_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32532_ ( .A({ _tmp_24, _09235_ }), .Y(_09234_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32533_ ( .A({ _09236_, _tmp_23[0], _tmp_23[33:32] }), .Y(_09235_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32534_ ( .A({ _09245_, _09244_, _09242_, _09237_ }), .Y(_09236_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32535_ ( .A({ _09241_, _09240_, _09239_, _09238_ }), .Y(_09237_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32536_ ( .A({ _tmp_23[24], _tmp_23[21], _tmp_23[19:18] }), .Y(_09238_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32537_ ( .A({ _tmp_23[31], _tmp_23[29:28], _tmp_23[25] }), .Y(_09239_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32538_ ( .A({ _tmp_23[7:6], _tmp_23[4], _tmp_23[1] }), .Y(_09240_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32539_ ( .A({ _tmp_23[16], _tmp_23[13], _tmp_23[11:10] }), .Y(_09241_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32540_ ( .A({ _09243_, _tmp_23[30], _tmp_23[27:26] }), .Y(_09242_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32541_ ( .A({ _tmp_23[23:22], _tmp_23[20], _tmp_23[17] }), .Y(_09243_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32542_ ( .A({ _tmp_23[8], _tmp_23[5], _tmp_23[3:2] }), .Y(_09244_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32543_ ( .A({ _tmp_23[15:14], _tmp_23[12], _tmp_23[9] }), .Y(_09245_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32544_ ( .A({ _wvalid_18, _05287_ }), .Y(_05288_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32545_ ( .A({ _dataflow_slice_valid_13, _09246_ }), .Y(_05290_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32546_ ( .A({ _tmp_26, _09247_ }), .Y(_09246_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32547_ ( .A({ _09248_, _tmp_25[0], _tmp_25[33:32] }), .Y(_09247_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32548_ ( .A({ _09257_, _09256_, _09254_, _09249_ }), .Y(_09248_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32549_ ( .A({ _09253_, _09252_, _09251_, _09250_ }), .Y(_09249_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32550_ ( .A({ _tmp_25[24], _tmp_25[21], _tmp_25[19:18] }), .Y(_09250_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32551_ ( .A({ _tmp_25[31], _tmp_25[29:28], _tmp_25[25] }), .Y(_09251_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32552_ ( .A({ _tmp_25[7:6], _tmp_25[4], _tmp_25[1] }), .Y(_09252_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32553_ ( .A({ _tmp_25[16], _tmp_25[13], _tmp_25[11:10] }), .Y(_09253_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32554_ ( .A({ _09255_, _tmp_25[30], _tmp_25[27:26] }), .Y(_09254_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32555_ ( .A({ _tmp_25[23:22], _tmp_25[20], _tmp_25[17] }), .Y(_09255_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32556_ ( .A({ _tmp_25[8], _tmp_25[5], _tmp_25[3:2] }), .Y(_09256_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32557_ ( .A({ _tmp_25[15:14], _tmp_25[12], _tmp_25[9] }), .Y(_09257_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32558_ ( .A({ _wvalid_18, _05290_ }), .Y(_05291_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _32559_ ( .A({ _dataflow_slice_valid_17, _tmp_34, _09258_ }), .Y(_05293_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32560_ ( .A({ _09259_, _tmp_33[0], _tmp_33[33:32] }), .Y(_09258_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32561_ ( .A({ _09268_, _09267_, _09265_, _09260_ }), .Y(_09259_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32562_ ( .A({ _09264_, _09263_, _09262_, _09261_ }), .Y(_09260_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32563_ ( .A({ _tmp_33[24], _tmp_33[21], _tmp_33[19:18] }), .Y(_09261_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32564_ ( .A({ _tmp_33[31], _tmp_33[29:28], _tmp_33[25] }), .Y(_09262_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32565_ ( .A({ _tmp_33[7:6], _tmp_33[4], _tmp_33[1] }), .Y(_09263_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32566_ ( .A({ _tmp_33[16], _tmp_33[13], _tmp_33[11:10] }), .Y(_09264_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32567_ ( .A({ _09266_, _tmp_33[30], _tmp_33[27:26] }), .Y(_09265_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32568_ ( .A({ _tmp_33[23:22], _tmp_33[20], _tmp_33[17] }), .Y(_09266_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32569_ ( .A({ _tmp_33[8], _tmp_33[5], _tmp_33[3:2] }), .Y(_09267_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32570_ ( .A({ _tmp_33[15:14], _tmp_33[12], _tmp_33[9] }), .Y(_09268_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32571_ ( .A({ _wvalid_31, _05293_ }), .Y(_05294_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _32572_ ( .A({ _dataflow_slice_valid_20, _tmp_65, _09269_ }), .Y(_05296_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32573_ ( .A({ _09270_, _tmp_64[0], _tmp_64[33:32] }), .Y(_09269_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32574_ ( .A({ _09279_, _09278_, _09276_, _09271_ }), .Y(_09270_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32575_ ( .A({ _09275_, _09274_, _09273_, _09272_ }), .Y(_09271_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32576_ ( .A({ _tmp_64[24], _tmp_64[21], _tmp_64[19:18] }), .Y(_09272_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32577_ ( .A({ _tmp_64[31], _tmp_64[29:28], _tmp_64[25] }), .Y(_09273_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32578_ ( .A({ _tmp_64[7:6], _tmp_64[4], _tmp_64[1] }), .Y(_09274_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32579_ ( .A({ _tmp_64[16], _tmp_64[13], _tmp_64[11:10] }), .Y(_09275_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32580_ ( .A({ _09277_, _tmp_64[30], _tmp_64[27:26] }), .Y(_09276_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32581_ ( .A({ _tmp_64[23:22], _tmp_64[20], _tmp_64[17] }), .Y(_09277_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32582_ ( .A({ _tmp_64[8], _tmp_64[5], _tmp_64[3:2] }), .Y(_09278_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32583_ ( .A({ _tmp_64[15:14], _tmp_64[12], _tmp_64[9] }), .Y(_09279_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32584_ ( .A({ _wvalid_31, _05296_ }), .Y(_05297_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _32585_ ( .A({ _dataflow_slice_valid_23, _tmp_96, _09280_ }), .Y(_05299_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32586_ ( .A({ _09281_, _tmp_95[0], _tmp_95[33:32] }), .Y(_09280_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32587_ ( .A({ _09290_, _09289_, _09287_, _09282_ }), .Y(_09281_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32588_ ( .A({ _09286_, _09285_, _09284_, _09283_ }), .Y(_09282_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32589_ ( .A({ _tmp_95[24], _tmp_95[21], _tmp_95[19:18] }), .Y(_09283_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32590_ ( .A({ _tmp_95[31], _tmp_95[29:28], _tmp_95[25] }), .Y(_09284_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32591_ ( .A({ _tmp_95[7:6], _tmp_95[4], _tmp_95[1] }), .Y(_09285_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32592_ ( .A({ _tmp_95[16], _tmp_95[13], _tmp_95[11:10] }), .Y(_09286_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32593_ ( .A({ _09288_, _tmp_95[30], _tmp_95[27:26] }), .Y(_09287_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32594_ ( .A({ _tmp_95[23:22], _tmp_95[20], _tmp_95[17] }), .Y(_09288_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32595_ ( .A({ _tmp_95[8], _tmp_95[5], _tmp_95[3:2] }), .Y(_09289_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32596_ ( .A({ _tmp_95[15:14], _tmp_95[12], _tmp_95[9] }), .Y(_09290_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32597_ ( .A({ _wvalid_31, _05299_ }), .Y(_05300_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _32598_ ( .A({ _dataflow_slice_valid_26, _tmp_127, _09291_ }), .Y(_05302_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32599_ ( .A({ _09292_, _tmp_126[0], _tmp_126[33:32] }), .Y(_09291_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32600_ ( .A({ _09301_, _09300_, _09298_, _09293_ }), .Y(_09292_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32601_ ( .A({ _09297_, _09296_, _09295_, _09294_ }), .Y(_09293_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32602_ ( .A({ _tmp_126[24], _tmp_126[21], _tmp_126[19:18] }), .Y(_09294_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32603_ ( .A({ _tmp_126[31], _tmp_126[29:28], _tmp_126[25] }), .Y(_09295_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32604_ ( .A({ _tmp_126[7:6], _tmp_126[4], _tmp_126[1] }), .Y(_09296_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32605_ ( .A({ _tmp_126[16], _tmp_126[13], _tmp_126[11:10] }), .Y(_09297_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32606_ ( .A({ _09299_, _tmp_126[30], _tmp_126[27:26] }), .Y(_09298_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32607_ ( .A({ _tmp_126[23:22], _tmp_126[20], _tmp_126[17] }), .Y(_09299_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32608_ ( .A({ _tmp_126[8], _tmp_126[5], _tmp_126[3:2] }), .Y(_09300_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32609_ ( .A({ _tmp_126[15:14], _tmp_126[12], _tmp_126[9] }), .Y(_09301_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32610_ ( .A({ _wvalid_31, _05302_ }), .Y(_05303_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32611_ ( .A({ _dataflow_slice_valid_30, _09302_ }), .Y(_05305_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32612_ ( .A({ _tmp_163, _09303_ }), .Y(_09302_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32613_ ( .A({ _09304_, _tmp_162[0], _tmp_162[33:32] }), .Y(_09303_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32614_ ( .A({ _09313_, _09312_, _09310_, _09305_ }), .Y(_09304_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32615_ ( .A({ _09309_, _09308_, _09307_, _09306_ }), .Y(_09305_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32616_ ( .A({ _tmp_162[24], _tmp_162[21], _tmp_162[19:18] }), .Y(_09306_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32617_ ( .A({ _tmp_162[31], _tmp_162[29:28], _tmp_162[25] }), .Y(_09307_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32618_ ( .A({ _tmp_162[7:6], _tmp_162[4], _tmp_162[1] }), .Y(_09308_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32619_ ( .A({ _tmp_162[16], _tmp_162[13], _tmp_162[11:10] }), .Y(_09309_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32620_ ( .A({ _09311_, _tmp_162[30], _tmp_162[27:26] }), .Y(_09310_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32621_ ( .A({ _tmp_162[23:22], _tmp_162[20], _tmp_162[17] }), .Y(_09311_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32622_ ( .A({ _tmp_162[8], _tmp_162[5], _tmp_162[3:2] }), .Y(_09312_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32623_ ( .A({ _tmp_162[15:14], _tmp_162[12], _tmp_162[9] }), .Y(_09313_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32624_ ( .A({ _wvalid_160, _05305_ }), .Y(_05306_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32625_ ( .A({ _dataflow_slice_valid_33, _09314_ }), .Y(_05308_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32626_ ( .A({ _tmp_176, _09315_ }), .Y(_09314_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32627_ ( .A({ _09316_, _tmp_175[0], _tmp_175[33:32] }), .Y(_09315_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32628_ ( .A({ _09325_, _09324_, _09322_, _09317_ }), .Y(_09316_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32629_ ( .A({ _09321_, _09320_, _09319_, _09318_ }), .Y(_09317_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32630_ ( .A({ _tmp_175[24], _tmp_175[21], _tmp_175[19:18] }), .Y(_09318_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32631_ ( .A({ _tmp_175[31], _tmp_175[29:28], _tmp_175[25] }), .Y(_09319_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32632_ ( .A({ _tmp_175[7:6], _tmp_175[4], _tmp_175[1] }), .Y(_09320_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32633_ ( .A({ _tmp_175[16], _tmp_175[13], _tmp_175[11:10] }), .Y(_09321_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32634_ ( .A({ _09323_, _tmp_175[30], _tmp_175[27:26] }), .Y(_09322_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32635_ ( .A({ _tmp_175[23:22], _tmp_175[20], _tmp_175[17] }), .Y(_09323_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32636_ ( .A({ _tmp_175[8], _tmp_175[5], _tmp_175[3:2] }), .Y(_09324_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32637_ ( .A({ _tmp_175[15:14], _tmp_175[12], _tmp_175[9] }), .Y(_09325_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32638_ ( .A({ _wvalid_160, _05308_ }), .Y(_05309_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32639_ ( .A({ _dataflow_slice_valid_36, _09326_ }), .Y(_05311_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32640_ ( .A({ _tmp_189, _09327_ }), .Y(_09326_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32641_ ( .A({ _09328_, _tmp_188[0], _tmp_188[33:32] }), .Y(_09327_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32642_ ( .A({ _09337_, _09336_, _09334_, _09329_ }), .Y(_09328_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32643_ ( .A({ _09333_, _09332_, _09331_, _09330_ }), .Y(_09329_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32644_ ( .A({ _tmp_188[24], _tmp_188[21], _tmp_188[19:18] }), .Y(_09330_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32645_ ( .A({ _tmp_188[31], _tmp_188[29:28], _tmp_188[25] }), .Y(_09331_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32646_ ( .A({ _tmp_188[7:6], _tmp_188[4], _tmp_188[1] }), .Y(_09332_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32647_ ( .A({ _tmp_188[16], _tmp_188[13], _tmp_188[11:10] }), .Y(_09333_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32648_ ( .A({ _09335_, _tmp_188[30], _tmp_188[27:26] }), .Y(_09334_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32649_ ( .A({ _tmp_188[23:22], _tmp_188[20], _tmp_188[17] }), .Y(_09335_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32650_ ( .A({ _tmp_188[8], _tmp_188[5], _tmp_188[3:2] }), .Y(_09336_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32651_ ( .A({ _tmp_188[15:14], _tmp_188[12], _tmp_188[9] }), .Y(_09337_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32652_ ( .A({ _wvalid_160, _05311_ }), .Y(_05312_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32653_ ( .A({ _dataflow_slice_valid_39, _09338_ }), .Y(_05314_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32654_ ( .A({ _tmp_202, _09339_ }), .Y(_09338_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32655_ ( .A({ _09340_, _tmp_201[0], _tmp_201[33:32] }), .Y(_09339_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32656_ ( .A({ _09349_, _09348_, _09346_, _09341_ }), .Y(_09340_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32657_ ( .A({ _09345_, _09344_, _09343_, _09342_ }), .Y(_09341_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32658_ ( .A({ _tmp_201[24], _tmp_201[21], _tmp_201[19:18] }), .Y(_09342_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32659_ ( .A({ _tmp_201[31], _tmp_201[29:28], _tmp_201[25] }), .Y(_09343_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32660_ ( .A({ _tmp_201[7:6], _tmp_201[4], _tmp_201[1] }), .Y(_09344_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32661_ ( .A({ _tmp_201[16], _tmp_201[13], _tmp_201[11:10] }), .Y(_09345_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32662_ ( .A({ _09347_, _tmp_201[30], _tmp_201[27:26] }), .Y(_09346_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32663_ ( .A({ _tmp_201[23:22], _tmp_201[20], _tmp_201[17] }), .Y(_09347_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32664_ ( .A({ _tmp_201[8], _tmp_201[5], _tmp_201[3:2] }), .Y(_09348_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32665_ ( .A({ _tmp_201[15:14], _tmp_201[12], _tmp_201[9] }), .Y(_09349_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32666_ ( .A({ _wvalid_160, _05314_ }), .Y(_05315_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32667_ ( .A({ _dataflow_slice_valid_43, _09350_ }), .Y(_05317_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32668_ ( .A({ _tmp_220, _09351_ }), .Y(_09350_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32669_ ( .A({ _09352_, _tmp_219[0], _tmp_219[33:32] }), .Y(_09351_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32670_ ( .A({ _09361_, _09360_, _09358_, _09353_ }), .Y(_09352_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32671_ ( .A({ _09357_, _09356_, _09355_, _09354_ }), .Y(_09353_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32672_ ( .A({ _tmp_219[24], _tmp_219[21], _tmp_219[19:18] }), .Y(_09354_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32673_ ( .A({ _tmp_219[31], _tmp_219[29:28], _tmp_219[25] }), .Y(_09355_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32674_ ( .A({ _tmp_219[7:6], _tmp_219[4], _tmp_219[1] }), .Y(_09356_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32675_ ( .A({ _tmp_219[16], _tmp_219[13], _tmp_219[11:10] }), .Y(_09357_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32676_ ( .A({ _09359_, _tmp_219[30], _tmp_219[27:26] }), .Y(_09358_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32677_ ( .A({ _tmp_219[23:22], _tmp_219[20], _tmp_219[17] }), .Y(_09359_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32678_ ( .A({ _tmp_219[8], _tmp_219[5], _tmp_219[3:2] }), .Y(_09360_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32679_ ( .A({ _tmp_219[15:14], _tmp_219[12], _tmp_219[9] }), .Y(_09361_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32680_ ( .A({ _wvalid_217, _05317_ }), .Y(_05318_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32681_ ( .A({ _dataflow_slice_valid_46, _09362_ }), .Y(_05320_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32682_ ( .A({ _tmp_233, _09363_ }), .Y(_09362_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32683_ ( .A({ _09364_, _tmp_232[0], _tmp_232[33:32] }), .Y(_09363_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32684_ ( .A({ _09373_, _09372_, _09370_, _09365_ }), .Y(_09364_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32685_ ( .A({ _09369_, _09368_, _09367_, _09366_ }), .Y(_09365_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32686_ ( .A({ _tmp_232[24], _tmp_232[21], _tmp_232[19:18] }), .Y(_09366_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32687_ ( .A({ _tmp_232[31], _tmp_232[29:28], _tmp_232[25] }), .Y(_09367_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32688_ ( .A({ _tmp_232[7:6], _tmp_232[4], _tmp_232[1] }), .Y(_09368_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32689_ ( .A({ _tmp_232[16], _tmp_232[13], _tmp_232[11:10] }), .Y(_09369_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32690_ ( .A({ _09371_, _tmp_232[30], _tmp_232[27:26] }), .Y(_09370_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32691_ ( .A({ _tmp_232[23:22], _tmp_232[20], _tmp_232[17] }), .Y(_09371_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32692_ ( .A({ _tmp_232[8], _tmp_232[5], _tmp_232[3:2] }), .Y(_09372_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32693_ ( .A({ _tmp_232[15:14], _tmp_232[12], _tmp_232[9] }), .Y(_09373_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32694_ ( .A({ _wvalid_217, _05320_ }), .Y(_05321_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32695_ ( .A({ _dataflow_slice_valid_49, _09374_ }), .Y(_05323_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32696_ ( .A({ _tmp_246, _09375_ }), .Y(_09374_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32697_ ( .A({ _09376_, _tmp_245[0], _tmp_245[33:32] }), .Y(_09375_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32698_ ( .A({ _09385_, _09384_, _09382_, _09377_ }), .Y(_09376_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32699_ ( .A({ _09381_, _09380_, _09379_, _09378_ }), .Y(_09377_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32700_ ( .A({ _tmp_245[24], _tmp_245[21], _tmp_245[19:18] }), .Y(_09378_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32701_ ( .A({ _tmp_245[31], _tmp_245[29:28], _tmp_245[25] }), .Y(_09379_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32702_ ( .A({ _tmp_245[7:6], _tmp_245[4], _tmp_245[1] }), .Y(_09380_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32703_ ( .A({ _tmp_245[16], _tmp_245[13], _tmp_245[11:10] }), .Y(_09381_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32704_ ( .A({ _09383_, _tmp_245[30], _tmp_245[27:26] }), .Y(_09382_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32705_ ( .A({ _tmp_245[23:22], _tmp_245[20], _tmp_245[17] }), .Y(_09383_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32706_ ( .A({ _tmp_245[8], _tmp_245[5], _tmp_245[3:2] }), .Y(_09384_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32707_ ( .A({ _tmp_245[15:14], _tmp_245[12], _tmp_245[9] }), .Y(_09385_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32708_ ( .A({ _wvalid_217, _05323_ }), .Y(_05324_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32709_ ( .A({ _dataflow_slice_valid_52, _09386_ }), .Y(_05326_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32710_ ( .A({ _tmp_259, _09387_ }), .Y(_09386_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32711_ ( .A({ _09388_, _tmp_258[0], _tmp_258[33:32] }), .Y(_09387_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32712_ ( .A({ _09397_, _09396_, _09394_, _09389_ }), .Y(_09388_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32713_ ( .A({ _09393_, _09392_, _09391_, _09390_ }), .Y(_09389_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32714_ ( .A({ _tmp_258[24], _tmp_258[21], _tmp_258[19:18] }), .Y(_09390_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32715_ ( .A({ _tmp_258[31], _tmp_258[29:28], _tmp_258[25] }), .Y(_09391_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32716_ ( .A({ _tmp_258[7:6], _tmp_258[4], _tmp_258[1] }), .Y(_09392_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32717_ ( .A({ _tmp_258[16], _tmp_258[13], _tmp_258[11:10] }), .Y(_09393_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32718_ ( .A({ _09395_, _tmp_258[30], _tmp_258[27:26] }), .Y(_09394_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32719_ ( .A({ _tmp_258[23:22], _tmp_258[20], _tmp_258[17] }), .Y(_09395_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32720_ ( .A({ _tmp_258[8], _tmp_258[5], _tmp_258[3:2] }), .Y(_09396_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32721_ ( .A({ _tmp_258[15:14], _tmp_258[12], _tmp_258[9] }), .Y(_09397_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32722_ ( .A({ _wvalid_217, _05326_ }), .Y(_05327_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32723_ ( .A({ _dataflow_slice_valid_56, _09398_ }), .Y(_05329_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32724_ ( .A({ _tmp_277, _09399_ }), .Y(_09398_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32725_ ( .A({ _09400_, _tmp_276[0], _tmp_276[33:32] }), .Y(_09399_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32726_ ( .A({ _09409_, _09408_, _09406_, _09401_ }), .Y(_09400_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32727_ ( .A({ _09405_, _09404_, _09403_, _09402_ }), .Y(_09401_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32728_ ( .A({ _tmp_276[24], _tmp_276[21], _tmp_276[19:18] }), .Y(_09402_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32729_ ( .A({ _tmp_276[31], _tmp_276[29:28], _tmp_276[25] }), .Y(_09403_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32730_ ( .A({ _tmp_276[7:6], _tmp_276[4], _tmp_276[1] }), .Y(_09404_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32731_ ( .A({ _tmp_276[16], _tmp_276[13], _tmp_276[11:10] }), .Y(_09405_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32732_ ( .A({ _09407_, _tmp_276[30], _tmp_276[27:26] }), .Y(_09406_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32733_ ( .A({ _tmp_276[23:22], _tmp_276[20], _tmp_276[17] }), .Y(_09407_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32734_ ( .A({ _tmp_276[8], _tmp_276[5], _tmp_276[3:2] }), .Y(_09408_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32735_ ( .A({ _tmp_276[15:14], _tmp_276[12], _tmp_276[9] }), .Y(_09409_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32736_ ( .A({ _wvalid_274, _05329_ }), .Y(_05330_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32737_ ( .A({ _dataflow_slice_valid_59, _09410_ }), .Y(_05332_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32738_ ( .A({ _tmp_290, _09411_ }), .Y(_09410_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32739_ ( .A({ _09412_, _tmp_289[0], _tmp_289[33:32] }), .Y(_09411_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32740_ ( .A({ _09421_, _09420_, _09418_, _09413_ }), .Y(_09412_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32741_ ( .A({ _09417_, _09416_, _09415_, _09414_ }), .Y(_09413_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32742_ ( .A({ _tmp_289[24], _tmp_289[21], _tmp_289[19:18] }), .Y(_09414_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32743_ ( .A({ _tmp_289[31], _tmp_289[29:28], _tmp_289[25] }), .Y(_09415_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32744_ ( .A({ _tmp_289[7:6], _tmp_289[4], _tmp_289[1] }), .Y(_09416_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32745_ ( .A({ _tmp_289[16], _tmp_289[13], _tmp_289[11:10] }), .Y(_09417_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32746_ ( .A({ _09419_, _tmp_289[30], _tmp_289[27:26] }), .Y(_09418_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32747_ ( .A({ _tmp_289[23:22], _tmp_289[20], _tmp_289[17] }), .Y(_09419_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32748_ ( .A({ _tmp_289[8], _tmp_289[5], _tmp_289[3:2] }), .Y(_09420_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32749_ ( .A({ _tmp_289[15:14], _tmp_289[12], _tmp_289[9] }), .Y(_09421_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32750_ ( .A({ _wvalid_274, _05332_ }), .Y(_05333_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32751_ ( .A({ _dataflow_slice_valid_62, _09422_ }), .Y(_05335_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32752_ ( .A({ _tmp_303, _09423_ }), .Y(_09422_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32753_ ( .A({ _09424_, _tmp_302[0], _tmp_302[33:32] }), .Y(_09423_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32754_ ( .A({ _09433_, _09432_, _09430_, _09425_ }), .Y(_09424_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32755_ ( .A({ _09429_, _09428_, _09427_, _09426_ }), .Y(_09425_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32756_ ( .A({ _tmp_302[24], _tmp_302[21], _tmp_302[19:18] }), .Y(_09426_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32757_ ( .A({ _tmp_302[31], _tmp_302[29:28], _tmp_302[25] }), .Y(_09427_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32758_ ( .A({ _tmp_302[7:6], _tmp_302[4], _tmp_302[1] }), .Y(_09428_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32759_ ( .A({ _tmp_302[16], _tmp_302[13], _tmp_302[11:10] }), .Y(_09429_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32760_ ( .A({ _09431_, _tmp_302[30], _tmp_302[27:26] }), .Y(_09430_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32761_ ( .A({ _tmp_302[23:22], _tmp_302[20], _tmp_302[17] }), .Y(_09431_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32762_ ( .A({ _tmp_302[8], _tmp_302[5], _tmp_302[3:2] }), .Y(_09432_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32763_ ( .A({ _tmp_302[15:14], _tmp_302[12], _tmp_302[9] }), .Y(_09433_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32764_ ( .A({ _wvalid_274, _05335_ }), .Y(_05336_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32765_ ( .A({ _dataflow_slice_valid_65, _09434_ }), .Y(_05338_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32766_ ( .A({ _tmp_316, _09435_ }), .Y(_09434_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32767_ ( .A({ _09436_, _tmp_315[0], _tmp_315[33:32] }), .Y(_09435_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32768_ ( .A({ _09445_, _09444_, _09442_, _09437_ }), .Y(_09436_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32769_ ( .A({ _09441_, _09440_, _09439_, _09438_ }), .Y(_09437_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32770_ ( .A({ _tmp_315[24], _tmp_315[21], _tmp_315[19:18] }), .Y(_09438_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32771_ ( .A({ _tmp_315[31], _tmp_315[29:28], _tmp_315[25] }), .Y(_09439_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32772_ ( .A({ _tmp_315[7:6], _tmp_315[4], _tmp_315[1] }), .Y(_09440_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32773_ ( .A({ _tmp_315[16], _tmp_315[13], _tmp_315[11:10] }), .Y(_09441_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32774_ ( .A({ _09443_, _tmp_315[30], _tmp_315[27:26] }), .Y(_09442_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32775_ ( .A({ _tmp_315[23:22], _tmp_315[20], _tmp_315[17] }), .Y(_09443_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32776_ ( .A({ _tmp_315[8], _tmp_315[5], _tmp_315[3:2] }), .Y(_09444_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32777_ ( .A({ _tmp_315[15:14], _tmp_315[12], _tmp_315[9] }), .Y(_09445_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32778_ ( .A({ _wvalid_274, _05338_ }), .Y(_05339_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32779_ ( .A({ _dataflow_slice_valid_78, _09446_ }), .Y(_05341_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32780_ ( .A({ _tmp_854, _09447_ }), .Y(_09446_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32781_ ( .A({ _09448_, _tmp_853[0], _tmp_853[33:32] }), .Y(_09447_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32782_ ( .A({ _09457_, _09456_, _09454_, _09449_ }), .Y(_09448_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32783_ ( .A({ _09453_, _09452_, _09451_, _09450_ }), .Y(_09449_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32784_ ( .A({ _tmp_853[24], _tmp_853[21], _tmp_853[19:18] }), .Y(_09450_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32785_ ( .A({ _tmp_853[31], _tmp_853[29:28], _tmp_853[25] }), .Y(_09451_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32786_ ( .A({ _tmp_853[7:6], _tmp_853[4], _tmp_853[1] }), .Y(_09452_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32787_ ( .A({ _tmp_853[16], _tmp_853[13], _tmp_853[11:10] }), .Y(_09453_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32788_ ( .A({ _09455_, _tmp_853[30], _tmp_853[27:26] }), .Y(_09454_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32789_ ( .A({ _tmp_853[23:22], _tmp_853[20], _tmp_853[17] }), .Y(_09455_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32790_ ( .A({ _tmp_853[8], _tmp_853[5], _tmp_853[3:2] }), .Y(_09456_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32791_ ( .A({ _tmp_853[15:14], _tmp_853[12], _tmp_853[9] }), .Y(_09457_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32792_ ( .A({ _wvalid_852, _05341_ }), .Y(_05342_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32793_ ( .A({ _dataflow_slice_valid_81, _09458_ }), .Y(_05344_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32794_ ( .A({ _tmp_856, _09459_ }), .Y(_09458_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32795_ ( .A({ _09460_, _tmp_855[0], _tmp_855[33:32] }), .Y(_09459_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32796_ ( .A({ _09469_, _09468_, _09466_, _09461_ }), .Y(_09460_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32797_ ( .A({ _09465_, _09464_, _09463_, _09462_ }), .Y(_09461_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32798_ ( .A({ _tmp_855[24], _tmp_855[21], _tmp_855[19:18] }), .Y(_09462_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32799_ ( .A({ _tmp_855[31], _tmp_855[29:28], _tmp_855[25] }), .Y(_09463_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32800_ ( .A({ _tmp_855[7:6], _tmp_855[4], _tmp_855[1] }), .Y(_09464_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32801_ ( .A({ _tmp_855[16], _tmp_855[13], _tmp_855[11:10] }), .Y(_09465_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32802_ ( .A({ _09467_, _tmp_855[30], _tmp_855[27:26] }), .Y(_09466_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32803_ ( .A({ _tmp_855[23:22], _tmp_855[20], _tmp_855[17] }), .Y(_09467_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32804_ ( .A({ _tmp_855[8], _tmp_855[5], _tmp_855[3:2] }), .Y(_09468_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32805_ ( .A({ _tmp_855[15:14], _tmp_855[12], _tmp_855[9] }), .Y(_09469_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32806_ ( .A({ _wvalid_852, _05344_ }), .Y(_05345_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32807_ ( .A({ _dataflow_slice_valid_84, _09470_ }), .Y(_05347_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32808_ ( .A({ _tmp_858, _09471_ }), .Y(_09470_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32809_ ( .A({ _09472_, _tmp_857[0], _tmp_857[33:32] }), .Y(_09471_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32810_ ( .A({ _09481_, _09480_, _09478_, _09473_ }), .Y(_09472_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32811_ ( .A({ _09477_, _09476_, _09475_, _09474_ }), .Y(_09473_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32812_ ( .A({ _tmp_857[24], _tmp_857[21], _tmp_857[19:18] }), .Y(_09474_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32813_ ( .A({ _tmp_857[31], _tmp_857[29:28], _tmp_857[25] }), .Y(_09475_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32814_ ( .A({ _tmp_857[7:6], _tmp_857[4], _tmp_857[1] }), .Y(_09476_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32815_ ( .A({ _tmp_857[16], _tmp_857[13], _tmp_857[11:10] }), .Y(_09477_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32816_ ( .A({ _09479_, _tmp_857[30], _tmp_857[27:26] }), .Y(_09478_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32817_ ( .A({ _tmp_857[23:22], _tmp_857[20], _tmp_857[17] }), .Y(_09479_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32818_ ( .A({ _tmp_857[8], _tmp_857[5], _tmp_857[3:2] }), .Y(_09480_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32819_ ( .A({ _tmp_857[15:14], _tmp_857[12], _tmp_857[9] }), .Y(_09481_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32820_ ( .A({ _wvalid_852, _05347_ }), .Y(_05348_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32821_ ( .A({ _dataflow_slice_valid_87, _09482_ }), .Y(_05350_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32822_ ( .A({ _tmp_860, _09483_ }), .Y(_09482_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32823_ ( .A({ _09484_, _tmp_859[0], _tmp_859[33:32] }), .Y(_09483_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32824_ ( .A({ _09493_, _09492_, _09490_, _09485_ }), .Y(_09484_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32825_ ( .A({ _09489_, _09488_, _09487_, _09486_ }), .Y(_09485_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32826_ ( .A({ _tmp_859[24], _tmp_859[21], _tmp_859[19:18] }), .Y(_09486_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32827_ ( .A({ _tmp_859[31], _tmp_859[29:28], _tmp_859[25] }), .Y(_09487_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32828_ ( .A({ _tmp_859[7:6], _tmp_859[4], _tmp_859[1] }), .Y(_09488_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32829_ ( .A({ _tmp_859[16], _tmp_859[13], _tmp_859[11:10] }), .Y(_09489_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32830_ ( .A({ _09491_, _tmp_859[30], _tmp_859[27:26] }), .Y(_09490_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32831_ ( .A({ _tmp_859[23:22], _tmp_859[20], _tmp_859[17] }), .Y(_09491_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32832_ ( .A({ _tmp_859[8], _tmp_859[5], _tmp_859[3:2] }), .Y(_09492_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32833_ ( .A({ _tmp_859[15:14], _tmp_859[12], _tmp_859[9] }), .Y(_09493_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32834_ ( .A({ _wvalid_852, _05350_ }), .Y(_05351_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32835_ ( .A({ _dataflow_slice_valid_100, _09494_ }), .Y(_05353_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32836_ ( .A({ _tmp_965, _09495_ }), .Y(_09494_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32837_ ( .A({ _09496_, _tmp_964[0], _tmp_964[33:32] }), .Y(_09495_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32838_ ( .A({ _09505_, _09504_, _09502_, _09497_ }), .Y(_09496_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32839_ ( .A({ _09501_, _09500_, _09499_, _09498_ }), .Y(_09497_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32840_ ( .A({ _tmp_964[24], _tmp_964[21], _tmp_964[19:18] }), .Y(_09498_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32841_ ( .A({ _tmp_964[31], _tmp_964[29:28], _tmp_964[25] }), .Y(_09499_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32842_ ( .A({ _tmp_964[7:6], _tmp_964[4], _tmp_964[1] }), .Y(_09500_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32843_ ( .A({ _tmp_964[16], _tmp_964[13], _tmp_964[11:10] }), .Y(_09501_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32844_ ( .A({ _09503_, _tmp_964[30], _tmp_964[27:26] }), .Y(_09502_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32845_ ( .A({ _tmp_964[23:22], _tmp_964[20], _tmp_964[17] }), .Y(_09503_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32846_ ( .A({ _tmp_964[8], _tmp_964[5], _tmp_964[3:2] }), .Y(_09504_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32847_ ( .A({ _tmp_964[15:14], _tmp_964[12], _tmp_964[9] }), .Y(_09505_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32848_ ( .A({ _wvalid_963, _05353_ }), .Y(_05354_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32849_ ( .A({ _dataflow_slice_valid_103, _09506_ }), .Y(_05356_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32850_ ( .A({ _tmp_967, _09507_ }), .Y(_09506_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32851_ ( .A({ _09508_, _tmp_966[0], _tmp_966[33:32] }), .Y(_09507_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32852_ ( .A({ _09517_, _09516_, _09514_, _09509_ }), .Y(_09508_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32853_ ( .A({ _09513_, _09512_, _09511_, _09510_ }), .Y(_09509_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32854_ ( .A({ _tmp_966[24], _tmp_966[21], _tmp_966[19:18] }), .Y(_09510_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32855_ ( .A({ _tmp_966[31], _tmp_966[29:28], _tmp_966[25] }), .Y(_09511_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32856_ ( .A({ _tmp_966[7:6], _tmp_966[4], _tmp_966[1] }), .Y(_09512_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32857_ ( .A({ _tmp_966[16], _tmp_966[13], _tmp_966[11:10] }), .Y(_09513_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32858_ ( .A({ _09515_, _tmp_966[30], _tmp_966[27:26] }), .Y(_09514_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32859_ ( .A({ _tmp_966[23:22], _tmp_966[20], _tmp_966[17] }), .Y(_09515_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32860_ ( .A({ _tmp_966[8], _tmp_966[5], _tmp_966[3:2] }), .Y(_09516_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32861_ ( .A({ _tmp_966[15:14], _tmp_966[12], _tmp_966[9] }), .Y(_09517_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32862_ ( .A({ _wvalid_963, _05356_ }), .Y(_05357_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32863_ ( .A({ _dataflow_slice_valid_106, _09518_ }), .Y(_05359_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32864_ ( .A({ _tmp_969, _09519_ }), .Y(_09518_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32865_ ( .A({ _09520_, _tmp_968[0], _tmp_968[33:32] }), .Y(_09519_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32866_ ( .A({ _09529_, _09528_, _09526_, _09521_ }), .Y(_09520_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32867_ ( .A({ _09525_, _09524_, _09523_, _09522_ }), .Y(_09521_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32868_ ( .A({ _tmp_968[24], _tmp_968[21], _tmp_968[19:18] }), .Y(_09522_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32869_ ( .A({ _tmp_968[31], _tmp_968[29:28], _tmp_968[25] }), .Y(_09523_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32870_ ( .A({ _tmp_968[7:6], _tmp_968[4], _tmp_968[1] }), .Y(_09524_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32871_ ( .A({ _tmp_968[16], _tmp_968[13], _tmp_968[11:10] }), .Y(_09525_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32872_ ( .A({ _09527_, _tmp_968[30], _tmp_968[27:26] }), .Y(_09526_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32873_ ( .A({ _tmp_968[23:22], _tmp_968[20], _tmp_968[17] }), .Y(_09527_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32874_ ( .A({ _tmp_968[8], _tmp_968[5], _tmp_968[3:2] }), .Y(_09528_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32875_ ( .A({ _tmp_968[15:14], _tmp_968[12], _tmp_968[9] }), .Y(_09529_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32876_ ( .A({ _wvalid_963, _05359_ }), .Y(_05360_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32877_ ( .A({ _dataflow_slice_valid_109, _09530_ }), .Y(_05362_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32878_ ( .A({ _tmp_971, _09531_ }), .Y(_09530_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32879_ ( .A({ _09532_, _tmp_970[0], _tmp_970[33:32] }), .Y(_09531_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32880_ ( .A({ _09541_, _09540_, _09538_, _09533_ }), .Y(_09532_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32881_ ( .A({ _09537_, _09536_, _09535_, _09534_ }), .Y(_09533_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32882_ ( .A({ _tmp_970[24], _tmp_970[21], _tmp_970[19:18] }), .Y(_09534_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32883_ ( .A({ _tmp_970[31], _tmp_970[29:28], _tmp_970[25] }), .Y(_09535_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32884_ ( .A({ _tmp_970[7:6], _tmp_970[4], _tmp_970[1] }), .Y(_09536_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32885_ ( .A({ _tmp_970[16], _tmp_970[13], _tmp_970[11:10] }), .Y(_09537_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32886_ ( .A({ _09539_, _tmp_970[30], _tmp_970[27:26] }), .Y(_09538_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32887_ ( .A({ _tmp_970[23:22], _tmp_970[20], _tmp_970[17] }), .Y(_09539_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32888_ ( .A({ _tmp_970[8], _tmp_970[5], _tmp_970[3:2] }), .Y(_09540_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32889_ ( .A({ _tmp_970[15:14], _tmp_970[12], _tmp_970[9] }), .Y(_09541_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32890_ ( .A({ _wvalid_963, _05362_ }), .Y(_05363_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32891_ ( .A({ _dataflow_slice_valid_113, _09542_ }), .Y(_05365_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32892_ ( .A({ _tmp_976, _09543_ }), .Y(_09542_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32893_ ( .A({ _09544_, _tmp_975[0], _tmp_975[33:32] }), .Y(_09543_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32894_ ( .A({ _09553_, _09552_, _09550_, _09545_ }), .Y(_09544_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32895_ ( .A({ _09549_, _09548_, _09547_, _09546_ }), .Y(_09545_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32896_ ( .A({ _tmp_975[24], _tmp_975[21], _tmp_975[19:18] }), .Y(_09546_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32897_ ( .A({ _tmp_975[31], _tmp_975[29:28], _tmp_975[25] }), .Y(_09547_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32898_ ( .A({ _tmp_975[7:6], _tmp_975[4], _tmp_975[1] }), .Y(_09548_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32899_ ( .A({ _tmp_975[16], _tmp_975[13], _tmp_975[11:10] }), .Y(_09549_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32900_ ( .A({ _09551_, _tmp_975[30], _tmp_975[27:26] }), .Y(_09550_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32901_ ( .A({ _tmp_975[23:22], _tmp_975[20], _tmp_975[17] }), .Y(_09551_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32902_ ( .A({ _tmp_975[8], _tmp_975[5], _tmp_975[3:2] }), .Y(_09552_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32903_ ( .A({ _tmp_975[15:14], _tmp_975[12], _tmp_975[9] }), .Y(_09553_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32904_ ( .A({ _wvalid_974, _05365_ }), .Y(_05366_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32905_ ( .A({ _dataflow_slice_valid_116, _09554_ }), .Y(_05368_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32906_ ( .A({ _tmp_978, _09555_ }), .Y(_09554_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32907_ ( .A({ _09556_, _tmp_977[0], _tmp_977[33:32] }), .Y(_09555_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32908_ ( .A({ _09565_, _09564_, _09562_, _09557_ }), .Y(_09556_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32909_ ( .A({ _09561_, _09560_, _09559_, _09558_ }), .Y(_09557_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32910_ ( .A({ _tmp_977[24], _tmp_977[21], _tmp_977[19:18] }), .Y(_09558_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32911_ ( .A({ _tmp_977[31], _tmp_977[29:28], _tmp_977[25] }), .Y(_09559_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32912_ ( .A({ _tmp_977[7:6], _tmp_977[4], _tmp_977[1] }), .Y(_09560_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32913_ ( .A({ _tmp_977[16], _tmp_977[13], _tmp_977[11:10] }), .Y(_09561_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32914_ ( .A({ _09563_, _tmp_977[30], _tmp_977[27:26] }), .Y(_09562_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32915_ ( .A({ _tmp_977[23:22], _tmp_977[20], _tmp_977[17] }), .Y(_09563_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32916_ ( .A({ _tmp_977[8], _tmp_977[5], _tmp_977[3:2] }), .Y(_09564_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32917_ ( .A({ _tmp_977[15:14], _tmp_977[12], _tmp_977[9] }), .Y(_09565_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32918_ ( .A({ _wvalid_974, _05368_ }), .Y(_05369_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32919_ ( .A({ _dataflow_slice_valid_119, _09566_ }), .Y(_05371_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32920_ ( .A({ _tmp_980, _09567_ }), .Y(_09566_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32921_ ( .A({ _09568_, _tmp_979[0], _tmp_979[33:32] }), .Y(_09567_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32922_ ( .A({ _09577_, _09576_, _09574_, _09569_ }), .Y(_09568_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32923_ ( .A({ _09573_, _09572_, _09571_, _09570_ }), .Y(_09569_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32924_ ( .A({ _tmp_979[24], _tmp_979[21], _tmp_979[19:18] }), .Y(_09570_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32925_ ( .A({ _tmp_979[31], _tmp_979[29:28], _tmp_979[25] }), .Y(_09571_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32926_ ( .A({ _tmp_979[7:6], _tmp_979[4], _tmp_979[1] }), .Y(_09572_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32927_ ( .A({ _tmp_979[16], _tmp_979[13], _tmp_979[11:10] }), .Y(_09573_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32928_ ( .A({ _09575_, _tmp_979[30], _tmp_979[27:26] }), .Y(_09574_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32929_ ( .A({ _tmp_979[23:22], _tmp_979[20], _tmp_979[17] }), .Y(_09575_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32930_ ( .A({ _tmp_979[8], _tmp_979[5], _tmp_979[3:2] }), .Y(_09576_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32931_ ( .A({ _tmp_979[15:14], _tmp_979[12], _tmp_979[9] }), .Y(_09577_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32932_ ( .A({ _wvalid_974, _05371_ }), .Y(_05372_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32933_ ( .A({ _dataflow_slice_valid_122, _09578_ }), .Y(_05374_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32934_ ( .A({ _tmp_982, _09579_ }), .Y(_09578_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32935_ ( .A({ _09580_, _tmp_981[0], _tmp_981[33:32] }), .Y(_09579_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32936_ ( .A({ _09589_, _09588_, _09586_, _09581_ }), .Y(_09580_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32937_ ( .A({ _09585_, _09584_, _09583_, _09582_ }), .Y(_09581_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32938_ ( .A({ _tmp_981[24], _tmp_981[21], _tmp_981[19:18] }), .Y(_09582_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32939_ ( .A({ _tmp_981[31], _tmp_981[29:28], _tmp_981[25] }), .Y(_09583_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32940_ ( .A({ _tmp_981[7:6], _tmp_981[4], _tmp_981[1] }), .Y(_09584_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32941_ ( .A({ _tmp_981[16], _tmp_981[13], _tmp_981[11:10] }), .Y(_09585_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32942_ ( .A({ _09587_, _tmp_981[30], _tmp_981[27:26] }), .Y(_09586_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32943_ ( .A({ _tmp_981[23:22], _tmp_981[20], _tmp_981[17] }), .Y(_09587_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32944_ ( .A({ _tmp_981[8], _tmp_981[5], _tmp_981[3:2] }), .Y(_09588_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32945_ ( .A({ _tmp_981[15:14], _tmp_981[12], _tmp_981[9] }), .Y(_09589_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32946_ ( .A({ _wvalid_974, _05374_ }), .Y(_05375_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32947_ ( .A({ _dataflow__delay_valid_132, _09590_ }), .Y(_05377_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32948_ ( .A({ _tmp_13, _09591_ }), .Y(_09590_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32949_ ( .A({ _09592_, _tmp_12[0], _tmp_12[33:32] }), .Y(_09591_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32950_ ( .A({ _09601_, _09600_, _09598_, _09593_ }), .Y(_09592_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32951_ ( .A({ _09597_, _09596_, _09595_, _09594_ }), .Y(_09593_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32952_ ( .A({ _tmp_12[24], _tmp_12[21], _tmp_12[19:18] }), .Y(_09594_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32953_ ( .A({ _tmp_12[31], _tmp_12[29:28], _tmp_12[25] }), .Y(_09595_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32954_ ( .A({ _tmp_12[7:6], _tmp_12[4], _tmp_12[1] }), .Y(_09596_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32955_ ( .A({ _tmp_12[16], _tmp_12[13], _tmp_12[11:10] }), .Y(_09597_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32956_ ( .A({ _09599_, _tmp_12[30], _tmp_12[27:26] }), .Y(_09598_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32957_ ( .A({ _tmp_12[23:22], _tmp_12[20], _tmp_12[17] }), .Y(_09599_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32958_ ( .A({ _tmp_12[8], _tmp_12[5], _tmp_12[3:2] }), .Y(_09600_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32959_ ( .A({ _tmp_12[15:14], _tmp_12[12], _tmp_12[9] }), .Y(_09601_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32960_ ( .A({ _wvalid_11, _05377_ }), .Y(_05378_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32961_ ( .A({ saxi_bready, saxi_bvalid }), .Y(_05380_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32962_ ( .A({ saxi_awvalid, saxi_awready }), .Y(_05382_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32963_ ( .A({ saxi_arvalid, saxi_arready }), .Y(_05383_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32964_ ( .A({ saxi_rvalid, saxi_rready }), .Y(_05385_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32965_ ( .A({ _tmp_7, _05384_, _04890_ }), .Y(_05386_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32966_ ( .A({ _saxi_register_fsm[0], _08047_, _05385_ }), .Y(_05384_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32967_ ( .A({ _tmp_7, _05384_, _04978_ }), .Y(_05387_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32968_ ( .A({ _tmp_7, _05384_, _04979_ }), .Y(_05388_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32969_ ( .A({ _tmp_7, _05384_, _04980_ }), .Y(_05389_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32970_ ( .A({ _tmp_7, _05384_, _04981_ }), .Y(_05390_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32971_ ( .A({ _tmp_7, _05384_, _04982_ }), .Y(_05391_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32972_ ( .A({ _tmp_7, _05384_, _04983_ }), .Y(_05392_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32973_ ( .A({ _tmp_7, _05384_, _04984_ }), .Y(_05393_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32974_ ( .A({ _tmp_7, _05384_, _04985_ }), .Y(_05394_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32975_ ( .A({ _tmp_7, _05384_, _04986_ }), .Y(_05395_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32976_ ( .A({ _tmp_7, _05384_, _04987_ }), .Y(_05396_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32977_ ( .A({ _tmp_7, _05384_, _04988_ }), .Y(_05397_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32978_ ( .A({ _tmp_7, _05384_, _04989_ }), .Y(_05398_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32979_ ( .A({ _tmp_7, _05384_, _04990_ }), .Y(_05399_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32980_ ( .A({ _05381_, _04890_ }), .Y(_05400_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32981_ ( .A({ saxi_wvalid, saxi_wready }), .Y(_05381_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32982_ ( .A({ _05381_, _04978_ }), .Y(_05401_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32983_ ( .A({ _05381_, _04979_ }), .Y(_05402_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32984_ ( .A({ _05381_, _04980_ }), .Y(_05403_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32985_ ( .A({ _05381_, _04981_ }), .Y(_05404_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32986_ ( .A({ _05381_, _04982_ }), .Y(_05405_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32987_ ( .A({ _05381_, _04983_ }), .Y(_05406_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32988_ ( .A({ _05381_, _04984_ }), .Y(_05407_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32989_ ( .A({ _05381_, _04985_ }), .Y(_05408_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32990_ ( .A({ _05381_, _04986_ }), .Y(_05409_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32991_ ( .A({ _05381_, _04987_ }), .Y(_05410_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32992_ ( .A({ _05381_, _04988_ }), .Y(_05411_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32993_ ( .A({ _05381_, _04989_ }), .Y(_05412_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32994_ ( .A({ _05381_, _04990_ }), .Y(_05413_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _32995_ ( .A({ _maxi_read_start, _09602_, _maxi_read_op_sel[1:0] }), .Y(_05414_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32996_ ( .A({ _maxi_read_op_sel[3], _09603_, _maxi_read_op_sel[2] }), .Y(_09602_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32997_ ( .A(_maxi_read_op_sel[7:4]), .Y(_09603_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32998_ ( .A({ _05414_, _09495_ }), .Y(_05415_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32999_ ( .A({ _dataflow_slice_valid_100, _09494_ }), .Y(_05355_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33000_ ( .A({ _09604_, _05355_ }), .Y(_05416_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33001_ ( .A({ _tmp_964[0], _09496_, _tmp_964[33:32] }), .Y(_09604_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33002_ ( .A({ _05414_, _09507_ }), .Y(_05417_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33003_ ( .A({ _dataflow_slice_valid_103, _09506_ }), .Y(_05358_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33004_ ( .A({ _09605_, _05358_ }), .Y(_05418_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33005_ ( .A({ _tmp_966[0], _09508_, _tmp_966[33:32] }), .Y(_09605_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33006_ ( .A({ _05414_, _09519_ }), .Y(_05419_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33007_ ( .A({ _dataflow_slice_valid_106, _09518_ }), .Y(_05361_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33008_ ( .A({ _09606_, _05361_ }), .Y(_05420_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33009_ ( .A({ _tmp_968[0], _09520_, _tmp_968[33:32] }), .Y(_09606_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33010_ ( .A({ _05414_, _09531_ }), .Y(_05421_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33011_ ( .A({ _dataflow_slice_valid_109, _09530_ }), .Y(_05364_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33012_ ( .A({ _09607_, _05364_ }), .Y(_05422_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33013_ ( .A({ _tmp_970[0], _09532_, _tmp_970[33:32] }), .Y(_09607_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33014_ ( .A({ _stream_matmul_15_source_20_source_ram_renable, _04991_ }), .Y(_tmp_1033) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _33015_ ( .A({ _maxi_read_start, _maxi_read_op_sel[1], _09608_, _maxi_read_op_sel[0] }), .Y(_05423_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33016_ ( .A({ _09603_, _maxi_read_op_sel[3:2] }), .Y(_09608_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33017_ ( .A({ _05423_, _09211_ }), .Y(_05424_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33018_ ( .A({ _dataflow_slice_valid_4, _09210_ }), .Y(_05283_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33019_ ( .A({ _09609_, _05283_ }), .Y(_05425_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33020_ ( .A({ _tmp_19[0], _09212_, _tmp_19[33:32] }), .Y(_09609_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33021_ ( .A({ _09610_, _stream_max_pool_serial_9_sink_3_sink_waddr[1] }), .Y(_05426_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33022_ ( .A({ _09611_, _stream_max_pool_serial_9_sink_3_sink_waddr[0] }), .Y(_09610_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33023_ ( .A({ _09613_, _09612_, _stream_max_pool_serial_9_sink_3_sink_ram_sel[2], _stream_max_pool_serial_9_sink_3_sink_ram_sel[0] }), .Y(_09611_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33024_ ( .A({ _stream_max_pool_serial_9_sink_3_sink_ram_sel[1], _stream_max_pool_serial_9_sink_3_sink_wenable, _stream_max_pool_serial_9_sink_3_sink_ram_sel[7] }), .Y(_09612_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33025_ ( .A(_stream_max_pool_serial_9_sink_3_sink_ram_sel[6:3]), .Y(_09613_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33026_ ( .A({ _tmp_910, _05434_ }), .Y(_tmp_915) );
  \$lut  #( .LUT(16'h8f00), .WIDTH(4) ) _33027_ ( .A({ _05433_, _dataflow_cat_valid_96, _09203_, _09208_ }), .Y(_05434_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33028_ ( .A({ _tmp_946, _tmp_934, _tmp_922, _tmp_910 }), .Y(_05433_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33029_ ( .A({ _tmp_918, _05434_, _tmp_910 }), .Y(_05427_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33030_ ( .A({ _tmp_917, _05434_, _tmp_910 }), .Y(_05428_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33031_ ( .A({ _maxi_write_start, _09208_ }), .Y(_05429_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33032_ ( .A({ _05429_, _09614_, _tmp_920, _tmp_919 }), .Y(_05430_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33033_ ( .A({ _09615_, _tmp_921[0] }), .Y(_09614_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33034_ ( .A({ _09625_, _09620_, _09618_, _09616_ }), .Y(_09615_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33035_ ( .A({ _09617_, _tmp_921[33:31] }), .Y(_09616_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33036_ ( .A({ _tmp_921[29:28], _tmp_921[26], _tmp_921[23] }), .Y(_09617_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33037_ ( .A({ _09619_, _tmp_921[2:1] }), .Y(_09618_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33038_ ( .A(_tmp_921[6:3]), .Y(_09619_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33039_ ( .A({ _09624_, _09623_, _09622_, _09621_ }), .Y(_09620_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33040_ ( .A(_tmp_921[14:11]), .Y(_09621_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33041_ ( .A(_tmp_921[10:7]), .Y(_09622_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33042_ ( .A(_tmp_921[22:19]), .Y(_09623_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33043_ ( .A(_tmp_921[18:15]), .Y(_09624_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33044_ ( .A({ _tmp_921[30], _tmp_921[27], _tmp_921[25:24] }), .Y(_09625_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33045_ ( .A({ _09614_, _05434_, _tmp_910 }), .Y(_05431_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33046_ ( .A({ _09615_, _tmp_921[0], _05434_, _tmp_910 }), .Y(_05432_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33047_ ( .A({ _05423_, _09223_ }), .Y(_05435_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33048_ ( .A({ _dataflow_slice_valid_7, _09222_ }), .Y(_05286_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33049_ ( .A({ _09626_, _05286_ }), .Y(_05436_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33050_ ( .A({ _tmp_21[0], _09224_, _tmp_21[33:32] }), .Y(_09626_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33051_ ( .A({ _09627_, _stream_max_pool_serial_9_sink_3_sink_waddr[1] }), .Y(_05437_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33052_ ( .A({ _stream_max_pool_serial_9_sink_3_sink_waddr[0], _09611_ }), .Y(_09627_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33053_ ( .A({ _tmp_922, _05434_ }), .Y(_tmp_927) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33054_ ( .A({ _tmp_930, _05434_, _tmp_922 }), .Y(_05438_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33055_ ( .A({ _tmp_929, _05434_, _tmp_922 }), .Y(_05439_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33056_ ( .A({ _05429_, _09628_, _tmp_932, _tmp_931 }), .Y(_05440_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33057_ ( .A({ _09629_, _tmp_933[0] }), .Y(_09628_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33058_ ( .A({ _09639_, _09634_, _09632_, _09630_ }), .Y(_09629_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33059_ ( .A({ _09631_, _tmp_933[33:31] }), .Y(_09630_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33060_ ( .A({ _tmp_933[29:28], _tmp_933[26], _tmp_933[23] }), .Y(_09631_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33061_ ( .A({ _09633_, _tmp_933[2:1] }), .Y(_09632_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33062_ ( .A(_tmp_933[6:3]), .Y(_09633_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33063_ ( .A({ _09638_, _09637_, _09636_, _09635_ }), .Y(_09634_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33064_ ( .A(_tmp_933[14:11]), .Y(_09635_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33065_ ( .A(_tmp_933[10:7]), .Y(_09636_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33066_ ( .A(_tmp_933[22:19]), .Y(_09637_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33067_ ( .A(_tmp_933[18:15]), .Y(_09638_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33068_ ( .A({ _tmp_933[30], _tmp_933[27], _tmp_933[25:24] }), .Y(_09639_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33069_ ( .A({ _09628_, _05434_, _tmp_922 }), .Y(_05441_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33070_ ( .A({ _09629_, _tmp_933[0], _05434_, _tmp_922 }), .Y(_05442_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33071_ ( .A({ _05423_, _09235_ }), .Y(_05443_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33072_ ( .A({ _dataflow_slice_valid_10, _09234_ }), .Y(_05289_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33073_ ( .A({ _09640_, _05289_ }), .Y(_05444_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33074_ ( .A({ _tmp_23[0], _09236_, _tmp_23[33:32] }), .Y(_09640_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33075_ ( .A({ _stream_max_pool_serial_9_sink_3_sink_waddr[1], _09610_ }), .Y(_05445_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33076_ ( .A({ _tmp_934, _05434_ }), .Y(_tmp_939) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33077_ ( .A({ _tmp_942, _05434_, _tmp_934 }), .Y(_05446_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33078_ ( .A({ _tmp_941, _05434_, _tmp_934 }), .Y(_05447_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33079_ ( .A({ _05429_, _09641_, _tmp_944, _tmp_943 }), .Y(_05448_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33080_ ( .A({ _09642_, _tmp_945[0] }), .Y(_09641_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33081_ ( .A({ _09652_, _09647_, _09645_, _09643_ }), .Y(_09642_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33082_ ( .A({ _09644_, _tmp_945[33:31] }), .Y(_09643_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33083_ ( .A({ _tmp_945[29:28], _tmp_945[26], _tmp_945[23] }), .Y(_09644_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33084_ ( .A({ _09646_, _tmp_945[2:1] }), .Y(_09645_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33085_ ( .A(_tmp_945[6:3]), .Y(_09646_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33086_ ( .A({ _09651_, _09650_, _09649_, _09648_ }), .Y(_09647_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33087_ ( .A(_tmp_945[14:11]), .Y(_09648_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33088_ ( .A(_tmp_945[10:7]), .Y(_09649_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33089_ ( .A(_tmp_945[22:19]), .Y(_09650_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33090_ ( .A(_tmp_945[18:15]), .Y(_09651_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33091_ ( .A({ _tmp_945[30], _tmp_945[27], _tmp_945[25:24] }), .Y(_09652_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33092_ ( .A({ _09641_, _05434_, _tmp_934 }), .Y(_05449_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33093_ ( .A({ _09642_, _tmp_945[0], _05434_, _tmp_934 }), .Y(_05450_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33094_ ( .A({ _05423_, _09247_ }), .Y(_05451_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33095_ ( .A({ _dataflow_slice_valid_13, _09246_ }), .Y(_05292_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33096_ ( .A({ _09653_, _05292_ }), .Y(_05452_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33097_ ( .A({ _tmp_25[0], _09248_, _tmp_25[33:32] }), .Y(_09653_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33098_ ( .A({ _stream_conv2d_8_source_8_source_ram_renable, _04992_ }), .Y(_tmp_347) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33099_ ( .A({ _stream_max_pool_serial_9_sink_3_sink_waddr[1], _09627_ }), .Y(_05453_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33100_ ( .A({ _tmp_946, _05434_ }), .Y(_tmp_951) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33101_ ( .A({ _tmp_954, _05434_, _tmp_946 }), .Y(_05454_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33102_ ( .A({ _tmp_953, _05434_, _tmp_946 }), .Y(_05455_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33103_ ( .A({ _05429_, _09654_, _tmp_956, _tmp_955 }), .Y(_05456_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33104_ ( .A({ _09655_, _tmp_957[0] }), .Y(_09654_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33105_ ( .A({ _09665_, _09660_, _09658_, _09656_ }), .Y(_09655_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33106_ ( .A({ _09657_, _tmp_957[33:31] }), .Y(_09656_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33107_ ( .A({ _tmp_957[29:28], _tmp_957[26], _tmp_957[23] }), .Y(_09657_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33108_ ( .A({ _09659_, _tmp_957[2:1] }), .Y(_09658_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33109_ ( .A(_tmp_957[6:3]), .Y(_09659_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33110_ ( .A({ _09664_, _09663_, _09662_, _09661_ }), .Y(_09660_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33111_ ( .A(_tmp_957[14:11]), .Y(_09661_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33112_ ( .A(_tmp_957[10:7]), .Y(_09662_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33113_ ( .A(_tmp_957[22:19]), .Y(_09663_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33114_ ( .A(_tmp_957[18:15]), .Y(_09664_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33115_ ( .A({ _tmp_957[30], _tmp_957[27], _tmp_957[25:24] }), .Y(_09665_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33116_ ( .A({ _09654_, _05434_, _tmp_946 }), .Y(_05457_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33117_ ( .A({ _09655_, _tmp_957[0], _05434_, _tmp_946 }), .Y(_05458_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33118_ ( .A({ _stream_matmul_15_source_8_source_ram_renable, _04993_ }), .Y(_tmp_1003) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33119_ ( .A({ _maxi_read_start, _maxi_read_op_sel[1:0], _09608_ }), .Y(_05459_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33120_ ( .A({ _05459_, _09258_ }), .Y(_05460_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33121_ ( .A({ _dataflow_slice_valid_17, _tmp_34, _09258_ }), .Y(_05295_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33122_ ( .A({ _09666_, _05295_ }), .Y(_05461_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33123_ ( .A({ _09668_, _09667_, _tmp_32[1:0] }), .Y(_09666_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33124_ ( .A(_tmp_32[9:6]), .Y(_09667_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33125_ ( .A(_tmp_32[5:2]), .Y(_09668_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33126_ ( .A({ _05152_, _05461_ }), .Y(_05462_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33127_ ( .A({ _05153_, _05295_ }), .Y(_05463_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33128_ ( .A({ _05154_, _05295_ }), .Y(_05464_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33129_ ( .A({ _05155_, _05295_ }), .Y(_05465_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33130_ ( .A({ _05156_, _05295_ }), .Y(_05466_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33131_ ( .A({ _05157_, _05295_ }), .Y(_05467_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33132_ ( .A({ _05158_, _05295_ }), .Y(_05468_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33133_ ( .A({ _05159_, _05295_ }), .Y(_05469_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33134_ ( .A({ _05160_, _05295_ }), .Y(_05470_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33135_ ( .A({ _05152_, _05295_ }), .Y(_05471_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33136_ ( .A({ _09669_, _05295_ }), .Y(_05472_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33137_ ( .A({ _09259_, _tmp_33[33:32] }), .Y(_09669_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33138_ ( .A({ _maxi_read_start, _maxi_read_op_sel[1:0], _09670_ }), .Y(_05473_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33139_ ( .A({ _09603_, _maxi_read_op_sel[2], _maxi_read_op_sel[3] }), .Y(_09670_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33140_ ( .A({ _05473_, _09447_ }), .Y(_05474_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33141_ ( .A({ _dataflow_slice_valid_78, _09446_ }), .Y(_05343_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33142_ ( .A({ _09671_, _05343_ }), .Y(_05475_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33143_ ( .A({ _tmp_853[0], _09448_, _tmp_853[33:32] }), .Y(_09671_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33144_ ( .A({ _09672_, _stream_matmul_15_sink_21_sink_waddr[1] }), .Y(_05476_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33145_ ( .A({ _09673_, _stream_matmul_15_sink_21_sink_waddr[0] }), .Y(_09672_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33146_ ( .A({ _09675_, _09674_, _stream_matmul_15_sink_21_sink_ram_sel[3], _stream_matmul_15_sink_21_sink_ram_sel[1] }), .Y(_09673_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33147_ ( .A({ _stream_matmul_15_sink_21_sink_ram_sel[2], _stream_matmul_15_sink_21_sink_ram_sel[0], _stream_matmul_15_sink_21_sink_wenable }), .Y(_09674_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33148_ ( .A(_stream_matmul_15_sink_21_sink_ram_sel[7:4]), .Y(_09675_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33149_ ( .A({ _tmp_1119, _05484_ }), .Y(_tmp_1124) );
  \$lut  #( .LUT(16'h8f00), .WIDTH(4) ) _33150_ ( .A({ _05483_, _dataflow_cat_valid_131, _09203_, _09209_ }), .Y(_05484_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33151_ ( .A({ _tmp_1155, _tmp_1143, _tmp_1131, _tmp_1119 }), .Y(_05483_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33152_ ( .A({ _tmp_1127, _05484_, _tmp_1119 }), .Y(_05477_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33153_ ( .A({ _tmp_1126, _05484_, _tmp_1119 }), .Y(_05478_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33154_ ( .A({ _maxi_write_start, _09209_ }), .Y(_05479_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33155_ ( .A({ _05479_, _09676_, _tmp_1129, _tmp_1128 }), .Y(_05480_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33156_ ( .A({ _09677_, _tmp_1130[0] }), .Y(_09676_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33157_ ( .A({ _09687_, _09682_, _09680_, _09678_ }), .Y(_09677_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33158_ ( .A({ _09679_, _tmp_1130[33:31] }), .Y(_09678_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33159_ ( .A({ _tmp_1130[29:28], _tmp_1130[26], _tmp_1130[23] }), .Y(_09679_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33160_ ( .A({ _09681_, _tmp_1130[2:1] }), .Y(_09680_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33161_ ( .A(_tmp_1130[6:3]), .Y(_09681_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33162_ ( .A({ _09686_, _09685_, _09684_, _09683_ }), .Y(_09682_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33163_ ( .A(_tmp_1130[14:11]), .Y(_09683_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33164_ ( .A(_tmp_1130[10:7]), .Y(_09684_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33165_ ( .A(_tmp_1130[22:19]), .Y(_09685_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33166_ ( .A(_tmp_1130[18:15]), .Y(_09686_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33167_ ( .A({ _tmp_1130[30], _tmp_1130[27], _tmp_1130[25:24] }), .Y(_09687_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33168_ ( .A({ _09676_, _05484_, _tmp_1119 }), .Y(_05481_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33169_ ( .A({ _09677_, _tmp_1130[0], _05484_, _tmp_1119 }), .Y(_05482_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33170_ ( .A({ _05459_, _09269_ }), .Y(_05485_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33171_ ( .A({ _dataflow_slice_valid_20, _tmp_65, _09269_ }), .Y(_05298_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33172_ ( .A({ _09688_, _05298_ }), .Y(_05486_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33173_ ( .A({ _09690_, _09689_, _tmp_63[1:0] }), .Y(_09688_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33174_ ( .A(_tmp_63[9:6]), .Y(_09689_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33175_ ( .A(_tmp_63[5:2]), .Y(_09690_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33176_ ( .A({ _05161_, _05486_ }), .Y(_05487_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33177_ ( .A({ _05162_, _05298_ }), .Y(_05488_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33178_ ( .A({ _05163_, _05298_ }), .Y(_05489_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33179_ ( .A({ _05164_, _05298_ }), .Y(_05490_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33180_ ( .A({ _05165_, _05298_ }), .Y(_05491_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33181_ ( .A({ _05166_, _05298_ }), .Y(_05492_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33182_ ( .A({ _05167_, _05298_ }), .Y(_05493_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33183_ ( .A({ _05168_, _05298_ }), .Y(_05494_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33184_ ( .A({ _05169_, _05298_ }), .Y(_05495_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33185_ ( .A({ _05161_, _05298_ }), .Y(_05496_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33186_ ( .A({ _09691_, _05298_ }), .Y(_05497_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33187_ ( .A({ _09270_, _tmp_64[33:32] }), .Y(_09691_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33188_ ( .A({ _05473_, _09459_ }), .Y(_05498_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33189_ ( .A({ _dataflow_slice_valid_81, _09458_ }), .Y(_05346_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33190_ ( .A({ _09692_, _05346_ }), .Y(_05499_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33191_ ( .A({ _tmp_855[0], _09460_, _tmp_855[33:32] }), .Y(_09692_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33192_ ( .A({ _09693_, _stream_matmul_15_sink_21_sink_waddr[1] }), .Y(_05500_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33193_ ( .A({ _stream_matmul_15_sink_21_sink_waddr[0], _09673_ }), .Y(_09693_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33194_ ( .A({ _tmp_1131, _05484_ }), .Y(_tmp_1136) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33195_ ( .A({ _tmp_1139, _05484_, _tmp_1131 }), .Y(_05501_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33196_ ( .A({ _tmp_1138, _05484_, _tmp_1131 }), .Y(_05502_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33197_ ( .A({ _05479_, _09694_, _tmp_1141, _tmp_1140 }), .Y(_05503_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33198_ ( .A({ _09695_, _tmp_1142[0] }), .Y(_09694_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33199_ ( .A({ _09705_, _09700_, _09698_, _09696_ }), .Y(_09695_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33200_ ( .A({ _09697_, _tmp_1142[33:31] }), .Y(_09696_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33201_ ( .A({ _tmp_1142[29:28], _tmp_1142[26], _tmp_1142[23] }), .Y(_09697_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33202_ ( .A({ _09699_, _tmp_1142[2:1] }), .Y(_09698_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33203_ ( .A(_tmp_1142[6:3]), .Y(_09699_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33204_ ( .A({ _09704_, _09703_, _09702_, _09701_ }), .Y(_09700_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33205_ ( .A(_tmp_1142[14:11]), .Y(_09701_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33206_ ( .A(_tmp_1142[10:7]), .Y(_09702_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33207_ ( .A(_tmp_1142[22:19]), .Y(_09703_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33208_ ( .A(_tmp_1142[18:15]), .Y(_09704_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33209_ ( .A({ _tmp_1142[30], _tmp_1142[27], _tmp_1142[25:24] }), .Y(_09705_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33210_ ( .A({ _09694_, _05484_, _tmp_1131 }), .Y(_05504_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33211_ ( .A({ _09695_, _tmp_1142[0], _05484_, _tmp_1131 }), .Y(_05505_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33212_ ( .A({ _05459_, _09280_ }), .Y(_05506_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33213_ ( .A({ _dataflow_slice_valid_23, _tmp_96, _09280_ }), .Y(_05301_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33214_ ( .A({ _09706_, _05301_ }), .Y(_05507_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33215_ ( .A({ _09708_, _09707_, _tmp_94[1:0] }), .Y(_09706_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33216_ ( .A(_tmp_94[9:6]), .Y(_09707_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33217_ ( .A(_tmp_94[5:2]), .Y(_09708_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33218_ ( .A({ _05170_, _05507_ }), .Y(_05508_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33219_ ( .A({ _05171_, _05301_ }), .Y(_05509_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33220_ ( .A({ _05172_, _05301_ }), .Y(_05510_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33221_ ( .A({ _05173_, _05301_ }), .Y(_05511_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33222_ ( .A({ _05174_, _05301_ }), .Y(_05512_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33223_ ( .A({ _05175_, _05301_ }), .Y(_05513_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33224_ ( .A({ _05176_, _05301_ }), .Y(_05514_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33225_ ( .A({ _05177_, _05301_ }), .Y(_05515_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33226_ ( .A({ _05178_, _05301_ }), .Y(_05516_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33227_ ( .A({ _05170_, _05301_ }), .Y(_05517_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33228_ ( .A({ _09709_, _05301_ }), .Y(_05518_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33229_ ( .A({ _09281_, _tmp_95[33:32] }), .Y(_09709_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33230_ ( .A({ _05473_, _09471_ }), .Y(_05519_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33231_ ( .A({ _dataflow_slice_valid_84, _09470_ }), .Y(_05349_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33232_ ( .A({ _09710_, _05349_ }), .Y(_05520_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33233_ ( .A({ _tmp_857[0], _09472_, _tmp_857[33:32] }), .Y(_09710_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33234_ ( .A({ _stream_matmul_15_sink_21_sink_waddr[1], _09672_ }), .Y(_05521_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33235_ ( .A({ _tmp_1143, _05484_ }), .Y(_tmp_1148) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33236_ ( .A({ _tmp_1151, _05484_, _tmp_1143 }), .Y(_05522_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33237_ ( .A({ _tmp_1150, _05484_, _tmp_1143 }), .Y(_05523_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33238_ ( .A({ _05479_, _09711_, _tmp_1153, _tmp_1152 }), .Y(_05524_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33239_ ( .A({ _09712_, _tmp_1154[0] }), .Y(_09711_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33240_ ( .A({ _09722_, _09717_, _09715_, _09713_ }), .Y(_09712_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33241_ ( .A({ _09714_, _tmp_1154[33:31] }), .Y(_09713_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33242_ ( .A({ _tmp_1154[29:28], _tmp_1154[26], _tmp_1154[23] }), .Y(_09714_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33243_ ( .A({ _09716_, _tmp_1154[2:1] }), .Y(_09715_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33244_ ( .A(_tmp_1154[6:3]), .Y(_09716_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33245_ ( .A({ _09721_, _09720_, _09719_, _09718_ }), .Y(_09717_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33246_ ( .A(_tmp_1154[14:11]), .Y(_09718_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33247_ ( .A(_tmp_1154[10:7]), .Y(_09719_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33248_ ( .A(_tmp_1154[22:19]), .Y(_09720_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33249_ ( .A(_tmp_1154[18:15]), .Y(_09721_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33250_ ( .A({ _tmp_1154[30], _tmp_1154[27], _tmp_1154[25:24] }), .Y(_09722_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33251_ ( .A({ _09711_, _05484_, _tmp_1143 }), .Y(_05525_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33252_ ( .A({ _09712_, _tmp_1154[0], _05484_, _tmp_1143 }), .Y(_05526_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33253_ ( .A({ _05459_, _09291_ }), .Y(_05527_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33254_ ( .A({ _dataflow_slice_valid_26, _tmp_127, _09291_ }), .Y(_05304_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33255_ ( .A({ _09723_, _05304_ }), .Y(_05528_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33256_ ( .A({ _09725_, _09724_, _tmp_125[1:0] }), .Y(_09723_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33257_ ( .A(_tmp_125[9:6]), .Y(_09724_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33258_ ( .A(_tmp_125[5:2]), .Y(_09725_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33259_ ( .A({ _05179_, _05528_ }), .Y(_05529_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33260_ ( .A({ _05180_, _05304_ }), .Y(_05530_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33261_ ( .A({ _05181_, _05304_ }), .Y(_05531_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33262_ ( .A({ _05182_, _05304_ }), .Y(_05532_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33263_ ( .A({ _05183_, _05304_ }), .Y(_05533_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33264_ ( .A({ _05184_, _05304_ }), .Y(_05534_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33265_ ( .A({ _05185_, _05304_ }), .Y(_05535_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33266_ ( .A({ _05186_, _05304_ }), .Y(_05536_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33267_ ( .A({ _05187_, _05304_ }), .Y(_05537_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33268_ ( .A({ _05179_, _05304_ }), .Y(_05538_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33269_ ( .A({ _09726_, _05304_ }), .Y(_05539_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33270_ ( .A({ _09292_, _tmp_126[33:32] }), .Y(_09726_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33271_ ( .A({ _stream_conv2d_8_source_28_source_ram_renable, _04994_ }), .Y(_tmp_457) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33272_ ( .A({ _05473_, _09483_ }), .Y(_05540_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33273_ ( .A({ _dataflow_slice_valid_87, _09482_ }), .Y(_05352_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33274_ ( .A({ _09727_, _05352_ }), .Y(_05541_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33275_ ( .A({ _tmp_859[0], _09484_, _tmp_859[33:32] }), .Y(_09727_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33276_ ( .A({ _stream_max_pool_serial_9_source_1_source_ram_renable, _04995_ }), .Y(_tmp_873) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33277_ ( .A({ _stream_matmul_15_sink_21_sink_waddr[1], _09693_ }), .Y(_05542_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33278_ ( .A({ _tmp_1155, _05484_ }), .Y(_tmp_1160) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33279_ ( .A({ _tmp_1163, _05484_, _tmp_1155 }), .Y(_05543_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33280_ ( .A({ _tmp_1162, _05484_, _tmp_1155 }), .Y(_05544_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33281_ ( .A({ _05479_, _09728_, _tmp_1165, _tmp_1164 }), .Y(_05545_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33282_ ( .A({ _09729_, _tmp_1166[0] }), .Y(_09728_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33283_ ( .A({ _09739_, _09734_, _09732_, _09730_ }), .Y(_09729_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33284_ ( .A({ _09731_, _tmp_1166[33:31] }), .Y(_09730_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33285_ ( .A({ _tmp_1166[29:28], _tmp_1166[26], _tmp_1166[23] }), .Y(_09731_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33286_ ( .A({ _09733_, _tmp_1166[2:1] }), .Y(_09732_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33287_ ( .A(_tmp_1166[6:3]), .Y(_09733_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33288_ ( .A({ _09738_, _09737_, _09736_, _09735_ }), .Y(_09734_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33289_ ( .A(_tmp_1166[14:11]), .Y(_09735_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33290_ ( .A(_tmp_1166[10:7]), .Y(_09736_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33291_ ( .A(_tmp_1166[22:19]), .Y(_09737_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33292_ ( .A(_tmp_1166[18:15]), .Y(_09738_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33293_ ( .A({ _tmp_1166[30], _tmp_1166[27], _tmp_1166[25:24] }), .Y(_09739_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33294_ ( .A({ _09728_, _05484_, _tmp_1155 }), .Y(_05546_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33295_ ( .A({ _09729_, _tmp_1166[0], _05484_, _tmp_1155 }), .Y(_05547_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _33296_ ( .A({ _maxi_read_start, _09602_, _maxi_read_op_sel[0], _maxi_read_op_sel[1] }), .Y(_05548_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33297_ ( .A({ _05548_, _09543_ }), .Y(_05549_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33298_ ( .A({ _dataflow_slice_valid_113, _09542_ }), .Y(_05367_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33299_ ( .A({ _09740_, _05367_ }), .Y(_05550_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33300_ ( .A({ _tmp_975[0], _09544_, _tmp_975[33:32] }), .Y(_09740_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33301_ ( .A({ _05548_, _09555_ }), .Y(_05551_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33302_ ( .A({ _dataflow_slice_valid_116, _09554_ }), .Y(_05370_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33303_ ( .A({ _09741_, _05370_ }), .Y(_05552_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33304_ ( .A({ _tmp_977[0], _09556_, _tmp_977[33:32] }), .Y(_09741_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33305_ ( .A({ _05548_, _09567_ }), .Y(_05553_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33306_ ( .A({ _dataflow_slice_valid_119, _09566_ }), .Y(_05373_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33307_ ( .A({ _09742_, _05373_ }), .Y(_05554_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33308_ ( .A({ _tmp_979[0], _09568_, _tmp_979[33:32] }), .Y(_09742_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33309_ ( .A({ _stream_conv2d_8_source_29_source_ram_renable, _04996_ }), .Y(_tmp_467) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33310_ ( .A({ _05548_, _09579_ }), .Y(_05555_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33311_ ( .A({ _dataflow_slice_valid_122, _09578_ }), .Y(_05376_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33312_ ( .A({ _09743_, _05376_ }), .Y(_05556_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33313_ ( .A({ _tmp_981[0], _09580_, _tmp_981[33:32] }), .Y(_09743_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33314_ ( .A({ _stream_matmul_15_source_19_source_ram_renable, _04997_ }), .Y(_tmp_1023) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33315_ ( .A({ _stream_conv2d_8_source_30_source_ram_renable, _04998_ }), .Y(_tmp_477) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33316_ ( .A({ _stream_conv2d_8_source_31_source_ram_renable, _04999_ }), .Y(_tmp_487) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33317_ ( .A({ _stream_conv2d_8_source_32_source_ram_renable, _05000_ }), .Y(_tmp_497) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33318_ ( .A({ _stream_conv2d_8_source_33_source_ram_renable, _05001_ }), .Y(_tmp_507) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33319_ ( .A({ _stream_conv2d_8_source_34_source_ram_renable, _05002_ }), .Y(_tmp_517) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33320_ ( .A({ _stream_conv2d_8_source_35_source_ram_renable, _05003_ }), .Y(_tmp_527) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33321_ ( .A({ _stream_conv2d_8_source_36_source_ram_renable, _05004_ }), .Y(_tmp_537) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33322_ ( .A({ _maxi_read_start, _09670_, _maxi_read_op_sel[1:0] }), .Y(_05557_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33323_ ( .A({ _05557_, _09303_ }), .Y(_05558_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33324_ ( .A({ _dataflow_slice_valid_30, _09302_ }), .Y(_05307_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33325_ ( .A({ _dataflow_slice_valid_30, _09744_, _09302_ }), .Y(_05559_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33326_ ( .A({ _09746_, _09745_, _tmp_161[1:0] }), .Y(_09744_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33327_ ( .A(_tmp_161[9:6]), .Y(_09745_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33328_ ( .A(_tmp_161[5:2]), .Y(_09746_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33329_ ( .A({ _05188_, _05559_ }), .Y(_05560_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33330_ ( .A({ _05189_, _05307_ }), .Y(_05561_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33331_ ( .A({ _05190_, _05307_ }), .Y(_05562_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33332_ ( .A({ _05188_, _05307_ }), .Y(_05563_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33333_ ( .A({ _09747_, _05307_ }), .Y(_05564_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33334_ ( .A({ _tmp_162[0], _09304_, _tmp_162[33:32] }), .Y(_09747_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33335_ ( .A({ _05557_, _09315_ }), .Y(_05565_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33336_ ( .A({ _dataflow_slice_valid_33, _09314_ }), .Y(_05310_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33337_ ( .A({ _dataflow_slice_valid_33, _09748_, _09314_ }), .Y(_05566_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33338_ ( .A({ _09750_, _09749_, _tmp_174[1:0] }), .Y(_09748_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33339_ ( .A(_tmp_174[9:6]), .Y(_09749_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33340_ ( .A(_tmp_174[5:2]), .Y(_09750_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33341_ ( .A({ _05191_, _05566_ }), .Y(_05567_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33342_ ( .A({ _05192_, _05310_ }), .Y(_05568_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33343_ ( .A({ _05193_, _05310_ }), .Y(_05569_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33344_ ( .A({ _05191_, _05310_ }), .Y(_05570_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33345_ ( .A({ _09751_, _05310_ }), .Y(_05571_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33346_ ( .A({ _tmp_175[0], _09316_, _tmp_175[33:32] }), .Y(_09751_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33347_ ( .A({ _05557_, _09327_ }), .Y(_05572_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33348_ ( .A({ _dataflow_slice_valid_36, _09326_ }), .Y(_05313_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33349_ ( .A({ _dataflow_slice_valid_36, _09752_, _09326_ }), .Y(_05573_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33350_ ( .A({ _09754_, _09753_, _tmp_187[1:0] }), .Y(_09752_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33351_ ( .A(_tmp_187[9:6]), .Y(_09753_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33352_ ( .A(_tmp_187[5:2]), .Y(_09754_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33353_ ( .A({ _05194_, _05573_ }), .Y(_05574_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33354_ ( .A({ _05195_, _05313_ }), .Y(_05575_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33355_ ( .A({ _05196_, _05313_ }), .Y(_05576_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33356_ ( .A({ _05194_, _05313_ }), .Y(_05577_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33357_ ( .A({ _09755_, _05313_ }), .Y(_05578_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33358_ ( .A({ _tmp_188[0], _09328_, _tmp_188[33:32] }), .Y(_09755_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33359_ ( .A({ _05557_, _09339_ }), .Y(_05579_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33360_ ( .A({ _dataflow_slice_valid_39, _09338_ }), .Y(_05316_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33361_ ( .A({ _dataflow_slice_valid_39, _09756_, _09338_ }), .Y(_05580_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33362_ ( .A({ _09758_, _09757_, _tmp_200[1:0] }), .Y(_09756_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33363_ ( .A(_tmp_200[9:6]), .Y(_09757_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33364_ ( .A(_tmp_200[5:2]), .Y(_09758_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33365_ ( .A({ _05197_, _05580_ }), .Y(_05581_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33366_ ( .A({ _05198_, _05316_ }), .Y(_05582_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33367_ ( .A({ _05199_, _05316_ }), .Y(_05583_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33368_ ( .A({ _05197_, _05316_ }), .Y(_05584_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33369_ ( .A({ _09759_, _05316_ }), .Y(_05585_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33370_ ( .A({ _tmp_201[0], _09340_, _tmp_201[33:32] }), .Y(_09759_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33371_ ( .A({ _stream_conv2d_8_source_19_source_ram_renable, _05005_ }), .Y(_tmp_367) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33372_ ( .A({ _stream_conv2d_8_source_20_source_ram_renable, _05006_ }), .Y(_tmp_377) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33373_ ( .A({ _stream_conv2d_8_source_21_source_ram_renable, _05007_ }), .Y(_tmp_387) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _33374_ ( .A({ _maxi_read_start, _09670_, _maxi_read_op_sel[0], _maxi_read_op_sel[1] }), .Y(_05586_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33375_ ( .A({ _05586_, _09351_ }), .Y(_05587_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33376_ ( .A({ _dataflow_slice_valid_43, _09350_ }), .Y(_05319_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33377_ ( .A({ _dataflow_slice_valid_43, _09760_, _09350_ }), .Y(_05588_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33378_ ( .A({ _09762_, _09761_, _tmp_218[1:0] }), .Y(_09760_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33379_ ( .A(_tmp_218[9:6]), .Y(_09761_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33380_ ( .A(_tmp_218[5:2]), .Y(_09762_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33381_ ( .A({ _05200_, _05588_ }), .Y(_05589_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33382_ ( .A({ _05201_, _05319_ }), .Y(_05590_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33383_ ( .A({ _05202_, _05319_ }), .Y(_05591_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33384_ ( .A({ _05200_, _05319_ }), .Y(_05592_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33385_ ( .A({ _09763_, _05319_ }), .Y(_05593_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33386_ ( .A({ _tmp_219[0], _09352_, _tmp_219[33:32] }), .Y(_09763_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33387_ ( .A({ _05586_, _09363_ }), .Y(_05594_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33388_ ( .A({ _dataflow_slice_valid_46, _09362_ }), .Y(_05322_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33389_ ( .A({ _dataflow_slice_valid_46, _09764_, _09362_ }), .Y(_05595_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33390_ ( .A({ _09766_, _09765_, _tmp_231[1:0] }), .Y(_09764_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33391_ ( .A(_tmp_231[9:6]), .Y(_09765_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33392_ ( .A(_tmp_231[5:2]), .Y(_09766_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33393_ ( .A({ _05203_, _05595_ }), .Y(_05596_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33394_ ( .A({ _05204_, _05322_ }), .Y(_05597_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33395_ ( .A({ _05205_, _05322_ }), .Y(_05598_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33396_ ( .A({ _05203_, _05322_ }), .Y(_05599_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33397_ ( .A({ _09767_, _05322_ }), .Y(_05600_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33398_ ( .A({ _tmp_232[0], _09364_, _tmp_232[33:32] }), .Y(_09767_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33399_ ( .A({ _05586_, _09375_ }), .Y(_05601_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33400_ ( .A({ _dataflow_slice_valid_49, _09374_ }), .Y(_05325_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33401_ ( .A({ _dataflow_slice_valid_49, _09768_, _09374_ }), .Y(_05602_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33402_ ( .A({ _09770_, _09769_, _tmp_244[1:0] }), .Y(_09768_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33403_ ( .A(_tmp_244[9:6]), .Y(_09769_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33404_ ( .A(_tmp_244[5:2]), .Y(_09770_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33405_ ( .A({ _05206_, _05602_ }), .Y(_05603_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33406_ ( .A({ _05207_, _05325_ }), .Y(_05604_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33407_ ( .A({ _05208_, _05325_ }), .Y(_05605_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33408_ ( .A({ _05206_, _05325_ }), .Y(_05606_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33409_ ( .A({ _09771_, _05325_ }), .Y(_05607_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33410_ ( .A({ _tmp_245[0], _09376_, _tmp_245[33:32] }), .Y(_09771_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33411_ ( .A({ _05586_, _09387_ }), .Y(_05608_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33412_ ( .A({ _dataflow_slice_valid_52, _09386_ }), .Y(_05328_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33413_ ( .A({ _dataflow_slice_valid_52, _09772_, _09386_ }), .Y(_05609_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33414_ ( .A({ _09774_, _09773_, _tmp_257[1:0] }), .Y(_09772_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33415_ ( .A(_tmp_257[9:6]), .Y(_09773_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33416_ ( .A(_tmp_257[5:2]), .Y(_09774_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33417_ ( .A({ _05209_, _05609_ }), .Y(_05610_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33418_ ( .A({ _05210_, _05328_ }), .Y(_05611_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33419_ ( .A({ _05211_, _05328_ }), .Y(_05612_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33420_ ( .A({ _05209_, _05328_ }), .Y(_05613_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33421_ ( .A({ _09775_, _05328_ }), .Y(_05614_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33422_ ( .A({ _tmp_258[0], _09388_, _tmp_258[33:32] }), .Y(_09775_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33423_ ( .A({ _stream_conv2d_8_source_22_source_ram_renable, _05008_ }), .Y(_tmp_397) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33424_ ( .A({ _stream_conv2d_8_source_23_source_ram_renable, _05009_ }), .Y(_tmp_407) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33425_ ( .A({ _stream_conv2d_8_source_24_source_ram_renable, _05010_ }), .Y(_tmp_417) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _33426_ ( .A({ _maxi_read_start, _maxi_read_op_sel[1], _09670_, _maxi_read_op_sel[0] }), .Y(_05615_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33427_ ( .A({ _05615_, _09399_ }), .Y(_05616_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33428_ ( .A({ _dataflow_slice_valid_56, _09398_ }), .Y(_05331_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33429_ ( .A({ _dataflow_slice_valid_56, _09776_, _09398_ }), .Y(_05617_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33430_ ( .A({ _09778_, _09777_, _tmp_275[1:0] }), .Y(_09776_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33431_ ( .A(_tmp_275[9:6]), .Y(_09777_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33432_ ( .A(_tmp_275[5:2]), .Y(_09778_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33433_ ( .A({ _05212_, _05617_ }), .Y(_05618_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33434_ ( .A({ _05213_, _05331_ }), .Y(_05619_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33435_ ( .A({ _05214_, _05331_ }), .Y(_05620_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33436_ ( .A({ _05212_, _05331_ }), .Y(_05621_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33437_ ( .A({ _09779_, _05331_ }), .Y(_05622_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33438_ ( .A({ _tmp_276[0], _09400_, _tmp_276[33:32] }), .Y(_09779_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33439_ ( .A({ _05615_, _09411_ }), .Y(_05623_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33440_ ( .A({ _dataflow_slice_valid_59, _09410_ }), .Y(_05334_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33441_ ( .A({ _dataflow_slice_valid_59, _09780_, _09410_ }), .Y(_05624_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33442_ ( .A({ _09782_, _09781_, _tmp_288[1:0] }), .Y(_09780_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33443_ ( .A(_tmp_288[9:6]), .Y(_09781_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33444_ ( .A(_tmp_288[5:2]), .Y(_09782_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33445_ ( .A({ _05215_, _05624_ }), .Y(_05625_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33446_ ( .A({ _05216_, _05334_ }), .Y(_05626_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33447_ ( .A({ _05217_, _05334_ }), .Y(_05627_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33448_ ( .A({ _05215_, _05334_ }), .Y(_05628_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33449_ ( .A({ _09783_, _05334_ }), .Y(_05629_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33450_ ( .A({ _tmp_289[0], _09412_, _tmp_289[33:32] }), .Y(_09783_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33451_ ( .A({ _05615_, _09423_ }), .Y(_05630_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33452_ ( .A({ _dataflow_slice_valid_62, _09422_ }), .Y(_05337_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33453_ ( .A({ _dataflow_slice_valid_62, _09784_, _09422_ }), .Y(_05631_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33454_ ( .A({ _09786_, _09785_, _tmp_301[1:0] }), .Y(_09784_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33455_ ( .A(_tmp_301[9:6]), .Y(_09785_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33456_ ( .A(_tmp_301[5:2]), .Y(_09786_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33457_ ( .A({ _05218_, _05631_ }), .Y(_05632_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33458_ ( .A({ _05219_, _05337_ }), .Y(_05633_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33459_ ( .A({ _05220_, _05337_ }), .Y(_05634_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33460_ ( .A({ _05218_, _05337_ }), .Y(_05635_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33461_ ( .A({ _09787_, _05337_ }), .Y(_05636_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33462_ ( .A({ _tmp_302[0], _09424_, _tmp_302[33:32] }), .Y(_09787_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33463_ ( .A({ _05615_, _09435_ }), .Y(_05637_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33464_ ( .A({ _dataflow_slice_valid_65, _09434_ }), .Y(_05340_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33465_ ( .A({ _dataflow_slice_valid_65, _09788_, _09434_ }), .Y(_05638_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33466_ ( .A({ _09790_, _09789_, _tmp_314[1:0] }), .Y(_09788_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33467_ ( .A(_tmp_314[9:6]), .Y(_09789_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33468_ ( .A(_tmp_314[5:2]), .Y(_09790_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33469_ ( .A({ _05221_, _05638_ }), .Y(_05639_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33470_ ( .A({ _05222_, _05340_ }), .Y(_05640_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33471_ ( .A({ _05223_, _05340_ }), .Y(_05641_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33472_ ( .A({ _05221_, _05340_ }), .Y(_05642_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33473_ ( .A({ _09791_, _05340_ }), .Y(_05643_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33474_ ( .A({ _tmp_315[0], _09436_, _tmp_315[33:32] }), .Y(_09791_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33475_ ( .A({ _stream_conv2d_8_source_25_source_ram_renable, _05011_ }), .Y(_tmp_427) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33476_ ( .A({ _stream_conv2d_8_source_26_source_ram_renable, _05012_ }), .Y(_tmp_437) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33477_ ( .A({ _stream_conv2d_8_source_27_source_ram_renable, _05013_ }), .Y(_tmp_447) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33478_ ( .A({ _09792_, _stream_conv2d_8_sink_37_sink_waddr[1] }), .Y(_05644_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33479_ ( .A({ _09793_, _stream_conv2d_8_sink_37_sink_waddr[0] }), .Y(_09792_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33480_ ( .A({ _09795_, _09794_, _stream_conv2d_8_sink_37_sink_ram_sel[3], _stream_conv2d_8_sink_37_sink_ram_sel[1] }), .Y(_09793_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33481_ ( .A({ _stream_conv2d_8_sink_37_sink_ram_sel[4], _stream_conv2d_8_sink_37_sink_ram_sel[2], _stream_conv2d_8_sink_37_sink_ram_sel[0] }), .Y(_09794_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33482_ ( .A({ _stream_conv2d_8_sink_37_sink_wenable, _stream_conv2d_8_sink_37_sink_ram_sel[7:5] }), .Y(_09795_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33483_ ( .A({ _tmp_799, _05652_ }), .Y(_tmp_804) );
  \$lut  #( .LUT(16'h8f00), .WIDTH(4) ) _33484_ ( .A({ _05651_, _dataflow_cat_valid_74, _09203_, _09204_ }), .Y(_05652_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33485_ ( .A({ _tmp_835, _tmp_823, _tmp_811, _tmp_799 }), .Y(_05651_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33486_ ( .A({ _tmp_807, _05652_, _tmp_799 }), .Y(_05645_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33487_ ( .A({ _tmp_806, _05652_, _tmp_799 }), .Y(_05646_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33488_ ( .A({ _maxi_write_start, _09204_ }), .Y(_05647_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33489_ ( .A({ _05647_, _09796_, _tmp_809, _tmp_808 }), .Y(_05648_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33490_ ( .A({ _09797_, _tmp_810[0] }), .Y(_09796_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33491_ ( .A({ _09807_, _09802_, _09800_, _09798_ }), .Y(_09797_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33492_ ( .A({ _09799_, _tmp_810[33:31] }), .Y(_09798_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33493_ ( .A({ _tmp_810[29:28], _tmp_810[26], _tmp_810[23] }), .Y(_09799_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33494_ ( .A({ _09801_, _tmp_810[2:1] }), .Y(_09800_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33495_ ( .A(_tmp_810[6:3]), .Y(_09801_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33496_ ( .A({ _09806_, _09805_, _09804_, _09803_ }), .Y(_09802_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33497_ ( .A(_tmp_810[14:11]), .Y(_09803_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33498_ ( .A(_tmp_810[10:7]), .Y(_09804_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33499_ ( .A(_tmp_810[22:19]), .Y(_09805_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33500_ ( .A(_tmp_810[18:15]), .Y(_09806_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33501_ ( .A({ _tmp_810[30], _tmp_810[27], _tmp_810[25:24] }), .Y(_09807_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33502_ ( .A({ _09796_, _05652_, _tmp_799 }), .Y(_05649_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33503_ ( .A({ _09797_, _tmp_810[0], _05652_, _tmp_799 }), .Y(_05650_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33504_ ( .A({ _09808_, _stream_conv2d_8_sink_37_sink_waddr[1] }), .Y(_05653_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33505_ ( .A({ _stream_conv2d_8_sink_37_sink_waddr[0], _09793_ }), .Y(_09808_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33506_ ( .A({ _tmp_811, _05652_ }), .Y(_tmp_816) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33507_ ( .A({ _tmp_819, _05652_, _tmp_811 }), .Y(_05654_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33508_ ( .A({ _tmp_818, _05652_, _tmp_811 }), .Y(_05655_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33509_ ( .A({ _05647_, _09809_, _tmp_821, _tmp_820 }), .Y(_05656_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33510_ ( .A({ _09810_, _tmp_822[0] }), .Y(_09809_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33511_ ( .A({ _09820_, _09815_, _09813_, _09811_ }), .Y(_09810_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33512_ ( .A({ _09812_, _tmp_822[33:31] }), .Y(_09811_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33513_ ( .A({ _tmp_822[29:28], _tmp_822[26], _tmp_822[23] }), .Y(_09812_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33514_ ( .A({ _09814_, _tmp_822[2:1] }), .Y(_09813_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33515_ ( .A(_tmp_822[6:3]), .Y(_09814_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33516_ ( .A({ _09819_, _09818_, _09817_, _09816_ }), .Y(_09815_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33517_ ( .A(_tmp_822[14:11]), .Y(_09816_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33518_ ( .A(_tmp_822[10:7]), .Y(_09817_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33519_ ( .A(_tmp_822[22:19]), .Y(_09818_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33520_ ( .A(_tmp_822[18:15]), .Y(_09819_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33521_ ( .A({ _tmp_822[30], _tmp_822[27], _tmp_822[25:24] }), .Y(_09820_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33522_ ( .A({ _09809_, _05652_, _tmp_811 }), .Y(_05657_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33523_ ( .A({ _09810_, _tmp_822[0], _05652_, _tmp_811 }), .Y(_05658_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33524_ ( .A({ _stream_conv2d_8_sink_37_sink_waddr[1], _09792_ }), .Y(_05659_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33525_ ( .A({ _tmp_823, _05652_ }), .Y(_tmp_828) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33526_ ( .A({ _tmp_831, _05652_, _tmp_823 }), .Y(_05660_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33527_ ( .A({ _tmp_830, _05652_, _tmp_823 }), .Y(_05661_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33528_ ( .A({ _05647_, _09821_, _tmp_833, _tmp_832 }), .Y(_05662_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33529_ ( .A({ _09822_, _tmp_834[0] }), .Y(_09821_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33530_ ( .A({ _09832_, _09827_, _09825_, _09823_ }), .Y(_09822_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33531_ ( .A({ _09824_, _tmp_834[33:31] }), .Y(_09823_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33532_ ( .A({ _tmp_834[29:28], _tmp_834[26], _tmp_834[23] }), .Y(_09824_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33533_ ( .A({ _09826_, _tmp_834[2:1] }), .Y(_09825_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33534_ ( .A(_tmp_834[6:3]), .Y(_09826_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33535_ ( .A({ _09831_, _09830_, _09829_, _09828_ }), .Y(_09827_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33536_ ( .A(_tmp_834[14:11]), .Y(_09828_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33537_ ( .A(_tmp_834[10:7]), .Y(_09829_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33538_ ( .A(_tmp_834[22:19]), .Y(_09830_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33539_ ( .A(_tmp_834[18:15]), .Y(_09831_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33540_ ( .A({ _tmp_834[30], _tmp_834[27], _tmp_834[25:24] }), .Y(_09832_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33541_ ( .A({ _09821_, _05652_, _tmp_823 }), .Y(_05663_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33542_ ( .A({ _09822_, _tmp_834[0], _05652_, _tmp_823 }), .Y(_05664_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33543_ ( .A({ _stream_conv2d_8_sink_37_sink_waddr[1], _09808_ }), .Y(_05665_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33544_ ( .A({ _tmp_835, _05652_ }), .Y(_tmp_840) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33545_ ( .A({ _tmp_843, _05652_, _tmp_835 }), .Y(_05666_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _33546_ ( .A({ _tmp_842, _05652_, _tmp_835 }), .Y(_05667_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33547_ ( .A({ _05647_, _09833_, _tmp_845, _tmp_844 }), .Y(_05668_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33548_ ( .A({ _09834_, _tmp_846[0] }), .Y(_09833_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33549_ ( .A({ _09844_, _09839_, _09837_, _09835_ }), .Y(_09834_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33550_ ( .A({ _09836_, _tmp_846[33:31] }), .Y(_09835_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33551_ ( .A({ _tmp_846[29:28], _tmp_846[26], _tmp_846[23] }), .Y(_09836_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33552_ ( .A({ _09838_, _tmp_846[2:1] }), .Y(_09837_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33553_ ( .A(_tmp_846[6:3]), .Y(_09838_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33554_ ( .A({ _09843_, _09842_, _09841_, _09840_ }), .Y(_09839_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33555_ ( .A(_tmp_846[14:11]), .Y(_09840_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33556_ ( .A(_tmp_846[10:7]), .Y(_09841_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33557_ ( .A(_tmp_846[22:19]), .Y(_09842_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33558_ ( .A(_tmp_846[18:15]), .Y(_09843_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33559_ ( .A({ _tmp_846[30], _tmp_846[27], _tmp_846[25:24] }), .Y(_09844_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33560_ ( .A({ _09833_, _05652_, _tmp_835 }), .Y(_05669_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33561_ ( .A({ _09834_, _tmp_846[0], _05652_, _tmp_835 }), .Y(_05670_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _33562_ ( .A({ _maxi_read_start, _09608_, _maxi_read_op_sel[0], _maxi_read_op_sel[1] }), .Y(_05671_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33563_ ( .A({ _05671_, _09591_ }), .Y(_05672_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33564_ ( .A({ _dataflow__delay_valid_132, _09590_ }), .Y(_05379_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33565_ ( .A({ _09845_, _05379_ }), .Y(_05673_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33566_ ( .A({ _tmp_12[0], _09592_, _tmp_12[33:32] }), .Y(_09845_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33567_ ( .A({ _stream_conv2d_8_source_6_source_ram_renable, _05014_ }), .Y(_tmp_336) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33568_ ( .A({ _stream_matmul_15_source_6_source_ram_renable, _05015_ }), .Y(_tmp_992) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33569_ ( .A({ _09846_, _05099_ }), .Y(_05675_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33570_ ( .A({ _09856_, _09851_, _09849_, _09847_ }), .Y(_09846_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33571_ ( .A({ _09848_, _source_stream_conv2d_8_source_6_pat_count_0[32:30] }), .Y(_09847_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33572_ ( .A({ _source_stream_conv2d_8_source_6_pat_count_0[28:27], _source_stream_conv2d_8_source_6_pat_count_0[25], _source_stream_conv2d_8_source_6_pat_count_0[22] }), .Y(_09848_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33573_ ( .A({ _09850_, _source_stream_conv2d_8_source_6_pat_count_0[1:0] }), .Y(_09849_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33574_ ( .A(_source_stream_conv2d_8_source_6_pat_count_0[5:2]), .Y(_09850_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33575_ ( .A({ _09855_, _09854_, _09853_, _09852_ }), .Y(_09851_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33576_ ( .A(_source_stream_conv2d_8_source_6_pat_count_0[13:10]), .Y(_09852_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33577_ ( .A(_source_stream_conv2d_8_source_6_pat_count_0[9:6]), .Y(_09853_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33578_ ( .A(_source_stream_conv2d_8_source_6_pat_count_0[21:18]), .Y(_09854_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33579_ ( .A(_source_stream_conv2d_8_source_6_pat_count_0[17:14]), .Y(_09855_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33580_ ( .A({ _source_stream_conv2d_8_source_6_pat_count_0[29], _source_stream_conv2d_8_source_6_pat_count_0[26], _source_stream_conv2d_8_source_6_pat_count_0[24:23] }), .Y(_09856_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33581_ ( .A({ _09857_, _05675_ }), .Y(_05676_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33582_ ( .A({ _09867_, _09865_, _09858_ }), .Y(_09857_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33583_ ( .A({ _09864_, _09859_, _source_stream_conv2d_8_source_6_pat_count_1[1:0] }), .Y(_09858_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33584_ ( .A({ _09863_, _09862_, _09861_, _09860_ }), .Y(_09859_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33585_ ( .A(_source_stream_conv2d_8_source_6_pat_count_1[13:10]), .Y(_09860_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33586_ ( .A(_source_stream_conv2d_8_source_6_pat_count_1[9:6]), .Y(_09861_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33587_ ( .A(_source_stream_conv2d_8_source_6_pat_count_1[21:18]), .Y(_09862_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33588_ ( .A(_source_stream_conv2d_8_source_6_pat_count_1[17:14]), .Y(_09863_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33589_ ( .A(_source_stream_conv2d_8_source_6_pat_count_1[5:2]), .Y(_09864_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33590_ ( .A({ _09866_, _source_stream_conv2d_8_source_6_pat_count_1[32:30] }), .Y(_09865_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33591_ ( .A({ _source_stream_conv2d_8_source_6_pat_count_1[28:27], _source_stream_conv2d_8_source_6_pat_count_1[25], _source_stream_conv2d_8_source_6_pat_count_1[22] }), .Y(_09866_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33592_ ( .A({ _source_stream_conv2d_8_source_6_pat_count_1[29], _source_stream_conv2d_8_source_6_pat_count_1[26], _source_stream_conv2d_8_source_6_pat_count_1[24:23] }), .Y(_09867_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33593_ ( .A({ _09868_, _09857_, _05675_ }), .Y(_05677_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33594_ ( .A({ _09878_, _09873_, _09871_, _09869_ }), .Y(_09868_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33595_ ( .A({ _09870_, _source_stream_conv2d_8_source_6_pat_count_2[32:30] }), .Y(_09869_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33596_ ( .A({ _source_stream_conv2d_8_source_6_pat_count_2[28:27], _source_stream_conv2d_8_source_6_pat_count_2[25], _source_stream_conv2d_8_source_6_pat_count_2[22] }), .Y(_09870_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33597_ ( .A({ _09872_, _source_stream_conv2d_8_source_6_pat_count_2[1:0] }), .Y(_09871_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33598_ ( .A(_source_stream_conv2d_8_source_6_pat_count_2[5:2]), .Y(_09872_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33599_ ( .A({ _09877_, _09876_, _09875_, _09874_ }), .Y(_09873_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33600_ ( .A(_source_stream_conv2d_8_source_6_pat_count_2[13:10]), .Y(_09874_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33601_ ( .A(_source_stream_conv2d_8_source_6_pat_count_2[9:6]), .Y(_09875_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33602_ ( .A(_source_stream_conv2d_8_source_6_pat_count_2[21:18]), .Y(_09876_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33603_ ( .A(_source_stream_conv2d_8_source_6_pat_count_2[17:14]), .Y(_09877_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33604_ ( .A({ _source_stream_conv2d_8_source_6_pat_count_2[29], _source_stream_conv2d_8_source_6_pat_count_2[26], _source_stream_conv2d_8_source_6_pat_count_2[24:23] }), .Y(_09878_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33605_ ( .A({ _05826_, _05099_ }), .Y(_05678_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33606_ ( .A({ _09879_, _09868_, _09846_, _09857_ }), .Y(_05826_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33607_ ( .A({ _09889_, _09884_, _09882_, _09880_ }), .Y(_09879_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33608_ ( .A({ _09881_, _source_stream_conv2d_8_source_6_pat_count_3[32:30] }), .Y(_09880_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33609_ ( .A({ _source_stream_conv2d_8_source_6_pat_count_3[28:27], _source_stream_conv2d_8_source_6_pat_count_3[25], _source_stream_conv2d_8_source_6_pat_count_3[22] }), .Y(_09881_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33610_ ( .A({ _09883_, _source_stream_conv2d_8_source_6_pat_count_3[1:0] }), .Y(_09882_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33611_ ( .A(_source_stream_conv2d_8_source_6_pat_count_3[5:2]), .Y(_09883_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33612_ ( .A({ _09888_, _09887_, _09886_, _09885_ }), .Y(_09884_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33613_ ( .A(_source_stream_conv2d_8_source_6_pat_count_3[13:10]), .Y(_09885_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33614_ ( .A(_source_stream_conv2d_8_source_6_pat_count_3[9:6]), .Y(_09886_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33615_ ( .A(_source_stream_conv2d_8_source_6_pat_count_3[21:18]), .Y(_09887_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33616_ ( .A(_source_stream_conv2d_8_source_6_pat_count_3[17:14]), .Y(_09888_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33617_ ( .A({ _source_stream_conv2d_8_source_6_pat_count_3[29], _source_stream_conv2d_8_source_6_pat_count_3[26], _source_stream_conv2d_8_source_6_pat_count_3[24:23] }), .Y(_09889_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33618_ ( .A({ _09890_, _05097_ }), .Y(_05680_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33619_ ( .A({ _09900_, _09895_, _09893_, _09891_ }), .Y(_09890_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33620_ ( .A({ _09892_, _source_stream_conv2d_8_source_8_pat_count_0[32:30] }), .Y(_09891_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33621_ ( .A({ _source_stream_conv2d_8_source_8_pat_count_0[28:27], _source_stream_conv2d_8_source_8_pat_count_0[25], _source_stream_conv2d_8_source_8_pat_count_0[22] }), .Y(_09892_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33622_ ( .A({ _09894_, _source_stream_conv2d_8_source_8_pat_count_0[1:0] }), .Y(_09893_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33623_ ( .A(_source_stream_conv2d_8_source_8_pat_count_0[5:2]), .Y(_09894_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33624_ ( .A({ _09899_, _09898_, _09897_, _09896_ }), .Y(_09895_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33625_ ( .A(_source_stream_conv2d_8_source_8_pat_count_0[13:10]), .Y(_09896_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33626_ ( .A(_source_stream_conv2d_8_source_8_pat_count_0[9:6]), .Y(_09897_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33627_ ( .A(_source_stream_conv2d_8_source_8_pat_count_0[21:18]), .Y(_09898_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33628_ ( .A(_source_stream_conv2d_8_source_8_pat_count_0[17:14]), .Y(_09899_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33629_ ( .A({ _source_stream_conv2d_8_source_8_pat_count_0[29], _source_stream_conv2d_8_source_8_pat_count_0[26], _source_stream_conv2d_8_source_8_pat_count_0[24:23] }), .Y(_09900_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33630_ ( .A({ _09901_, _05680_ }), .Y(_05681_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33631_ ( .A({ _09911_, _09909_, _09902_ }), .Y(_09901_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33632_ ( .A({ _09908_, _09903_, _source_stream_conv2d_8_source_8_pat_count_1[1:0] }), .Y(_09902_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33633_ ( .A({ _09907_, _09906_, _09905_, _09904_ }), .Y(_09903_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33634_ ( .A(_source_stream_conv2d_8_source_8_pat_count_1[13:10]), .Y(_09904_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33635_ ( .A(_source_stream_conv2d_8_source_8_pat_count_1[9:6]), .Y(_09905_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33636_ ( .A(_source_stream_conv2d_8_source_8_pat_count_1[21:18]), .Y(_09906_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33637_ ( .A(_source_stream_conv2d_8_source_8_pat_count_1[17:14]), .Y(_09907_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33638_ ( .A(_source_stream_conv2d_8_source_8_pat_count_1[5:2]), .Y(_09908_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33639_ ( .A({ _09910_, _source_stream_conv2d_8_source_8_pat_count_1[32:30] }), .Y(_09909_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33640_ ( .A({ _source_stream_conv2d_8_source_8_pat_count_1[28:27], _source_stream_conv2d_8_source_8_pat_count_1[25], _source_stream_conv2d_8_source_8_pat_count_1[22] }), .Y(_09910_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33641_ ( .A({ _source_stream_conv2d_8_source_8_pat_count_1[29], _source_stream_conv2d_8_source_8_pat_count_1[26], _source_stream_conv2d_8_source_8_pat_count_1[24:23] }), .Y(_09911_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33642_ ( .A({ _09890_, _09912_, _05097_ }), .Y(_05682_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33643_ ( .A({ _09913_, _09901_ }), .Y(_09912_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33644_ ( .A({ _09923_, _09918_, _09916_, _09914_ }), .Y(_09913_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33645_ ( .A({ _09915_, _source_stream_conv2d_8_source_8_pat_count_2[32:30] }), .Y(_09914_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33646_ ( .A({ _source_stream_conv2d_8_source_8_pat_count_2[28:27], _source_stream_conv2d_8_source_8_pat_count_2[25], _source_stream_conv2d_8_source_8_pat_count_2[22] }), .Y(_09915_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33647_ ( .A({ _09917_, _source_stream_conv2d_8_source_8_pat_count_2[1:0] }), .Y(_09916_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33648_ ( .A(_source_stream_conv2d_8_source_8_pat_count_2[5:2]), .Y(_09917_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33649_ ( .A({ _09922_, _09921_, _09920_, _09919_ }), .Y(_09918_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33650_ ( .A(_source_stream_conv2d_8_source_8_pat_count_2[13:10]), .Y(_09919_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33651_ ( .A(_source_stream_conv2d_8_source_8_pat_count_2[9:6]), .Y(_09920_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33652_ ( .A(_source_stream_conv2d_8_source_8_pat_count_2[21:18]), .Y(_09921_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33653_ ( .A(_source_stream_conv2d_8_source_8_pat_count_2[17:14]), .Y(_09922_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33654_ ( .A({ _source_stream_conv2d_8_source_8_pat_count_2[29], _source_stream_conv2d_8_source_8_pat_count_2[26], _source_stream_conv2d_8_source_8_pat_count_2[24:23] }), .Y(_09923_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33655_ ( .A({ _09924_, _05682_ }), .Y(_05683_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33656_ ( .A({ _09934_, _09932_, _09925_ }), .Y(_09924_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33657_ ( .A({ _09931_, _09926_, _source_stream_conv2d_8_source_8_pat_count_3[1:0] }), .Y(_09925_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33658_ ( .A({ _09930_, _09929_, _09928_, _09927_ }), .Y(_09926_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33659_ ( .A(_source_stream_conv2d_8_source_8_pat_count_3[13:10]), .Y(_09927_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33660_ ( .A(_source_stream_conv2d_8_source_8_pat_count_3[9:6]), .Y(_09928_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33661_ ( .A(_source_stream_conv2d_8_source_8_pat_count_3[21:18]), .Y(_09929_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33662_ ( .A(_source_stream_conv2d_8_source_8_pat_count_3[17:14]), .Y(_09930_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33663_ ( .A(_source_stream_conv2d_8_source_8_pat_count_3[5:2]), .Y(_09931_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33664_ ( .A({ _09933_, _source_stream_conv2d_8_source_8_pat_count_3[32:30] }), .Y(_09932_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33665_ ( .A({ _source_stream_conv2d_8_source_8_pat_count_3[28:27], _source_stream_conv2d_8_source_8_pat_count_3[25], _source_stream_conv2d_8_source_8_pat_count_3[22] }), .Y(_09933_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33666_ ( .A({ _source_stream_conv2d_8_source_8_pat_count_3[29], _source_stream_conv2d_8_source_8_pat_count_3[26], _source_stream_conv2d_8_source_8_pat_count_3[24:23] }), .Y(_09934_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33667_ ( .A({ _09935_, _05095_ }), .Y(_05685_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33668_ ( .A({ _09945_, _09940_, _09938_, _09936_ }), .Y(_09935_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33669_ ( .A({ _09937_, _source_stream_conv2d_8_source_19_pat_count_0[32:30] }), .Y(_09936_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33670_ ( .A({ _source_stream_conv2d_8_source_19_pat_count_0[28:27], _source_stream_conv2d_8_source_19_pat_count_0[25], _source_stream_conv2d_8_source_19_pat_count_0[22] }), .Y(_09937_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33671_ ( .A({ _09939_, _source_stream_conv2d_8_source_19_pat_count_0[1:0] }), .Y(_09938_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33672_ ( .A(_source_stream_conv2d_8_source_19_pat_count_0[5:2]), .Y(_09939_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33673_ ( .A({ _09944_, _09943_, _09942_, _09941_ }), .Y(_09940_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33674_ ( .A(_source_stream_conv2d_8_source_19_pat_count_0[13:10]), .Y(_09941_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33675_ ( .A(_source_stream_conv2d_8_source_19_pat_count_0[9:6]), .Y(_09942_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33676_ ( .A(_source_stream_conv2d_8_source_19_pat_count_0[21:18]), .Y(_09943_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33677_ ( .A(_source_stream_conv2d_8_source_19_pat_count_0[17:14]), .Y(_09944_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33678_ ( .A({ _source_stream_conv2d_8_source_19_pat_count_0[29], _source_stream_conv2d_8_source_19_pat_count_0[26], _source_stream_conv2d_8_source_19_pat_count_0[24:23] }), .Y(_09945_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33679_ ( .A({ _09946_, _05685_ }), .Y(_05686_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33680_ ( .A({ _09956_, _09954_, _09947_ }), .Y(_09946_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33681_ ( .A({ _09953_, _09948_, _source_stream_conv2d_8_source_19_pat_count_1[1:0] }), .Y(_09947_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33682_ ( .A({ _09952_, _09951_, _09950_, _09949_ }), .Y(_09948_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33683_ ( .A(_source_stream_conv2d_8_source_19_pat_count_1[13:10]), .Y(_09949_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33684_ ( .A(_source_stream_conv2d_8_source_19_pat_count_1[9:6]), .Y(_09950_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33685_ ( .A(_source_stream_conv2d_8_source_19_pat_count_1[21:18]), .Y(_09951_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33686_ ( .A(_source_stream_conv2d_8_source_19_pat_count_1[17:14]), .Y(_09952_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33687_ ( .A(_source_stream_conv2d_8_source_19_pat_count_1[5:2]), .Y(_09953_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33688_ ( .A({ _09955_, _source_stream_conv2d_8_source_19_pat_count_1[32:30] }), .Y(_09954_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33689_ ( .A({ _source_stream_conv2d_8_source_19_pat_count_1[28:27], _source_stream_conv2d_8_source_19_pat_count_1[25], _source_stream_conv2d_8_source_19_pat_count_1[22] }), .Y(_09955_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33690_ ( .A({ _source_stream_conv2d_8_source_19_pat_count_1[29], _source_stream_conv2d_8_source_19_pat_count_1[26], _source_stream_conv2d_8_source_19_pat_count_1[24:23] }), .Y(_09956_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33691_ ( .A({ _09935_, _09957_, _05095_ }), .Y(_05687_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33692_ ( .A({ _09958_, _09946_ }), .Y(_09957_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33693_ ( .A({ _09968_, _09963_, _09961_, _09959_ }), .Y(_09958_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33694_ ( .A({ _09960_, _source_stream_conv2d_8_source_19_pat_count_2[32:30] }), .Y(_09959_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33695_ ( .A({ _source_stream_conv2d_8_source_19_pat_count_2[28:27], _source_stream_conv2d_8_source_19_pat_count_2[25], _source_stream_conv2d_8_source_19_pat_count_2[22] }), .Y(_09960_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33696_ ( .A({ _09962_, _source_stream_conv2d_8_source_19_pat_count_2[1:0] }), .Y(_09961_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33697_ ( .A(_source_stream_conv2d_8_source_19_pat_count_2[5:2]), .Y(_09962_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33698_ ( .A({ _09967_, _09966_, _09965_, _09964_ }), .Y(_09963_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33699_ ( .A(_source_stream_conv2d_8_source_19_pat_count_2[13:10]), .Y(_09964_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33700_ ( .A(_source_stream_conv2d_8_source_19_pat_count_2[9:6]), .Y(_09965_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33701_ ( .A(_source_stream_conv2d_8_source_19_pat_count_2[21:18]), .Y(_09966_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33702_ ( .A(_source_stream_conv2d_8_source_19_pat_count_2[17:14]), .Y(_09967_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33703_ ( .A({ _source_stream_conv2d_8_source_19_pat_count_2[29], _source_stream_conv2d_8_source_19_pat_count_2[26], _source_stream_conv2d_8_source_19_pat_count_2[24:23] }), .Y(_09968_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33704_ ( .A({ _09969_, _05687_ }), .Y(_05688_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33705_ ( .A({ _09979_, _09977_, _09970_ }), .Y(_09969_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33706_ ( .A({ _09976_, _09971_, _source_stream_conv2d_8_source_19_pat_count_3[1:0] }), .Y(_09970_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33707_ ( .A({ _09975_, _09974_, _09973_, _09972_ }), .Y(_09971_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33708_ ( .A(_source_stream_conv2d_8_source_19_pat_count_3[13:10]), .Y(_09972_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33709_ ( .A(_source_stream_conv2d_8_source_19_pat_count_3[9:6]), .Y(_09973_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33710_ ( .A(_source_stream_conv2d_8_source_19_pat_count_3[21:18]), .Y(_09974_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33711_ ( .A(_source_stream_conv2d_8_source_19_pat_count_3[17:14]), .Y(_09975_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33712_ ( .A(_source_stream_conv2d_8_source_19_pat_count_3[5:2]), .Y(_09976_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33713_ ( .A({ _09978_, _source_stream_conv2d_8_source_19_pat_count_3[32:30] }), .Y(_09977_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33714_ ( .A({ _source_stream_conv2d_8_source_19_pat_count_3[28:27], _source_stream_conv2d_8_source_19_pat_count_3[25], _source_stream_conv2d_8_source_19_pat_count_3[22] }), .Y(_09978_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33715_ ( .A({ _source_stream_conv2d_8_source_19_pat_count_3[29], _source_stream_conv2d_8_source_19_pat_count_3[26], _source_stream_conv2d_8_source_19_pat_count_3[24:23] }), .Y(_09979_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33716_ ( .A({ _09980_, _05093_ }), .Y(_05690_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33717_ ( .A({ _09990_, _09985_, _09983_, _09981_ }), .Y(_09980_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33718_ ( .A({ _09982_, _source_stream_conv2d_8_source_20_pat_count_0[32:30] }), .Y(_09981_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33719_ ( .A({ _source_stream_conv2d_8_source_20_pat_count_0[28:27], _source_stream_conv2d_8_source_20_pat_count_0[25], _source_stream_conv2d_8_source_20_pat_count_0[22] }), .Y(_09982_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33720_ ( .A({ _09984_, _source_stream_conv2d_8_source_20_pat_count_0[1:0] }), .Y(_09983_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33721_ ( .A(_source_stream_conv2d_8_source_20_pat_count_0[5:2]), .Y(_09984_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33722_ ( .A({ _09989_, _09988_, _09987_, _09986_ }), .Y(_09985_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33723_ ( .A(_source_stream_conv2d_8_source_20_pat_count_0[13:10]), .Y(_09986_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33724_ ( .A(_source_stream_conv2d_8_source_20_pat_count_0[9:6]), .Y(_09987_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33725_ ( .A(_source_stream_conv2d_8_source_20_pat_count_0[21:18]), .Y(_09988_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33726_ ( .A(_source_stream_conv2d_8_source_20_pat_count_0[17:14]), .Y(_09989_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33727_ ( .A({ _source_stream_conv2d_8_source_20_pat_count_0[29], _source_stream_conv2d_8_source_20_pat_count_0[26], _source_stream_conv2d_8_source_20_pat_count_0[24:23] }), .Y(_09990_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33728_ ( .A({ _09991_, _05690_ }), .Y(_05691_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33729_ ( .A({ _10001_, _09999_, _09992_ }), .Y(_09991_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33730_ ( .A({ _09998_, _09993_, _source_stream_conv2d_8_source_20_pat_count_1[1:0] }), .Y(_09992_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33731_ ( .A({ _09997_, _09996_, _09995_, _09994_ }), .Y(_09993_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33732_ ( .A(_source_stream_conv2d_8_source_20_pat_count_1[13:10]), .Y(_09994_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33733_ ( .A(_source_stream_conv2d_8_source_20_pat_count_1[9:6]), .Y(_09995_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33734_ ( .A(_source_stream_conv2d_8_source_20_pat_count_1[21:18]), .Y(_09996_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33735_ ( .A(_source_stream_conv2d_8_source_20_pat_count_1[17:14]), .Y(_09997_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33736_ ( .A(_source_stream_conv2d_8_source_20_pat_count_1[5:2]), .Y(_09998_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33737_ ( .A({ _10000_, _source_stream_conv2d_8_source_20_pat_count_1[32:30] }), .Y(_09999_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33738_ ( .A({ _source_stream_conv2d_8_source_20_pat_count_1[28:27], _source_stream_conv2d_8_source_20_pat_count_1[25], _source_stream_conv2d_8_source_20_pat_count_1[22] }), .Y(_10000_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33739_ ( .A({ _source_stream_conv2d_8_source_20_pat_count_1[29], _source_stream_conv2d_8_source_20_pat_count_1[26], _source_stream_conv2d_8_source_20_pat_count_1[24:23] }), .Y(_10001_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33740_ ( .A({ _10002_, _09991_, _05690_ }), .Y(_05692_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33741_ ( .A({ _10012_, _10007_, _10005_, _10003_ }), .Y(_10002_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33742_ ( .A({ _10004_, _source_stream_conv2d_8_source_20_pat_count_2[32:30] }), .Y(_10003_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33743_ ( .A({ _source_stream_conv2d_8_source_20_pat_count_2[28:27], _source_stream_conv2d_8_source_20_pat_count_2[25], _source_stream_conv2d_8_source_20_pat_count_2[22] }), .Y(_10004_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33744_ ( .A({ _10006_, _source_stream_conv2d_8_source_20_pat_count_2[1:0] }), .Y(_10005_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33745_ ( .A(_source_stream_conv2d_8_source_20_pat_count_2[5:2]), .Y(_10006_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33746_ ( .A({ _10011_, _10010_, _10009_, _10008_ }), .Y(_10007_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33747_ ( .A(_source_stream_conv2d_8_source_20_pat_count_2[13:10]), .Y(_10008_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33748_ ( .A(_source_stream_conv2d_8_source_20_pat_count_2[9:6]), .Y(_10009_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33749_ ( .A(_source_stream_conv2d_8_source_20_pat_count_2[21:18]), .Y(_10010_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33750_ ( .A(_source_stream_conv2d_8_source_20_pat_count_2[17:14]), .Y(_10011_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33751_ ( .A({ _source_stream_conv2d_8_source_20_pat_count_2[29], _source_stream_conv2d_8_source_20_pat_count_2[26], _source_stream_conv2d_8_source_20_pat_count_2[24:23] }), .Y(_10012_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33752_ ( .A({ _05829_, _05093_ }), .Y(_05693_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33753_ ( .A({ _10013_, _10002_, _09980_, _09991_ }), .Y(_05829_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33754_ ( .A({ _10023_, _10018_, _10016_, _10014_ }), .Y(_10013_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33755_ ( .A({ _10015_, _source_stream_conv2d_8_source_20_pat_count_3[32:30] }), .Y(_10014_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33756_ ( .A({ _source_stream_conv2d_8_source_20_pat_count_3[28:27], _source_stream_conv2d_8_source_20_pat_count_3[25], _source_stream_conv2d_8_source_20_pat_count_3[22] }), .Y(_10015_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33757_ ( .A({ _10017_, _source_stream_conv2d_8_source_20_pat_count_3[1:0] }), .Y(_10016_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33758_ ( .A(_source_stream_conv2d_8_source_20_pat_count_3[5:2]), .Y(_10017_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33759_ ( .A({ _10022_, _10021_, _10020_, _10019_ }), .Y(_10018_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33760_ ( .A(_source_stream_conv2d_8_source_20_pat_count_3[13:10]), .Y(_10019_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33761_ ( .A(_source_stream_conv2d_8_source_20_pat_count_3[9:6]), .Y(_10020_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33762_ ( .A(_source_stream_conv2d_8_source_20_pat_count_3[21:18]), .Y(_10021_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33763_ ( .A(_source_stream_conv2d_8_source_20_pat_count_3[17:14]), .Y(_10022_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33764_ ( .A({ _source_stream_conv2d_8_source_20_pat_count_3[29], _source_stream_conv2d_8_source_20_pat_count_3[26], _source_stream_conv2d_8_source_20_pat_count_3[24:23] }), .Y(_10023_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33765_ ( .A({ _10024_, _05091_ }), .Y(_05695_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33766_ ( .A({ _10034_, _10029_, _10027_, _10025_ }), .Y(_10024_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33767_ ( .A({ _10026_, _source_stream_conv2d_8_source_21_pat_count_0[32:30] }), .Y(_10025_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33768_ ( .A({ _source_stream_conv2d_8_source_21_pat_count_0[28:27], _source_stream_conv2d_8_source_21_pat_count_0[25], _source_stream_conv2d_8_source_21_pat_count_0[22] }), .Y(_10026_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33769_ ( .A({ _10028_, _source_stream_conv2d_8_source_21_pat_count_0[1:0] }), .Y(_10027_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33770_ ( .A(_source_stream_conv2d_8_source_21_pat_count_0[5:2]), .Y(_10028_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33771_ ( .A({ _10033_, _10032_, _10031_, _10030_ }), .Y(_10029_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33772_ ( .A(_source_stream_conv2d_8_source_21_pat_count_0[13:10]), .Y(_10030_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33773_ ( .A(_source_stream_conv2d_8_source_21_pat_count_0[9:6]), .Y(_10031_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33774_ ( .A(_source_stream_conv2d_8_source_21_pat_count_0[21:18]), .Y(_10032_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33775_ ( .A(_source_stream_conv2d_8_source_21_pat_count_0[17:14]), .Y(_10033_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33776_ ( .A({ _source_stream_conv2d_8_source_21_pat_count_0[29], _source_stream_conv2d_8_source_21_pat_count_0[26], _source_stream_conv2d_8_source_21_pat_count_0[24:23] }), .Y(_10034_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33777_ ( .A({ _10035_, _05695_ }), .Y(_05696_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33778_ ( .A({ _10045_, _10043_, _10036_ }), .Y(_10035_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33779_ ( .A({ _10042_, _10037_, _source_stream_conv2d_8_source_21_pat_count_1[1:0] }), .Y(_10036_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33780_ ( .A({ _10041_, _10040_, _10039_, _10038_ }), .Y(_10037_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33781_ ( .A(_source_stream_conv2d_8_source_21_pat_count_1[13:10]), .Y(_10038_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33782_ ( .A(_source_stream_conv2d_8_source_21_pat_count_1[9:6]), .Y(_10039_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33783_ ( .A(_source_stream_conv2d_8_source_21_pat_count_1[21:18]), .Y(_10040_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33784_ ( .A(_source_stream_conv2d_8_source_21_pat_count_1[17:14]), .Y(_10041_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33785_ ( .A(_source_stream_conv2d_8_source_21_pat_count_1[5:2]), .Y(_10042_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33786_ ( .A({ _10044_, _source_stream_conv2d_8_source_21_pat_count_1[32:30] }), .Y(_10043_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33787_ ( .A({ _source_stream_conv2d_8_source_21_pat_count_1[28:27], _source_stream_conv2d_8_source_21_pat_count_1[25], _source_stream_conv2d_8_source_21_pat_count_1[22] }), .Y(_10044_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33788_ ( .A({ _source_stream_conv2d_8_source_21_pat_count_1[29], _source_stream_conv2d_8_source_21_pat_count_1[26], _source_stream_conv2d_8_source_21_pat_count_1[24:23] }), .Y(_10045_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33789_ ( .A({ _10046_, _10035_, _05695_ }), .Y(_05697_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33790_ ( .A({ _10056_, _10051_, _10049_, _10047_ }), .Y(_10046_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33791_ ( .A({ _10048_, _source_stream_conv2d_8_source_21_pat_count_2[32:30] }), .Y(_10047_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33792_ ( .A({ _source_stream_conv2d_8_source_21_pat_count_2[28:27], _source_stream_conv2d_8_source_21_pat_count_2[25], _source_stream_conv2d_8_source_21_pat_count_2[22] }), .Y(_10048_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33793_ ( .A({ _10050_, _source_stream_conv2d_8_source_21_pat_count_2[1:0] }), .Y(_10049_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33794_ ( .A(_source_stream_conv2d_8_source_21_pat_count_2[5:2]), .Y(_10050_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33795_ ( .A({ _10055_, _10054_, _10053_, _10052_ }), .Y(_10051_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33796_ ( .A(_source_stream_conv2d_8_source_21_pat_count_2[13:10]), .Y(_10052_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33797_ ( .A(_source_stream_conv2d_8_source_21_pat_count_2[9:6]), .Y(_10053_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33798_ ( .A(_source_stream_conv2d_8_source_21_pat_count_2[21:18]), .Y(_10054_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33799_ ( .A(_source_stream_conv2d_8_source_21_pat_count_2[17:14]), .Y(_10055_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33800_ ( .A({ _source_stream_conv2d_8_source_21_pat_count_2[29], _source_stream_conv2d_8_source_21_pat_count_2[26], _source_stream_conv2d_8_source_21_pat_count_2[24:23] }), .Y(_10056_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33801_ ( .A({ _05830_, _05091_ }), .Y(_05698_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33802_ ( .A({ _10057_, _10046_, _10024_, _10035_ }), .Y(_05830_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33803_ ( .A({ _10067_, _10062_, _10060_, _10058_ }), .Y(_10057_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33804_ ( .A({ _10059_, _source_stream_conv2d_8_source_21_pat_count_3[32:30] }), .Y(_10058_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33805_ ( .A({ _source_stream_conv2d_8_source_21_pat_count_3[28:27], _source_stream_conv2d_8_source_21_pat_count_3[25], _source_stream_conv2d_8_source_21_pat_count_3[22] }), .Y(_10059_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33806_ ( .A({ _10061_, _source_stream_conv2d_8_source_21_pat_count_3[1:0] }), .Y(_10060_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33807_ ( .A(_source_stream_conv2d_8_source_21_pat_count_3[5:2]), .Y(_10061_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33808_ ( .A({ _10066_, _10065_, _10064_, _10063_ }), .Y(_10062_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33809_ ( .A(_source_stream_conv2d_8_source_21_pat_count_3[13:10]), .Y(_10063_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33810_ ( .A(_source_stream_conv2d_8_source_21_pat_count_3[9:6]), .Y(_10064_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33811_ ( .A(_source_stream_conv2d_8_source_21_pat_count_3[21:18]), .Y(_10065_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33812_ ( .A(_source_stream_conv2d_8_source_21_pat_count_3[17:14]), .Y(_10066_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33813_ ( .A({ _source_stream_conv2d_8_source_21_pat_count_3[29], _source_stream_conv2d_8_source_21_pat_count_3[26], _source_stream_conv2d_8_source_21_pat_count_3[24:23] }), .Y(_10067_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33814_ ( .A({ _10068_, _05089_ }), .Y(_05700_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33815_ ( .A({ _10078_, _10073_, _10071_, _10069_ }), .Y(_10068_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33816_ ( .A({ _10070_, _source_stream_conv2d_8_source_22_pat_count_0[32:30] }), .Y(_10069_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33817_ ( .A({ _source_stream_conv2d_8_source_22_pat_count_0[28:27], _source_stream_conv2d_8_source_22_pat_count_0[25], _source_stream_conv2d_8_source_22_pat_count_0[22] }), .Y(_10070_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33818_ ( .A({ _10072_, _source_stream_conv2d_8_source_22_pat_count_0[1:0] }), .Y(_10071_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33819_ ( .A(_source_stream_conv2d_8_source_22_pat_count_0[5:2]), .Y(_10072_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33820_ ( .A({ _10077_, _10076_, _10075_, _10074_ }), .Y(_10073_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33821_ ( .A(_source_stream_conv2d_8_source_22_pat_count_0[13:10]), .Y(_10074_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33822_ ( .A(_source_stream_conv2d_8_source_22_pat_count_0[9:6]), .Y(_10075_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33823_ ( .A(_source_stream_conv2d_8_source_22_pat_count_0[21:18]), .Y(_10076_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33824_ ( .A(_source_stream_conv2d_8_source_22_pat_count_0[17:14]), .Y(_10077_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33825_ ( .A({ _source_stream_conv2d_8_source_22_pat_count_0[29], _source_stream_conv2d_8_source_22_pat_count_0[26], _source_stream_conv2d_8_source_22_pat_count_0[24:23] }), .Y(_10078_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33826_ ( .A({ _10079_, _05700_ }), .Y(_05701_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33827_ ( .A({ _10089_, _10087_, _10080_ }), .Y(_10079_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33828_ ( .A({ _10086_, _10081_, _source_stream_conv2d_8_source_22_pat_count_1[1:0] }), .Y(_10080_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33829_ ( .A({ _10085_, _10084_, _10083_, _10082_ }), .Y(_10081_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33830_ ( .A(_source_stream_conv2d_8_source_22_pat_count_1[13:10]), .Y(_10082_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33831_ ( .A(_source_stream_conv2d_8_source_22_pat_count_1[9:6]), .Y(_10083_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33832_ ( .A(_source_stream_conv2d_8_source_22_pat_count_1[21:18]), .Y(_10084_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33833_ ( .A(_source_stream_conv2d_8_source_22_pat_count_1[17:14]), .Y(_10085_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33834_ ( .A(_source_stream_conv2d_8_source_22_pat_count_1[5:2]), .Y(_10086_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33835_ ( .A({ _10088_, _source_stream_conv2d_8_source_22_pat_count_1[32:30] }), .Y(_10087_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33836_ ( .A({ _source_stream_conv2d_8_source_22_pat_count_1[28:27], _source_stream_conv2d_8_source_22_pat_count_1[25], _source_stream_conv2d_8_source_22_pat_count_1[22] }), .Y(_10088_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33837_ ( .A({ _source_stream_conv2d_8_source_22_pat_count_1[29], _source_stream_conv2d_8_source_22_pat_count_1[26], _source_stream_conv2d_8_source_22_pat_count_1[24:23] }), .Y(_10089_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33838_ ( .A({ _10090_, _10079_, _05700_ }), .Y(_05702_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33839_ ( .A({ _10100_, _10095_, _10093_, _10091_ }), .Y(_10090_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33840_ ( .A({ _10092_, _source_stream_conv2d_8_source_22_pat_count_2[32:30] }), .Y(_10091_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33841_ ( .A({ _source_stream_conv2d_8_source_22_pat_count_2[28:27], _source_stream_conv2d_8_source_22_pat_count_2[25], _source_stream_conv2d_8_source_22_pat_count_2[22] }), .Y(_10092_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33842_ ( .A({ _10094_, _source_stream_conv2d_8_source_22_pat_count_2[1:0] }), .Y(_10093_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33843_ ( .A(_source_stream_conv2d_8_source_22_pat_count_2[5:2]), .Y(_10094_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33844_ ( .A({ _10099_, _10098_, _10097_, _10096_ }), .Y(_10095_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33845_ ( .A(_source_stream_conv2d_8_source_22_pat_count_2[13:10]), .Y(_10096_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33846_ ( .A(_source_stream_conv2d_8_source_22_pat_count_2[9:6]), .Y(_10097_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33847_ ( .A(_source_stream_conv2d_8_source_22_pat_count_2[21:18]), .Y(_10098_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33848_ ( .A(_source_stream_conv2d_8_source_22_pat_count_2[17:14]), .Y(_10099_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33849_ ( .A({ _source_stream_conv2d_8_source_22_pat_count_2[29], _source_stream_conv2d_8_source_22_pat_count_2[26], _source_stream_conv2d_8_source_22_pat_count_2[24:23] }), .Y(_10100_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33850_ ( .A({ _05831_, _05089_ }), .Y(_05703_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33851_ ( .A({ _10101_, _10090_, _10068_, _10079_ }), .Y(_05831_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33852_ ( .A({ _10111_, _10106_, _10104_, _10102_ }), .Y(_10101_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33853_ ( .A({ _10103_, _source_stream_conv2d_8_source_22_pat_count_3[32:30] }), .Y(_10102_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33854_ ( .A({ _source_stream_conv2d_8_source_22_pat_count_3[28:27], _source_stream_conv2d_8_source_22_pat_count_3[25], _source_stream_conv2d_8_source_22_pat_count_3[22] }), .Y(_10103_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33855_ ( .A({ _10105_, _source_stream_conv2d_8_source_22_pat_count_3[1:0] }), .Y(_10104_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33856_ ( .A(_source_stream_conv2d_8_source_22_pat_count_3[5:2]), .Y(_10105_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33857_ ( .A({ _10110_, _10109_, _10108_, _10107_ }), .Y(_10106_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33858_ ( .A(_source_stream_conv2d_8_source_22_pat_count_3[13:10]), .Y(_10107_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33859_ ( .A(_source_stream_conv2d_8_source_22_pat_count_3[9:6]), .Y(_10108_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33860_ ( .A(_source_stream_conv2d_8_source_22_pat_count_3[21:18]), .Y(_10109_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33861_ ( .A(_source_stream_conv2d_8_source_22_pat_count_3[17:14]), .Y(_10110_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33862_ ( .A({ _source_stream_conv2d_8_source_22_pat_count_3[29], _source_stream_conv2d_8_source_22_pat_count_3[26], _source_stream_conv2d_8_source_22_pat_count_3[24:23] }), .Y(_10111_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33863_ ( .A({ _10112_, _05087_ }), .Y(_05705_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33864_ ( .A({ _10122_, _10117_, _10115_, _10113_ }), .Y(_10112_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33865_ ( .A({ _10114_, _source_stream_conv2d_8_source_23_pat_count_0[32:30] }), .Y(_10113_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33866_ ( .A({ _source_stream_conv2d_8_source_23_pat_count_0[28:27], _source_stream_conv2d_8_source_23_pat_count_0[25], _source_stream_conv2d_8_source_23_pat_count_0[22] }), .Y(_10114_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33867_ ( .A({ _10116_, _source_stream_conv2d_8_source_23_pat_count_0[1:0] }), .Y(_10115_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33868_ ( .A(_source_stream_conv2d_8_source_23_pat_count_0[5:2]), .Y(_10116_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33869_ ( .A({ _10121_, _10120_, _10119_, _10118_ }), .Y(_10117_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33870_ ( .A(_source_stream_conv2d_8_source_23_pat_count_0[13:10]), .Y(_10118_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33871_ ( .A(_source_stream_conv2d_8_source_23_pat_count_0[9:6]), .Y(_10119_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33872_ ( .A(_source_stream_conv2d_8_source_23_pat_count_0[21:18]), .Y(_10120_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33873_ ( .A(_source_stream_conv2d_8_source_23_pat_count_0[17:14]), .Y(_10121_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33874_ ( .A({ _source_stream_conv2d_8_source_23_pat_count_0[29], _source_stream_conv2d_8_source_23_pat_count_0[26], _source_stream_conv2d_8_source_23_pat_count_0[24:23] }), .Y(_10122_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33875_ ( .A({ _10123_, _05705_ }), .Y(_05706_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33876_ ( .A({ _10133_, _10131_, _10124_ }), .Y(_10123_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33877_ ( .A({ _10130_, _10125_, _source_stream_conv2d_8_source_23_pat_count_1[1:0] }), .Y(_10124_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33878_ ( .A({ _10129_, _10128_, _10127_, _10126_ }), .Y(_10125_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33879_ ( .A(_source_stream_conv2d_8_source_23_pat_count_1[13:10]), .Y(_10126_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33880_ ( .A(_source_stream_conv2d_8_source_23_pat_count_1[9:6]), .Y(_10127_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33881_ ( .A(_source_stream_conv2d_8_source_23_pat_count_1[21:18]), .Y(_10128_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33882_ ( .A(_source_stream_conv2d_8_source_23_pat_count_1[17:14]), .Y(_10129_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33883_ ( .A(_source_stream_conv2d_8_source_23_pat_count_1[5:2]), .Y(_10130_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33884_ ( .A({ _10132_, _source_stream_conv2d_8_source_23_pat_count_1[32:30] }), .Y(_10131_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33885_ ( .A({ _source_stream_conv2d_8_source_23_pat_count_1[28:27], _source_stream_conv2d_8_source_23_pat_count_1[25], _source_stream_conv2d_8_source_23_pat_count_1[22] }), .Y(_10132_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33886_ ( .A({ _source_stream_conv2d_8_source_23_pat_count_1[29], _source_stream_conv2d_8_source_23_pat_count_1[26], _source_stream_conv2d_8_source_23_pat_count_1[24:23] }), .Y(_10133_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33887_ ( .A({ _10134_, _10123_, _05705_ }), .Y(_05707_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33888_ ( .A({ _10144_, _10139_, _10137_, _10135_ }), .Y(_10134_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33889_ ( .A({ _10136_, _source_stream_conv2d_8_source_23_pat_count_2[32:30] }), .Y(_10135_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33890_ ( .A({ _source_stream_conv2d_8_source_23_pat_count_2[28:27], _source_stream_conv2d_8_source_23_pat_count_2[25], _source_stream_conv2d_8_source_23_pat_count_2[22] }), .Y(_10136_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33891_ ( .A({ _10138_, _source_stream_conv2d_8_source_23_pat_count_2[1:0] }), .Y(_10137_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33892_ ( .A(_source_stream_conv2d_8_source_23_pat_count_2[5:2]), .Y(_10138_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33893_ ( .A({ _10143_, _10142_, _10141_, _10140_ }), .Y(_10139_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33894_ ( .A(_source_stream_conv2d_8_source_23_pat_count_2[13:10]), .Y(_10140_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33895_ ( .A(_source_stream_conv2d_8_source_23_pat_count_2[9:6]), .Y(_10141_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33896_ ( .A(_source_stream_conv2d_8_source_23_pat_count_2[21:18]), .Y(_10142_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33897_ ( .A(_source_stream_conv2d_8_source_23_pat_count_2[17:14]), .Y(_10143_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33898_ ( .A({ _source_stream_conv2d_8_source_23_pat_count_2[29], _source_stream_conv2d_8_source_23_pat_count_2[26], _source_stream_conv2d_8_source_23_pat_count_2[24:23] }), .Y(_10144_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33899_ ( .A({ _05832_, _05087_ }), .Y(_05708_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33900_ ( .A({ _10145_, _10134_, _10112_, _10123_ }), .Y(_05832_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33901_ ( .A({ _10155_, _10150_, _10148_, _10146_ }), .Y(_10145_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33902_ ( .A({ _10147_, _source_stream_conv2d_8_source_23_pat_count_3[32:30] }), .Y(_10146_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33903_ ( .A({ _source_stream_conv2d_8_source_23_pat_count_3[28:27], _source_stream_conv2d_8_source_23_pat_count_3[25], _source_stream_conv2d_8_source_23_pat_count_3[22] }), .Y(_10147_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33904_ ( .A({ _10149_, _source_stream_conv2d_8_source_23_pat_count_3[1:0] }), .Y(_10148_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33905_ ( .A(_source_stream_conv2d_8_source_23_pat_count_3[5:2]), .Y(_10149_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33906_ ( .A({ _10154_, _10153_, _10152_, _10151_ }), .Y(_10150_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33907_ ( .A(_source_stream_conv2d_8_source_23_pat_count_3[13:10]), .Y(_10151_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33908_ ( .A(_source_stream_conv2d_8_source_23_pat_count_3[9:6]), .Y(_10152_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33909_ ( .A(_source_stream_conv2d_8_source_23_pat_count_3[21:18]), .Y(_10153_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33910_ ( .A(_source_stream_conv2d_8_source_23_pat_count_3[17:14]), .Y(_10154_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33911_ ( .A({ _source_stream_conv2d_8_source_23_pat_count_3[29], _source_stream_conv2d_8_source_23_pat_count_3[26], _source_stream_conv2d_8_source_23_pat_count_3[24:23] }), .Y(_10155_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33912_ ( .A({ _10156_, _05085_ }), .Y(_05710_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33913_ ( .A({ _10166_, _10161_, _10159_, _10157_ }), .Y(_10156_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33914_ ( .A({ _10158_, _source_stream_conv2d_8_source_24_pat_count_0[32:30] }), .Y(_10157_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33915_ ( .A({ _source_stream_conv2d_8_source_24_pat_count_0[28:27], _source_stream_conv2d_8_source_24_pat_count_0[25], _source_stream_conv2d_8_source_24_pat_count_0[22] }), .Y(_10158_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33916_ ( .A({ _10160_, _source_stream_conv2d_8_source_24_pat_count_0[1:0] }), .Y(_10159_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33917_ ( .A(_source_stream_conv2d_8_source_24_pat_count_0[5:2]), .Y(_10160_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33918_ ( .A({ _10165_, _10164_, _10163_, _10162_ }), .Y(_10161_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33919_ ( .A(_source_stream_conv2d_8_source_24_pat_count_0[13:10]), .Y(_10162_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33920_ ( .A(_source_stream_conv2d_8_source_24_pat_count_0[9:6]), .Y(_10163_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33921_ ( .A(_source_stream_conv2d_8_source_24_pat_count_0[21:18]), .Y(_10164_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33922_ ( .A(_source_stream_conv2d_8_source_24_pat_count_0[17:14]), .Y(_10165_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33923_ ( .A({ _source_stream_conv2d_8_source_24_pat_count_0[29], _source_stream_conv2d_8_source_24_pat_count_0[26], _source_stream_conv2d_8_source_24_pat_count_0[24:23] }), .Y(_10166_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33924_ ( .A({ _10167_, _05710_ }), .Y(_05711_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33925_ ( .A({ _10177_, _10175_, _10168_ }), .Y(_10167_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33926_ ( .A({ _10174_, _10169_, _source_stream_conv2d_8_source_24_pat_count_1[1:0] }), .Y(_10168_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33927_ ( .A({ _10173_, _10172_, _10171_, _10170_ }), .Y(_10169_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33928_ ( .A(_source_stream_conv2d_8_source_24_pat_count_1[13:10]), .Y(_10170_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33929_ ( .A(_source_stream_conv2d_8_source_24_pat_count_1[9:6]), .Y(_10171_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33930_ ( .A(_source_stream_conv2d_8_source_24_pat_count_1[21:18]), .Y(_10172_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33931_ ( .A(_source_stream_conv2d_8_source_24_pat_count_1[17:14]), .Y(_10173_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33932_ ( .A(_source_stream_conv2d_8_source_24_pat_count_1[5:2]), .Y(_10174_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33933_ ( .A({ _10176_, _source_stream_conv2d_8_source_24_pat_count_1[32:30] }), .Y(_10175_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33934_ ( .A({ _source_stream_conv2d_8_source_24_pat_count_1[28:27], _source_stream_conv2d_8_source_24_pat_count_1[25], _source_stream_conv2d_8_source_24_pat_count_1[22] }), .Y(_10176_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33935_ ( .A({ _source_stream_conv2d_8_source_24_pat_count_1[29], _source_stream_conv2d_8_source_24_pat_count_1[26], _source_stream_conv2d_8_source_24_pat_count_1[24:23] }), .Y(_10177_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33936_ ( .A({ _10178_, _10167_, _05710_ }), .Y(_05712_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33937_ ( .A({ _10188_, _10183_, _10181_, _10179_ }), .Y(_10178_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33938_ ( .A({ _10180_, _source_stream_conv2d_8_source_24_pat_count_2[32:30] }), .Y(_10179_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33939_ ( .A({ _source_stream_conv2d_8_source_24_pat_count_2[28:27], _source_stream_conv2d_8_source_24_pat_count_2[25], _source_stream_conv2d_8_source_24_pat_count_2[22] }), .Y(_10180_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33940_ ( .A({ _10182_, _source_stream_conv2d_8_source_24_pat_count_2[1:0] }), .Y(_10181_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33941_ ( .A(_source_stream_conv2d_8_source_24_pat_count_2[5:2]), .Y(_10182_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33942_ ( .A({ _10187_, _10186_, _10185_, _10184_ }), .Y(_10183_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33943_ ( .A(_source_stream_conv2d_8_source_24_pat_count_2[13:10]), .Y(_10184_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33944_ ( .A(_source_stream_conv2d_8_source_24_pat_count_2[9:6]), .Y(_10185_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33945_ ( .A(_source_stream_conv2d_8_source_24_pat_count_2[21:18]), .Y(_10186_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33946_ ( .A(_source_stream_conv2d_8_source_24_pat_count_2[17:14]), .Y(_10187_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33947_ ( .A({ _source_stream_conv2d_8_source_24_pat_count_2[29], _source_stream_conv2d_8_source_24_pat_count_2[26], _source_stream_conv2d_8_source_24_pat_count_2[24:23] }), .Y(_10188_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33948_ ( .A({ _05833_, _05085_ }), .Y(_05713_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33949_ ( .A({ _10189_, _10178_, _10156_, _10167_ }), .Y(_05833_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33950_ ( .A({ _10199_, _10194_, _10192_, _10190_ }), .Y(_10189_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33951_ ( .A({ _10191_, _source_stream_conv2d_8_source_24_pat_count_3[32:30] }), .Y(_10190_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33952_ ( .A({ _source_stream_conv2d_8_source_24_pat_count_3[28:27], _source_stream_conv2d_8_source_24_pat_count_3[25], _source_stream_conv2d_8_source_24_pat_count_3[22] }), .Y(_10191_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33953_ ( .A({ _10193_, _source_stream_conv2d_8_source_24_pat_count_3[1:0] }), .Y(_10192_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33954_ ( .A(_source_stream_conv2d_8_source_24_pat_count_3[5:2]), .Y(_10193_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33955_ ( .A({ _10198_, _10197_, _10196_, _10195_ }), .Y(_10194_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33956_ ( .A(_source_stream_conv2d_8_source_24_pat_count_3[13:10]), .Y(_10195_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33957_ ( .A(_source_stream_conv2d_8_source_24_pat_count_3[9:6]), .Y(_10196_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33958_ ( .A(_source_stream_conv2d_8_source_24_pat_count_3[21:18]), .Y(_10197_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33959_ ( .A(_source_stream_conv2d_8_source_24_pat_count_3[17:14]), .Y(_10198_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33960_ ( .A({ _source_stream_conv2d_8_source_24_pat_count_3[29], _source_stream_conv2d_8_source_24_pat_count_3[26], _source_stream_conv2d_8_source_24_pat_count_3[24:23] }), .Y(_10199_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33961_ ( .A({ _10200_, _05083_ }), .Y(_05715_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33962_ ( .A({ _10210_, _10205_, _10203_, _10201_ }), .Y(_10200_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33963_ ( .A({ _10202_, _source_stream_conv2d_8_source_25_pat_count_0[32:30] }), .Y(_10201_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33964_ ( .A({ _source_stream_conv2d_8_source_25_pat_count_0[28:27], _source_stream_conv2d_8_source_25_pat_count_0[25], _source_stream_conv2d_8_source_25_pat_count_0[22] }), .Y(_10202_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33965_ ( .A({ _10204_, _source_stream_conv2d_8_source_25_pat_count_0[1:0] }), .Y(_10203_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33966_ ( .A(_source_stream_conv2d_8_source_25_pat_count_0[5:2]), .Y(_10204_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33967_ ( .A({ _10209_, _10208_, _10207_, _10206_ }), .Y(_10205_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33968_ ( .A(_source_stream_conv2d_8_source_25_pat_count_0[13:10]), .Y(_10206_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33969_ ( .A(_source_stream_conv2d_8_source_25_pat_count_0[9:6]), .Y(_10207_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33970_ ( .A(_source_stream_conv2d_8_source_25_pat_count_0[21:18]), .Y(_10208_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33971_ ( .A(_source_stream_conv2d_8_source_25_pat_count_0[17:14]), .Y(_10209_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33972_ ( .A({ _source_stream_conv2d_8_source_25_pat_count_0[29], _source_stream_conv2d_8_source_25_pat_count_0[26], _source_stream_conv2d_8_source_25_pat_count_0[24:23] }), .Y(_10210_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33973_ ( .A({ _10211_, _05715_ }), .Y(_05716_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33974_ ( .A({ _10221_, _10219_, _10212_ }), .Y(_10211_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33975_ ( .A({ _10218_, _10213_, _source_stream_conv2d_8_source_25_pat_count_1[1:0] }), .Y(_10212_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33976_ ( .A({ _10217_, _10216_, _10215_, _10214_ }), .Y(_10213_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33977_ ( .A(_source_stream_conv2d_8_source_25_pat_count_1[13:10]), .Y(_10214_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33978_ ( .A(_source_stream_conv2d_8_source_25_pat_count_1[9:6]), .Y(_10215_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33979_ ( .A(_source_stream_conv2d_8_source_25_pat_count_1[21:18]), .Y(_10216_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33980_ ( .A(_source_stream_conv2d_8_source_25_pat_count_1[17:14]), .Y(_10217_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33981_ ( .A(_source_stream_conv2d_8_source_25_pat_count_1[5:2]), .Y(_10218_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33982_ ( .A({ _10220_, _source_stream_conv2d_8_source_25_pat_count_1[32:30] }), .Y(_10219_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33983_ ( .A({ _source_stream_conv2d_8_source_25_pat_count_1[28:27], _source_stream_conv2d_8_source_25_pat_count_1[25], _source_stream_conv2d_8_source_25_pat_count_1[22] }), .Y(_10220_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33984_ ( .A({ _source_stream_conv2d_8_source_25_pat_count_1[29], _source_stream_conv2d_8_source_25_pat_count_1[26], _source_stream_conv2d_8_source_25_pat_count_1[24:23] }), .Y(_10221_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33985_ ( .A({ _10222_, _10211_, _05715_ }), .Y(_05717_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33986_ ( .A({ _10232_, _10227_, _10225_, _10223_ }), .Y(_10222_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33987_ ( .A({ _10224_, _source_stream_conv2d_8_source_25_pat_count_2[32:30] }), .Y(_10223_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33988_ ( .A({ _source_stream_conv2d_8_source_25_pat_count_2[28:27], _source_stream_conv2d_8_source_25_pat_count_2[25], _source_stream_conv2d_8_source_25_pat_count_2[22] }), .Y(_10224_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33989_ ( .A({ _10226_, _source_stream_conv2d_8_source_25_pat_count_2[1:0] }), .Y(_10225_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33990_ ( .A(_source_stream_conv2d_8_source_25_pat_count_2[5:2]), .Y(_10226_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33991_ ( .A({ _10231_, _10230_, _10229_, _10228_ }), .Y(_10227_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33992_ ( .A(_source_stream_conv2d_8_source_25_pat_count_2[13:10]), .Y(_10228_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33993_ ( .A(_source_stream_conv2d_8_source_25_pat_count_2[9:6]), .Y(_10229_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33994_ ( .A(_source_stream_conv2d_8_source_25_pat_count_2[21:18]), .Y(_10230_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33995_ ( .A(_source_stream_conv2d_8_source_25_pat_count_2[17:14]), .Y(_10231_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33996_ ( .A({ _source_stream_conv2d_8_source_25_pat_count_2[29], _source_stream_conv2d_8_source_25_pat_count_2[26], _source_stream_conv2d_8_source_25_pat_count_2[24:23] }), .Y(_10232_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33997_ ( .A({ _05834_, _05083_ }), .Y(_05718_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33998_ ( .A({ _10222_, _10233_, _10211_ }), .Y(_05834_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33999_ ( .A({ _10243_, _10241_, _10234_, _10200_ }), .Y(_10233_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34000_ ( .A({ _10240_, _10235_, _source_stream_conv2d_8_source_25_pat_count_3[1:0] }), .Y(_10234_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34001_ ( .A({ _10239_, _10238_, _10237_, _10236_ }), .Y(_10235_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34002_ ( .A(_source_stream_conv2d_8_source_25_pat_count_3[13:10]), .Y(_10236_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34003_ ( .A(_source_stream_conv2d_8_source_25_pat_count_3[9:6]), .Y(_10237_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34004_ ( .A(_source_stream_conv2d_8_source_25_pat_count_3[21:18]), .Y(_10238_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34005_ ( .A(_source_stream_conv2d_8_source_25_pat_count_3[17:14]), .Y(_10239_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34006_ ( .A(_source_stream_conv2d_8_source_25_pat_count_3[5:2]), .Y(_10240_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34007_ ( .A({ _10242_, _source_stream_conv2d_8_source_25_pat_count_3[32:30] }), .Y(_10241_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34008_ ( .A({ _source_stream_conv2d_8_source_25_pat_count_3[28:27], _source_stream_conv2d_8_source_25_pat_count_3[25], _source_stream_conv2d_8_source_25_pat_count_3[22] }), .Y(_10242_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34009_ ( .A({ _source_stream_conv2d_8_source_25_pat_count_3[29], _source_stream_conv2d_8_source_25_pat_count_3[26], _source_stream_conv2d_8_source_25_pat_count_3[24:23] }), .Y(_10243_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34010_ ( .A({ _10244_, _05081_ }), .Y(_05720_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34011_ ( .A({ _10254_, _10253_, _10252_, _10245_ }), .Y(_10244_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34012_ ( .A({ _10251_, _10246_, _source_stream_conv2d_8_source_26_pat_count_0[1:0] }), .Y(_10245_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34013_ ( .A({ _10250_, _10249_, _10248_, _10247_ }), .Y(_10246_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34014_ ( .A(_source_stream_conv2d_8_source_26_pat_count_0[13:10]), .Y(_10247_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34015_ ( .A(_source_stream_conv2d_8_source_26_pat_count_0[9:6]), .Y(_10248_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34016_ ( .A(_source_stream_conv2d_8_source_26_pat_count_0[21:18]), .Y(_10249_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34017_ ( .A(_source_stream_conv2d_8_source_26_pat_count_0[17:14]), .Y(_10250_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34018_ ( .A(_source_stream_conv2d_8_source_26_pat_count_0[5:2]), .Y(_10251_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34019_ ( .A(_source_stream_conv2d_8_source_26_pat_count_0[32:30]), .Y(_10252_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34020_ ( .A(_source_stream_conv2d_8_source_26_pat_count_0[29:26]), .Y(_10253_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34021_ ( .A(_source_stream_conv2d_8_source_26_pat_count_0[25:22]), .Y(_10254_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34022_ ( .A({ _10255_, _05720_ }), .Y(_05721_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34023_ ( .A({ _10265_, _10263_, _10256_ }), .Y(_10255_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34024_ ( .A({ _10262_, _10257_, _source_stream_conv2d_8_source_26_pat_count_1[1:0] }), .Y(_10256_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34025_ ( .A({ _10261_, _10260_, _10259_, _10258_ }), .Y(_10257_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34026_ ( .A(_source_stream_conv2d_8_source_26_pat_count_1[13:10]), .Y(_10258_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34027_ ( .A(_source_stream_conv2d_8_source_26_pat_count_1[9:6]), .Y(_10259_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34028_ ( .A(_source_stream_conv2d_8_source_26_pat_count_1[21:18]), .Y(_10260_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34029_ ( .A(_source_stream_conv2d_8_source_26_pat_count_1[17:14]), .Y(_10261_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34030_ ( .A(_source_stream_conv2d_8_source_26_pat_count_1[5:2]), .Y(_10262_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34031_ ( .A({ _10264_, _source_stream_conv2d_8_source_26_pat_count_1[32:30] }), .Y(_10263_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34032_ ( .A({ _source_stream_conv2d_8_source_26_pat_count_1[28:27], _source_stream_conv2d_8_source_26_pat_count_1[25], _source_stream_conv2d_8_source_26_pat_count_1[22] }), .Y(_10264_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34033_ ( .A({ _source_stream_conv2d_8_source_26_pat_count_1[29], _source_stream_conv2d_8_source_26_pat_count_1[26], _source_stream_conv2d_8_source_26_pat_count_1[24:23] }), .Y(_10265_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34034_ ( .A({ _10266_, _10255_, _05720_ }), .Y(_05722_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34035_ ( .A({ _10276_, _10271_, _10269_, _10267_ }), .Y(_10266_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34036_ ( .A({ _10268_, _source_stream_conv2d_8_source_26_pat_count_2[32:30] }), .Y(_10267_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34037_ ( .A({ _source_stream_conv2d_8_source_26_pat_count_2[28:27], _source_stream_conv2d_8_source_26_pat_count_2[25], _source_stream_conv2d_8_source_26_pat_count_2[22] }), .Y(_10268_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34038_ ( .A({ _10270_, _source_stream_conv2d_8_source_26_pat_count_2[1:0] }), .Y(_10269_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34039_ ( .A(_source_stream_conv2d_8_source_26_pat_count_2[5:2]), .Y(_10270_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34040_ ( .A({ _10275_, _10274_, _10273_, _10272_ }), .Y(_10271_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34041_ ( .A(_source_stream_conv2d_8_source_26_pat_count_2[13:10]), .Y(_10272_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34042_ ( .A(_source_stream_conv2d_8_source_26_pat_count_2[9:6]), .Y(_10273_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34043_ ( .A(_source_stream_conv2d_8_source_26_pat_count_2[21:18]), .Y(_10274_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34044_ ( .A(_source_stream_conv2d_8_source_26_pat_count_2[17:14]), .Y(_10275_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34045_ ( .A({ _source_stream_conv2d_8_source_26_pat_count_2[29], _source_stream_conv2d_8_source_26_pat_count_2[26], _source_stream_conv2d_8_source_26_pat_count_2[24:23] }), .Y(_10276_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34046_ ( .A({ _05835_, _05081_ }), .Y(_05723_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34047_ ( .A({ _10277_, _10266_, _10255_, _10244_ }), .Y(_05835_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34048_ ( .A({ _10287_, _10282_, _10280_, _10278_ }), .Y(_10277_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34049_ ( .A({ _10279_, _source_stream_conv2d_8_source_26_pat_count_3[32:30] }), .Y(_10278_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34050_ ( .A({ _source_stream_conv2d_8_source_26_pat_count_3[28:27], _source_stream_conv2d_8_source_26_pat_count_3[25], _source_stream_conv2d_8_source_26_pat_count_3[22] }), .Y(_10279_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34051_ ( .A({ _10281_, _source_stream_conv2d_8_source_26_pat_count_3[1:0] }), .Y(_10280_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34052_ ( .A(_source_stream_conv2d_8_source_26_pat_count_3[5:2]), .Y(_10281_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34053_ ( .A({ _10286_, _10285_, _10284_, _10283_ }), .Y(_10282_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34054_ ( .A(_source_stream_conv2d_8_source_26_pat_count_3[13:10]), .Y(_10283_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34055_ ( .A(_source_stream_conv2d_8_source_26_pat_count_3[9:6]), .Y(_10284_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34056_ ( .A(_source_stream_conv2d_8_source_26_pat_count_3[21:18]), .Y(_10285_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34057_ ( .A(_source_stream_conv2d_8_source_26_pat_count_3[17:14]), .Y(_10286_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34058_ ( .A({ _source_stream_conv2d_8_source_26_pat_count_3[29], _source_stream_conv2d_8_source_26_pat_count_3[26], _source_stream_conv2d_8_source_26_pat_count_3[24:23] }), .Y(_10287_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34059_ ( .A({ _10288_, _05079_ }), .Y(_05725_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34060_ ( .A({ _10298_, _10293_, _10291_, _10289_ }), .Y(_10288_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34061_ ( .A({ _10290_, _source_stream_conv2d_8_source_27_pat_count_0[32:30] }), .Y(_10289_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34062_ ( .A({ _source_stream_conv2d_8_source_27_pat_count_0[28:27], _source_stream_conv2d_8_source_27_pat_count_0[25], _source_stream_conv2d_8_source_27_pat_count_0[22] }), .Y(_10290_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34063_ ( .A({ _10292_, _source_stream_conv2d_8_source_27_pat_count_0[1:0] }), .Y(_10291_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34064_ ( .A(_source_stream_conv2d_8_source_27_pat_count_0[5:2]), .Y(_10292_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34065_ ( .A({ _10297_, _10296_, _10295_, _10294_ }), .Y(_10293_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34066_ ( .A(_source_stream_conv2d_8_source_27_pat_count_0[13:10]), .Y(_10294_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34067_ ( .A(_source_stream_conv2d_8_source_27_pat_count_0[9:6]), .Y(_10295_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34068_ ( .A(_source_stream_conv2d_8_source_27_pat_count_0[21:18]), .Y(_10296_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34069_ ( .A(_source_stream_conv2d_8_source_27_pat_count_0[17:14]), .Y(_10297_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34070_ ( .A({ _source_stream_conv2d_8_source_27_pat_count_0[29], _source_stream_conv2d_8_source_27_pat_count_0[26], _source_stream_conv2d_8_source_27_pat_count_0[24:23] }), .Y(_10298_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34071_ ( .A({ _10299_, _05725_ }), .Y(_05726_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34072_ ( .A({ _10309_, _10307_, _10300_ }), .Y(_10299_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34073_ ( .A({ _10306_, _10301_, _source_stream_conv2d_8_source_27_pat_count_1[1:0] }), .Y(_10300_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34074_ ( .A({ _10305_, _10304_, _10303_, _10302_ }), .Y(_10301_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34075_ ( .A(_source_stream_conv2d_8_source_27_pat_count_1[13:10]), .Y(_10302_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34076_ ( .A(_source_stream_conv2d_8_source_27_pat_count_1[9:6]), .Y(_10303_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34077_ ( .A(_source_stream_conv2d_8_source_27_pat_count_1[21:18]), .Y(_10304_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34078_ ( .A(_source_stream_conv2d_8_source_27_pat_count_1[17:14]), .Y(_10305_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34079_ ( .A(_source_stream_conv2d_8_source_27_pat_count_1[5:2]), .Y(_10306_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34080_ ( .A({ _10308_, _source_stream_conv2d_8_source_27_pat_count_1[32:30] }), .Y(_10307_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34081_ ( .A({ _source_stream_conv2d_8_source_27_pat_count_1[28:27], _source_stream_conv2d_8_source_27_pat_count_1[25], _source_stream_conv2d_8_source_27_pat_count_1[22] }), .Y(_10308_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34082_ ( .A({ _source_stream_conv2d_8_source_27_pat_count_1[29], _source_stream_conv2d_8_source_27_pat_count_1[26], _source_stream_conv2d_8_source_27_pat_count_1[24:23] }), .Y(_10309_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34083_ ( .A({ _10310_, _10299_, _05725_ }), .Y(_05727_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34084_ ( .A({ _10320_, _10315_, _10313_, _10311_ }), .Y(_10310_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34085_ ( .A({ _10312_, _source_stream_conv2d_8_source_27_pat_count_2[32:30] }), .Y(_10311_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34086_ ( .A({ _source_stream_conv2d_8_source_27_pat_count_2[28:27], _source_stream_conv2d_8_source_27_pat_count_2[25], _source_stream_conv2d_8_source_27_pat_count_2[22] }), .Y(_10312_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34087_ ( .A({ _10314_, _source_stream_conv2d_8_source_27_pat_count_2[1:0] }), .Y(_10313_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34088_ ( .A(_source_stream_conv2d_8_source_27_pat_count_2[5:2]), .Y(_10314_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34089_ ( .A({ _10319_, _10318_, _10317_, _10316_ }), .Y(_10315_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34090_ ( .A(_source_stream_conv2d_8_source_27_pat_count_2[13:10]), .Y(_10316_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34091_ ( .A(_source_stream_conv2d_8_source_27_pat_count_2[9:6]), .Y(_10317_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34092_ ( .A(_source_stream_conv2d_8_source_27_pat_count_2[21:18]), .Y(_10318_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34093_ ( .A(_source_stream_conv2d_8_source_27_pat_count_2[17:14]), .Y(_10319_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34094_ ( .A({ _source_stream_conv2d_8_source_27_pat_count_2[29], _source_stream_conv2d_8_source_27_pat_count_2[26], _source_stream_conv2d_8_source_27_pat_count_2[24:23] }), .Y(_10320_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34095_ ( .A({ _05836_, _05079_ }), .Y(_05728_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34096_ ( .A({ _10321_, _10310_, _10288_, _10299_ }), .Y(_05836_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34097_ ( .A({ _10331_, _10326_, _10324_, _10322_ }), .Y(_10321_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34098_ ( .A({ _10323_, _source_stream_conv2d_8_source_27_pat_count_3[32:30] }), .Y(_10322_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34099_ ( .A({ _source_stream_conv2d_8_source_27_pat_count_3[28:27], _source_stream_conv2d_8_source_27_pat_count_3[25], _source_stream_conv2d_8_source_27_pat_count_3[22] }), .Y(_10323_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34100_ ( .A({ _10325_, _source_stream_conv2d_8_source_27_pat_count_3[1:0] }), .Y(_10324_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34101_ ( .A(_source_stream_conv2d_8_source_27_pat_count_3[5:2]), .Y(_10325_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34102_ ( .A({ _10330_, _10329_, _10328_, _10327_ }), .Y(_10326_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34103_ ( .A(_source_stream_conv2d_8_source_27_pat_count_3[13:10]), .Y(_10327_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34104_ ( .A(_source_stream_conv2d_8_source_27_pat_count_3[9:6]), .Y(_10328_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34105_ ( .A(_source_stream_conv2d_8_source_27_pat_count_3[21:18]), .Y(_10329_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34106_ ( .A(_source_stream_conv2d_8_source_27_pat_count_3[17:14]), .Y(_10330_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34107_ ( .A({ _source_stream_conv2d_8_source_27_pat_count_3[29], _source_stream_conv2d_8_source_27_pat_count_3[26], _source_stream_conv2d_8_source_27_pat_count_3[24:23] }), .Y(_10331_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34108_ ( .A({ _10332_, _05077_ }), .Y(_05730_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34109_ ( .A({ _10342_, _10337_, _10335_, _10333_ }), .Y(_10332_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34110_ ( .A({ _10334_, _source_stream_conv2d_8_source_28_pat_count_0[32:30] }), .Y(_10333_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34111_ ( .A({ _source_stream_conv2d_8_source_28_pat_count_0[28:27], _source_stream_conv2d_8_source_28_pat_count_0[25], _source_stream_conv2d_8_source_28_pat_count_0[22] }), .Y(_10334_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34112_ ( .A({ _10336_, _source_stream_conv2d_8_source_28_pat_count_0[1:0] }), .Y(_10335_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34113_ ( .A(_source_stream_conv2d_8_source_28_pat_count_0[5:2]), .Y(_10336_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34114_ ( .A({ _10341_, _10340_, _10339_, _10338_ }), .Y(_10337_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34115_ ( .A(_source_stream_conv2d_8_source_28_pat_count_0[13:10]), .Y(_10338_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34116_ ( .A(_source_stream_conv2d_8_source_28_pat_count_0[9:6]), .Y(_10339_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34117_ ( .A(_source_stream_conv2d_8_source_28_pat_count_0[21:18]), .Y(_10340_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34118_ ( .A(_source_stream_conv2d_8_source_28_pat_count_0[17:14]), .Y(_10341_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34119_ ( .A({ _source_stream_conv2d_8_source_28_pat_count_0[29], _source_stream_conv2d_8_source_28_pat_count_0[26], _source_stream_conv2d_8_source_28_pat_count_0[24:23] }), .Y(_10342_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34120_ ( .A({ _10343_, _05730_ }), .Y(_05731_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34121_ ( .A({ _10353_, _10351_, _10344_ }), .Y(_10343_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34122_ ( .A({ _10350_, _10345_, _source_stream_conv2d_8_source_28_pat_count_1[1:0] }), .Y(_10344_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34123_ ( .A({ _10349_, _10348_, _10347_, _10346_ }), .Y(_10345_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34124_ ( .A(_source_stream_conv2d_8_source_28_pat_count_1[13:10]), .Y(_10346_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34125_ ( .A(_source_stream_conv2d_8_source_28_pat_count_1[9:6]), .Y(_10347_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34126_ ( .A(_source_stream_conv2d_8_source_28_pat_count_1[21:18]), .Y(_10348_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34127_ ( .A(_source_stream_conv2d_8_source_28_pat_count_1[17:14]), .Y(_10349_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34128_ ( .A(_source_stream_conv2d_8_source_28_pat_count_1[5:2]), .Y(_10350_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34129_ ( .A({ _10352_, _source_stream_conv2d_8_source_28_pat_count_1[32:30] }), .Y(_10351_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34130_ ( .A({ _source_stream_conv2d_8_source_28_pat_count_1[28:27], _source_stream_conv2d_8_source_28_pat_count_1[25], _source_stream_conv2d_8_source_28_pat_count_1[22] }), .Y(_10352_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34131_ ( .A({ _source_stream_conv2d_8_source_28_pat_count_1[29], _source_stream_conv2d_8_source_28_pat_count_1[26], _source_stream_conv2d_8_source_28_pat_count_1[24:23] }), .Y(_10353_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34132_ ( .A({ _10354_, _10343_, _05730_ }), .Y(_05732_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34133_ ( .A({ _10364_, _10359_, _10357_, _10355_ }), .Y(_10354_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34134_ ( .A({ _10356_, _source_stream_conv2d_8_source_28_pat_count_2[32:30] }), .Y(_10355_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34135_ ( .A({ _source_stream_conv2d_8_source_28_pat_count_2[28:27], _source_stream_conv2d_8_source_28_pat_count_2[25], _source_stream_conv2d_8_source_28_pat_count_2[22] }), .Y(_10356_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34136_ ( .A({ _10358_, _source_stream_conv2d_8_source_28_pat_count_2[1:0] }), .Y(_10357_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34137_ ( .A(_source_stream_conv2d_8_source_28_pat_count_2[5:2]), .Y(_10358_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34138_ ( .A({ _10363_, _10362_, _10361_, _10360_ }), .Y(_10359_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34139_ ( .A(_source_stream_conv2d_8_source_28_pat_count_2[13:10]), .Y(_10360_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34140_ ( .A(_source_stream_conv2d_8_source_28_pat_count_2[9:6]), .Y(_10361_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34141_ ( .A(_source_stream_conv2d_8_source_28_pat_count_2[21:18]), .Y(_10362_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34142_ ( .A(_source_stream_conv2d_8_source_28_pat_count_2[17:14]), .Y(_10363_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34143_ ( .A({ _source_stream_conv2d_8_source_28_pat_count_2[29], _source_stream_conv2d_8_source_28_pat_count_2[26], _source_stream_conv2d_8_source_28_pat_count_2[24:23] }), .Y(_10364_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34144_ ( .A({ _05837_, _05077_ }), .Y(_05733_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34145_ ( .A({ _10365_, _10354_, _10332_, _10343_ }), .Y(_05837_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34146_ ( .A({ _10375_, _10370_, _10368_, _10366_ }), .Y(_10365_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34147_ ( .A({ _10367_, _source_stream_conv2d_8_source_28_pat_count_3[32:30] }), .Y(_10366_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34148_ ( .A({ _source_stream_conv2d_8_source_28_pat_count_3[28:27], _source_stream_conv2d_8_source_28_pat_count_3[25], _source_stream_conv2d_8_source_28_pat_count_3[22] }), .Y(_10367_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34149_ ( .A({ _10369_, _source_stream_conv2d_8_source_28_pat_count_3[1:0] }), .Y(_10368_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34150_ ( .A(_source_stream_conv2d_8_source_28_pat_count_3[5:2]), .Y(_10369_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34151_ ( .A({ _10374_, _10373_, _10372_, _10371_ }), .Y(_10370_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34152_ ( .A(_source_stream_conv2d_8_source_28_pat_count_3[13:10]), .Y(_10371_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34153_ ( .A(_source_stream_conv2d_8_source_28_pat_count_3[9:6]), .Y(_10372_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34154_ ( .A(_source_stream_conv2d_8_source_28_pat_count_3[21:18]), .Y(_10373_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34155_ ( .A(_source_stream_conv2d_8_source_28_pat_count_3[17:14]), .Y(_10374_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34156_ ( .A({ _source_stream_conv2d_8_source_28_pat_count_3[29], _source_stream_conv2d_8_source_28_pat_count_3[26], _source_stream_conv2d_8_source_28_pat_count_3[24:23] }), .Y(_10375_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34157_ ( .A({ _10376_, _05075_ }), .Y(_05735_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34158_ ( .A({ _10386_, _10381_, _10379_, _10377_ }), .Y(_10376_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34159_ ( .A({ _10378_, _source_stream_conv2d_8_source_29_pat_count_0[32:30] }), .Y(_10377_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34160_ ( .A({ _source_stream_conv2d_8_source_29_pat_count_0[28:27], _source_stream_conv2d_8_source_29_pat_count_0[25], _source_stream_conv2d_8_source_29_pat_count_0[22] }), .Y(_10378_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34161_ ( .A({ _10380_, _source_stream_conv2d_8_source_29_pat_count_0[1:0] }), .Y(_10379_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34162_ ( .A(_source_stream_conv2d_8_source_29_pat_count_0[5:2]), .Y(_10380_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34163_ ( .A({ _10385_, _10384_, _10383_, _10382_ }), .Y(_10381_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34164_ ( .A(_source_stream_conv2d_8_source_29_pat_count_0[13:10]), .Y(_10382_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34165_ ( .A(_source_stream_conv2d_8_source_29_pat_count_0[9:6]), .Y(_10383_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34166_ ( .A(_source_stream_conv2d_8_source_29_pat_count_0[21:18]), .Y(_10384_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34167_ ( .A(_source_stream_conv2d_8_source_29_pat_count_0[17:14]), .Y(_10385_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34168_ ( .A({ _source_stream_conv2d_8_source_29_pat_count_0[29], _source_stream_conv2d_8_source_29_pat_count_0[26], _source_stream_conv2d_8_source_29_pat_count_0[24:23] }), .Y(_10386_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34169_ ( .A({ _10387_, _05735_ }), .Y(_05736_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34170_ ( .A({ _10397_, _10395_, _10388_ }), .Y(_10387_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34171_ ( .A({ _10394_, _10389_, _source_stream_conv2d_8_source_29_pat_count_1[1:0] }), .Y(_10388_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34172_ ( .A({ _10393_, _10392_, _10391_, _10390_ }), .Y(_10389_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34173_ ( .A(_source_stream_conv2d_8_source_29_pat_count_1[13:10]), .Y(_10390_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34174_ ( .A(_source_stream_conv2d_8_source_29_pat_count_1[9:6]), .Y(_10391_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34175_ ( .A(_source_stream_conv2d_8_source_29_pat_count_1[21:18]), .Y(_10392_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34176_ ( .A(_source_stream_conv2d_8_source_29_pat_count_1[17:14]), .Y(_10393_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34177_ ( .A(_source_stream_conv2d_8_source_29_pat_count_1[5:2]), .Y(_10394_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34178_ ( .A({ _10396_, _source_stream_conv2d_8_source_29_pat_count_1[32:30] }), .Y(_10395_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34179_ ( .A({ _source_stream_conv2d_8_source_29_pat_count_1[28:27], _source_stream_conv2d_8_source_29_pat_count_1[25], _source_stream_conv2d_8_source_29_pat_count_1[22] }), .Y(_10396_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34180_ ( .A({ _source_stream_conv2d_8_source_29_pat_count_1[29], _source_stream_conv2d_8_source_29_pat_count_1[26], _source_stream_conv2d_8_source_29_pat_count_1[24:23] }), .Y(_10397_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34181_ ( .A({ _10398_, _10387_, _05735_ }), .Y(_05737_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34182_ ( .A({ _10408_, _10403_, _10401_, _10399_ }), .Y(_10398_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34183_ ( .A({ _10400_, _source_stream_conv2d_8_source_29_pat_count_2[32:30] }), .Y(_10399_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34184_ ( .A({ _source_stream_conv2d_8_source_29_pat_count_2[28:27], _source_stream_conv2d_8_source_29_pat_count_2[25], _source_stream_conv2d_8_source_29_pat_count_2[22] }), .Y(_10400_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34185_ ( .A({ _10402_, _source_stream_conv2d_8_source_29_pat_count_2[1:0] }), .Y(_10401_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34186_ ( .A(_source_stream_conv2d_8_source_29_pat_count_2[5:2]), .Y(_10402_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34187_ ( .A({ _10407_, _10406_, _10405_, _10404_ }), .Y(_10403_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34188_ ( .A(_source_stream_conv2d_8_source_29_pat_count_2[13:10]), .Y(_10404_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34189_ ( .A(_source_stream_conv2d_8_source_29_pat_count_2[9:6]), .Y(_10405_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34190_ ( .A(_source_stream_conv2d_8_source_29_pat_count_2[21:18]), .Y(_10406_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34191_ ( .A(_source_stream_conv2d_8_source_29_pat_count_2[17:14]), .Y(_10407_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34192_ ( .A({ _source_stream_conv2d_8_source_29_pat_count_2[29], _source_stream_conv2d_8_source_29_pat_count_2[26], _source_stream_conv2d_8_source_29_pat_count_2[24:23] }), .Y(_10408_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34193_ ( .A({ _05838_, _05075_ }), .Y(_05738_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34194_ ( .A({ _10398_, _10409_, _10387_ }), .Y(_05838_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34195_ ( .A({ _10419_, _10417_, _10410_, _10376_ }), .Y(_10409_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34196_ ( .A({ _10416_, _10411_, _source_stream_conv2d_8_source_29_pat_count_3[1:0] }), .Y(_10410_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34197_ ( .A({ _10415_, _10414_, _10413_, _10412_ }), .Y(_10411_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34198_ ( .A(_source_stream_conv2d_8_source_29_pat_count_3[13:10]), .Y(_10412_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34199_ ( .A(_source_stream_conv2d_8_source_29_pat_count_3[9:6]), .Y(_10413_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34200_ ( .A(_source_stream_conv2d_8_source_29_pat_count_3[21:18]), .Y(_10414_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34201_ ( .A(_source_stream_conv2d_8_source_29_pat_count_3[17:14]), .Y(_10415_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34202_ ( .A(_source_stream_conv2d_8_source_29_pat_count_3[5:2]), .Y(_10416_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34203_ ( .A({ _10418_, _source_stream_conv2d_8_source_29_pat_count_3[32:30] }), .Y(_10417_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34204_ ( .A({ _source_stream_conv2d_8_source_29_pat_count_3[28:27], _source_stream_conv2d_8_source_29_pat_count_3[25], _source_stream_conv2d_8_source_29_pat_count_3[22] }), .Y(_10418_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34205_ ( .A({ _source_stream_conv2d_8_source_29_pat_count_3[29], _source_stream_conv2d_8_source_29_pat_count_3[26], _source_stream_conv2d_8_source_29_pat_count_3[24:23] }), .Y(_10419_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34206_ ( .A({ _10420_, _05073_ }), .Y(_05740_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34207_ ( .A({ _10430_, _10425_, _10423_, _10421_ }), .Y(_10420_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34208_ ( .A({ _10422_, _source_stream_conv2d_8_source_30_pat_count_0[32:30] }), .Y(_10421_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34209_ ( .A({ _source_stream_conv2d_8_source_30_pat_count_0[28:27], _source_stream_conv2d_8_source_30_pat_count_0[25], _source_stream_conv2d_8_source_30_pat_count_0[22] }), .Y(_10422_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34210_ ( .A({ _10424_, _source_stream_conv2d_8_source_30_pat_count_0[1:0] }), .Y(_10423_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34211_ ( .A(_source_stream_conv2d_8_source_30_pat_count_0[5:2]), .Y(_10424_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34212_ ( .A({ _10429_, _10428_, _10427_, _10426_ }), .Y(_10425_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34213_ ( .A(_source_stream_conv2d_8_source_30_pat_count_0[13:10]), .Y(_10426_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34214_ ( .A(_source_stream_conv2d_8_source_30_pat_count_0[9:6]), .Y(_10427_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34215_ ( .A(_source_stream_conv2d_8_source_30_pat_count_0[21:18]), .Y(_10428_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34216_ ( .A(_source_stream_conv2d_8_source_30_pat_count_0[17:14]), .Y(_10429_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34217_ ( .A({ _source_stream_conv2d_8_source_30_pat_count_0[29], _source_stream_conv2d_8_source_30_pat_count_0[26], _source_stream_conv2d_8_source_30_pat_count_0[24:23] }), .Y(_10430_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34218_ ( .A({ _10431_, _05740_ }), .Y(_05741_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34219_ ( .A({ _10441_, _10439_, _10432_ }), .Y(_10431_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34220_ ( .A({ _10438_, _10433_, _source_stream_conv2d_8_source_30_pat_count_1[1:0] }), .Y(_10432_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34221_ ( .A({ _10437_, _10436_, _10435_, _10434_ }), .Y(_10433_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34222_ ( .A(_source_stream_conv2d_8_source_30_pat_count_1[13:10]), .Y(_10434_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34223_ ( .A(_source_stream_conv2d_8_source_30_pat_count_1[9:6]), .Y(_10435_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34224_ ( .A(_source_stream_conv2d_8_source_30_pat_count_1[21:18]), .Y(_10436_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34225_ ( .A(_source_stream_conv2d_8_source_30_pat_count_1[17:14]), .Y(_10437_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34226_ ( .A(_source_stream_conv2d_8_source_30_pat_count_1[5:2]), .Y(_10438_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34227_ ( .A({ _10440_, _source_stream_conv2d_8_source_30_pat_count_1[32:30] }), .Y(_10439_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34228_ ( .A({ _source_stream_conv2d_8_source_30_pat_count_1[28:27], _source_stream_conv2d_8_source_30_pat_count_1[25], _source_stream_conv2d_8_source_30_pat_count_1[22] }), .Y(_10440_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34229_ ( .A({ _source_stream_conv2d_8_source_30_pat_count_1[29], _source_stream_conv2d_8_source_30_pat_count_1[26], _source_stream_conv2d_8_source_30_pat_count_1[24:23] }), .Y(_10441_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34230_ ( .A({ _10442_, _10431_, _05740_ }), .Y(_05742_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34231_ ( .A({ _10452_, _10447_, _10445_, _10443_ }), .Y(_10442_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34232_ ( .A({ _10444_, _source_stream_conv2d_8_source_30_pat_count_2[32:30] }), .Y(_10443_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34233_ ( .A({ _source_stream_conv2d_8_source_30_pat_count_2[28:27], _source_stream_conv2d_8_source_30_pat_count_2[25], _source_stream_conv2d_8_source_30_pat_count_2[22] }), .Y(_10444_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34234_ ( .A({ _10446_, _source_stream_conv2d_8_source_30_pat_count_2[1:0] }), .Y(_10445_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34235_ ( .A(_source_stream_conv2d_8_source_30_pat_count_2[5:2]), .Y(_10446_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34236_ ( .A({ _10451_, _10450_, _10449_, _10448_ }), .Y(_10447_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34237_ ( .A(_source_stream_conv2d_8_source_30_pat_count_2[13:10]), .Y(_10448_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34238_ ( .A(_source_stream_conv2d_8_source_30_pat_count_2[9:6]), .Y(_10449_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34239_ ( .A(_source_stream_conv2d_8_source_30_pat_count_2[21:18]), .Y(_10450_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34240_ ( .A(_source_stream_conv2d_8_source_30_pat_count_2[17:14]), .Y(_10451_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34241_ ( .A({ _source_stream_conv2d_8_source_30_pat_count_2[29], _source_stream_conv2d_8_source_30_pat_count_2[26], _source_stream_conv2d_8_source_30_pat_count_2[24:23] }), .Y(_10452_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34242_ ( .A({ _05839_, _05073_ }), .Y(_05743_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34243_ ( .A({ _10442_, _10453_, _10431_ }), .Y(_05839_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34244_ ( .A({ _10463_, _10461_, _10454_, _10420_ }), .Y(_10453_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34245_ ( .A({ _10460_, _10455_, _source_stream_conv2d_8_source_30_pat_count_3[1:0] }), .Y(_10454_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34246_ ( .A({ _10459_, _10458_, _10457_, _10456_ }), .Y(_10455_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34247_ ( .A(_source_stream_conv2d_8_source_30_pat_count_3[13:10]), .Y(_10456_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34248_ ( .A(_source_stream_conv2d_8_source_30_pat_count_3[9:6]), .Y(_10457_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34249_ ( .A(_source_stream_conv2d_8_source_30_pat_count_3[21:18]), .Y(_10458_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34250_ ( .A(_source_stream_conv2d_8_source_30_pat_count_3[17:14]), .Y(_10459_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34251_ ( .A(_source_stream_conv2d_8_source_30_pat_count_3[5:2]), .Y(_10460_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34252_ ( .A({ _10462_, _source_stream_conv2d_8_source_30_pat_count_3[32:30] }), .Y(_10461_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34253_ ( .A({ _source_stream_conv2d_8_source_30_pat_count_3[28:27], _source_stream_conv2d_8_source_30_pat_count_3[25], _source_stream_conv2d_8_source_30_pat_count_3[22] }), .Y(_10462_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34254_ ( .A({ _source_stream_conv2d_8_source_30_pat_count_3[29], _source_stream_conv2d_8_source_30_pat_count_3[26], _source_stream_conv2d_8_source_30_pat_count_3[24:23] }), .Y(_10463_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34255_ ( .A({ _10464_, _05071_ }), .Y(_05745_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34256_ ( .A({ _10474_, _10473_, _10472_, _10465_ }), .Y(_10464_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34257_ ( .A({ _10471_, _10466_, _source_stream_conv2d_8_source_31_pat_count_0[1:0] }), .Y(_10465_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34258_ ( .A({ _10470_, _10469_, _10468_, _10467_ }), .Y(_10466_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34259_ ( .A(_source_stream_conv2d_8_source_31_pat_count_0[13:10]), .Y(_10467_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34260_ ( .A(_source_stream_conv2d_8_source_31_pat_count_0[9:6]), .Y(_10468_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34261_ ( .A(_source_stream_conv2d_8_source_31_pat_count_0[21:18]), .Y(_10469_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34262_ ( .A(_source_stream_conv2d_8_source_31_pat_count_0[17:14]), .Y(_10470_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34263_ ( .A(_source_stream_conv2d_8_source_31_pat_count_0[5:2]), .Y(_10471_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34264_ ( .A(_source_stream_conv2d_8_source_31_pat_count_0[32:30]), .Y(_10472_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34265_ ( .A(_source_stream_conv2d_8_source_31_pat_count_0[29:26]), .Y(_10473_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34266_ ( .A(_source_stream_conv2d_8_source_31_pat_count_0[25:22]), .Y(_10474_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34267_ ( .A({ _10475_, _05745_ }), .Y(_05746_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34268_ ( .A({ _10485_, _10483_, _10476_ }), .Y(_10475_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34269_ ( .A({ _10482_, _10477_, _source_stream_conv2d_8_source_31_pat_count_1[1:0] }), .Y(_10476_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34270_ ( .A({ _10481_, _10480_, _10479_, _10478_ }), .Y(_10477_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34271_ ( .A(_source_stream_conv2d_8_source_31_pat_count_1[13:10]), .Y(_10478_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34272_ ( .A(_source_stream_conv2d_8_source_31_pat_count_1[9:6]), .Y(_10479_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34273_ ( .A(_source_stream_conv2d_8_source_31_pat_count_1[21:18]), .Y(_10480_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34274_ ( .A(_source_stream_conv2d_8_source_31_pat_count_1[17:14]), .Y(_10481_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34275_ ( .A(_source_stream_conv2d_8_source_31_pat_count_1[5:2]), .Y(_10482_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34276_ ( .A({ _10484_, _source_stream_conv2d_8_source_31_pat_count_1[32:30] }), .Y(_10483_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34277_ ( .A({ _source_stream_conv2d_8_source_31_pat_count_1[28:27], _source_stream_conv2d_8_source_31_pat_count_1[25], _source_stream_conv2d_8_source_31_pat_count_1[22] }), .Y(_10484_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34278_ ( .A({ _source_stream_conv2d_8_source_31_pat_count_1[29], _source_stream_conv2d_8_source_31_pat_count_1[26], _source_stream_conv2d_8_source_31_pat_count_1[24:23] }), .Y(_10485_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34279_ ( .A({ _10486_, _05745_ }), .Y(_05747_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34280_ ( .A({ _10496_, _10493_, _10487_, _10475_ }), .Y(_10486_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34281_ ( .A({ _10492_, _10490_, _10488_ }), .Y(_10487_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34282_ ( .A({ _10489_, _source_stream_conv2d_8_source_31_pat_count_2[17], _source_stream_conv2d_8_source_31_pat_count_2[14], _source_stream_conv2d_8_source_31_pat_count_2[4] }), .Y(_10488_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34283_ ( .A({ _source_stream_conv2d_8_source_31_pat_count_2[21], _source_stream_conv2d_8_source_31_pat_count_2[18], _source_stream_conv2d_8_source_31_pat_count_2[16:15] }), .Y(_10489_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34284_ ( .A({ _10491_, _source_stream_conv2d_8_source_31_pat_count_2[10], _source_stream_conv2d_8_source_31_pat_count_2[5] }), .Y(_10490_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34285_ ( .A({ _source_stream_conv2d_8_source_31_pat_count_2[13], _source_stream_conv2d_8_source_31_pat_count_2[8:7] }), .Y(_10491_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34286_ ( .A({ _source_stream_conv2d_8_source_31_pat_count_2[12:11], _source_stream_conv2d_8_source_31_pat_count_2[9], _source_stream_conv2d_8_source_31_pat_count_2[6] }), .Y(_10492_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34287_ ( .A({ _10494_, _source_stream_conv2d_8_source_31_pat_count_2[2], _source_stream_conv2d_8_source_31_pat_count_2[0] }), .Y(_10493_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34288_ ( .A({ _10495_, _source_stream_conv2d_8_source_31_pat_count_2[29], _source_stream_conv2d_8_source_31_pat_count_2[26] }), .Y(_10494_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34289_ ( .A(_source_stream_conv2d_8_source_31_pat_count_2[32:30]), .Y(_10495_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34290_ ( .A({ _10497_, _source_stream_conv2d_8_source_31_pat_count_2[25:23] }), .Y(_10496_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34291_ ( .A({ _10498_, _source_stream_conv2d_8_source_31_pat_count_2[27], _source_stream_conv2d_8_source_31_pat_count_2[20], _source_stream_conv2d_8_source_31_pat_count_2[1] }), .Y(_10497_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34292_ ( .A({ _source_stream_conv2d_8_source_31_pat_count_2[28], _source_stream_conv2d_8_source_31_pat_count_2[22], _source_stream_conv2d_8_source_31_pat_count_2[19], _source_stream_conv2d_8_source_31_pat_count_2[3] }), .Y(_10498_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34293_ ( .A({ _10499_, _05747_ }), .Y(_05748_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34294_ ( .A({ _10509_, _10507_, _10500_ }), .Y(_10499_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34295_ ( .A({ _10506_, _10501_, _source_stream_conv2d_8_source_31_pat_count_3[1:0] }), .Y(_10500_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34296_ ( .A({ _10505_, _10504_, _10503_, _10502_ }), .Y(_10501_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34297_ ( .A(_source_stream_conv2d_8_source_31_pat_count_3[13:10]), .Y(_10502_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34298_ ( .A(_source_stream_conv2d_8_source_31_pat_count_3[9:6]), .Y(_10503_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34299_ ( .A(_source_stream_conv2d_8_source_31_pat_count_3[21:18]), .Y(_10504_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34300_ ( .A(_source_stream_conv2d_8_source_31_pat_count_3[17:14]), .Y(_10505_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34301_ ( .A(_source_stream_conv2d_8_source_31_pat_count_3[5:2]), .Y(_10506_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34302_ ( .A({ _10508_, _source_stream_conv2d_8_source_31_pat_count_3[32:30] }), .Y(_10507_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34303_ ( .A({ _source_stream_conv2d_8_source_31_pat_count_3[28:27], _source_stream_conv2d_8_source_31_pat_count_3[25], _source_stream_conv2d_8_source_31_pat_count_3[22] }), .Y(_10508_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34304_ ( .A({ _source_stream_conv2d_8_source_31_pat_count_3[29], _source_stream_conv2d_8_source_31_pat_count_3[26], _source_stream_conv2d_8_source_31_pat_count_3[24:23] }), .Y(_10509_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34305_ ( .A({ _10510_, _05069_ }), .Y(_05750_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34306_ ( .A({ _10520_, _10515_, _10513_, _10511_ }), .Y(_10510_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34307_ ( .A({ _10512_, _source_stream_conv2d_8_source_32_pat_count_0[32:30] }), .Y(_10511_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34308_ ( .A({ _source_stream_conv2d_8_source_32_pat_count_0[28:27], _source_stream_conv2d_8_source_32_pat_count_0[25], _source_stream_conv2d_8_source_32_pat_count_0[22] }), .Y(_10512_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34309_ ( .A({ _10514_, _source_stream_conv2d_8_source_32_pat_count_0[1:0] }), .Y(_10513_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34310_ ( .A(_source_stream_conv2d_8_source_32_pat_count_0[5:2]), .Y(_10514_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34311_ ( .A({ _10519_, _10518_, _10517_, _10516_ }), .Y(_10515_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34312_ ( .A(_source_stream_conv2d_8_source_32_pat_count_0[13:10]), .Y(_10516_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34313_ ( .A(_source_stream_conv2d_8_source_32_pat_count_0[9:6]), .Y(_10517_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34314_ ( .A(_source_stream_conv2d_8_source_32_pat_count_0[21:18]), .Y(_10518_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34315_ ( .A(_source_stream_conv2d_8_source_32_pat_count_0[17:14]), .Y(_10519_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34316_ ( .A({ _source_stream_conv2d_8_source_32_pat_count_0[29], _source_stream_conv2d_8_source_32_pat_count_0[26], _source_stream_conv2d_8_source_32_pat_count_0[24:23] }), .Y(_10520_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34317_ ( .A({ _10521_, _05750_ }), .Y(_05751_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34318_ ( .A({ _10531_, _10529_, _10522_ }), .Y(_10521_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34319_ ( .A({ _10528_, _10523_, _source_stream_conv2d_8_source_32_pat_count_1[1:0] }), .Y(_10522_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34320_ ( .A({ _10527_, _10526_, _10525_, _10524_ }), .Y(_10523_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34321_ ( .A(_source_stream_conv2d_8_source_32_pat_count_1[13:10]), .Y(_10524_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34322_ ( .A(_source_stream_conv2d_8_source_32_pat_count_1[9:6]), .Y(_10525_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34323_ ( .A(_source_stream_conv2d_8_source_32_pat_count_1[21:18]), .Y(_10526_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34324_ ( .A(_source_stream_conv2d_8_source_32_pat_count_1[17:14]), .Y(_10527_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34325_ ( .A(_source_stream_conv2d_8_source_32_pat_count_1[5:2]), .Y(_10528_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34326_ ( .A({ _10530_, _source_stream_conv2d_8_source_32_pat_count_1[32:30] }), .Y(_10529_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34327_ ( .A({ _source_stream_conv2d_8_source_32_pat_count_1[28:27], _source_stream_conv2d_8_source_32_pat_count_1[25], _source_stream_conv2d_8_source_32_pat_count_1[22] }), .Y(_10530_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34328_ ( .A({ _source_stream_conv2d_8_source_32_pat_count_1[29], _source_stream_conv2d_8_source_32_pat_count_1[26], _source_stream_conv2d_8_source_32_pat_count_1[24:23] }), .Y(_10531_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34329_ ( .A({ _10532_, _05750_ }), .Y(_05752_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34330_ ( .A({ _10533_, _10521_ }), .Y(_10532_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34331_ ( .A({ _10543_, _10538_, _10536_, _10534_ }), .Y(_10533_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34332_ ( .A({ _10535_, _source_stream_conv2d_8_source_32_pat_count_2[32:30] }), .Y(_10534_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34333_ ( .A({ _source_stream_conv2d_8_source_32_pat_count_2[28:27], _source_stream_conv2d_8_source_32_pat_count_2[25], _source_stream_conv2d_8_source_32_pat_count_2[22] }), .Y(_10535_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34334_ ( .A({ _10537_, _source_stream_conv2d_8_source_32_pat_count_2[1:0] }), .Y(_10536_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34335_ ( .A(_source_stream_conv2d_8_source_32_pat_count_2[5:2]), .Y(_10537_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34336_ ( .A({ _10542_, _10541_, _10540_, _10539_ }), .Y(_10538_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34337_ ( .A(_source_stream_conv2d_8_source_32_pat_count_2[13:10]), .Y(_10539_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34338_ ( .A(_source_stream_conv2d_8_source_32_pat_count_2[9:6]), .Y(_10540_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34339_ ( .A(_source_stream_conv2d_8_source_32_pat_count_2[21:18]), .Y(_10541_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34340_ ( .A(_source_stream_conv2d_8_source_32_pat_count_2[17:14]), .Y(_10542_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34341_ ( .A({ _source_stream_conv2d_8_source_32_pat_count_2[29], _source_stream_conv2d_8_source_32_pat_count_2[26], _source_stream_conv2d_8_source_32_pat_count_2[24:23] }), .Y(_10543_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34342_ ( .A({ _10544_, _05752_ }), .Y(_05753_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34343_ ( .A({ _10554_, _10552_, _10545_ }), .Y(_10544_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34344_ ( .A({ _10551_, _10546_, _source_stream_conv2d_8_source_32_pat_count_3[1:0] }), .Y(_10545_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34345_ ( .A({ _10550_, _10549_, _10548_, _10547_ }), .Y(_10546_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34346_ ( .A(_source_stream_conv2d_8_source_32_pat_count_3[13:10]), .Y(_10547_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34347_ ( .A(_source_stream_conv2d_8_source_32_pat_count_3[9:6]), .Y(_10548_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34348_ ( .A(_source_stream_conv2d_8_source_32_pat_count_3[21:18]), .Y(_10549_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34349_ ( .A(_source_stream_conv2d_8_source_32_pat_count_3[17:14]), .Y(_10550_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34350_ ( .A(_source_stream_conv2d_8_source_32_pat_count_3[5:2]), .Y(_10551_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34351_ ( .A({ _10553_, _source_stream_conv2d_8_source_32_pat_count_3[32:30] }), .Y(_10552_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34352_ ( .A({ _source_stream_conv2d_8_source_32_pat_count_3[28:27], _source_stream_conv2d_8_source_32_pat_count_3[25], _source_stream_conv2d_8_source_32_pat_count_3[22] }), .Y(_10553_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34353_ ( .A({ _source_stream_conv2d_8_source_32_pat_count_3[29], _source_stream_conv2d_8_source_32_pat_count_3[26], _source_stream_conv2d_8_source_32_pat_count_3[24:23] }), .Y(_10554_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34354_ ( .A({ _10555_, _05067_ }), .Y(_05755_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34355_ ( .A({ _10565_, _10564_, _10563_, _10556_ }), .Y(_10555_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34356_ ( .A({ _10562_, _10557_, _source_stream_conv2d_8_source_33_pat_count_0[1:0] }), .Y(_10556_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34357_ ( .A({ _10561_, _10560_, _10559_, _10558_ }), .Y(_10557_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34358_ ( .A(_source_stream_conv2d_8_source_33_pat_count_0[13:10]), .Y(_10558_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34359_ ( .A(_source_stream_conv2d_8_source_33_pat_count_0[9:6]), .Y(_10559_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34360_ ( .A(_source_stream_conv2d_8_source_33_pat_count_0[21:18]), .Y(_10560_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34361_ ( .A(_source_stream_conv2d_8_source_33_pat_count_0[17:14]), .Y(_10561_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34362_ ( .A(_source_stream_conv2d_8_source_33_pat_count_0[5:2]), .Y(_10562_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34363_ ( .A(_source_stream_conv2d_8_source_33_pat_count_0[32:30]), .Y(_10563_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34364_ ( .A(_source_stream_conv2d_8_source_33_pat_count_0[29:26]), .Y(_10564_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34365_ ( .A(_source_stream_conv2d_8_source_33_pat_count_0[25:22]), .Y(_10565_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34366_ ( .A({ _10566_, _05755_ }), .Y(_05756_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34367_ ( .A({ _10576_, _10574_, _10567_ }), .Y(_10566_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34368_ ( .A({ _10573_, _10568_, _source_stream_conv2d_8_source_33_pat_count_1[1:0] }), .Y(_10567_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34369_ ( .A({ _10572_, _10571_, _10570_, _10569_ }), .Y(_10568_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34370_ ( .A(_source_stream_conv2d_8_source_33_pat_count_1[13:10]), .Y(_10569_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34371_ ( .A(_source_stream_conv2d_8_source_33_pat_count_1[9:6]), .Y(_10570_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34372_ ( .A(_source_stream_conv2d_8_source_33_pat_count_1[21:18]), .Y(_10571_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34373_ ( .A(_source_stream_conv2d_8_source_33_pat_count_1[17:14]), .Y(_10572_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34374_ ( .A(_source_stream_conv2d_8_source_33_pat_count_1[5:2]), .Y(_10573_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34375_ ( .A({ _10575_, _source_stream_conv2d_8_source_33_pat_count_1[32:30] }), .Y(_10574_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34376_ ( .A({ _source_stream_conv2d_8_source_33_pat_count_1[28:27], _source_stream_conv2d_8_source_33_pat_count_1[25], _source_stream_conv2d_8_source_33_pat_count_1[22] }), .Y(_10575_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34377_ ( .A({ _source_stream_conv2d_8_source_33_pat_count_1[29], _source_stream_conv2d_8_source_33_pat_count_1[26], _source_stream_conv2d_8_source_33_pat_count_1[24:23] }), .Y(_10576_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34378_ ( .A({ _10577_, _05755_ }), .Y(_05757_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34379_ ( .A({ _10584_, _10578_, _10566_ }), .Y(_10577_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34380_ ( .A({ _10583_, _10581_, _10579_ }), .Y(_10578_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34381_ ( .A({ _10580_, _source_stream_conv2d_8_source_33_pat_count_2[17], _source_stream_conv2d_8_source_33_pat_count_2[14], _source_stream_conv2d_8_source_33_pat_count_2[4] }), .Y(_10579_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34382_ ( .A({ _source_stream_conv2d_8_source_33_pat_count_2[21], _source_stream_conv2d_8_source_33_pat_count_2[18], _source_stream_conv2d_8_source_33_pat_count_2[16:15] }), .Y(_10580_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34383_ ( .A({ _10582_, _source_stream_conv2d_8_source_33_pat_count_2[27], _source_stream_conv2d_8_source_33_pat_count_2[20], _source_stream_conv2d_8_source_33_pat_count_2[1] }), .Y(_10581_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34384_ ( .A({ _source_stream_conv2d_8_source_33_pat_count_2[28], _source_stream_conv2d_8_source_33_pat_count_2[22], _source_stream_conv2d_8_source_33_pat_count_2[19], _source_stream_conv2d_8_source_33_pat_count_2[3] }), .Y(_10582_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34385_ ( .A({ _source_stream_conv2d_8_source_33_pat_count_2[12:11], _source_stream_conv2d_8_source_33_pat_count_2[9], _source_stream_conv2d_8_source_33_pat_count_2[6] }), .Y(_10583_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34386_ ( .A({ _10588_, _10585_, _source_stream_conv2d_8_source_33_pat_count_2[2], _source_stream_conv2d_8_source_33_pat_count_2[0] }), .Y(_10584_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34387_ ( .A({ _10587_, _10586_, _source_stream_conv2d_8_source_33_pat_count_2[10], _source_stream_conv2d_8_source_33_pat_count_2[5] }), .Y(_10585_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34388_ ( .A(_source_stream_conv2d_8_source_33_pat_count_2[25:23]), .Y(_10586_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34389_ ( .A({ _source_stream_conv2d_8_source_33_pat_count_2[13], _source_stream_conv2d_8_source_33_pat_count_2[8:7] }), .Y(_10587_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34390_ ( .A({ _10589_, _source_stream_conv2d_8_source_33_pat_count_2[29], _source_stream_conv2d_8_source_33_pat_count_2[26] }), .Y(_10588_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34391_ ( .A(_source_stream_conv2d_8_source_33_pat_count_2[32:30]), .Y(_10589_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34392_ ( .A({ _10590_, _05757_ }), .Y(_05758_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34393_ ( .A({ _10600_, _10598_, _10591_ }), .Y(_10590_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34394_ ( .A({ _10597_, _10592_, _source_stream_conv2d_8_source_33_pat_count_3[1:0] }), .Y(_10591_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34395_ ( .A({ _10596_, _10595_, _10594_, _10593_ }), .Y(_10592_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34396_ ( .A(_source_stream_conv2d_8_source_33_pat_count_3[13:10]), .Y(_10593_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34397_ ( .A(_source_stream_conv2d_8_source_33_pat_count_3[9:6]), .Y(_10594_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34398_ ( .A(_source_stream_conv2d_8_source_33_pat_count_3[21:18]), .Y(_10595_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34399_ ( .A(_source_stream_conv2d_8_source_33_pat_count_3[17:14]), .Y(_10596_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34400_ ( .A(_source_stream_conv2d_8_source_33_pat_count_3[5:2]), .Y(_10597_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34401_ ( .A({ _10599_, _source_stream_conv2d_8_source_33_pat_count_3[32:30] }), .Y(_10598_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34402_ ( .A({ _source_stream_conv2d_8_source_33_pat_count_3[28:27], _source_stream_conv2d_8_source_33_pat_count_3[25], _source_stream_conv2d_8_source_33_pat_count_3[22] }), .Y(_10599_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34403_ ( .A({ _source_stream_conv2d_8_source_33_pat_count_3[29], _source_stream_conv2d_8_source_33_pat_count_3[26], _source_stream_conv2d_8_source_33_pat_count_3[24:23] }), .Y(_10600_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34404_ ( .A({ _10601_, _05066_ }), .Y(_05760_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34405_ ( .A({ _10611_, _10610_, _10609_, _10602_ }), .Y(_10601_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34406_ ( .A({ _10608_, _10603_, _source_stream_conv2d_8_source_34_pat_count_0[1:0] }), .Y(_10602_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34407_ ( .A({ _10607_, _10606_, _10605_, _10604_ }), .Y(_10603_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34408_ ( .A(_source_stream_conv2d_8_source_34_pat_count_0[13:10]), .Y(_10604_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34409_ ( .A(_source_stream_conv2d_8_source_34_pat_count_0[9:6]), .Y(_10605_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34410_ ( .A(_source_stream_conv2d_8_source_34_pat_count_0[21:18]), .Y(_10606_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34411_ ( .A(_source_stream_conv2d_8_source_34_pat_count_0[17:14]), .Y(_10607_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34412_ ( .A(_source_stream_conv2d_8_source_34_pat_count_0[5:2]), .Y(_10608_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34413_ ( .A(_source_stream_conv2d_8_source_34_pat_count_0[32:30]), .Y(_10609_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34414_ ( .A(_source_stream_conv2d_8_source_34_pat_count_0[29:26]), .Y(_10610_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34415_ ( .A(_source_stream_conv2d_8_source_34_pat_count_0[25:22]), .Y(_10611_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34416_ ( .A({ _10612_, _05760_ }), .Y(_05761_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34417_ ( .A({ _10622_, _10620_, _10613_ }), .Y(_10612_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34418_ ( .A({ _10619_, _10614_, _source_stream_conv2d_8_source_34_pat_count_1[1:0] }), .Y(_10613_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34419_ ( .A({ _10618_, _10617_, _10616_, _10615_ }), .Y(_10614_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34420_ ( .A(_source_stream_conv2d_8_source_34_pat_count_1[13:10]), .Y(_10615_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34421_ ( .A(_source_stream_conv2d_8_source_34_pat_count_1[9:6]), .Y(_10616_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34422_ ( .A(_source_stream_conv2d_8_source_34_pat_count_1[21:18]), .Y(_10617_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34423_ ( .A(_source_stream_conv2d_8_source_34_pat_count_1[17:14]), .Y(_10618_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34424_ ( .A(_source_stream_conv2d_8_source_34_pat_count_1[5:2]), .Y(_10619_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34425_ ( .A({ _10621_, _source_stream_conv2d_8_source_34_pat_count_1[32:30] }), .Y(_10620_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34426_ ( .A({ _source_stream_conv2d_8_source_34_pat_count_1[28:27], _source_stream_conv2d_8_source_34_pat_count_1[25], _source_stream_conv2d_8_source_34_pat_count_1[22] }), .Y(_10621_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34427_ ( .A({ _source_stream_conv2d_8_source_34_pat_count_1[29], _source_stream_conv2d_8_source_34_pat_count_1[26], _source_stream_conv2d_8_source_34_pat_count_1[24:23] }), .Y(_10622_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34428_ ( .A({ _10623_, _05760_ }), .Y(_05762_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34429_ ( .A({ _10633_, _10630_, _10624_, _10612_ }), .Y(_10623_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34430_ ( .A({ _10629_, _10627_, _10625_ }), .Y(_10624_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34431_ ( .A({ _10626_, _source_stream_conv2d_8_source_34_pat_count_2[17], _source_stream_conv2d_8_source_34_pat_count_2[14], _source_stream_conv2d_8_source_34_pat_count_2[4] }), .Y(_10625_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34432_ ( .A({ _source_stream_conv2d_8_source_34_pat_count_2[21], _source_stream_conv2d_8_source_34_pat_count_2[18], _source_stream_conv2d_8_source_34_pat_count_2[16:15] }), .Y(_10626_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34433_ ( .A({ _10628_, _source_stream_conv2d_8_source_34_pat_count_2[10], _source_stream_conv2d_8_source_34_pat_count_2[5] }), .Y(_10627_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34434_ ( .A({ _source_stream_conv2d_8_source_34_pat_count_2[13], _source_stream_conv2d_8_source_34_pat_count_2[8:7] }), .Y(_10628_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34435_ ( .A({ _source_stream_conv2d_8_source_34_pat_count_2[12:11], _source_stream_conv2d_8_source_34_pat_count_2[9], _source_stream_conv2d_8_source_34_pat_count_2[6] }), .Y(_10629_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34436_ ( .A({ _10631_, _source_stream_conv2d_8_source_34_pat_count_2[2], _source_stream_conv2d_8_source_34_pat_count_2[0] }), .Y(_10630_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34437_ ( .A({ _10632_, _source_stream_conv2d_8_source_34_pat_count_2[29], _source_stream_conv2d_8_source_34_pat_count_2[26] }), .Y(_10631_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34438_ ( .A(_source_stream_conv2d_8_source_34_pat_count_2[32:30]), .Y(_10632_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34439_ ( .A({ _10634_, _source_stream_conv2d_8_source_34_pat_count_2[25:23] }), .Y(_10633_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34440_ ( .A({ _10635_, _source_stream_conv2d_8_source_34_pat_count_2[27], _source_stream_conv2d_8_source_34_pat_count_2[20], _source_stream_conv2d_8_source_34_pat_count_2[1] }), .Y(_10634_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34441_ ( .A({ _source_stream_conv2d_8_source_34_pat_count_2[28], _source_stream_conv2d_8_source_34_pat_count_2[22], _source_stream_conv2d_8_source_34_pat_count_2[19], _source_stream_conv2d_8_source_34_pat_count_2[3] }), .Y(_10635_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34442_ ( .A({ _10636_, _05762_ }), .Y(_05763_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34443_ ( .A({ _10646_, _10644_, _10637_ }), .Y(_10636_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34444_ ( .A({ _10643_, _10638_, _source_stream_conv2d_8_source_34_pat_count_3[1:0] }), .Y(_10637_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34445_ ( .A({ _10642_, _10641_, _10640_, _10639_ }), .Y(_10638_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34446_ ( .A(_source_stream_conv2d_8_source_34_pat_count_3[13:10]), .Y(_10639_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34447_ ( .A(_source_stream_conv2d_8_source_34_pat_count_3[9:6]), .Y(_10640_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34448_ ( .A(_source_stream_conv2d_8_source_34_pat_count_3[21:18]), .Y(_10641_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34449_ ( .A(_source_stream_conv2d_8_source_34_pat_count_3[17:14]), .Y(_10642_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34450_ ( .A(_source_stream_conv2d_8_source_34_pat_count_3[5:2]), .Y(_10643_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34451_ ( .A({ _10645_, _source_stream_conv2d_8_source_34_pat_count_3[32:30] }), .Y(_10644_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34452_ ( .A({ _source_stream_conv2d_8_source_34_pat_count_3[28:27], _source_stream_conv2d_8_source_34_pat_count_3[25], _source_stream_conv2d_8_source_34_pat_count_3[22] }), .Y(_10645_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34453_ ( .A({ _source_stream_conv2d_8_source_34_pat_count_3[29], _source_stream_conv2d_8_source_34_pat_count_3[26], _source_stream_conv2d_8_source_34_pat_count_3[24:23] }), .Y(_10646_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34454_ ( .A({ _10647_, _05064_ }), .Y(_05765_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34455_ ( .A({ _10657_, _10656_, _10655_, _10648_ }), .Y(_10647_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34456_ ( .A({ _10654_, _10649_, _source_stream_conv2d_8_source_35_pat_count_0[1:0] }), .Y(_10648_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34457_ ( .A({ _10653_, _10652_, _10651_, _10650_ }), .Y(_10649_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34458_ ( .A(_source_stream_conv2d_8_source_35_pat_count_0[13:10]), .Y(_10650_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34459_ ( .A(_source_stream_conv2d_8_source_35_pat_count_0[9:6]), .Y(_10651_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34460_ ( .A(_source_stream_conv2d_8_source_35_pat_count_0[21:18]), .Y(_10652_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34461_ ( .A(_source_stream_conv2d_8_source_35_pat_count_0[17:14]), .Y(_10653_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34462_ ( .A(_source_stream_conv2d_8_source_35_pat_count_0[5:2]), .Y(_10654_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34463_ ( .A(_source_stream_conv2d_8_source_35_pat_count_0[32:30]), .Y(_10655_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34464_ ( .A(_source_stream_conv2d_8_source_35_pat_count_0[29:26]), .Y(_10656_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34465_ ( .A(_source_stream_conv2d_8_source_35_pat_count_0[25:22]), .Y(_10657_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34466_ ( .A({ _10658_, _05765_ }), .Y(_05766_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34467_ ( .A({ _10668_, _10666_, _10659_ }), .Y(_10658_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34468_ ( .A({ _10665_, _10660_, _source_stream_conv2d_8_source_35_pat_count_1[1:0] }), .Y(_10659_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34469_ ( .A({ _10664_, _10663_, _10662_, _10661_ }), .Y(_10660_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34470_ ( .A(_source_stream_conv2d_8_source_35_pat_count_1[13:10]), .Y(_10661_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34471_ ( .A(_source_stream_conv2d_8_source_35_pat_count_1[9:6]), .Y(_10662_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34472_ ( .A(_source_stream_conv2d_8_source_35_pat_count_1[21:18]), .Y(_10663_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34473_ ( .A(_source_stream_conv2d_8_source_35_pat_count_1[17:14]), .Y(_10664_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34474_ ( .A(_source_stream_conv2d_8_source_35_pat_count_1[5:2]), .Y(_10665_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34475_ ( .A({ _10667_, _source_stream_conv2d_8_source_35_pat_count_1[32:30] }), .Y(_10666_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34476_ ( .A({ _source_stream_conv2d_8_source_35_pat_count_1[28:27], _source_stream_conv2d_8_source_35_pat_count_1[25], _source_stream_conv2d_8_source_35_pat_count_1[22] }), .Y(_10667_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34477_ ( .A({ _source_stream_conv2d_8_source_35_pat_count_1[29], _source_stream_conv2d_8_source_35_pat_count_1[26], _source_stream_conv2d_8_source_35_pat_count_1[24:23] }), .Y(_10668_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34478_ ( .A({ _10669_, _05765_ }), .Y(_05767_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34479_ ( .A({ _10679_, _10676_, _10670_, _10658_ }), .Y(_10669_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34480_ ( .A({ _10675_, _10673_, _10671_ }), .Y(_10670_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34481_ ( .A({ _10672_, _source_stream_conv2d_8_source_35_pat_count_2[17], _source_stream_conv2d_8_source_35_pat_count_2[14], _source_stream_conv2d_8_source_35_pat_count_2[4] }), .Y(_10671_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34482_ ( .A({ _source_stream_conv2d_8_source_35_pat_count_2[21], _source_stream_conv2d_8_source_35_pat_count_2[18], _source_stream_conv2d_8_source_35_pat_count_2[16:15] }), .Y(_10672_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34483_ ( .A({ _10674_, _source_stream_conv2d_8_source_35_pat_count_2[10], _source_stream_conv2d_8_source_35_pat_count_2[5] }), .Y(_10673_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34484_ ( .A({ _source_stream_conv2d_8_source_35_pat_count_2[13], _source_stream_conv2d_8_source_35_pat_count_2[8:7] }), .Y(_10674_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34485_ ( .A({ _source_stream_conv2d_8_source_35_pat_count_2[12:11], _source_stream_conv2d_8_source_35_pat_count_2[9], _source_stream_conv2d_8_source_35_pat_count_2[6] }), .Y(_10675_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34486_ ( .A({ _10677_, _source_stream_conv2d_8_source_35_pat_count_2[2], _source_stream_conv2d_8_source_35_pat_count_2[0] }), .Y(_10676_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34487_ ( .A({ _10678_, _source_stream_conv2d_8_source_35_pat_count_2[29], _source_stream_conv2d_8_source_35_pat_count_2[26] }), .Y(_10677_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34488_ ( .A(_source_stream_conv2d_8_source_35_pat_count_2[32:30]), .Y(_10678_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34489_ ( .A({ _10680_, _source_stream_conv2d_8_source_35_pat_count_2[25:23] }), .Y(_10679_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34490_ ( .A({ _10681_, _source_stream_conv2d_8_source_35_pat_count_2[27], _source_stream_conv2d_8_source_35_pat_count_2[20], _source_stream_conv2d_8_source_35_pat_count_2[1] }), .Y(_10680_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34491_ ( .A({ _source_stream_conv2d_8_source_35_pat_count_2[28], _source_stream_conv2d_8_source_35_pat_count_2[22], _source_stream_conv2d_8_source_35_pat_count_2[19], _source_stream_conv2d_8_source_35_pat_count_2[3] }), .Y(_10681_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34492_ ( .A({ _10682_, _05767_ }), .Y(_05768_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34493_ ( .A({ _10692_, _10690_, _10683_ }), .Y(_10682_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34494_ ( .A({ _10689_, _10684_, _source_stream_conv2d_8_source_35_pat_count_3[1:0] }), .Y(_10683_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34495_ ( .A({ _10688_, _10687_, _10686_, _10685_ }), .Y(_10684_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34496_ ( .A(_source_stream_conv2d_8_source_35_pat_count_3[13:10]), .Y(_10685_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34497_ ( .A(_source_stream_conv2d_8_source_35_pat_count_3[9:6]), .Y(_10686_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34498_ ( .A(_source_stream_conv2d_8_source_35_pat_count_3[21:18]), .Y(_10687_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34499_ ( .A(_source_stream_conv2d_8_source_35_pat_count_3[17:14]), .Y(_10688_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34500_ ( .A(_source_stream_conv2d_8_source_35_pat_count_3[5:2]), .Y(_10689_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34501_ ( .A({ _10691_, _source_stream_conv2d_8_source_35_pat_count_3[32:30] }), .Y(_10690_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34502_ ( .A({ _source_stream_conv2d_8_source_35_pat_count_3[28:27], _source_stream_conv2d_8_source_35_pat_count_3[25], _source_stream_conv2d_8_source_35_pat_count_3[22] }), .Y(_10691_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34503_ ( .A({ _source_stream_conv2d_8_source_35_pat_count_3[29], _source_stream_conv2d_8_source_35_pat_count_3[26], _source_stream_conv2d_8_source_35_pat_count_3[24:23] }), .Y(_10692_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34504_ ( .A({ _10693_, _05061_ }), .Y(_05770_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34505_ ( .A({ _10703_, _10702_, _10701_, _10694_ }), .Y(_10693_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34506_ ( .A({ _10700_, _10695_, _source_stream_conv2d_8_source_36_pat_count_0[1:0] }), .Y(_10694_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34507_ ( .A({ _10699_, _10698_, _10697_, _10696_ }), .Y(_10695_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34508_ ( .A(_source_stream_conv2d_8_source_36_pat_count_0[13:10]), .Y(_10696_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34509_ ( .A(_source_stream_conv2d_8_source_36_pat_count_0[9:6]), .Y(_10697_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34510_ ( .A(_source_stream_conv2d_8_source_36_pat_count_0[21:18]), .Y(_10698_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34511_ ( .A(_source_stream_conv2d_8_source_36_pat_count_0[17:14]), .Y(_10699_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34512_ ( .A(_source_stream_conv2d_8_source_36_pat_count_0[5:2]), .Y(_10700_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34513_ ( .A(_source_stream_conv2d_8_source_36_pat_count_0[32:30]), .Y(_10701_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34514_ ( .A(_source_stream_conv2d_8_source_36_pat_count_0[29:26]), .Y(_10702_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34515_ ( .A(_source_stream_conv2d_8_source_36_pat_count_0[25:22]), .Y(_10703_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34516_ ( .A({ _10704_, _05061_ }), .Y(_05771_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34517_ ( .A({ _10714_, _10712_, _10705_, _10693_ }), .Y(_10704_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34518_ ( .A({ _10711_, _10706_, _source_stream_conv2d_8_source_36_pat_count_1[1:0] }), .Y(_10705_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34519_ ( .A({ _10710_, _10709_, _10708_, _10707_ }), .Y(_10706_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34520_ ( .A(_source_stream_conv2d_8_source_36_pat_count_1[13:10]), .Y(_10707_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34521_ ( .A(_source_stream_conv2d_8_source_36_pat_count_1[9:6]), .Y(_10708_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34522_ ( .A(_source_stream_conv2d_8_source_36_pat_count_1[21:18]), .Y(_10709_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34523_ ( .A(_source_stream_conv2d_8_source_36_pat_count_1[17:14]), .Y(_10710_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34524_ ( .A(_source_stream_conv2d_8_source_36_pat_count_1[5:2]), .Y(_10711_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34525_ ( .A({ _10713_, _source_stream_conv2d_8_source_36_pat_count_1[32:30] }), .Y(_10712_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34526_ ( .A({ _source_stream_conv2d_8_source_36_pat_count_1[28:27], _source_stream_conv2d_8_source_36_pat_count_1[25], _source_stream_conv2d_8_source_36_pat_count_1[22] }), .Y(_10713_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34527_ ( .A({ _source_stream_conv2d_8_source_36_pat_count_1[29], _source_stream_conv2d_8_source_36_pat_count_1[26], _source_stream_conv2d_8_source_36_pat_count_1[24:23] }), .Y(_10714_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34528_ ( .A({ _10715_, _05771_ }), .Y(_05772_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34529_ ( .A({ _10725_, _10720_, _10718_, _10716_ }), .Y(_10715_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34530_ ( .A({ _10717_, _source_stream_conv2d_8_source_36_pat_count_2[32:30] }), .Y(_10716_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34531_ ( .A({ _source_stream_conv2d_8_source_36_pat_count_2[28:27], _source_stream_conv2d_8_source_36_pat_count_2[25], _source_stream_conv2d_8_source_36_pat_count_2[22] }), .Y(_10717_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34532_ ( .A({ _10719_, _source_stream_conv2d_8_source_36_pat_count_2[1:0] }), .Y(_10718_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34533_ ( .A(_source_stream_conv2d_8_source_36_pat_count_2[5:2]), .Y(_10719_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34534_ ( .A({ _10724_, _10723_, _10722_, _10721_ }), .Y(_10720_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34535_ ( .A(_source_stream_conv2d_8_source_36_pat_count_2[13:10]), .Y(_10721_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34536_ ( .A(_source_stream_conv2d_8_source_36_pat_count_2[9:6]), .Y(_10722_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34537_ ( .A(_source_stream_conv2d_8_source_36_pat_count_2[21:18]), .Y(_10723_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34538_ ( .A(_source_stream_conv2d_8_source_36_pat_count_2[17:14]), .Y(_10724_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34539_ ( .A({ _source_stream_conv2d_8_source_36_pat_count_2[29], _source_stream_conv2d_8_source_36_pat_count_2[26], _source_stream_conv2d_8_source_36_pat_count_2[24:23] }), .Y(_10725_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34540_ ( .A({ _10726_, _05771_ }), .Y(_05773_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34541_ ( .A({ _10737_, _10736_, _10715_, _10727_ }), .Y(_10726_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34542_ ( .A({ _10735_, _10733_, _10728_ }), .Y(_10727_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34543_ ( .A({ _10732_, _10731_, _10729_ }), .Y(_10728_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34544_ ( .A({ _10730_, _source_stream_conv2d_8_source_36_pat_count_3[1:0] }), .Y(_10729_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34545_ ( .A(_source_stream_conv2d_8_source_36_pat_count_3[5:2]), .Y(_10730_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34546_ ( .A({ _source_stream_conv2d_8_source_36_pat_count_3[13], _source_stream_conv2d_8_source_36_pat_count_3[10], _source_stream_conv2d_8_source_36_pat_count_3[8:7] }), .Y(_10731_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34547_ ( .A({ _source_stream_conv2d_8_source_36_pat_count_3[20:19], _source_stream_conv2d_8_source_36_pat_count_3[17], _source_stream_conv2d_8_source_36_pat_count_3[14] }), .Y(_10732_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34548_ ( .A({ _10734_, _source_stream_conv2d_8_source_36_pat_count_3[32:30] }), .Y(_10733_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34549_ ( .A({ _source_stream_conv2d_8_source_36_pat_count_3[28:27], _source_stream_conv2d_8_source_36_pat_count_3[25], _source_stream_conv2d_8_source_36_pat_count_3[22] }), .Y(_10734_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34550_ ( .A({ _source_stream_conv2d_8_source_36_pat_count_3[29], _source_stream_conv2d_8_source_36_pat_count_3[26], _source_stream_conv2d_8_source_36_pat_count_3[24:23] }), .Y(_10735_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34551_ ( .A({ _source_stream_conv2d_8_source_36_pat_count_3[12:11], _source_stream_conv2d_8_source_36_pat_count_3[9], _source_stream_conv2d_8_source_36_pat_count_3[6] }), .Y(_10736_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34552_ ( .A({ _source_stream_conv2d_8_source_36_pat_count_3[21], _source_stream_conv2d_8_source_36_pat_count_3[18], _source_stream_conv2d_8_source_36_pat_count_3[16:15] }), .Y(_10737_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34553_ ( .A({ __delay_data_1371, _stream_conv2d_8_sink_37_sink_fsm_20[0], _21900_ }), .Y(_05775_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34554_ ( .A({ _stream_conv2d_8_start_flag, _04903_ }), .Y(_tmp_541) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34555_ ( .A({ _10738_, _05043_ }), .Y(_05777_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34556_ ( .A({ _10748_, _10747_, _10746_, _10739_ }), .Y(_10738_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34557_ ( .A({ _10745_, _10740_, _source_stream_max_pool_serial_9_source_1_pat_count_0[1:0] }), .Y(_10739_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34558_ ( .A({ _10744_, _10743_, _10742_, _10741_ }), .Y(_10740_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34559_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_0[13:10]), .Y(_10741_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34560_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_0[9:6]), .Y(_10742_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34561_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_0[21:18]), .Y(_10743_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34562_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_0[17:14]), .Y(_10744_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34563_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_0[5:2]), .Y(_10745_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34564_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_0[32:30]), .Y(_10746_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34565_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_0[29:26]), .Y(_10747_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34566_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_0[25:22]), .Y(_10748_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34567_ ( .A({ _10749_, _05777_ }), .Y(_05778_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34568_ ( .A({ _10759_, _10757_, _10750_ }), .Y(_10749_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34569_ ( .A({ _10756_, _10751_, _source_stream_max_pool_serial_9_source_1_pat_count_1[1:0] }), .Y(_10750_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34570_ ( .A({ _10755_, _10754_, _10753_, _10752_ }), .Y(_10751_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34571_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_1[13:10]), .Y(_10752_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34572_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_1[9:6]), .Y(_10753_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34573_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_1[21:18]), .Y(_10754_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34574_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_1[17:14]), .Y(_10755_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34575_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_1[5:2]), .Y(_10756_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34576_ ( .A({ _10758_, _source_stream_max_pool_serial_9_source_1_pat_count_1[32:30] }), .Y(_10757_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34577_ ( .A({ _source_stream_max_pool_serial_9_source_1_pat_count_1[28:27], _source_stream_max_pool_serial_9_source_1_pat_count_1[25], _source_stream_max_pool_serial_9_source_1_pat_count_1[22] }), .Y(_10758_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34578_ ( .A({ _source_stream_max_pool_serial_9_source_1_pat_count_1[29], _source_stream_max_pool_serial_9_source_1_pat_count_1[26], _source_stream_max_pool_serial_9_source_1_pat_count_1[24:23] }), .Y(_10759_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34579_ ( .A({ _10760_, _05777_ }), .Y(_05779_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34580_ ( .A({ _10761_, _10749_ }), .Y(_10760_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34581_ ( .A({ _10771_, _10770_, _10769_, _10762_ }), .Y(_10761_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34582_ ( .A({ _10768_, _10763_, _source_stream_max_pool_serial_9_source_1_pat_count_2[1:0] }), .Y(_10762_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34583_ ( .A({ _10767_, _10766_, _10765_, _10764_ }), .Y(_10763_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34584_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_2[13:10]), .Y(_10764_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34585_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_2[9:6]), .Y(_10765_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34586_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_2[21:18]), .Y(_10766_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34587_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_2[17:14]), .Y(_10767_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34588_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_2[5:2]), .Y(_10768_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34589_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_2[32:30]), .Y(_10769_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34590_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_2[29:26]), .Y(_10770_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34591_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_2[25:22]), .Y(_10771_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34592_ ( .A({ _10772_, _05779_ }), .Y(_05780_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34593_ ( .A({ _10782_, _10780_, _10773_ }), .Y(_10772_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34594_ ( .A({ _10779_, _10774_, _source_stream_max_pool_serial_9_source_1_pat_count_3[1:0] }), .Y(_10773_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34595_ ( .A({ _10778_, _10777_, _10776_, _10775_ }), .Y(_10774_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34596_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_3[13:10]), .Y(_10775_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34597_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_3[9:6]), .Y(_10776_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34598_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_3[21:18]), .Y(_10777_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34599_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_3[17:14]), .Y(_10778_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34600_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_3[5:2]), .Y(_10779_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34601_ ( .A({ _10781_, _source_stream_max_pool_serial_9_source_1_pat_count_3[32:30] }), .Y(_10780_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34602_ ( .A({ _source_stream_max_pool_serial_9_source_1_pat_count_3[28:27], _source_stream_max_pool_serial_9_source_1_pat_count_3[25], _source_stream_max_pool_serial_9_source_1_pat_count_3[22] }), .Y(_10781_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34603_ ( .A({ _source_stream_max_pool_serial_9_source_1_pat_count_3[29], _source_stream_max_pool_serial_9_source_1_pat_count_3[26], _source_stream_max_pool_serial_9_source_1_pat_count_3[24:23] }), .Y(_10782_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34604_ ( .A({ __substreamoutput_data_774, _stream_max_pool_serial_9_sink_3_sink_fsm_1[0], _21891_ }), .Y(_05782_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34605_ ( .A({ _stream_max_pool_serial_9_start_flag, _04902_ }), .Y(_tmp_878) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34606_ ( .A({ _10783_, _05023_ }), .Y(_05784_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34607_ ( .A({ _10793_, _10792_, _10791_, _10784_ }), .Y(_10783_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34608_ ( .A({ _10790_, _10785_, _source_stream_matmul_15_source_6_pat_count_0[1:0] }), .Y(_10784_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34609_ ( .A({ _10789_, _10788_, _10787_, _10786_ }), .Y(_10785_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34610_ ( .A(_source_stream_matmul_15_source_6_pat_count_0[13:10]), .Y(_10786_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34611_ ( .A(_source_stream_matmul_15_source_6_pat_count_0[9:6]), .Y(_10787_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34612_ ( .A(_source_stream_matmul_15_source_6_pat_count_0[21:18]), .Y(_10788_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34613_ ( .A(_source_stream_matmul_15_source_6_pat_count_0[17:14]), .Y(_10789_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34614_ ( .A(_source_stream_matmul_15_source_6_pat_count_0[5:2]), .Y(_10790_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34615_ ( .A(_source_stream_matmul_15_source_6_pat_count_0[32:30]), .Y(_10791_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34616_ ( .A(_source_stream_matmul_15_source_6_pat_count_0[29:26]), .Y(_10792_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34617_ ( .A(_source_stream_matmul_15_source_6_pat_count_0[25:22]), .Y(_10793_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34618_ ( .A({ _10794_, _05784_ }), .Y(_05785_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34619_ ( .A({ _10804_, _10802_, _10795_ }), .Y(_10794_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34620_ ( .A({ _10801_, _10796_, _source_stream_matmul_15_source_6_pat_count_1[1:0] }), .Y(_10795_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34621_ ( .A({ _10800_, _10799_, _10798_, _10797_ }), .Y(_10796_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34622_ ( .A(_source_stream_matmul_15_source_6_pat_count_1[13:10]), .Y(_10797_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34623_ ( .A(_source_stream_matmul_15_source_6_pat_count_1[9:6]), .Y(_10798_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34624_ ( .A(_source_stream_matmul_15_source_6_pat_count_1[21:18]), .Y(_10799_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34625_ ( .A(_source_stream_matmul_15_source_6_pat_count_1[17:14]), .Y(_10800_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34626_ ( .A(_source_stream_matmul_15_source_6_pat_count_1[5:2]), .Y(_10801_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34627_ ( .A({ _10803_, _source_stream_matmul_15_source_6_pat_count_1[32:30] }), .Y(_10802_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34628_ ( .A({ _source_stream_matmul_15_source_6_pat_count_1[28:27], _source_stream_matmul_15_source_6_pat_count_1[25], _source_stream_matmul_15_source_6_pat_count_1[22] }), .Y(_10803_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34629_ ( .A({ _source_stream_matmul_15_source_6_pat_count_1[29], _source_stream_matmul_15_source_6_pat_count_1[26], _source_stream_matmul_15_source_6_pat_count_1[24:23] }), .Y(_10804_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34630_ ( .A({ _10805_, _05785_ }), .Y(_05786_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34631_ ( .A({ _10815_, _10810_, _10808_, _10806_ }), .Y(_10805_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34632_ ( .A({ _10807_, _source_stream_matmul_15_source_6_pat_count_2[32:30] }), .Y(_10806_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34633_ ( .A({ _source_stream_matmul_15_source_6_pat_count_2[28:27], _source_stream_matmul_15_source_6_pat_count_2[25], _source_stream_matmul_15_source_6_pat_count_2[22] }), .Y(_10807_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34634_ ( .A({ _10809_, _source_stream_matmul_15_source_6_pat_count_2[1:0] }), .Y(_10808_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34635_ ( .A(_source_stream_matmul_15_source_6_pat_count_2[5:2]), .Y(_10809_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34636_ ( .A({ _10814_, _10813_, _10812_, _10811_ }), .Y(_10810_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34637_ ( .A(_source_stream_matmul_15_source_6_pat_count_2[13:10]), .Y(_10811_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34638_ ( .A(_source_stream_matmul_15_source_6_pat_count_2[9:6]), .Y(_10812_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34639_ ( .A(_source_stream_matmul_15_source_6_pat_count_2[21:18]), .Y(_10813_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34640_ ( .A(_source_stream_matmul_15_source_6_pat_count_2[17:14]), .Y(_10814_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34641_ ( .A({ _source_stream_matmul_15_source_6_pat_count_2[29], _source_stream_matmul_15_source_6_pat_count_2[26], _source_stream_matmul_15_source_6_pat_count_2[24:23] }), .Y(_10815_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34642_ ( .A({ _05858_, _05023_ }), .Y(_05787_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34643_ ( .A({ _10816_, _10805_, _10794_, _10783_ }), .Y(_05858_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34644_ ( .A({ _10826_, _10821_, _10819_, _10817_ }), .Y(_10816_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34645_ ( .A({ _10818_, _source_stream_matmul_15_source_6_pat_count_3[32:30] }), .Y(_10817_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34646_ ( .A({ _source_stream_matmul_15_source_6_pat_count_3[28:27], _source_stream_matmul_15_source_6_pat_count_3[25], _source_stream_matmul_15_source_6_pat_count_3[22] }), .Y(_10818_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34647_ ( .A({ _10820_, _source_stream_matmul_15_source_6_pat_count_3[1:0] }), .Y(_10819_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34648_ ( .A(_source_stream_matmul_15_source_6_pat_count_3[5:2]), .Y(_10820_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34649_ ( .A({ _10825_, _10824_, _10823_, _10822_ }), .Y(_10821_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34650_ ( .A(_source_stream_matmul_15_source_6_pat_count_3[13:10]), .Y(_10822_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34651_ ( .A(_source_stream_matmul_15_source_6_pat_count_3[9:6]), .Y(_10823_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34652_ ( .A(_source_stream_matmul_15_source_6_pat_count_3[21:18]), .Y(_10824_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34653_ ( .A(_source_stream_matmul_15_source_6_pat_count_3[17:14]), .Y(_10825_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34654_ ( .A({ _source_stream_matmul_15_source_6_pat_count_3[29], _source_stream_matmul_15_source_6_pat_count_3[26], _source_stream_matmul_15_source_6_pat_count_3[24:23] }), .Y(_10826_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34655_ ( .A({ _10827_, _05025_ }), .Y(_05789_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34656_ ( .A({ _10837_, _10836_, _10835_, _10828_ }), .Y(_10827_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34657_ ( .A({ _10834_, _10829_, _source_stream_matmul_15_source_8_pat_count_0[1:0] }), .Y(_10828_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34658_ ( .A({ _10833_, _10832_, _10831_, _10830_ }), .Y(_10829_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34659_ ( .A(_source_stream_matmul_15_source_8_pat_count_0[13:10]), .Y(_10830_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34660_ ( .A(_source_stream_matmul_15_source_8_pat_count_0[9:6]), .Y(_10831_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34661_ ( .A(_source_stream_matmul_15_source_8_pat_count_0[21:18]), .Y(_10832_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34662_ ( .A(_source_stream_matmul_15_source_8_pat_count_0[17:14]), .Y(_10833_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34663_ ( .A(_source_stream_matmul_15_source_8_pat_count_0[5:2]), .Y(_10834_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34664_ ( .A(_source_stream_matmul_15_source_8_pat_count_0[32:30]), .Y(_10835_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34665_ ( .A(_source_stream_matmul_15_source_8_pat_count_0[29:26]), .Y(_10836_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34666_ ( .A(_source_stream_matmul_15_source_8_pat_count_0[25:22]), .Y(_10837_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34667_ ( .A({ _10838_, _05789_ }), .Y(_05790_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34668_ ( .A({ _10848_, _10846_, _10839_ }), .Y(_10838_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34669_ ( .A({ _10845_, _10840_, _source_stream_matmul_15_source_8_pat_count_1[1:0] }), .Y(_10839_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34670_ ( .A({ _10844_, _10843_, _10842_, _10841_ }), .Y(_10840_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34671_ ( .A(_source_stream_matmul_15_source_8_pat_count_1[13:10]), .Y(_10841_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34672_ ( .A(_source_stream_matmul_15_source_8_pat_count_1[9:6]), .Y(_10842_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34673_ ( .A(_source_stream_matmul_15_source_8_pat_count_1[21:18]), .Y(_10843_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34674_ ( .A(_source_stream_matmul_15_source_8_pat_count_1[17:14]), .Y(_10844_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34675_ ( .A(_source_stream_matmul_15_source_8_pat_count_1[5:2]), .Y(_10845_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34676_ ( .A({ _10847_, _source_stream_matmul_15_source_8_pat_count_1[32:30] }), .Y(_10846_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34677_ ( .A({ _source_stream_matmul_15_source_8_pat_count_1[28:27], _source_stream_matmul_15_source_8_pat_count_1[25], _source_stream_matmul_15_source_8_pat_count_1[22] }), .Y(_10847_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34678_ ( .A({ _source_stream_matmul_15_source_8_pat_count_1[29], _source_stream_matmul_15_source_8_pat_count_1[26], _source_stream_matmul_15_source_8_pat_count_1[24:23] }), .Y(_10848_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34679_ ( .A({ _10849_, _05789_ }), .Y(_05791_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34680_ ( .A({ _10859_, _10853_, _10850_, _10838_ }), .Y(_10849_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34681_ ( .A({ _10851_, _source_stream_matmul_15_source_8_pat_count_2[32], _source_stream_matmul_15_source_8_pat_count_2[12], _source_stream_matmul_15_source_8_pat_count_2[6] }), .Y(_10850_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34682_ ( .A({ _10852_, _source_stream_matmul_15_source_8_pat_count_2[17], _source_stream_matmul_15_source_8_pat_count_2[14], _source_stream_matmul_15_source_8_pat_count_2[4] }), .Y(_10851_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34683_ ( .A({ _source_stream_matmul_15_source_8_pat_count_2[21], _source_stream_matmul_15_source_8_pat_count_2[18], _source_stream_matmul_15_source_8_pat_count_2[16:15] }), .Y(_10852_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34684_ ( .A({ _10857_, _10854_, _source_stream_matmul_15_source_8_pat_count_2[2], _source_stream_matmul_15_source_8_pat_count_2[0] }), .Y(_10853_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34685_ ( .A({ _10856_, _10855_, _source_stream_matmul_15_source_8_pat_count_2[10], _source_stream_matmul_15_source_8_pat_count_2[5] }), .Y(_10854_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34686_ ( .A(_source_stream_matmul_15_source_8_pat_count_2[25:23]), .Y(_10855_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34687_ ( .A({ _source_stream_matmul_15_source_8_pat_count_2[13], _source_stream_matmul_15_source_8_pat_count_2[8:7] }), .Y(_10856_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34688_ ( .A({ _10858_, _source_stream_matmul_15_source_8_pat_count_2[29], _source_stream_matmul_15_source_8_pat_count_2[26] }), .Y(_10857_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34689_ ( .A({ _source_stream_matmul_15_source_8_pat_count_2[31:30], _source_stream_matmul_15_source_8_pat_count_2[11], _source_stream_matmul_15_source_8_pat_count_2[9] }), .Y(_10858_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34690_ ( .A({ _10860_, _source_stream_matmul_15_source_8_pat_count_2[27], _source_stream_matmul_15_source_8_pat_count_2[20], _source_stream_matmul_15_source_8_pat_count_2[1] }), .Y(_10859_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34691_ ( .A({ _source_stream_matmul_15_source_8_pat_count_2[28], _source_stream_matmul_15_source_8_pat_count_2[22], _source_stream_matmul_15_source_8_pat_count_2[19], _source_stream_matmul_15_source_8_pat_count_2[3] }), .Y(_10860_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34692_ ( .A({ _10861_, _05791_ }), .Y(_05792_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34693_ ( .A({ _10871_, _10869_, _10862_ }), .Y(_10861_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34694_ ( .A({ _10868_, _10863_, _source_stream_matmul_15_source_8_pat_count_3[1:0] }), .Y(_10862_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34695_ ( .A({ _10867_, _10866_, _10865_, _10864_ }), .Y(_10863_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34696_ ( .A(_source_stream_matmul_15_source_8_pat_count_3[13:10]), .Y(_10864_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34697_ ( .A(_source_stream_matmul_15_source_8_pat_count_3[9:6]), .Y(_10865_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34698_ ( .A(_source_stream_matmul_15_source_8_pat_count_3[21:18]), .Y(_10866_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34699_ ( .A(_source_stream_matmul_15_source_8_pat_count_3[17:14]), .Y(_10867_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34700_ ( .A(_source_stream_matmul_15_source_8_pat_count_3[5:2]), .Y(_10868_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34701_ ( .A({ _10870_, _source_stream_matmul_15_source_8_pat_count_3[32:30] }), .Y(_10869_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34702_ ( .A({ _source_stream_matmul_15_source_8_pat_count_3[28:27], _source_stream_matmul_15_source_8_pat_count_3[25], _source_stream_matmul_15_source_8_pat_count_3[22] }), .Y(_10870_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34703_ ( .A({ _source_stream_matmul_15_source_8_pat_count_3[29], _source_stream_matmul_15_source_8_pat_count_3[26], _source_stream_matmul_15_source_8_pat_count_3[24:23] }), .Y(_10871_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34704_ ( .A({ _10872_, _05021_ }), .Y(_05794_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34705_ ( .A({ _10882_, _10881_, _10880_, _10873_ }), .Y(_10872_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34706_ ( .A({ _10879_, _10874_, _source_stream_matmul_15_source_19_pat_count_0[1:0] }), .Y(_10873_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34707_ ( .A({ _10878_, _10877_, _10876_, _10875_ }), .Y(_10874_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34708_ ( .A(_source_stream_matmul_15_source_19_pat_count_0[13:10]), .Y(_10875_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34709_ ( .A(_source_stream_matmul_15_source_19_pat_count_0[9:6]), .Y(_10876_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34710_ ( .A(_source_stream_matmul_15_source_19_pat_count_0[21:18]), .Y(_10877_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34711_ ( .A(_source_stream_matmul_15_source_19_pat_count_0[17:14]), .Y(_10878_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34712_ ( .A(_source_stream_matmul_15_source_19_pat_count_0[5:2]), .Y(_10879_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34713_ ( .A(_source_stream_matmul_15_source_19_pat_count_0[32:30]), .Y(_10880_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34714_ ( .A(_source_stream_matmul_15_source_19_pat_count_0[29:26]), .Y(_10881_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34715_ ( .A(_source_stream_matmul_15_source_19_pat_count_0[25:22]), .Y(_10882_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34716_ ( .A({ _10883_, _05021_ }), .Y(_05795_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34717_ ( .A({ _10893_, _10891_, _10884_, _10872_ }), .Y(_10883_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34718_ ( .A({ _10890_, _10885_, _source_stream_matmul_15_source_19_pat_count_1[1:0] }), .Y(_10884_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34719_ ( .A({ _10889_, _10888_, _10887_, _10886_ }), .Y(_10885_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34720_ ( .A(_source_stream_matmul_15_source_19_pat_count_1[13:10]), .Y(_10886_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34721_ ( .A(_source_stream_matmul_15_source_19_pat_count_1[9:6]), .Y(_10887_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34722_ ( .A(_source_stream_matmul_15_source_19_pat_count_1[21:18]), .Y(_10888_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34723_ ( .A(_source_stream_matmul_15_source_19_pat_count_1[17:14]), .Y(_10889_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34724_ ( .A(_source_stream_matmul_15_source_19_pat_count_1[5:2]), .Y(_10890_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34725_ ( .A({ _10892_, _source_stream_matmul_15_source_19_pat_count_1[32:30] }), .Y(_10891_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34726_ ( .A({ _source_stream_matmul_15_source_19_pat_count_1[28:27], _source_stream_matmul_15_source_19_pat_count_1[25], _source_stream_matmul_15_source_19_pat_count_1[22] }), .Y(_10892_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34727_ ( .A({ _source_stream_matmul_15_source_19_pat_count_1[29], _source_stream_matmul_15_source_19_pat_count_1[26], _source_stream_matmul_15_source_19_pat_count_1[24:23] }), .Y(_10893_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34728_ ( .A({ _10894_, _05795_ }), .Y(_05796_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34729_ ( .A({ _10904_, _10899_, _10897_, _10895_ }), .Y(_10894_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34730_ ( .A({ _10896_, _source_stream_matmul_15_source_19_pat_count_2[32:30] }), .Y(_10895_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34731_ ( .A({ _source_stream_matmul_15_source_19_pat_count_2[28:27], _source_stream_matmul_15_source_19_pat_count_2[25], _source_stream_matmul_15_source_19_pat_count_2[22] }), .Y(_10896_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34732_ ( .A({ _10898_, _source_stream_matmul_15_source_19_pat_count_2[1:0] }), .Y(_10897_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34733_ ( .A(_source_stream_matmul_15_source_19_pat_count_2[5:2]), .Y(_10898_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34734_ ( .A({ _10903_, _10902_, _10901_, _10900_ }), .Y(_10899_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34735_ ( .A(_source_stream_matmul_15_source_19_pat_count_2[13:10]), .Y(_10900_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34736_ ( .A(_source_stream_matmul_15_source_19_pat_count_2[9:6]), .Y(_10901_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34737_ ( .A(_source_stream_matmul_15_source_19_pat_count_2[21:18]), .Y(_10902_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34738_ ( .A(_source_stream_matmul_15_source_19_pat_count_2[17:14]), .Y(_10903_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34739_ ( .A({ _source_stream_matmul_15_source_19_pat_count_2[29], _source_stream_matmul_15_source_19_pat_count_2[26], _source_stream_matmul_15_source_19_pat_count_2[24:23] }), .Y(_10904_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34740_ ( .A({ _10905_, _05795_ }), .Y(_05797_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34741_ ( .A({ _10916_, _10915_, _10894_, _10906_ }), .Y(_10905_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34742_ ( .A({ _10914_, _10912_, _10907_ }), .Y(_10906_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34743_ ( .A({ _10911_, _10910_, _10908_ }), .Y(_10907_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34744_ ( .A({ _10909_, _source_stream_matmul_15_source_19_pat_count_3[1:0] }), .Y(_10908_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34745_ ( .A(_source_stream_matmul_15_source_19_pat_count_3[5:2]), .Y(_10909_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34746_ ( .A({ _source_stream_matmul_15_source_19_pat_count_3[13], _source_stream_matmul_15_source_19_pat_count_3[10], _source_stream_matmul_15_source_19_pat_count_3[8:7] }), .Y(_10910_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34747_ ( .A({ _source_stream_matmul_15_source_19_pat_count_3[20:19], _source_stream_matmul_15_source_19_pat_count_3[17], _source_stream_matmul_15_source_19_pat_count_3[14] }), .Y(_10911_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34748_ ( .A({ _10913_, _source_stream_matmul_15_source_19_pat_count_3[32:30] }), .Y(_10912_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34749_ ( .A({ _source_stream_matmul_15_source_19_pat_count_3[28:27], _source_stream_matmul_15_source_19_pat_count_3[25], _source_stream_matmul_15_source_19_pat_count_3[22] }), .Y(_10913_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34750_ ( .A({ _source_stream_matmul_15_source_19_pat_count_3[29], _source_stream_matmul_15_source_19_pat_count_3[26], _source_stream_matmul_15_source_19_pat_count_3[24:23] }), .Y(_10914_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34751_ ( .A({ _source_stream_matmul_15_source_19_pat_count_3[12:11], _source_stream_matmul_15_source_19_pat_count_3[9], _source_stream_matmul_15_source_19_pat_count_3[6] }), .Y(_10915_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34752_ ( .A({ _source_stream_matmul_15_source_19_pat_count_3[21], _source_stream_matmul_15_source_19_pat_count_3[18], _source_stream_matmul_15_source_19_pat_count_3[16:15] }), .Y(_10916_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34753_ ( .A({ _10917_, _05020_ }), .Y(_05799_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34754_ ( .A({ _10927_, _10926_, _10925_, _10918_ }), .Y(_10917_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34755_ ( .A({ _10924_, _10919_, _source_stream_matmul_15_source_20_pat_count_0[1:0] }), .Y(_10918_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34756_ ( .A({ _10923_, _10922_, _10921_, _10920_ }), .Y(_10919_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34757_ ( .A(_source_stream_matmul_15_source_20_pat_count_0[13:10]), .Y(_10920_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34758_ ( .A(_source_stream_matmul_15_source_20_pat_count_0[9:6]), .Y(_10921_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34759_ ( .A(_source_stream_matmul_15_source_20_pat_count_0[21:18]), .Y(_10922_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34760_ ( .A(_source_stream_matmul_15_source_20_pat_count_0[17:14]), .Y(_10923_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34761_ ( .A(_source_stream_matmul_15_source_20_pat_count_0[5:2]), .Y(_10924_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34762_ ( .A(_source_stream_matmul_15_source_20_pat_count_0[32:30]), .Y(_10925_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34763_ ( .A(_source_stream_matmul_15_source_20_pat_count_0[29:26]), .Y(_10926_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34764_ ( .A(_source_stream_matmul_15_source_20_pat_count_0[25:22]), .Y(_10927_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34765_ ( .A({ _10928_, _05799_ }), .Y(_05800_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34766_ ( .A({ _10938_, _10936_, _10929_ }), .Y(_10928_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34767_ ( .A({ _10935_, _10930_, _source_stream_matmul_15_source_20_pat_count_1[1:0] }), .Y(_10929_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34768_ ( .A({ _10934_, _10933_, _10932_, _10931_ }), .Y(_10930_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34769_ ( .A(_source_stream_matmul_15_source_20_pat_count_1[13:10]), .Y(_10931_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34770_ ( .A(_source_stream_matmul_15_source_20_pat_count_1[9:6]), .Y(_10932_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34771_ ( .A(_source_stream_matmul_15_source_20_pat_count_1[21:18]), .Y(_10933_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34772_ ( .A(_source_stream_matmul_15_source_20_pat_count_1[17:14]), .Y(_10934_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34773_ ( .A(_source_stream_matmul_15_source_20_pat_count_1[5:2]), .Y(_10935_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34774_ ( .A({ _10937_, _source_stream_matmul_15_source_20_pat_count_1[32:30] }), .Y(_10936_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34775_ ( .A({ _source_stream_matmul_15_source_20_pat_count_1[28:27], _source_stream_matmul_15_source_20_pat_count_1[25], _source_stream_matmul_15_source_20_pat_count_1[22] }), .Y(_10937_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34776_ ( .A({ _source_stream_matmul_15_source_20_pat_count_1[29], _source_stream_matmul_15_source_20_pat_count_1[26], _source_stream_matmul_15_source_20_pat_count_1[24:23] }), .Y(_10938_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34777_ ( .A({ _10939_, _05799_ }), .Y(_05801_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34778_ ( .A({ _10940_, _10928_ }), .Y(_10939_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34779_ ( .A({ _10950_, _10949_, _10948_, _10941_ }), .Y(_10940_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34780_ ( .A({ _10947_, _10942_, _source_stream_matmul_15_source_20_pat_count_2[1:0] }), .Y(_10941_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34781_ ( .A({ _10946_, _10945_, _10944_, _10943_ }), .Y(_10942_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34782_ ( .A(_source_stream_matmul_15_source_20_pat_count_2[13:10]), .Y(_10943_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34783_ ( .A(_source_stream_matmul_15_source_20_pat_count_2[9:6]), .Y(_10944_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34784_ ( .A(_source_stream_matmul_15_source_20_pat_count_2[21:18]), .Y(_10945_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34785_ ( .A(_source_stream_matmul_15_source_20_pat_count_2[17:14]), .Y(_10946_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34786_ ( .A(_source_stream_matmul_15_source_20_pat_count_2[5:2]), .Y(_10947_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34787_ ( .A(_source_stream_matmul_15_source_20_pat_count_2[32:30]), .Y(_10948_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34788_ ( .A(_source_stream_matmul_15_source_20_pat_count_2[29:26]), .Y(_10949_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34789_ ( .A(_source_stream_matmul_15_source_20_pat_count_2[25:22]), .Y(_10950_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34790_ ( .A({ _10951_, _05801_ }), .Y(_05802_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34791_ ( .A({ _10961_, _10959_, _10952_ }), .Y(_10951_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34792_ ( .A({ _10958_, _10953_, _source_stream_matmul_15_source_20_pat_count_3[1:0] }), .Y(_10952_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34793_ ( .A({ _10957_, _10956_, _10955_, _10954_ }), .Y(_10953_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34794_ ( .A(_source_stream_matmul_15_source_20_pat_count_3[13:10]), .Y(_10954_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34795_ ( .A(_source_stream_matmul_15_source_20_pat_count_3[9:6]), .Y(_10955_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34796_ ( .A(_source_stream_matmul_15_source_20_pat_count_3[21:18]), .Y(_10956_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34797_ ( .A(_source_stream_matmul_15_source_20_pat_count_3[17:14]), .Y(_10957_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34798_ ( .A(_source_stream_matmul_15_source_20_pat_count_3[5:2]), .Y(_10958_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34799_ ( .A({ _10960_, _source_stream_matmul_15_source_20_pat_count_3[32:30] }), .Y(_10959_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34800_ ( .A({ _source_stream_matmul_15_source_20_pat_count_3[28:27], _source_stream_matmul_15_source_20_pat_count_3[25], _source_stream_matmul_15_source_20_pat_count_3[22] }), .Y(_10960_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34801_ ( .A({ _source_stream_matmul_15_source_20_pat_count_3[29], _source_stream_matmul_15_source_20_pat_count_3[26], _source_stream_matmul_15_source_20_pat_count_3[24:23] }), .Y(_10961_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34802_ ( .A({ __delay_data_1498, _stream_matmul_15_sink_21_sink_fsm_4[0], _21881_ }), .Y(_05804_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34803_ ( .A({ _stream_matmul_15_start_flag, _04901_ }), .Y(_tmp_1037) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34804_ ( .A({ conv2d_8_mux_dma_flag_0, conv2d_8_mux_dma_pad_mask_0 }), .Y(_05868_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34805_ ( .A({ conv2d_8_mux_dma_flag_1, conv2d_8_mux_dma_pad_mask_1 }), .Y(_05869_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34806_ ( .A({ conv2d_8_mux_dma_flag_2, conv2d_8_mux_dma_pad_mask_2 }), .Y(_05870_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _34807_ ( .A({ conv2d_8_update_filter, _10962_, _03964_, _10969_ }), .Y(_05805_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34808_ ( .A({ _10968_, _10963_ }), .Y(_10962_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34809_ ( .A({ _10967_, _10966_, _10965_, _10964_ }), .Y(_10963_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34810_ ( .A({ _03972_, _03971_, _03970_, _03969_ }), .Y(_10964_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34811_ ( .A({ _03968_, _03967_, _03966_, _03965_ }), .Y(_10965_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34812_ ( .A({ _03986_, _03985_, _03983_, _03982_ }), .Y(_10966_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34813_ ( .A({ _03980_, _03979_, _03977_, _03974_ }), .Y(_10967_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34814_ ( .A({ _03981_, _03978_, _03976_, _03975_ }), .Y(_10968_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34815_ ( .A({ _10972_, _10971_, _10970_ }), .Y(_10969_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34816_ ( .A({ _03963_, _03993_, _03992_ }), .Y(_10970_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34817_ ( .A({ _03991_, _03990_, _03989_, _03988_ }), .Y(_10971_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34818_ ( .A({ _03987_, _03984_, _03973_, _03962_ }), .Y(_10972_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34819_ ( .A({ conv2d_8_mux_next_dma_flag_0, _10973_ }), .Y(_05806_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34820_ ( .A({ _10983_, _10982_, _10978_, _10974_ }), .Y(_10973_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _34821_ ( .A({ _04028_, _10975_, _10977_ }), .Y(_10974_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34822_ ( .A({ _10976_, _04027_, _04057_, _04056_ }), .Y(_10975_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34823_ ( .A({ _04055_, _04052_, _04048_, _04037_ }), .Y(_10976_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34824_ ( .A({ _04054_, _04053_, _04051_, _04026_ }), .Y(_10977_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34825_ ( .A({ _10981_, _10980_, _10979_ }), .Y(_10978_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34826_ ( .A({ _04050_, _04049_, _04047_, _04046_ }), .Y(_10979_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34827_ ( .A({ _04045_, _04044_, _04043_, _04042_ }), .Y(_10980_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34828_ ( .A({ _04041_, _04040_, _04039_, _04038_ }), .Y(_10981_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34829_ ( .A({ _04036_, _04033_, _04031_, _04030_ }), .Y(_10982_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34830_ ( .A({ _04035_, _04034_, _04032_, _04029_ }), .Y(_10983_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _34831_ ( .A({ conv2d_8_mux_next_dma_flag_1, _10984_, _04060_, _10991_ }), .Y(_05807_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34832_ ( .A({ _10990_, _10989_, _10985_ }), .Y(_10984_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34833_ ( .A({ _10988_, _10987_, _10986_ }), .Y(_10985_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34834_ ( .A({ _04082_, _04081_, _04079_, _04078_ }), .Y(_10986_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34835_ ( .A({ _04077_, _04076_, _04075_, _04074_ }), .Y(_10987_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34836_ ( .A({ _04073_, _04072_, _04071_, _04070_ }), .Y(_10988_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34837_ ( .A({ _04068_, _04067_, _04066_, _04065_ }), .Y(_10989_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34838_ ( .A({ _04064_, _04063_, _04062_, _04061_ }), .Y(_10990_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34839_ ( .A({ _10994_, _10993_, _10992_ }), .Y(_10991_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34840_ ( .A({ _04059_, _04089_, _04088_ }), .Y(_10992_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34841_ ( .A({ _04087_, _04086_, _04085_, _04084_ }), .Y(_10993_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34842_ ( .A({ _04083_, _04080_, _04069_, _04058_ }), .Y(_10994_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _34843_ ( .A({ conv2d_8_mux_next_dma_flag_2, _10995_, _04092_, _11002_ }), .Y(_05808_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34844_ ( .A({ _11001_, _11000_, _10996_ }), .Y(_10995_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34845_ ( .A({ _10999_, _10998_, _10997_ }), .Y(_10996_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34846_ ( .A({ _04114_, _04113_, _04111_, _04110_ }), .Y(_10997_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34847_ ( .A({ _04109_, _04108_, _04107_, _04106_ }), .Y(_10998_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34848_ ( .A({ _04105_, _04104_, _04103_, _04102_ }), .Y(_10999_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34849_ ( .A({ _04100_, _04099_, _04098_, _04097_ }), .Y(_11000_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34850_ ( .A({ _04096_, _04095_, _04094_, _04093_ }), .Y(_11001_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34851_ ( .A({ _11005_, _11004_, _11003_ }), .Y(_11002_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34852_ ( .A({ _04091_, _04121_, _04120_ }), .Y(_11003_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34853_ ( .A({ _04119_, _04118_, _04117_, _04116_ }), .Y(_11004_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34854_ ( .A({ _04115_, _04112_, _04101_, _04090_ }), .Y(_11005_) );
  \$lut  #( .LUT(16'h00bf), .WIDTH(4) ) _34855_ ( .A({ conv2d_8_skip_write_out, _11008_, _11016_, _11284_ }), .Y(_05809_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _34856_ ( .A({ cparam_conv2d_8_max_col_count[2], conv2d_8_prev_row_count[2], _11007_ }), .Y(_11006_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _34857_ ( .A({ cparam_conv2d_8_max_col_count[0], cparam_conv2d_8_max_col_count[1], conv2d_8_prev_row_count[0], conv2d_8_prev_row_count[1] }), .Y(_11007_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34858_ ( .A({ _11015_, _11014_, _11009_ }), .Y(_11008_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34859_ ( .A({ _11013_, _11012_, _11011_, _11010_ }), .Y(_11009_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34860_ ( .A(conv2d_8_prev_row_count[23:20]), .Y(_11010_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34861_ ( .A(conv2d_8_prev_row_count[19:16]), .Y(_11011_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34862_ ( .A(conv2d_8_prev_row_count[31:28]), .Y(_11012_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34863_ ( .A(conv2d_8_prev_row_count[27:24]), .Y(_11013_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34864_ ( .A(conv2d_8_prev_row_count[15:12]), .Y(_11014_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34865_ ( .A(conv2d_8_prev_row_count[11:8]), .Y(_11015_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34866_ ( .A(conv2d_8_prev_row_count[7:5]), .Y(_11016_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34867_ ( .A({ _11031_, _11017_, _11008_ }), .Y(_05810_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34868_ ( .A({ _11026_, _11021_, _11018_ }), .Y(_11017_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34869_ ( .A({ _11020_, _11019_, _11016_ }), .Y(_11018_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34870_ ( .A({ conv2d_8_skip_write_out, conv2d_8_prev_och_count[31:29] }), .Y(_11019_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34871_ ( .A(conv2d_8_prev_och_count[28:25]), .Y(_11020_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34872_ ( .A({ _11025_, _11024_, _11023_, _11022_ }), .Y(_11021_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34873_ ( .A(conv2d_8_prev_och_count[16:13]), .Y(_11022_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34874_ ( .A(conv2d_8_prev_och_count[12:9]), .Y(_11023_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34875_ ( .A(conv2d_8_prev_och_count[24:21]), .Y(_11024_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34876_ ( .A(conv2d_8_prev_och_count[20:17]), .Y(_11025_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34877_ ( .A({ _11030_, _11029_, _11028_, _11027_ }), .Y(_11026_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34878_ ( .A({ conv2d_8_prev_och_count[0], conv2d_8_prev_bat_count[31:29] }), .Y(_11027_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34879_ ( .A(conv2d_8_prev_bat_count[28:25]), .Y(_11028_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34880_ ( .A(conv2d_8_prev_och_count[8:5]), .Y(_11029_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34881_ ( .A(conv2d_8_prev_och_count[4:1]), .Y(_11030_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34882_ ( .A({ _11040_, _11039_, _11037_, _11032_ }), .Y(_11031_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34883_ ( .A({ _11036_, _11035_, _11034_, _11033_ }), .Y(_11032_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34884_ ( .A({ conv2d_8_prev_bat_count[16], conv2d_8_prev_bat_count[13], conv2d_8_prev_bat_count[11:10] }), .Y(_11033_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34885_ ( .A({ conv2d_8_prev_bat_count[23:22], conv2d_8_prev_bat_count[20], conv2d_8_prev_bat_count[17] }), .Y(_11034_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34886_ ( .A({ conv2d_8_prev_bat_count[0], conv2d_8_prev_row_count[2:0] }), .Y(_11035_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34887_ ( .A({ conv2d_8_prev_bat_count[8], conv2d_8_prev_bat_count[5], conv2d_8_prev_bat_count[3:2] }), .Y(_11036_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34888_ ( .A({ _11038_, conv2d_8_prev_row_count[4:3] }), .Y(_11037_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34889_ ( .A({ conv2d_8_prev_bat_count[7:6], conv2d_8_prev_bat_count[4], conv2d_8_prev_bat_count[1] }), .Y(_11038_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34890_ ( .A({ conv2d_8_prev_bat_count[15:14], conv2d_8_prev_bat_count[12], conv2d_8_prev_bat_count[9] }), .Y(_11039_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34891_ ( .A({ conv2d_8_prev_bat_count[24], conv2d_8_prev_bat_count[21], conv2d_8_prev_bat_count[19:18] }), .Y(_11040_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34892_ ( .A({ _05262_, _11041_ }), .Y(_05811_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34893_ ( .A({ _11047_, _11046_, _11044_, _11042_ }), .Y(_11041_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34894_ ( .A({ _11043_, _04126_, _04125_ }), .Y(_11042_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34895_ ( .A({ _04130_, _04129_, _04128_, _04127_ }), .Y(_11043_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34896_ ( .A({ _11045_, _04147_, _04146_, _04145_ }), .Y(_11044_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34897_ ( .A({ _04143_, _04142_, _04141_, _04140_ }), .Y(_11045_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34898_ ( .A({ _04139_, _04138_, _04137_, _04136_ }), .Y(_11046_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34899_ ( .A({ _04135_, _04134_, _04132_, _04131_ }), .Y(_11047_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34900_ ( .A({ _09188_, _maxi_read_op_sel[0], _09608_, _maxi_read_op_sel[1] }), .Y(_05812_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34901_ ( .A({ _maxi_read_op_sel[1], _09188_, _09608_, _maxi_read_op_sel[0] }), .Y(_05814_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34902_ ( .A({ _maxi_read_op_sel[1:0], _09608_, _09188_ }), .Y(_05815_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34903_ ( .A({ _09188_, _maxi_read_op_sel[0], _09670_, _maxi_read_op_sel[1] }), .Y(_05817_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34904_ ( .A({ _09670_, _09188_, _maxi_read_op_sel[1:0] }), .Y(_05816_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34905_ ( .A({ _maxi_read_op_sel[1], _09188_, _09670_, _maxi_read_op_sel[0] }), .Y(_05818_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34906_ ( .A({ _maxi_read_op_sel[1:0], _09670_, _09188_ }), .Y(_05819_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34907_ ( .A({ _09602_, _09188_, _maxi_read_op_sel[1:0] }), .Y(_05820_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34908_ ( .A({ _09188_, _maxi_read_op_sel[0], _09602_, _maxi_read_op_sel[1] }), .Y(_05821_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34909_ ( .A({ maxi_rlast, _09188_ }), .Y(_05813_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34910_ ( .A({ _05813_, _11048_ }), .Y(_05822_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34911_ ( .A({ _07419_, _07428_, _07425_, _maxi_read_rest_size[8] }), .Y(_11048_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34912_ ( .A({ _11048_, _05813_ }), .Y(_05823_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34913_ ( .A({ _05902_, conv2d_8_skip_comp }), .Y(_05824_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34914_ ( .A({ cparam_conv2d_8_pad_col_left, _05242_ }), .Y(_05825_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34915_ ( .A({ _stream_conv2d_8_source_6_source_mode[1], _stream_conv2d_8_start }), .Y(_05674_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34916_ ( .A({ _stream_conv2d_8_source_8_source_mode[1], _stream_conv2d_8_start }), .Y(_05679_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34917_ ( .A({ _09890_, _09924_, _09912_ }), .Y(_05827_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34918_ ( .A({ _stream_conv2d_8_source_19_source_mode[1], _stream_conv2d_8_start }), .Y(_05684_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34919_ ( .A({ _09935_, _09969_, _09957_ }), .Y(_05828_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34920_ ( .A({ _stream_conv2d_8_source_20_source_mode[1], _stream_conv2d_8_start }), .Y(_05689_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34921_ ( .A({ _stream_conv2d_8_source_21_source_mode[1], _stream_conv2d_8_start }), .Y(_05694_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34922_ ( .A({ _stream_conv2d_8_source_22_source_mode[1], _stream_conv2d_8_start }), .Y(_05699_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34923_ ( .A({ _stream_conv2d_8_source_23_source_mode[1], _stream_conv2d_8_start }), .Y(_05704_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34924_ ( .A({ _stream_conv2d_8_source_24_source_mode[1], _stream_conv2d_8_start }), .Y(_05709_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34925_ ( .A({ _stream_conv2d_8_source_25_source_mode[1], _stream_conv2d_8_start }), .Y(_05714_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34926_ ( .A({ _stream_conv2d_8_source_26_source_mode[1], _stream_conv2d_8_start }), .Y(_05719_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34927_ ( .A({ _stream_conv2d_8_source_27_source_mode[1], _stream_conv2d_8_start }), .Y(_05724_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34928_ ( .A({ _stream_conv2d_8_source_28_source_mode[1], _stream_conv2d_8_start }), .Y(_05729_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34929_ ( .A({ _stream_conv2d_8_source_29_source_mode[1], _stream_conv2d_8_start }), .Y(_05734_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34930_ ( .A({ _stream_conv2d_8_source_30_source_mode[1], _stream_conv2d_8_start }), .Y(_05739_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34931_ ( .A({ _stream_conv2d_8_source_31_source_mode[1], _stream_conv2d_8_start }), .Y(_05744_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34932_ ( .A({ _10499_, _10464_, _10486_ }), .Y(_05840_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34933_ ( .A({ _stream_conv2d_8_source_32_source_mode[1], _stream_conv2d_8_start }), .Y(_05749_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34934_ ( .A({ _10510_, _10544_, _10532_ }), .Y(_05841_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34935_ ( .A({ _stream_conv2d_8_source_33_source_mode[1], _stream_conv2d_8_start }), .Y(_05754_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34936_ ( .A({ _10590_, _10555_, _10577_ }), .Y(_05842_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34937_ ( .A({ _stream_conv2d_8_source_34_source_mode[1], _stream_conv2d_8_start }), .Y(_05759_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34938_ ( .A({ _10636_, _10601_, _10623_ }), .Y(_05843_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34939_ ( .A({ _stream_conv2d_8_source_35_source_mode[1], _stream_conv2d_8_start }), .Y(_05764_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34940_ ( .A({ _10682_, _10647_, _10669_ }), .Y(_05844_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34941_ ( .A({ _stream_conv2d_8_source_36_source_mode[1], _stream_conv2d_8_start }), .Y(_05769_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34942_ ( .A({ _10726_, _10704_ }), .Y(_05845_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34943_ ( .A({ _stream_conv2d_8_sink_37_sink_mode[0], __stream_conv2d_8_start_46 }), .Y(_05774_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34944_ ( .A({ _11058_, _11057_, _11056_, _11049_ }), .Y(_05846_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34945_ ( .A({ _11055_, _11050_, _stream_conv2d_8_sink_37_sink_count[2:1] }), .Y(_11049_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34946_ ( .A({ _11054_, _11053_, _11052_, _11051_ }), .Y(_11050_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34947_ ( .A(_stream_conv2d_8_sink_37_sink_count[14:11]), .Y(_11051_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34948_ ( .A(_stream_conv2d_8_sink_37_sink_count[10:7]), .Y(_11052_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34949_ ( .A(_stream_conv2d_8_sink_37_sink_count[22:19]), .Y(_11053_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34950_ ( .A(_stream_conv2d_8_sink_37_sink_count[18:15]), .Y(_11054_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34951_ ( .A(_stream_conv2d_8_sink_37_sink_count[6:3]), .Y(_11055_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34952_ ( .A({ _stream_conv2d_8_sink_37_sink_count[0], __delay_data_1371, _stream_conv2d_8_sink_37_sink_count[32:31] }), .Y(_11056_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34953_ ( .A(_stream_conv2d_8_sink_37_sink_count[30:27]), .Y(_11057_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34954_ ( .A(_stream_conv2d_8_sink_37_sink_count[26:23]), .Y(_11058_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34955_ ( .A({ _05263_, _11059_ }), .Y(_05847_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34956_ ( .A({ _11065_, _11064_, _11062_, _11060_ }), .Y(_11059_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34957_ ( .A({ _11061_, _04223_, _04222_ }), .Y(_11060_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34958_ ( .A({ _04227_, _04226_, _04225_, _04224_ }), .Y(_11061_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34959_ ( .A({ _11063_, _04244_, _04243_, _04242_ }), .Y(_11062_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34960_ ( .A({ _04240_, _04239_, _04238_, _04237_ }), .Y(_11063_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34961_ ( .A({ _04236_, _04235_, _04234_, _04233_ }), .Y(_11064_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34962_ ( .A({ _04232_, _04231_, _04229_, _04228_ }), .Y(_11065_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34963_ ( .A({ _maxi_write_data_done, _11066_ }), .Y(_05848_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34964_ ( .A({ _07309_, _07318_, _07315_, _maxi_write_rest_size[8] }), .Y(_11066_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34965_ ( .A({ _maxi_write_data_done, _11066_ }), .Y(_05849_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34966_ ( .A({ _11081_, _11067_ }), .Y(_05851_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34967_ ( .A({ _11080_, _11079_, _11078_, _11068_ }), .Y(_11067_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34968_ ( .A({ _11077_, _11076_, _11074_, _11069_ }), .Y(_11068_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34969_ ( .A({ _11073_, _11072_, _11071_, _11070_ }), .Y(_11069_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34970_ ( .A(max_pool_serial_9_prev_bat_count[16:13]), .Y(_11070_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34971_ ( .A(max_pool_serial_9_prev_bat_count[12:9]), .Y(_11071_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34972_ ( .A(max_pool_serial_9_prev_bat_count[24:21]), .Y(_11072_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34973_ ( .A(max_pool_serial_9_prev_bat_count[20:17]), .Y(_11073_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34974_ ( .A({ _11075_, max_pool_serial_9_prev_row_count[1:0] }), .Y(_11074_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34975_ ( .A({ max_pool_serial_9_prev_bat_count[0], max_pool_serial_9_prev_row_count[4:2] }), .Y(_11075_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34976_ ( .A(max_pool_serial_9_prev_bat_count[8:5]), .Y(_11076_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34977_ ( .A(max_pool_serial_9_prev_bat_count[4:1]), .Y(_11077_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _34978_ ( .A(max_pool_serial_9_prev_row_count[7:5]), .Y(_11078_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34979_ ( .A({ max_pool_serial_9_skip_write_out, max_pool_serial_9_prev_bat_count[31:29] }), .Y(_11079_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34980_ ( .A(max_pool_serial_9_prev_bat_count[28:25]), .Y(_11080_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34981_ ( .A({ _11088_, _11087_, _11082_ }), .Y(_11081_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34982_ ( .A({ _11086_, _11085_, _11084_, _11083_ }), .Y(_11082_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34983_ ( .A(max_pool_serial_9_prev_row_count[23:20]), .Y(_11083_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34984_ ( .A(max_pool_serial_9_prev_row_count[19:16]), .Y(_11084_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34985_ ( .A(max_pool_serial_9_prev_row_count[31:28]), .Y(_11085_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34986_ ( .A(max_pool_serial_9_prev_row_count[27:24]), .Y(_11086_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34987_ ( .A(max_pool_serial_9_prev_row_count[15:12]), .Y(_11087_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34988_ ( .A(max_pool_serial_9_prev_row_count[11:8]), .Y(_11088_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _34989_ ( .A({ max_pool_serial_9_prev_row_count[3], cparam_max_pool_serial_9_max_col_count[3], max_pool_serial_9_prev_row_count[4], cparam_max_pool_serial_9_max_col_count[4] }), .Y(_11089_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _34990_ ( .A({ cparam_max_pool_serial_9_max_col_count[0], cparam_max_pool_serial_9_max_col_count[1], max_pool_serial_9_prev_row_count[0], max_pool_serial_9_prev_row_count[1] }), .Y(_11090_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _34991_ ( .A({ cparam_max_pool_serial_9_max_col_count[2], max_pool_serial_9_prev_row_count[2], cparam_max_pool_serial_9_max_col_count[3], max_pool_serial_9_prev_row_count[3] }), .Y(_11091_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34992_ ( .A({ _08312_, max_pool_serial_9_skip_comp }), .Y(_05852_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34993_ ( .A({ _stream_max_pool_serial_9_source_1_source_mode[1], _stream_max_pool_serial_9_start }), .Y(_05776_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34994_ ( .A({ _stream_max_pool_serial_9_sink_3_sink_mode[0], __stream_max_pool_serial_9_start_10 }), .Y(_05781_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34995_ ( .A({ _10772_, _10738_, _10760_ }), .Y(_05853_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34996_ ( .A({ _11101_, _11100_, _11099_, _11092_ }), .Y(_05854_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34997_ ( .A({ _11098_, _11093_, _stream_max_pool_serial_9_sink_3_sink_count[2:1] }), .Y(_11092_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34998_ ( .A({ _11097_, _11096_, _11095_, _11094_ }), .Y(_11093_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34999_ ( .A(_stream_max_pool_serial_9_sink_3_sink_count[14:11]), .Y(_11094_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35000_ ( .A(_stream_max_pool_serial_9_sink_3_sink_count[10:7]), .Y(_11095_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35001_ ( .A(_stream_max_pool_serial_9_sink_3_sink_count[22:19]), .Y(_11096_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35002_ ( .A(_stream_max_pool_serial_9_sink_3_sink_count[18:15]), .Y(_11097_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35003_ ( .A(_stream_max_pool_serial_9_sink_3_sink_count[6:3]), .Y(_11098_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35004_ ( .A({ _stream_max_pool_serial_9_sink_3_sink_count[0], __substreamoutput_data_774, _stream_max_pool_serial_9_sink_3_sink_count[32:31] }), .Y(_11099_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35005_ ( .A(_stream_max_pool_serial_9_sink_3_sink_count[30:27]), .Y(_11100_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35006_ ( .A(_stream_max_pool_serial_9_sink_3_sink_count[26:23]), .Y(_11101_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _35007_ ( .A({ matmul_15_mux_dma_flag_0, matmul_15_mux_dma_pad_mask_0 }), .Y(_05871_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35008_ ( .A({ _11129_, _11124_, _11116_, _11102_ }), .Y(_05855_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35009_ ( .A({ _11115_, _11110_, _11108_, _11103_ }), .Y(_11102_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35010_ ( .A({ _11107_, _11106_, _11105_, _11104_ }), .Y(_11103_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35011_ ( .A(matmul_15_prev_och_count[23:20]), .Y(_11104_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35012_ ( .A(matmul_15_prev_och_count[19:16]), .Y(_11105_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35013_ ( .A(matmul_15_prev_och_count[31:28]), .Y(_11106_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35014_ ( .A(matmul_15_prev_och_count[27:24]), .Y(_11107_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35015_ ( .A({ matmul_15_skip_write_out, _11109_, matmul_15_prev_och_count[3:2] }), .Y(_11108_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35016_ ( .A({ matmul_15_prev_och_count[1:0], matmul_15_prev_bat_count[31:30] }), .Y(_11109_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35017_ ( .A({ _11114_, _11113_, _11112_, _11111_ }), .Y(_11110_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35018_ ( .A(matmul_15_prev_bat_count[21:18]), .Y(_11111_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35019_ ( .A(matmul_15_prev_bat_count[17:14]), .Y(_11112_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35020_ ( .A(matmul_15_prev_bat_count[29:26]), .Y(_11113_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35021_ ( .A(matmul_15_prev_bat_count[25:22]), .Y(_11114_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35022_ ( .A(matmul_15_prev_och_count[7:4]), .Y(_11115_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35023_ ( .A({ _11123_, _11122_, _11120_, _11117_ }), .Y(_11116_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35024_ ( .A({ _11119_, _11118_ }), .Y(_11117_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35025_ ( .A(matmul_15_prev_och_count[15:12]), .Y(_11118_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35026_ ( .A(matmul_15_prev_och_count[11:8]), .Y(_11119_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _35027_ ( .A({ _11121_, matmul_15_prev_row_count[1:0] }), .Y(_11120_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35028_ ( .A(matmul_15_prev_row_count[5:2]), .Y(_11121_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35029_ ( .A(matmul_15_prev_row_count[13:10]), .Y(_11122_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35030_ ( .A(matmul_15_prev_row_count[9:6]), .Y(_11123_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35031_ ( .A({ _11128_, _11127_, _11126_, _11125_ }), .Y(_11124_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35032_ ( .A(matmul_15_prev_bat_count[5:2]), .Y(_11125_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35033_ ( .A({ matmul_15_prev_bat_count[1:0], matmul_15_prev_row_count[31:30] }), .Y(_11126_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35034_ ( .A(matmul_15_prev_bat_count[13:10]), .Y(_11127_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35035_ ( .A(matmul_15_prev_bat_count[9:6]), .Y(_11128_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35036_ ( .A({ _11133_, _11132_, _11131_, _11130_ }), .Y(_11129_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35037_ ( .A(matmul_15_prev_row_count[21:18]), .Y(_11130_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35038_ ( .A(matmul_15_prev_row_count[17:14]), .Y(_11131_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35039_ ( .A(matmul_15_prev_row_count[29:26]), .Y(_11132_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35040_ ( .A(matmul_15_prev_row_count[25:22]), .Y(_11133_) );
  \$lut  #( .LUT(16'h007f), .WIDTH(4) ) _35041_ ( .A({ matmul_15_skip_write_out, _11134_, _11117_, _11103_ }), .Y(_05856_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _35042_ ( .A({ _11115_, matmul_15_prev_och_count[3], matmul_15_prev_och_count[1], matmul_15_prev_och_count[2] }), .Y(_11134_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35043_ ( .A({ _06622_, matmul_15_skip_comp }), .Y(_05857_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35044_ ( .A({ _stream_matmul_15_source_6_source_mode[1], _stream_matmul_15_start }), .Y(_05783_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35045_ ( .A({ _stream_matmul_15_source_8_source_mode[1], _stream_matmul_15_start }), .Y(_05788_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35046_ ( .A({ _10861_, _10827_, _10849_ }), .Y(_05859_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35047_ ( .A({ _stream_matmul_15_source_19_source_mode[1], _stream_matmul_15_start }), .Y(_05793_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35048_ ( .A({ _10905_, _10883_ }), .Y(_05860_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35049_ ( .A({ _stream_matmul_15_source_20_source_mode[1], _stream_matmul_15_start }), .Y(_05798_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35050_ ( .A({ _10951_, _10917_, _10939_ }), .Y(_05861_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35051_ ( .A({ _stream_matmul_15_sink_21_sink_mode[0], __stream_matmul_15_start_38 }), .Y(_05803_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35052_ ( .A({ _11144_, _11143_, _11142_, _11135_ }), .Y(_05862_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35053_ ( .A({ _11141_, _11136_, _stream_matmul_15_sink_21_sink_count[2:1] }), .Y(_11135_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35054_ ( .A({ _11140_, _11139_, _11138_, _11137_ }), .Y(_11136_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35055_ ( .A(_stream_matmul_15_sink_21_sink_count[14:11]), .Y(_11137_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35056_ ( .A(_stream_matmul_15_sink_21_sink_count[10:7]), .Y(_11138_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35057_ ( .A(_stream_matmul_15_sink_21_sink_count[22:19]), .Y(_11139_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35058_ ( .A(_stream_matmul_15_sink_21_sink_count[18:15]), .Y(_11140_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35059_ ( .A(_stream_matmul_15_sink_21_sink_count[6:3]), .Y(_11141_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35060_ ( .A({ _stream_matmul_15_sink_21_sink_count[0], __delay_data_1498, _stream_matmul_15_sink_21_sink_count[32:31] }), .Y(_11142_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35061_ ( .A(_stream_matmul_15_sink_21_sink_count[30:27]), .Y(_11143_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35062_ ( .A(_stream_matmul_15_sink_21_sink_count[26:23]), .Y(_11144_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _35063_ ( .A(__variable_wdata_174), .Y(_05259_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _35064_ ( .A(__variable_wdata_159), .Y(_05258_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _35065_ ( .A(__variable_wdata_144), .Y(_05257_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _35066_ ( .A(__variable_wdata_129), .Y(_05256_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _35067_ ( .A(__variable_wdata_114), .Y(_05255_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _35068_ ( .A(__variable_wdata_99), .Y(_05254_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _35069_ ( .A(__variable_wdata_84), .Y(_05253_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _35070_ ( .A(__variable_wdata_69), .Y(_05252_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _35071_ ( .A(__variable_wdata_54), .Y(_05251_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _35072_ ( .A({ _11145_, __variable_wdata_1[1:0] }), .Y(_05249_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35073_ ( .A(__variable_wdata_1[5:2]), .Y(_11145_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35074_ ( .A({ _14119_, _06012_ }), .Y(_14120_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35075_ ( .A({ _14079_, _06012_ }), .Y(_14111_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35076_ ( .A({ _14055_, _06012_ }), .Y(_14087_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35077_ ( .A({ _14066_, _06012_ }), .Y(_14098_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35078_ ( .A({ _14077_, _06012_ }), .Y(_14109_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35079_ ( .A({ _14080_, _06012_ }), .Y(_14112_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35080_ ( .A({ _14081_, _06012_ }), .Y(_14113_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35081_ ( .A({ _14082_, _06012_ }), .Y(_14114_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35082_ ( .A({ _14083_, _06012_ }), .Y(_14115_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35083_ ( .A({ _14084_, _06012_ }), .Y(_14116_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35084_ ( .A({ _14085_, _06012_ }), .Y(_14117_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35085_ ( .A({ _14086_, _06012_ }), .Y(_14118_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35086_ ( .A({ _14056_, _06012_ }), .Y(_14088_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35087_ ( .A({ _14057_, _06012_ }), .Y(_14089_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35088_ ( .A({ _14058_, _06012_ }), .Y(_14090_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35089_ ( .A({ _14059_, _06012_ }), .Y(_14091_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35090_ ( .A({ _14060_, _06012_ }), .Y(_14092_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35091_ ( .A({ _14061_, _06012_ }), .Y(_14093_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35092_ ( .A({ _14062_, _06012_ }), .Y(_14094_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35093_ ( .A({ _14063_, _06012_ }), .Y(_14095_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35094_ ( .A({ _14064_, _06012_ }), .Y(_14096_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35095_ ( .A({ _14065_, _06012_ }), .Y(_14097_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35096_ ( .A({ _14067_, _06012_ }), .Y(_14099_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35097_ ( .A({ _14068_, _06012_ }), .Y(_14100_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35098_ ( .A({ _14069_, _06012_ }), .Y(_14101_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35099_ ( .A({ _14070_, _06012_ }), .Y(_14102_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35100_ ( .A({ _14071_, _06012_ }), .Y(_14103_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35101_ ( .A({ _14072_, _06012_ }), .Y(_14104_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35102_ ( .A({ _14073_, _06012_ }), .Y(_14105_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35103_ ( .A({ _14074_, _06012_ }), .Y(_14106_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35104_ ( .A({ _14075_, _06012_ }), .Y(_14107_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35105_ ( .A({ _14076_, _06012_ }), .Y(_14108_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35106_ ( .A({ _14078_, _06012_ }), .Y(_14110_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35107_ ( .A({ _13989_, _06012_ }), .Y(_14021_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35108_ ( .A({ _14000_, _06012_ }), .Y(_14032_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35109_ ( .A({ _14011_, _06012_ }), .Y(_14043_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35110_ ( .A({ _14014_, _06012_ }), .Y(_14046_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35111_ ( .A({ _14015_, _06012_ }), .Y(_14047_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35112_ ( .A({ _14016_, _06012_ }), .Y(_14048_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35113_ ( .A({ _14017_, _06012_ }), .Y(_14049_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35114_ ( .A({ _14018_, _06012_ }), .Y(_14050_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35115_ ( .A({ _14019_, _06012_ }), .Y(_14051_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35116_ ( .A({ _14020_, _06012_ }), .Y(_14052_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35117_ ( .A({ _13990_, _06012_ }), .Y(_14022_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35118_ ( .A({ _13991_, _06012_ }), .Y(_14023_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35119_ ( .A({ _13992_, _06012_ }), .Y(_14024_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35120_ ( .A({ _13993_, _06012_ }), .Y(_14025_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35121_ ( .A({ _13994_, _06012_ }), .Y(_14026_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35122_ ( .A({ _13995_, _06012_ }), .Y(_14027_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35123_ ( .A({ _13996_, _06012_ }), .Y(_14028_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35124_ ( .A({ _13997_, _06012_ }), .Y(_14029_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35125_ ( .A({ _13998_, _06012_ }), .Y(_14030_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35126_ ( .A({ _13999_, _06012_ }), .Y(_14031_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35127_ ( .A({ _14001_, _06012_ }), .Y(_14033_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35128_ ( .A({ _14002_, _06012_ }), .Y(_14034_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35129_ ( .A({ _14003_, _06012_ }), .Y(_14035_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35130_ ( .A({ _14004_, _06012_ }), .Y(_14036_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35131_ ( .A({ _14005_, _06012_ }), .Y(_14037_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35132_ ( .A({ _14006_, _06012_ }), .Y(_14038_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35133_ ( .A({ _14007_, _06012_ }), .Y(_14039_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35134_ ( .A({ _14008_, _06012_ }), .Y(_14040_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35135_ ( .A({ _14009_, _06012_ }), .Y(_14041_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35136_ ( .A({ _14010_, _06012_ }), .Y(_14042_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35137_ ( .A({ _14012_, _06012_ }), .Y(_14044_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35138_ ( .A({ _14013_, _06012_ }), .Y(_14045_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35139_ ( .A({ _14053_, _06012_ }), .Y(_14054_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35140_ ( .A({ _13925_, _06012_ }), .Y(_13957_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35141_ ( .A({ _13936_, _06012_ }), .Y(_13968_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35142_ ( .A({ _13947_, _06012_ }), .Y(_13979_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35143_ ( .A({ _13950_, _06012_ }), .Y(_13982_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35144_ ( .A({ _13951_, _06012_ }), .Y(_13983_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35145_ ( .A({ _13952_, _06012_ }), .Y(_13984_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35146_ ( .A({ _13953_, _06012_ }), .Y(_13985_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35147_ ( .A({ _13954_, _06012_ }), .Y(_13986_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35148_ ( .A({ _13955_, _06012_ }), .Y(_13987_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35149_ ( .A({ _13956_, _06012_ }), .Y(_13988_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35150_ ( .A({ _13926_, _06012_ }), .Y(_13958_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35151_ ( .A({ _13927_, _06012_ }), .Y(_13959_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35152_ ( .A({ _13928_, _06012_ }), .Y(_13960_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35153_ ( .A({ _13929_, _06012_ }), .Y(_13961_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35154_ ( .A({ _13930_, _06012_ }), .Y(_13962_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35155_ ( .A({ _13931_, _06012_ }), .Y(_13963_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35156_ ( .A({ _13932_, _06012_ }), .Y(_13964_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35157_ ( .A({ _13933_, _06012_ }), .Y(_13965_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35158_ ( .A({ _13934_, _06012_ }), .Y(_13966_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35159_ ( .A({ _13935_, _06012_ }), .Y(_13967_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35160_ ( .A({ _13937_, _06012_ }), .Y(_13969_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35161_ ( .A({ _13938_, _06012_ }), .Y(_13970_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35162_ ( .A({ _13939_, _06012_ }), .Y(_13971_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35163_ ( .A({ _13940_, _06012_ }), .Y(_13972_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35164_ ( .A({ _13941_, _06012_ }), .Y(_13973_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35165_ ( .A({ _13942_, _06012_ }), .Y(_13974_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35166_ ( .A({ _13943_, _06012_ }), .Y(_13975_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35167_ ( .A({ _13944_, _06012_ }), .Y(_13976_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35168_ ( .A({ _13945_, _06012_ }), .Y(_13977_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35169_ ( .A({ _13946_, _06012_ }), .Y(_13978_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35170_ ( .A({ _13948_, _06012_ }), .Y(_13980_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35171_ ( .A({ _13949_, _06012_ }), .Y(_13981_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35172_ ( .A({ _18880_, _05909_ }), .Y(_18912_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35173_ ( .A({ _18891_, _05909_ }), .Y(_18923_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35174_ ( .A({ _18902_, _05909_ }), .Y(_18934_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35175_ ( .A({ _18905_, _05909_ }), .Y(_18937_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35176_ ( .A({ _18906_, _05909_ }), .Y(_18938_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35177_ ( .A({ _18907_, _05909_ }), .Y(_18939_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35178_ ( .A({ _18908_, _05909_ }), .Y(_18940_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35179_ ( .A({ _18909_, _05909_ }), .Y(_18941_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35180_ ( .A({ _18910_, _05909_ }), .Y(_18942_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35181_ ( .A({ _18911_, _05909_ }), .Y(_18943_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35182_ ( .A({ _18881_, _05909_ }), .Y(_18913_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35183_ ( .A({ _18882_, _05909_ }), .Y(_18914_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35184_ ( .A({ _18883_, _05909_ }), .Y(_18915_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35185_ ( .A({ _18884_, _05909_ }), .Y(_18916_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35186_ ( .A({ _18885_, _05909_ }), .Y(_18917_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35187_ ( .A({ _18886_, _05909_ }), .Y(_18918_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35188_ ( .A({ _18887_, _05909_ }), .Y(_18919_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35189_ ( .A({ _18888_, _05909_ }), .Y(_18920_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35190_ ( .A({ _18889_, _05909_ }), .Y(_18921_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35191_ ( .A({ _18890_, _05909_ }), .Y(_18922_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35192_ ( .A({ _18892_, _05909_ }), .Y(_18924_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35193_ ( .A({ _18893_, _05909_ }), .Y(_18925_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35194_ ( .A({ _18894_, _05909_ }), .Y(_18926_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35195_ ( .A({ _18895_, _05909_ }), .Y(_18927_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35196_ ( .A({ _18896_, _05909_ }), .Y(_18928_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35197_ ( .A({ _18897_, _05909_ }), .Y(_18929_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35198_ ( .A({ _18898_, _05909_ }), .Y(_18930_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35199_ ( .A({ _18899_, _05909_ }), .Y(_18931_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35200_ ( .A({ _18900_, _05909_ }), .Y(_18932_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35201_ ( .A({ _18901_, _05909_ }), .Y(_18933_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35202_ ( .A({ _18903_, _05909_ }), .Y(_18935_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35203_ ( .A({ _18904_, _05909_ }), .Y(_18936_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35204_ ( .A({ _13921_, _06012_ }), .Y(_13922_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35205_ ( .A({ _13923_, _06012_ }), .Y(_13924_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35206_ ( .A({ _04284_, _05874_ }), .Y(_13887_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35207_ ( .A({ _04295_, _05874_ }), .Y(_13898_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35208_ ( .A({ _04306_, _05874_ }), .Y(_13909_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35209_ ( .A({ _04309_, _05874_ }), .Y(_13912_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35210_ ( .A({ _04310_, _05874_ }), .Y(_13913_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35211_ ( .A({ _04311_, _05874_ }), .Y(_13914_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35212_ ( .A({ _04312_, _05874_ }), .Y(_13915_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35213_ ( .A({ _04313_, _05874_ }), .Y(_13916_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35214_ ( .A({ _04314_, _05874_ }), .Y(_13917_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35215_ ( .A({ _04315_, _05874_ }), .Y(_13918_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35216_ ( .A({ _04285_, _05874_ }), .Y(_13888_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35217_ ( .A({ _04286_, _05874_ }), .Y(_13889_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35218_ ( .A({ _04287_, _05874_ }), .Y(_13890_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35219_ ( .A({ _04288_, _05874_ }), .Y(_13891_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35220_ ( .A({ _04289_, _05874_ }), .Y(_13892_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35221_ ( .A({ _04290_, _05874_ }), .Y(_13893_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35222_ ( .A({ _04291_, _05874_ }), .Y(_13894_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35223_ ( .A({ _04292_, _05874_ }), .Y(_13895_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35224_ ( .A({ _04293_, _05874_ }), .Y(_13896_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35225_ ( .A({ _04294_, _05874_ }), .Y(_13897_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35226_ ( .A({ _04296_, _05874_ }), .Y(_13899_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35227_ ( .A({ _04297_, _05874_ }), .Y(_13900_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35228_ ( .A({ _04298_, _05874_ }), .Y(_13901_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35229_ ( .A({ _04299_, _05874_ }), .Y(_13902_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35230_ ( .A({ _04300_, _05874_ }), .Y(_13903_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35231_ ( .A({ _04301_, _05874_ }), .Y(_13904_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35232_ ( .A({ _04302_, _05874_ }), .Y(_13905_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35233_ ( .A({ _04303_, _05874_ }), .Y(_13906_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35234_ ( .A({ _04304_, _05874_ }), .Y(_13907_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35235_ ( .A({ _04305_, _05874_ }), .Y(_13908_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35236_ ( .A({ _04307_, _05874_ }), .Y(_13910_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35237_ ( .A({ _04308_, _05874_ }), .Y(_13911_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35238_ ( .A({ _13823_, _06479_ }), .Y(_13855_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35239_ ( .A({ _13834_, _06479_ }), .Y(_13866_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35240_ ( .A({ _13845_, _06479_ }), .Y(_13877_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35241_ ( .A({ _13848_, _06479_ }), .Y(_13880_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35242_ ( .A({ _13849_, _06479_ }), .Y(_13881_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35243_ ( .A({ _13850_, _06479_ }), .Y(_13882_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35244_ ( .A({ _13851_, _06479_ }), .Y(_13883_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35245_ ( .A({ _13852_, _06479_ }), .Y(_13884_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35246_ ( .A({ _13853_, _06479_ }), .Y(_13885_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35247_ ( .A({ _13854_, _06479_ }), .Y(_13886_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35248_ ( .A({ _13824_, _06479_ }), .Y(_13856_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35249_ ( .A({ _13825_, _06479_ }), .Y(_13857_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35250_ ( .A({ _13826_, _06479_ }), .Y(_13858_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35251_ ( .A({ _13827_, _06479_ }), .Y(_13859_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35252_ ( .A({ _13828_, _06479_ }), .Y(_13860_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35253_ ( .A({ _13829_, _06479_ }), .Y(_13861_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35254_ ( .A({ _13830_, _06479_ }), .Y(_13862_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35255_ ( .A({ _13831_, _06479_ }), .Y(_13863_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35256_ ( .A({ _13832_, _06479_ }), .Y(_13864_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35257_ ( .A({ _13833_, _06479_ }), .Y(_13865_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35258_ ( .A({ _13835_, _06479_ }), .Y(_13867_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35259_ ( .A({ _13836_, _06479_ }), .Y(_13868_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35260_ ( .A({ _13837_, _06479_ }), .Y(_13869_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35261_ ( .A({ _13838_, _06479_ }), .Y(_13870_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35262_ ( .A({ _13839_, _06479_ }), .Y(_13871_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35263_ ( .A({ _13840_, _06479_ }), .Y(_13872_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35264_ ( .A({ _13841_, _06479_ }), .Y(_13873_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35265_ ( .A({ _13842_, _06479_ }), .Y(_13874_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35266_ ( .A({ _13843_, _06479_ }), .Y(_13875_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35267_ ( .A({ _13844_, _06479_ }), .Y(_13876_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35268_ ( .A({ _13846_, _06479_ }), .Y(_13878_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35269_ ( .A({ _13847_, _06479_ }), .Y(_13879_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35270_ ( .A({ _13695_, _06479_ }), .Y(_13727_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35271_ ( .A({ _13706_, _06479_ }), .Y(_13738_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35272_ ( .A({ _13717_, _06479_ }), .Y(_13749_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35273_ ( .A({ _13720_, _06479_ }), .Y(_13752_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35274_ ( .A({ _13721_, _06479_ }), .Y(_13753_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35275_ ( .A({ _13722_, _06479_ }), .Y(_13754_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35276_ ( .A({ _13723_, _06479_ }), .Y(_13755_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35277_ ( .A({ _13724_, _06479_ }), .Y(_13756_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35278_ ( .A({ _13725_, _06479_ }), .Y(_13757_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35279_ ( .A({ _13726_, _06479_ }), .Y(_13758_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35280_ ( .A({ _13696_, _06479_ }), .Y(_13728_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35281_ ( .A({ _13697_, _06479_ }), .Y(_13729_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35282_ ( .A({ _13698_, _06479_ }), .Y(_13730_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35283_ ( .A({ _13699_, _06479_ }), .Y(_13731_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35284_ ( .A({ _13700_, _06479_ }), .Y(_13732_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35285_ ( .A({ _13701_, _06479_ }), .Y(_13733_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35286_ ( .A({ _13702_, _06479_ }), .Y(_13734_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35287_ ( .A({ _13703_, _06479_ }), .Y(_13735_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35288_ ( .A({ _13704_, _06479_ }), .Y(_13736_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35289_ ( .A({ _13705_, _06479_ }), .Y(_13737_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35290_ ( .A({ _13707_, _06479_ }), .Y(_13739_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35291_ ( .A({ _13708_, _06479_ }), .Y(_13740_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35292_ ( .A({ _13709_, _06479_ }), .Y(_13741_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35293_ ( .A({ _13710_, _06479_ }), .Y(_13742_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35294_ ( .A({ _13711_, _06479_ }), .Y(_13743_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35295_ ( .A({ _13712_, _06479_ }), .Y(_13744_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35296_ ( .A({ _13713_, _06479_ }), .Y(_13745_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35297_ ( .A({ _13714_, _06479_ }), .Y(_13746_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35298_ ( .A({ _13715_, _06479_ }), .Y(_13747_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35299_ ( .A({ _13716_, _06479_ }), .Y(_13748_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35300_ ( .A({ _13718_, _06479_ }), .Y(_13750_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35301_ ( .A({ _13719_, _06479_ }), .Y(_13751_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35302_ ( .A({ _18944_, _05909_ }), .Y(_18976_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35303_ ( .A({ _18955_, _05909_ }), .Y(_18987_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35304_ ( .A({ _18966_, _05909_ }), .Y(_18998_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35305_ ( .A({ _18969_, _05909_ }), .Y(_19001_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35306_ ( .A({ _18970_, _05909_ }), .Y(_19002_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35307_ ( .A({ _18971_, _05909_ }), .Y(_19003_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35308_ ( .A({ _18972_, _05909_ }), .Y(_19004_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35309_ ( .A({ _18973_, _05909_ }), .Y(_19005_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35310_ ( .A({ _18974_, _05909_ }), .Y(_19006_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35311_ ( .A({ _18975_, _05909_ }), .Y(_19007_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35312_ ( .A({ _18945_, _05909_ }), .Y(_18977_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35313_ ( .A({ _18946_, _05909_ }), .Y(_18978_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35314_ ( .A({ _18947_, _05909_ }), .Y(_18979_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35315_ ( .A({ _18948_, _05909_ }), .Y(_18980_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35316_ ( .A({ _18949_, _05909_ }), .Y(_18981_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35317_ ( .A({ _18950_, _05909_ }), .Y(_18982_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35318_ ( .A({ _18951_, _05909_ }), .Y(_18983_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35319_ ( .A({ _18952_, _05909_ }), .Y(_18984_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35320_ ( .A({ _18953_, _05909_ }), .Y(_18985_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35321_ ( .A({ _18954_, _05909_ }), .Y(_18986_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35322_ ( .A({ _18956_, _05909_ }), .Y(_18988_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35323_ ( .A({ _18957_, _05909_ }), .Y(_18989_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35324_ ( .A({ _18958_, _05909_ }), .Y(_18990_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35325_ ( .A({ _18959_, _05909_ }), .Y(_18991_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35326_ ( .A({ _18960_, _05909_ }), .Y(_18992_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35327_ ( .A({ _18961_, _05909_ }), .Y(_18993_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35328_ ( .A({ _18962_, _05909_ }), .Y(_18994_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35329_ ( .A({ _18963_, _05909_ }), .Y(_18995_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35330_ ( .A({ _18964_, _05909_ }), .Y(_18996_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35331_ ( .A({ _18965_, _05909_ }), .Y(_18997_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35332_ ( .A({ _18967_, _05909_ }), .Y(_18999_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35333_ ( .A({ _18968_, _05909_ }), .Y(_19000_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35334_ ( .A({ _13759_, _06479_ }), .Y(_13791_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35335_ ( .A({ _13770_, _06479_ }), .Y(_13802_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35336_ ( .A({ _13781_, _06479_ }), .Y(_13813_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35337_ ( .A({ _13784_, _06479_ }), .Y(_13816_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35338_ ( .A({ _13785_, _06479_ }), .Y(_13817_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35339_ ( .A({ _13786_, _06479_ }), .Y(_13818_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35340_ ( .A({ _13787_, _06479_ }), .Y(_13819_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35341_ ( .A({ _13788_, _06479_ }), .Y(_13820_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35342_ ( .A({ _13789_, _06479_ }), .Y(_13821_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35343_ ( .A({ _13790_, _06479_ }), .Y(_13822_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35344_ ( .A({ _13760_, _06479_ }), .Y(_13792_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35345_ ( .A({ _13761_, _06479_ }), .Y(_13793_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35346_ ( .A({ _13762_, _06479_ }), .Y(_13794_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35347_ ( .A({ _13763_, _06479_ }), .Y(_13795_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35348_ ( .A({ _13764_, _06479_ }), .Y(_13796_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35349_ ( .A({ _13765_, _06479_ }), .Y(_13797_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35350_ ( .A({ _13766_, _06479_ }), .Y(_13798_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35351_ ( .A({ _13767_, _06479_ }), .Y(_13799_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35352_ ( .A({ _13768_, _06479_ }), .Y(_13800_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35353_ ( .A({ _13769_, _06479_ }), .Y(_13801_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35354_ ( .A({ _13771_, _06479_ }), .Y(_13803_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35355_ ( .A({ _13772_, _06479_ }), .Y(_13804_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35356_ ( .A({ _13773_, _06479_ }), .Y(_13805_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35357_ ( .A({ _13774_, _06479_ }), .Y(_13806_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35358_ ( .A({ _13775_, _06479_ }), .Y(_13807_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35359_ ( .A({ _13776_, _06479_ }), .Y(_13808_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35360_ ( .A({ _13777_, _06479_ }), .Y(_13809_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35361_ ( .A({ _13778_, _06479_ }), .Y(_13810_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35362_ ( .A({ _13779_, _06479_ }), .Y(_13811_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35363_ ( .A({ _13780_, _06479_ }), .Y(_13812_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35364_ ( .A({ _13782_, _06479_ }), .Y(_13814_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35365_ ( .A({ _13783_, _06479_ }), .Y(_13815_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35366_ ( .A({ _19008_, _05909_ }), .Y(_19040_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35367_ ( .A({ _19019_, _05909_ }), .Y(_19051_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35368_ ( .A({ _19030_, _05909_ }), .Y(_19062_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35369_ ( .A({ _19033_, _05909_ }), .Y(_19065_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35370_ ( .A({ _19034_, _05909_ }), .Y(_19066_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35371_ ( .A({ _19035_, _05909_ }), .Y(_19067_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35372_ ( .A({ _19036_, _05909_ }), .Y(_19068_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35373_ ( .A({ _19037_, _05909_ }), .Y(_19069_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35374_ ( .A({ _19038_, _05909_ }), .Y(_19070_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35375_ ( .A({ _19039_, _05909_ }), .Y(_19071_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35376_ ( .A({ _19009_, _05909_ }), .Y(_19041_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35377_ ( .A({ _19010_, _05909_ }), .Y(_19042_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35378_ ( .A({ _19011_, _05909_ }), .Y(_19043_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35379_ ( .A({ _19012_, _05909_ }), .Y(_19044_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35380_ ( .A({ _19013_, _05909_ }), .Y(_19045_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35381_ ( .A({ _19014_, _05909_ }), .Y(_19046_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35382_ ( .A({ _19015_, _05909_ }), .Y(_19047_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35383_ ( .A({ _19016_, _05909_ }), .Y(_19048_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35384_ ( .A({ _19017_, _05909_ }), .Y(_19049_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35385_ ( .A({ _19018_, _05909_ }), .Y(_19050_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35386_ ( .A({ _19020_, _05909_ }), .Y(_19052_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35387_ ( .A({ _19021_, _05909_ }), .Y(_19053_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35388_ ( .A({ _19022_, _05909_ }), .Y(_19054_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35389_ ( .A({ _19023_, _05909_ }), .Y(_19055_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35390_ ( .A({ _19024_, _05909_ }), .Y(_19056_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35391_ ( .A({ _19025_, _05909_ }), .Y(_19057_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35392_ ( .A({ _19026_, _05909_ }), .Y(_19058_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35393_ ( .A({ _19027_, _05909_ }), .Y(_19059_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35394_ ( .A({ _19028_, _05909_ }), .Y(_19060_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35395_ ( .A({ _19029_, _05909_ }), .Y(_19061_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35396_ ( .A({ _19031_, _05909_ }), .Y(_19063_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35397_ ( .A({ _19032_, _05909_ }), .Y(_19064_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35398_ ( .A({ _19072_, _05909_ }), .Y(_19104_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35399_ ( .A({ _19083_, _05909_ }), .Y(_19115_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35400_ ( .A({ _19094_, _05909_ }), .Y(_19126_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35401_ ( .A({ _19097_, _05909_ }), .Y(_19129_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35402_ ( .A({ _19098_, _05909_ }), .Y(_19130_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35403_ ( .A({ _19099_, _05909_ }), .Y(_19131_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35404_ ( .A({ _19100_, _05909_ }), .Y(_19132_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35405_ ( .A({ _19101_, _05909_ }), .Y(_19133_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35406_ ( .A({ _19102_, _05909_ }), .Y(_19134_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35407_ ( .A({ _19103_, _05909_ }), .Y(_19135_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35408_ ( .A({ _19073_, _05909_ }), .Y(_19105_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35409_ ( .A({ _19074_, _05909_ }), .Y(_19106_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35410_ ( .A({ _19075_, _05909_ }), .Y(_19107_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35411_ ( .A({ _19076_, _05909_ }), .Y(_19108_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35412_ ( .A({ _19077_, _05909_ }), .Y(_19109_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35413_ ( .A({ _19078_, _05909_ }), .Y(_19110_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35414_ ( .A({ _19079_, _05909_ }), .Y(_19111_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35415_ ( .A({ _19080_, _05909_ }), .Y(_19112_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35416_ ( .A({ _19081_, _05909_ }), .Y(_19113_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35417_ ( .A({ _19082_, _05909_ }), .Y(_19114_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35418_ ( .A({ _19084_, _05909_ }), .Y(_19116_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35419_ ( .A({ _19085_, _05909_ }), .Y(_19117_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35420_ ( .A({ _19086_, _05909_ }), .Y(_19118_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35421_ ( .A({ _19087_, _05909_ }), .Y(_19119_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35422_ ( .A({ _19088_, _05909_ }), .Y(_19120_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35423_ ( .A({ _19089_, _05909_ }), .Y(_19121_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35424_ ( .A({ _19090_, _05909_ }), .Y(_19122_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35425_ ( .A({ _19091_, _05909_ }), .Y(_19123_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35426_ ( .A({ _19092_, _05909_ }), .Y(_19124_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35427_ ( .A({ _19093_, _05909_ }), .Y(_19125_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35428_ ( .A({ _19095_, _05909_ }), .Y(_19127_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35429_ ( .A({ _19096_, _05909_ }), .Y(_19128_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35430_ ( .A({ _19136_, _05909_ }), .Y(_19168_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35431_ ( .A({ _19147_, _05909_ }), .Y(_19179_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35432_ ( .A({ _19158_, _05909_ }), .Y(_19190_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35433_ ( .A({ _19161_, _05909_ }), .Y(_19193_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35434_ ( .A({ _19162_, _05909_ }), .Y(_19194_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35435_ ( .A({ _19163_, _05909_ }), .Y(_19195_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35436_ ( .A({ _19164_, _05909_ }), .Y(_19196_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35437_ ( .A({ _19165_, _05909_ }), .Y(_19197_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35438_ ( .A({ _19166_, _05909_ }), .Y(_19198_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35439_ ( .A({ _19167_, _05909_ }), .Y(_19199_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35440_ ( .A({ _19137_, _05909_ }), .Y(_19169_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35441_ ( .A({ _19138_, _05909_ }), .Y(_19170_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35442_ ( .A({ _19139_, _05909_ }), .Y(_19171_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35443_ ( .A({ _19140_, _05909_ }), .Y(_19172_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35444_ ( .A({ _19141_, _05909_ }), .Y(_19173_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35445_ ( .A({ _19142_, _05909_ }), .Y(_19174_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35446_ ( .A({ _19143_, _05909_ }), .Y(_19175_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35447_ ( .A({ _19144_, _05909_ }), .Y(_19176_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35448_ ( .A({ _19145_, _05909_ }), .Y(_19177_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35449_ ( .A({ _19146_, _05909_ }), .Y(_19178_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35450_ ( .A({ _19148_, _05909_ }), .Y(_19180_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35451_ ( .A({ _19149_, _05909_ }), .Y(_19181_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35452_ ( .A({ _19150_, _05909_ }), .Y(_19182_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35453_ ( .A({ _19151_, _05909_ }), .Y(_19183_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35454_ ( .A({ _19152_, _05909_ }), .Y(_19184_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35455_ ( .A({ _19153_, _05909_ }), .Y(_19185_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35456_ ( .A({ _19154_, _05909_ }), .Y(_19186_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35457_ ( .A({ _19155_, _05909_ }), .Y(_19187_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35458_ ( .A({ _19156_, _05909_ }), .Y(_19188_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35459_ ( .A({ _19157_, _05909_ }), .Y(_19189_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35460_ ( .A({ _19159_, _05909_ }), .Y(_19191_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35461_ ( .A({ _19160_, _05909_ }), .Y(_19192_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35462_ ( .A({ _19200_, _05909_ }), .Y(_19232_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35463_ ( .A({ _19211_, _05909_ }), .Y(_19243_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35464_ ( .A({ _19222_, _05909_ }), .Y(_19254_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35465_ ( .A({ _19225_, _05909_ }), .Y(_19257_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35466_ ( .A({ _19226_, _05909_ }), .Y(_19258_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35467_ ( .A({ _19227_, _05909_ }), .Y(_19259_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35468_ ( .A({ _19228_, _05909_ }), .Y(_19260_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35469_ ( .A({ _19229_, _05909_ }), .Y(_19261_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35470_ ( .A({ _19230_, _05909_ }), .Y(_19262_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35471_ ( .A({ _19231_, _05909_ }), .Y(_19263_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35472_ ( .A({ _19201_, _05909_ }), .Y(_19233_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35473_ ( .A({ _19202_, _05909_ }), .Y(_19234_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35474_ ( .A({ _19203_, _05909_ }), .Y(_19235_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35475_ ( .A({ _19204_, _05909_ }), .Y(_19236_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35476_ ( .A({ _19205_, _05909_ }), .Y(_19237_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35477_ ( .A({ _19206_, _05909_ }), .Y(_19238_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35478_ ( .A({ _19207_, _05909_ }), .Y(_19239_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35479_ ( .A({ _19208_, _05909_ }), .Y(_19240_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35480_ ( .A({ _19209_, _05909_ }), .Y(_19241_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35481_ ( .A({ _19210_, _05909_ }), .Y(_19242_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35482_ ( .A({ _19212_, _05909_ }), .Y(_19244_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35483_ ( .A({ _19213_, _05909_ }), .Y(_19245_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35484_ ( .A({ _19214_, _05909_ }), .Y(_19246_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35485_ ( .A({ _19215_, _05909_ }), .Y(_19247_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35486_ ( .A({ _19216_, _05909_ }), .Y(_19248_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35487_ ( .A({ _19217_, _05909_ }), .Y(_19249_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35488_ ( .A({ _19218_, _05909_ }), .Y(_19250_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35489_ ( .A({ _19219_, _05909_ }), .Y(_19251_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35490_ ( .A({ _19220_, _05909_ }), .Y(_19252_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35491_ ( .A({ _19221_, _05909_ }), .Y(_19253_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35492_ ( .A({ _19223_, _05909_ }), .Y(_19255_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35493_ ( .A({ _19224_, _05909_ }), .Y(_19256_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35494_ ( .A({ _19264_, _05909_ }), .Y(_19266_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35495_ ( .A({ _19265_, _05909_ }), .Y(_19267_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35496_ ( .A({ _04380_, _11896_ }), .Y(_12767_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35497_ ( .A({ _04391_, _11896_ }), .Y(_12778_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35498_ ( .A({ _04402_, _11896_ }), .Y(_12789_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35499_ ( .A({ _04405_, _11896_ }), .Y(_12792_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35500_ ( .A({ _04406_, _11896_ }), .Y(_12793_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35501_ ( .A({ _04407_, _11896_ }), .Y(_12794_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35502_ ( .A({ _04408_, _11896_ }), .Y(_12795_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35503_ ( .A({ _04409_, _11896_ }), .Y(_12796_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35504_ ( .A({ _04410_, _11896_ }), .Y(_12797_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35505_ ( .A({ _04411_, _11896_ }), .Y(_12798_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35506_ ( .A({ _04381_, _11896_ }), .Y(_12768_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35507_ ( .A({ _04382_, _11896_ }), .Y(_12769_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35508_ ( .A({ _04383_, _11896_ }), .Y(_12770_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35509_ ( .A({ _04384_, _11896_ }), .Y(_12771_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35510_ ( .A({ _04385_, _11896_ }), .Y(_12772_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35511_ ( .A({ _04386_, _11896_ }), .Y(_12773_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35512_ ( .A({ _04387_, _11896_ }), .Y(_12774_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35513_ ( .A({ _04388_, _11896_ }), .Y(_12775_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35514_ ( .A({ _04389_, _11896_ }), .Y(_12776_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35515_ ( .A({ _04390_, _11896_ }), .Y(_12777_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35516_ ( .A({ _04392_, _11896_ }), .Y(_12779_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35517_ ( .A({ _04393_, _11896_ }), .Y(_12780_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35518_ ( .A({ _04394_, _11896_ }), .Y(_12781_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35519_ ( .A({ _04395_, _11896_ }), .Y(_12782_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35520_ ( .A({ _04396_, _11896_ }), .Y(_12783_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35521_ ( .A({ _04397_, _11896_ }), .Y(_12784_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35522_ ( .A({ _04398_, _11896_ }), .Y(_12785_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35523_ ( .A({ _04399_, _11896_ }), .Y(_12786_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35524_ ( .A({ _04400_, _11896_ }), .Y(_12787_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35525_ ( .A({ _04401_, _11896_ }), .Y(_12788_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35526_ ( .A({ _04403_, _11896_ }), .Y(_12790_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35527_ ( .A({ _04404_, _11896_ }), .Y(_12791_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35528_ ( .A({ conv2d_8_och_count[0], _05909_ }), .Y(_19268_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35529_ ( .A({ conv2d_8_och_count[1], _05909_ }), .Y(_19279_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35530_ ( .A({ conv2d_8_och_count[2], _05909_ }), .Y(_19290_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35531_ ( .A({ conv2d_8_och_count[3], _05909_ }), .Y(_19293_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35532_ ( .A({ conv2d_8_och_count[4], _05909_ }), .Y(_19294_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35533_ ( .A({ conv2d_8_och_count[5], _05909_ }), .Y(_19295_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35534_ ( .A({ conv2d_8_och_count[6], _05909_ }), .Y(_19296_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35535_ ( .A({ conv2d_8_och_count[7], _05909_ }), .Y(_19297_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35536_ ( .A({ conv2d_8_och_count[8], _05909_ }), .Y(_19298_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35537_ ( .A({ conv2d_8_och_count[9], _05909_ }), .Y(_19299_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35538_ ( .A({ conv2d_8_och_count[10], _05909_ }), .Y(_19269_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35539_ ( .A({ conv2d_8_och_count[11], _05909_ }), .Y(_19270_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35540_ ( .A({ conv2d_8_och_count[12], _05909_ }), .Y(_19271_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35541_ ( .A({ conv2d_8_och_count[13], _05909_ }), .Y(_19272_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35542_ ( .A({ conv2d_8_och_count[14], _05909_ }), .Y(_19273_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35543_ ( .A({ conv2d_8_och_count[15], _05909_ }), .Y(_19274_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35544_ ( .A({ conv2d_8_och_count[16], _05909_ }), .Y(_19275_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35545_ ( .A({ conv2d_8_och_count[17], _05909_ }), .Y(_19276_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35546_ ( .A({ conv2d_8_och_count[18], _05909_ }), .Y(_19277_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35547_ ( .A({ conv2d_8_och_count[19], _05909_ }), .Y(_19278_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35548_ ( .A({ conv2d_8_och_count[20], _05909_ }), .Y(_19280_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35549_ ( .A({ conv2d_8_och_count[21], _05909_ }), .Y(_19281_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35550_ ( .A({ conv2d_8_och_count[22], _05909_ }), .Y(_19282_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35551_ ( .A({ conv2d_8_och_count[23], _05909_ }), .Y(_19283_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35552_ ( .A({ conv2d_8_och_count[24], _05909_ }), .Y(_19284_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35553_ ( .A({ conv2d_8_och_count[25], _05909_ }), .Y(_19285_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35554_ ( .A({ conv2d_8_och_count[26], _05909_ }), .Y(_19286_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35555_ ( .A({ conv2d_8_och_count[27], _05909_ }), .Y(_19287_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35556_ ( .A({ conv2d_8_och_count[28], _05909_ }), .Y(_19288_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35557_ ( .A({ conv2d_8_och_count[29], _05909_ }), .Y(_19289_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35558_ ( .A({ conv2d_8_och_count[30], _05909_ }), .Y(_19291_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35559_ ( .A({ conv2d_8_och_count[31], _05909_ }), .Y(_19292_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35560_ ( .A({ _12607_, _11896_ }), .Y(_12639_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35561_ ( .A({ _12618_, _11896_ }), .Y(_12650_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35562_ ( .A({ _12629_, _11896_ }), .Y(_12661_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35563_ ( .A({ _12632_, _11896_ }), .Y(_12664_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35564_ ( .A({ _12633_, _11896_ }), .Y(_12665_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35565_ ( .A({ _12634_, _11896_ }), .Y(_12666_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35566_ ( .A({ _12635_, _11896_ }), .Y(_12667_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35567_ ( .A({ _12636_, _11896_ }), .Y(_12668_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35568_ ( .A({ _12637_, _11896_ }), .Y(_12669_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35569_ ( .A({ _12638_, _11896_ }), .Y(_12670_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35570_ ( .A({ _12608_, _11896_ }), .Y(_12640_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35571_ ( .A({ _12609_, _11896_ }), .Y(_12641_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35572_ ( .A({ _12610_, _11896_ }), .Y(_12642_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35573_ ( .A({ _12611_, _11896_ }), .Y(_12643_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35574_ ( .A({ _12612_, _11896_ }), .Y(_12644_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35575_ ( .A({ _12613_, _11896_ }), .Y(_12645_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35576_ ( .A({ _12614_, _11896_ }), .Y(_12646_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35577_ ( .A({ _12615_, _11896_ }), .Y(_12647_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35578_ ( .A({ _12616_, _11896_ }), .Y(_12648_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35579_ ( .A({ _12617_, _11896_ }), .Y(_12649_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35580_ ( .A({ _12619_, _11896_ }), .Y(_12651_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35581_ ( .A({ _12620_, _11896_ }), .Y(_12652_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35582_ ( .A({ _12621_, _11896_ }), .Y(_12653_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35583_ ( .A({ _12622_, _11896_ }), .Y(_12654_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35584_ ( .A({ _12623_, _11896_ }), .Y(_12655_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35585_ ( .A({ _12624_, _11896_ }), .Y(_12656_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35586_ ( .A({ _12625_, _11896_ }), .Y(_12657_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35587_ ( .A({ _12626_, _11896_ }), .Y(_12658_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35588_ ( .A({ _12627_, _11896_ }), .Y(_12659_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35589_ ( .A({ _12628_, _11896_ }), .Y(_12660_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35590_ ( .A({ _12630_, _11896_ }), .Y(_12662_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35591_ ( .A({ _12631_, _11896_ }), .Y(_12663_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35592_ ( .A({ _12671_, _11896_ }), .Y(_12703_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35593_ ( .A({ _12682_, _11896_ }), .Y(_12714_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35594_ ( .A({ _12693_, _11896_ }), .Y(_12725_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35595_ ( .A({ _12696_, _11896_ }), .Y(_12728_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35596_ ( .A({ _12697_, _11896_ }), .Y(_12729_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35597_ ( .A({ _12698_, _11896_ }), .Y(_12730_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35598_ ( .A({ _12699_, _11896_ }), .Y(_12731_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35599_ ( .A({ _12700_, _11896_ }), .Y(_12732_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35600_ ( .A({ _12701_, _11896_ }), .Y(_12733_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35601_ ( .A({ _12702_, _11896_ }), .Y(_12734_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35602_ ( .A({ _12672_, _11896_ }), .Y(_12704_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35603_ ( .A({ _12673_, _11896_ }), .Y(_12705_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35604_ ( .A({ _12674_, _11896_ }), .Y(_12706_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35605_ ( .A({ _12675_, _11896_ }), .Y(_12707_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35606_ ( .A({ _12676_, _11896_ }), .Y(_12708_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35607_ ( .A({ _12677_, _11896_ }), .Y(_12709_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35608_ ( .A({ _12678_, _11896_ }), .Y(_12710_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35609_ ( .A({ _12679_, _11896_ }), .Y(_12711_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35610_ ( .A({ _12680_, _11896_ }), .Y(_12712_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35611_ ( .A({ _12681_, _11896_ }), .Y(_12713_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35612_ ( .A({ _12683_, _11896_ }), .Y(_12715_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35613_ ( .A({ _12684_, _11896_ }), .Y(_12716_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35614_ ( .A({ _12685_, _11896_ }), .Y(_12717_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35615_ ( .A({ _12686_, _11896_ }), .Y(_12718_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35616_ ( .A({ _12687_, _11896_ }), .Y(_12719_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35617_ ( .A({ _12688_, _11896_ }), .Y(_12720_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35618_ ( .A({ _12689_, _11896_ }), .Y(_12721_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35619_ ( .A({ _12690_, _11896_ }), .Y(_12722_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35620_ ( .A({ _12691_, _11896_ }), .Y(_12723_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35621_ ( .A({ _12692_, _11896_ }), .Y(_12724_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35622_ ( .A({ _12694_, _11896_ }), .Y(_12726_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35623_ ( .A({ _12695_, _11896_ }), .Y(_12727_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35624_ ( .A({ conv2d_8_bat_count[0], _05909_ }), .Y(_19300_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35625_ ( .A({ conv2d_8_bat_count[1], _05909_ }), .Y(_19311_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35626_ ( .A({ conv2d_8_bat_count[2], _05909_ }), .Y(_19322_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35627_ ( .A({ conv2d_8_bat_count[3], _05909_ }), .Y(_19325_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35628_ ( .A({ conv2d_8_bat_count[4], _05909_ }), .Y(_19326_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35629_ ( .A({ conv2d_8_bat_count[5], _05909_ }), .Y(_19327_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35630_ ( .A({ conv2d_8_bat_count[6], _05909_ }), .Y(_19328_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35631_ ( .A({ conv2d_8_bat_count[7], _05909_ }), .Y(_19329_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35632_ ( .A({ conv2d_8_bat_count[8], _05909_ }), .Y(_19330_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35633_ ( .A({ conv2d_8_bat_count[9], _05909_ }), .Y(_19331_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35634_ ( .A({ conv2d_8_bat_count[10], _05909_ }), .Y(_19301_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35635_ ( .A({ conv2d_8_bat_count[11], _05909_ }), .Y(_19302_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35636_ ( .A({ conv2d_8_bat_count[12], _05909_ }), .Y(_19303_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35637_ ( .A({ conv2d_8_bat_count[13], _05909_ }), .Y(_19304_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35638_ ( .A({ conv2d_8_bat_count[14], _05909_ }), .Y(_19305_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35639_ ( .A({ conv2d_8_bat_count[15], _05909_ }), .Y(_19306_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35640_ ( .A({ conv2d_8_bat_count[16], _05909_ }), .Y(_19307_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35641_ ( .A({ conv2d_8_bat_count[17], _05909_ }), .Y(_19308_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35642_ ( .A({ conv2d_8_bat_count[18], _05909_ }), .Y(_19309_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35643_ ( .A({ conv2d_8_bat_count[19], _05909_ }), .Y(_19310_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35644_ ( .A({ conv2d_8_bat_count[20], _05909_ }), .Y(_19312_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35645_ ( .A({ conv2d_8_bat_count[21], _05909_ }), .Y(_19313_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35646_ ( .A({ conv2d_8_bat_count[22], _05909_ }), .Y(_19314_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35647_ ( .A({ conv2d_8_bat_count[23], _05909_ }), .Y(_19315_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35648_ ( .A({ conv2d_8_bat_count[24], _05909_ }), .Y(_19316_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35649_ ( .A({ conv2d_8_bat_count[25], _05909_ }), .Y(_19317_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35650_ ( .A({ conv2d_8_bat_count[26], _05909_ }), .Y(_19318_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35651_ ( .A({ conv2d_8_bat_count[27], _05909_ }), .Y(_19319_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35652_ ( .A({ conv2d_8_bat_count[28], _05909_ }), .Y(_19320_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35653_ ( .A({ conv2d_8_bat_count[29], _05909_ }), .Y(_19321_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35654_ ( .A({ conv2d_8_bat_count[30], _05909_ }), .Y(_19323_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35655_ ( .A({ conv2d_8_bat_count[31], _05909_ }), .Y(_19324_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35656_ ( .A({ _12543_, _11896_ }), .Y(_12575_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35657_ ( .A({ _12554_, _11896_ }), .Y(_12586_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35658_ ( .A({ _12565_, _11896_ }), .Y(_12597_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35659_ ( .A({ _12568_, _11896_ }), .Y(_12600_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35660_ ( .A({ _12569_, _11896_ }), .Y(_12601_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35661_ ( .A({ _12570_, _11896_ }), .Y(_12602_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35662_ ( .A({ _12571_, _11896_ }), .Y(_12603_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35663_ ( .A({ _12572_, _11896_ }), .Y(_12604_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35664_ ( .A({ _12573_, _11896_ }), .Y(_12605_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35665_ ( .A({ _12574_, _11896_ }), .Y(_12606_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35666_ ( .A({ _12544_, _11896_ }), .Y(_12576_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35667_ ( .A({ _12545_, _11896_ }), .Y(_12577_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35668_ ( .A({ _12546_, _11896_ }), .Y(_12578_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35669_ ( .A({ _12547_, _11896_ }), .Y(_12579_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35670_ ( .A({ _12548_, _11896_ }), .Y(_12580_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35671_ ( .A({ _12549_, _11896_ }), .Y(_12581_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35672_ ( .A({ _12550_, _11896_ }), .Y(_12582_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35673_ ( .A({ _12551_, _11896_ }), .Y(_12583_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35674_ ( .A({ _12552_, _11896_ }), .Y(_12584_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35675_ ( .A({ _12553_, _11896_ }), .Y(_12585_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35676_ ( .A({ _12555_, _11896_ }), .Y(_12587_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35677_ ( .A({ _12556_, _11896_ }), .Y(_12588_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35678_ ( .A({ _12557_, _11896_ }), .Y(_12589_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35679_ ( .A({ _12558_, _11896_ }), .Y(_12590_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35680_ ( .A({ _12559_, _11896_ }), .Y(_12591_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35681_ ( .A({ _12560_, _11896_ }), .Y(_12592_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35682_ ( .A({ _12561_, _11896_ }), .Y(_12593_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35683_ ( .A({ _12562_, _11896_ }), .Y(_12594_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35684_ ( .A({ _12563_, _11896_ }), .Y(_12595_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35685_ ( .A({ _12564_, _11896_ }), .Y(_12596_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35686_ ( .A({ _12566_, _11896_ }), .Y(_12598_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35687_ ( .A({ _12567_, _11896_ }), .Y(_12599_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35688_ ( .A({ _18552_, _05909_ }), .Y(_18553_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35689_ ( .A({ _12479_, _06611_ }), .Y(_12511_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35690_ ( .A({ _12490_, _06611_ }), .Y(_12522_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35691_ ( .A({ _12501_, _06611_ }), .Y(_12533_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35692_ ( .A({ _12504_, _06611_ }), .Y(_12536_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35693_ ( .A({ _12505_, _06611_ }), .Y(_12537_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35694_ ( .A({ _12506_, _06611_ }), .Y(_12538_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35695_ ( .A({ _12507_, _06611_ }), .Y(_12539_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35696_ ( .A({ _12508_, _06611_ }), .Y(_12540_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35697_ ( .A({ _12509_, _06611_ }), .Y(_12541_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35698_ ( .A({ _12510_, _06611_ }), .Y(_12542_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35699_ ( .A({ _12480_, _06611_ }), .Y(_12512_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35700_ ( .A({ _12481_, _06611_ }), .Y(_12513_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35701_ ( .A({ _12482_, _06611_ }), .Y(_12514_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35702_ ( .A({ _12483_, _06611_ }), .Y(_12515_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35703_ ( .A({ _12484_, _06611_ }), .Y(_12516_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35704_ ( .A({ _12485_, _06611_ }), .Y(_12517_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35705_ ( .A({ _12486_, _06611_ }), .Y(_12518_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35706_ ( .A({ _12487_, _06611_ }), .Y(_12519_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35707_ ( .A({ _12488_, _06611_ }), .Y(_12520_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35708_ ( .A({ _12489_, _06611_ }), .Y(_12521_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35709_ ( .A({ _12491_, _06611_ }), .Y(_12523_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35710_ ( .A({ _12492_, _06611_ }), .Y(_12524_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35711_ ( .A({ _12493_, _06611_ }), .Y(_12525_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35712_ ( .A({ _12494_, _06611_ }), .Y(_12526_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35713_ ( .A({ _12495_, _06611_ }), .Y(_12527_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35714_ ( .A({ _12496_, _06611_ }), .Y(_12528_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35715_ ( .A({ _12497_, _06611_ }), .Y(_12529_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35716_ ( .A({ _12498_, _06611_ }), .Y(_12530_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35717_ ( .A({ _12499_, _06611_ }), .Y(_12531_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35718_ ( .A({ _12500_, _06611_ }), .Y(_12532_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35719_ ( .A({ _12502_, _06611_ }), .Y(_12534_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35720_ ( .A({ _12503_, _06611_ }), .Y(_12535_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35721_ ( .A({ _04412_, _11896_ }), .Y(_12447_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35722_ ( .A({ _04423_, _11896_ }), .Y(_12458_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35723_ ( .A({ _04434_, _11896_ }), .Y(_12469_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35724_ ( .A({ _04437_, _11896_ }), .Y(_12472_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35725_ ( .A({ _04438_, _11896_ }), .Y(_12473_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35726_ ( .A({ _04439_, _11896_ }), .Y(_12474_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35727_ ( .A({ _04440_, _11896_ }), .Y(_12475_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35728_ ( .A({ _04441_, _11896_ }), .Y(_12476_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35729_ ( .A({ _04442_, _11896_ }), .Y(_12477_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35730_ ( .A({ _04443_, _11896_ }), .Y(_12478_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35731_ ( .A({ _04413_, _11896_ }), .Y(_12448_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35732_ ( .A({ _04414_, _11896_ }), .Y(_12449_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35733_ ( .A({ _04415_, _11896_ }), .Y(_12450_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35734_ ( .A({ _04416_, _11896_ }), .Y(_12451_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35735_ ( .A({ _04417_, _11896_ }), .Y(_12452_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35736_ ( .A({ _04418_, _11896_ }), .Y(_12453_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35737_ ( .A({ _04419_, _11896_ }), .Y(_12454_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35738_ ( .A({ _04420_, _11896_ }), .Y(_12455_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35739_ ( .A({ _04421_, _11896_ }), .Y(_12456_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35740_ ( .A({ _04422_, _11896_ }), .Y(_12457_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35741_ ( .A({ _04424_, _11896_ }), .Y(_12459_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35742_ ( .A({ _04425_, _11896_ }), .Y(_12460_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35743_ ( .A({ _04426_, _11896_ }), .Y(_12461_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35744_ ( .A({ _04427_, _11896_ }), .Y(_12462_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35745_ ( .A({ _04428_, _11896_ }), .Y(_12463_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35746_ ( .A({ _04429_, _11896_ }), .Y(_12464_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35747_ ( .A({ _04430_, _11896_ }), .Y(_12465_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35748_ ( .A({ _04431_, _11896_ }), .Y(_12466_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35749_ ( .A({ _04432_, _11896_ }), .Y(_12467_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35750_ ( .A({ _04433_, _11896_ }), .Y(_12468_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35751_ ( .A({ _04435_, _11896_ }), .Y(_12470_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35752_ ( .A({ _04436_, _11896_ }), .Y(_12471_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35753_ ( .A({ _12383_, _11896_ }), .Y(_12415_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35754_ ( .A({ _12394_, _11896_ }), .Y(_12426_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35755_ ( .A({ _12405_, _11896_ }), .Y(_12437_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35756_ ( .A({ _12408_, _11896_ }), .Y(_12440_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35757_ ( .A({ _12409_, _11896_ }), .Y(_12441_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35758_ ( .A({ _12410_, _11896_ }), .Y(_12442_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35759_ ( .A({ _12411_, _11896_ }), .Y(_12443_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35760_ ( .A({ _12412_, _11896_ }), .Y(_12444_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35761_ ( .A({ _12413_, _11896_ }), .Y(_12445_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35762_ ( .A({ _12414_, _11896_ }), .Y(_12446_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35763_ ( .A({ _12384_, _11896_ }), .Y(_12416_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35764_ ( .A({ _12385_, _11896_ }), .Y(_12417_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35765_ ( .A({ _12386_, _11896_ }), .Y(_12418_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35766_ ( .A({ _12387_, _11896_ }), .Y(_12419_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35767_ ( .A({ _12388_, _11896_ }), .Y(_12420_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35768_ ( .A({ _12389_, _11896_ }), .Y(_12421_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35769_ ( .A({ _12390_, _11896_ }), .Y(_12422_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35770_ ( .A({ _12391_, _11896_ }), .Y(_12423_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35771_ ( .A({ _12392_, _11896_ }), .Y(_12424_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35772_ ( .A({ _12393_, _11896_ }), .Y(_12425_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35773_ ( .A({ _12395_, _11896_ }), .Y(_12427_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35774_ ( .A({ _12396_, _11896_ }), .Y(_12428_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35775_ ( .A({ _12397_, _11896_ }), .Y(_12429_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35776_ ( .A({ _12398_, _11896_ }), .Y(_12430_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35777_ ( .A({ _12399_, _11896_ }), .Y(_12431_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35778_ ( .A({ _12400_, _11896_ }), .Y(_12432_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35779_ ( .A({ _12401_, _11896_ }), .Y(_12433_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35780_ ( .A({ _12402_, _11896_ }), .Y(_12434_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35781_ ( .A({ _12403_, _11896_ }), .Y(_12435_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35782_ ( .A({ _12404_, _11896_ }), .Y(_12436_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35783_ ( .A({ _12406_, _11896_ }), .Y(_12438_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35784_ ( .A({ _12407_, _11896_ }), .Y(_12439_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35785_ ( .A({ matmul_15_row_count[0], _11896_ }), .Y(_12287_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35786_ ( .A({ matmul_15_row_count[1], _11896_ }), .Y(_12298_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35787_ ( .A({ matmul_15_row_count[2], _11896_ }), .Y(_12309_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35788_ ( .A({ matmul_15_row_count[3], _11896_ }), .Y(_12312_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35789_ ( .A({ matmul_15_row_count[4], _11896_ }), .Y(_12313_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35790_ ( .A({ matmul_15_row_count[5], _11896_ }), .Y(_12314_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35791_ ( .A({ matmul_15_row_count[6], _11896_ }), .Y(_12315_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35792_ ( .A({ matmul_15_row_count[7], _11896_ }), .Y(_12316_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35793_ ( .A({ matmul_15_row_count[8], _11896_ }), .Y(_12317_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35794_ ( .A({ matmul_15_row_count[9], _11896_ }), .Y(_12318_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35795_ ( .A({ matmul_15_row_count[10], _11896_ }), .Y(_12288_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35796_ ( .A({ matmul_15_row_count[11], _11896_ }), .Y(_12289_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35797_ ( .A({ matmul_15_row_count[12], _11896_ }), .Y(_12290_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35798_ ( .A({ matmul_15_row_count[13], _11896_ }), .Y(_12291_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35799_ ( .A({ matmul_15_row_count[14], _11896_ }), .Y(_12292_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35800_ ( .A({ matmul_15_row_count[15], _11896_ }), .Y(_12293_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35801_ ( .A({ matmul_15_row_count[16], _11896_ }), .Y(_12294_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35802_ ( .A({ matmul_15_row_count[17], _11896_ }), .Y(_12295_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35803_ ( .A({ matmul_15_row_count[18], _11896_ }), .Y(_12296_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35804_ ( .A({ matmul_15_row_count[19], _11896_ }), .Y(_12297_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35805_ ( .A({ matmul_15_row_count[20], _11896_ }), .Y(_12299_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35806_ ( .A({ matmul_15_row_count[21], _11896_ }), .Y(_12300_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35807_ ( .A({ matmul_15_row_count[22], _11896_ }), .Y(_12301_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35808_ ( .A({ matmul_15_row_count[23], _11896_ }), .Y(_12302_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35809_ ( .A({ matmul_15_row_count[24], _11896_ }), .Y(_12303_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35810_ ( .A({ matmul_15_row_count[25], _11896_ }), .Y(_12304_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35811_ ( .A({ matmul_15_row_count[26], _11896_ }), .Y(_12305_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35812_ ( .A({ matmul_15_row_count[27], _11896_ }), .Y(_12306_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35813_ ( .A({ matmul_15_row_count[28], _11896_ }), .Y(_12307_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35814_ ( .A({ matmul_15_row_count[29], _11896_ }), .Y(_12308_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35815_ ( .A({ matmul_15_row_count[30], _11896_ }), .Y(_12310_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35816_ ( .A({ matmul_15_row_count[31], _11896_ }), .Y(_12311_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35817_ ( .A({ matmul_15_och_count[0], _11896_ }), .Y(_12223_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35818_ ( .A({ matmul_15_och_count[1], _11896_ }), .Y(_12234_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35819_ ( .A({ matmul_15_och_count[2], _11896_ }), .Y(_12245_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35820_ ( .A({ matmul_15_och_count[3], _11896_ }), .Y(_12248_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35821_ ( .A({ matmul_15_och_count[4], _11896_ }), .Y(_12249_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35822_ ( .A({ matmul_15_och_count[5], _11896_ }), .Y(_12250_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35823_ ( .A({ matmul_15_och_count[6], _11896_ }), .Y(_12251_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35824_ ( .A({ matmul_15_och_count[7], _11896_ }), .Y(_12252_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35825_ ( .A({ matmul_15_och_count[8], _11896_ }), .Y(_12253_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35826_ ( .A({ matmul_15_och_count[9], _11896_ }), .Y(_12254_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35827_ ( .A({ matmul_15_och_count[10], _11896_ }), .Y(_12224_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35828_ ( .A({ matmul_15_och_count[11], _11896_ }), .Y(_12225_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35829_ ( .A({ matmul_15_och_count[12], _11896_ }), .Y(_12226_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35830_ ( .A({ matmul_15_och_count[13], _11896_ }), .Y(_12227_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35831_ ( .A({ matmul_15_och_count[14], _11896_ }), .Y(_12228_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35832_ ( .A({ matmul_15_och_count[15], _11896_ }), .Y(_12229_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35833_ ( .A({ matmul_15_och_count[16], _11896_ }), .Y(_12230_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35834_ ( .A({ matmul_15_och_count[17], _11896_ }), .Y(_12231_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35835_ ( .A({ matmul_15_och_count[18], _11896_ }), .Y(_12232_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35836_ ( .A({ matmul_15_och_count[19], _11896_ }), .Y(_12233_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35837_ ( .A({ matmul_15_och_count[20], _11896_ }), .Y(_12235_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35838_ ( .A({ matmul_15_och_count[21], _11896_ }), .Y(_12236_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35839_ ( .A({ matmul_15_och_count[22], _11896_ }), .Y(_12237_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35840_ ( .A({ matmul_15_och_count[23], _11896_ }), .Y(_12238_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35841_ ( .A({ matmul_15_och_count[24], _11896_ }), .Y(_12239_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35842_ ( .A({ matmul_15_och_count[25], _11896_ }), .Y(_12240_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35843_ ( .A({ matmul_15_och_count[26], _11896_ }), .Y(_12241_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35844_ ( .A({ matmul_15_och_count[27], _11896_ }), .Y(_12242_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35845_ ( .A({ matmul_15_och_count[28], _11896_ }), .Y(_12243_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35846_ ( .A({ matmul_15_och_count[29], _11896_ }), .Y(_12244_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35847_ ( .A({ matmul_15_och_count[30], _11896_ }), .Y(_12246_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35848_ ( .A({ matmul_15_och_count[31], _11896_ }), .Y(_12247_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35849_ ( .A({ conv2d_8_row_count[0], _05909_ }), .Y(_19332_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35850_ ( .A({ conv2d_8_row_count[1], _05909_ }), .Y(_19343_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35851_ ( .A({ conv2d_8_row_count[2], _05909_ }), .Y(_19354_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35852_ ( .A({ conv2d_8_row_count[3], _05909_ }), .Y(_19357_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35853_ ( .A({ conv2d_8_row_count[4], _05909_ }), .Y(_19358_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35854_ ( .A({ conv2d_8_row_count[5], _05909_ }), .Y(_19359_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35855_ ( .A({ conv2d_8_row_count[6], _05909_ }), .Y(_19360_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35856_ ( .A({ conv2d_8_row_count[7], _05909_ }), .Y(_19361_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35857_ ( .A({ conv2d_8_row_count[8], _05909_ }), .Y(_19362_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35858_ ( .A({ conv2d_8_row_count[9], _05909_ }), .Y(_19363_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35859_ ( .A({ conv2d_8_row_count[10], _05909_ }), .Y(_19333_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35860_ ( .A({ conv2d_8_row_count[11], _05909_ }), .Y(_19334_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35861_ ( .A({ conv2d_8_row_count[12], _05909_ }), .Y(_19335_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35862_ ( .A({ conv2d_8_row_count[13], _05909_ }), .Y(_19336_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35863_ ( .A({ conv2d_8_row_count[14], _05909_ }), .Y(_19337_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35864_ ( .A({ conv2d_8_row_count[15], _05909_ }), .Y(_19338_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35865_ ( .A({ conv2d_8_row_count[16], _05909_ }), .Y(_19339_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35866_ ( .A({ conv2d_8_row_count[17], _05909_ }), .Y(_19340_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35867_ ( .A({ conv2d_8_row_count[18], _05909_ }), .Y(_19341_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35868_ ( .A({ conv2d_8_row_count[19], _05909_ }), .Y(_19342_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35869_ ( .A({ conv2d_8_row_count[20], _05909_ }), .Y(_19344_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35870_ ( .A({ conv2d_8_row_count[21], _05909_ }), .Y(_19345_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35871_ ( .A({ conv2d_8_row_count[22], _05909_ }), .Y(_19346_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35872_ ( .A({ conv2d_8_row_count[23], _05909_ }), .Y(_19347_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35873_ ( .A({ conv2d_8_row_count[24], _05909_ }), .Y(_19348_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35874_ ( .A({ conv2d_8_row_count[25], _05909_ }), .Y(_19349_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35875_ ( .A({ conv2d_8_row_count[26], _05909_ }), .Y(_19350_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35876_ ( .A({ conv2d_8_row_count[27], _05909_ }), .Y(_19351_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35877_ ( .A({ conv2d_8_row_count[28], _05909_ }), .Y(_19352_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35878_ ( .A({ conv2d_8_row_count[29], _05909_ }), .Y(_19353_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35879_ ( .A({ conv2d_8_row_count[30], _05909_ }), .Y(_19355_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35880_ ( .A({ conv2d_8_row_count[31], _05909_ }), .Y(_19356_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35881_ ( .A({ matmul_15_bat_count[0], _11896_ }), .Y(_12255_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35882_ ( .A({ matmul_15_bat_count[1], _11896_ }), .Y(_12266_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35883_ ( .A({ matmul_15_bat_count[2], _11896_ }), .Y(_12277_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35884_ ( .A({ matmul_15_bat_count[3], _11896_ }), .Y(_12280_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35885_ ( .A({ matmul_15_bat_count[4], _11896_ }), .Y(_12281_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35886_ ( .A({ matmul_15_bat_count[5], _11896_ }), .Y(_12282_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35887_ ( .A({ matmul_15_bat_count[6], _11896_ }), .Y(_12283_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35888_ ( .A({ matmul_15_bat_count[7], _11896_ }), .Y(_12284_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35889_ ( .A({ matmul_15_bat_count[8], _11896_ }), .Y(_12285_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35890_ ( .A({ matmul_15_bat_count[9], _11896_ }), .Y(_12286_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35891_ ( .A({ matmul_15_bat_count[10], _11896_ }), .Y(_12256_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35892_ ( .A({ matmul_15_bat_count[11], _11896_ }), .Y(_12257_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35893_ ( .A({ matmul_15_bat_count[12], _11896_ }), .Y(_12258_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35894_ ( .A({ matmul_15_bat_count[13], _11896_ }), .Y(_12259_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35895_ ( .A({ matmul_15_bat_count[14], _11896_ }), .Y(_12260_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35896_ ( .A({ matmul_15_bat_count[15], _11896_ }), .Y(_12261_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35897_ ( .A({ matmul_15_bat_count[16], _11896_ }), .Y(_12262_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35898_ ( .A({ matmul_15_bat_count[17], _11896_ }), .Y(_12263_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35899_ ( .A({ matmul_15_bat_count[18], _11896_ }), .Y(_12264_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35900_ ( .A({ matmul_15_bat_count[19], _11896_ }), .Y(_12265_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35901_ ( .A({ matmul_15_bat_count[20], _11896_ }), .Y(_12267_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35902_ ( .A({ matmul_15_bat_count[21], _11896_ }), .Y(_12268_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35903_ ( .A({ matmul_15_bat_count[22], _11896_ }), .Y(_12269_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35904_ ( .A({ matmul_15_bat_count[23], _11896_ }), .Y(_12270_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35905_ ( .A({ matmul_15_bat_count[24], _11896_ }), .Y(_12271_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35906_ ( .A({ matmul_15_bat_count[25], _11896_ }), .Y(_12272_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35907_ ( .A({ matmul_15_bat_count[26], _11896_ }), .Y(_12273_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35908_ ( .A({ matmul_15_bat_count[27], _11896_ }), .Y(_12274_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35909_ ( .A({ matmul_15_bat_count[28], _11896_ }), .Y(_12275_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35910_ ( .A({ matmul_15_bat_count[29], _11896_ }), .Y(_12276_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35911_ ( .A({ matmul_15_bat_count[30], _11896_ }), .Y(_12278_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35912_ ( .A({ matmul_15_bat_count[31], _11896_ }), .Y(_12279_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35913_ ( .A({ _18554_, _05909_ }), .Y(_18555_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35914_ ( .A({ _12095_, _11896_ }), .Y(_12127_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35915_ ( .A({ _12106_, _11896_ }), .Y(_12138_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35916_ ( .A({ _12117_, _11896_ }), .Y(_12149_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35917_ ( .A({ _12120_, _11896_ }), .Y(_12152_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35918_ ( .A({ _12121_, _11896_ }), .Y(_12153_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35919_ ( .A({ _12122_, _11896_ }), .Y(_12154_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35920_ ( .A({ _12123_, _11896_ }), .Y(_12155_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35921_ ( .A({ _12124_, _11896_ }), .Y(_12156_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35922_ ( .A({ _12125_, _11896_ }), .Y(_12157_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35923_ ( .A({ _12126_, _11896_ }), .Y(_12158_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35924_ ( .A({ _12096_, _11896_ }), .Y(_12128_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35925_ ( .A({ _12097_, _11896_ }), .Y(_12129_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35926_ ( .A({ _12098_, _11896_ }), .Y(_12130_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35927_ ( .A({ _12099_, _11896_ }), .Y(_12131_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35928_ ( .A({ _12100_, _11896_ }), .Y(_12132_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35929_ ( .A({ _12101_, _11896_ }), .Y(_12133_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35930_ ( .A({ _12102_, _11896_ }), .Y(_12134_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35931_ ( .A({ _12103_, _11896_ }), .Y(_12135_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35932_ ( .A({ _12104_, _11896_ }), .Y(_12136_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35933_ ( .A({ _12105_, _11896_ }), .Y(_12137_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35934_ ( .A({ _12107_, _11896_ }), .Y(_12139_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35935_ ( .A({ _12108_, _11896_ }), .Y(_12140_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35936_ ( .A({ _12109_, _11896_ }), .Y(_12141_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35937_ ( .A({ _12110_, _11896_ }), .Y(_12142_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35938_ ( .A({ _12111_, _11896_ }), .Y(_12143_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35939_ ( .A({ _12112_, _11896_ }), .Y(_12144_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35940_ ( .A({ _12113_, _11896_ }), .Y(_12145_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35941_ ( .A({ _12114_, _11896_ }), .Y(_12146_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35942_ ( .A({ _12115_, _11896_ }), .Y(_12147_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35943_ ( .A({ _12116_, _11896_ }), .Y(_12148_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35944_ ( .A({ _12118_, _11896_ }), .Y(_12150_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35945_ ( .A({ _12119_, _11896_ }), .Y(_12151_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35946_ ( .A({ _12093_, _11896_ }), .Y(_12094_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35947_ ( .A({ _12159_, _11896_ }), .Y(_12191_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35948_ ( .A({ _12170_, _11896_ }), .Y(_12202_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35949_ ( .A({ _12181_, _11896_ }), .Y(_12213_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35950_ ( .A({ _12184_, _11896_ }), .Y(_12216_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35951_ ( .A({ _12185_, _11896_ }), .Y(_12217_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35952_ ( .A({ _12186_, _11896_ }), .Y(_12218_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35953_ ( .A({ _12187_, _11896_ }), .Y(_12219_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35954_ ( .A({ _12188_, _11896_ }), .Y(_12220_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35955_ ( .A({ _12189_, _11896_ }), .Y(_12221_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35956_ ( .A({ _12190_, _11896_ }), .Y(_12222_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35957_ ( .A({ _12160_, _11896_ }), .Y(_12192_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35958_ ( .A({ _12161_, _11896_ }), .Y(_12193_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35959_ ( .A({ _12162_, _11896_ }), .Y(_12194_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35960_ ( .A({ _12163_, _11896_ }), .Y(_12195_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35961_ ( .A({ _12164_, _11896_ }), .Y(_12196_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35962_ ( .A({ _12165_, _11896_ }), .Y(_12197_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35963_ ( .A({ _12166_, _11896_ }), .Y(_12198_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35964_ ( .A({ _12167_, _11896_ }), .Y(_12199_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35965_ ( .A({ _12168_, _11896_ }), .Y(_12200_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35966_ ( .A({ _12169_, _11896_ }), .Y(_12201_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35967_ ( .A({ _12171_, _11896_ }), .Y(_12203_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35968_ ( .A({ _12172_, _11896_ }), .Y(_12204_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35969_ ( .A({ _12173_, _11896_ }), .Y(_12205_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35970_ ( .A({ _12174_, _11896_ }), .Y(_12206_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35971_ ( .A({ _12175_, _11896_ }), .Y(_12207_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35972_ ( .A({ _12176_, _11896_ }), .Y(_12208_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35973_ ( .A({ _12177_, _11896_ }), .Y(_12209_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35974_ ( .A({ _12178_, _11896_ }), .Y(_12210_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35975_ ( .A({ _12179_, _11896_ }), .Y(_12211_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35976_ ( .A({ _12180_, _11896_ }), .Y(_12212_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35977_ ( .A({ _12182_, _11896_ }), .Y(_12214_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35978_ ( .A({ _12183_, _11896_ }), .Y(_12215_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35979_ ( .A({ _17839_, _07122_ }), .Y(_17871_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35980_ ( .A({ _17850_, _07122_ }), .Y(_17882_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35981_ ( .A({ _17861_, _07122_ }), .Y(_17893_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35982_ ( .A({ _17864_, _07122_ }), .Y(_17896_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35983_ ( .A({ _17865_, _07122_ }), .Y(_17897_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35984_ ( .A({ _17866_, _07122_ }), .Y(_17898_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35985_ ( .A({ _17867_, _07122_ }), .Y(_17899_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35986_ ( .A({ _17868_, _07122_ }), .Y(_17900_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35987_ ( .A({ _17869_, _07122_ }), .Y(_17901_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35988_ ( .A({ _17870_, _07122_ }), .Y(_17902_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35989_ ( .A({ _17840_, _07122_ }), .Y(_17872_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35990_ ( .A({ _17841_, _07122_ }), .Y(_17873_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35991_ ( .A({ _17842_, _07122_ }), .Y(_17874_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35992_ ( .A({ _17843_, _07122_ }), .Y(_17875_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35993_ ( .A({ _17844_, _07122_ }), .Y(_17876_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35994_ ( .A({ _17845_, _07122_ }), .Y(_17877_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35995_ ( .A({ _17846_, _07122_ }), .Y(_17878_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35996_ ( .A({ _17847_, _07122_ }), .Y(_17879_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35997_ ( .A({ _17848_, _07122_ }), .Y(_17880_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35998_ ( .A({ _17849_, _07122_ }), .Y(_17881_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35999_ ( .A({ _17851_, _07122_ }), .Y(_17883_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36000_ ( .A({ _17852_, _07122_ }), .Y(_17884_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36001_ ( .A({ _17853_, _07122_ }), .Y(_17885_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36002_ ( .A({ _17854_, _07122_ }), .Y(_17886_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36003_ ( .A({ _17855_, _07122_ }), .Y(_17887_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36004_ ( .A({ _17856_, _07122_ }), .Y(_17888_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36005_ ( .A({ _17857_, _07122_ }), .Y(_17889_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36006_ ( .A({ _17858_, _07122_ }), .Y(_17890_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36007_ ( .A({ _17859_, _07122_ }), .Y(_17891_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36008_ ( .A({ _17860_, _07122_ }), .Y(_17892_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36009_ ( .A({ _17862_, _07122_ }), .Y(_17894_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36010_ ( .A({ _17863_, _07122_ }), .Y(_17895_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36011_ ( .A({ _12029_, _11896_ }), .Y(_12061_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36012_ ( .A({ _12040_, _11896_ }), .Y(_12072_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36013_ ( .A({ _12051_, _11896_ }), .Y(_12083_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36014_ ( .A({ _12054_, _11896_ }), .Y(_12086_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36015_ ( .A({ _12055_, _11896_ }), .Y(_12087_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36016_ ( .A({ _12056_, _11896_ }), .Y(_12088_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36017_ ( .A({ _12057_, _11896_ }), .Y(_12089_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36018_ ( .A({ _12058_, _11896_ }), .Y(_12090_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36019_ ( .A({ _12059_, _11896_ }), .Y(_12091_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36020_ ( .A({ _12060_, _11896_ }), .Y(_12092_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36021_ ( .A({ _12030_, _11896_ }), .Y(_12062_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36022_ ( .A({ _12031_, _11896_ }), .Y(_12063_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36023_ ( .A({ _12032_, _11896_ }), .Y(_12064_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36024_ ( .A({ _12033_, _11896_ }), .Y(_12065_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36025_ ( .A({ _12034_, _11896_ }), .Y(_12066_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36026_ ( .A({ _12035_, _11896_ }), .Y(_12067_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36027_ ( .A({ _12036_, _11896_ }), .Y(_12068_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36028_ ( .A({ _12037_, _11896_ }), .Y(_12069_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36029_ ( .A({ _12038_, _11896_ }), .Y(_12070_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36030_ ( .A({ _12039_, _11896_ }), .Y(_12071_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36031_ ( .A({ _12041_, _11896_ }), .Y(_12073_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36032_ ( .A({ _12042_, _11896_ }), .Y(_12074_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36033_ ( .A({ _12043_, _11896_ }), .Y(_12075_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36034_ ( .A({ _12044_, _11896_ }), .Y(_12076_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36035_ ( .A({ _12045_, _11896_ }), .Y(_12077_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36036_ ( .A({ _12046_, _11896_ }), .Y(_12078_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36037_ ( .A({ _12047_, _11896_ }), .Y(_12079_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36038_ ( .A({ _12048_, _11896_ }), .Y(_12080_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36039_ ( .A({ _12049_, _11896_ }), .Y(_12081_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36040_ ( .A({ _12050_, _11896_ }), .Y(_12082_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36041_ ( .A({ _12052_, _11896_ }), .Y(_12084_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36042_ ( .A({ _12053_, _11896_ }), .Y(_12085_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36043_ ( .A({ _11965_, _11896_ }), .Y(_11997_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36044_ ( .A({ _11976_, _11896_ }), .Y(_12008_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36045_ ( .A({ _11987_, _11896_ }), .Y(_12019_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36046_ ( .A({ _11990_, _11896_ }), .Y(_12022_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36047_ ( .A({ _11991_, _11896_ }), .Y(_12023_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36048_ ( .A({ _11992_, _11896_ }), .Y(_12024_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36049_ ( .A({ _11993_, _11896_ }), .Y(_12025_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36050_ ( .A({ _11994_, _11896_ }), .Y(_12026_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36051_ ( .A({ _11995_, _11896_ }), .Y(_12027_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36052_ ( .A({ _11996_, _11896_ }), .Y(_12028_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36053_ ( .A({ _11966_, _11896_ }), .Y(_11998_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36054_ ( .A({ _11967_, _11896_ }), .Y(_11999_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36055_ ( .A({ _11968_, _11896_ }), .Y(_12000_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36056_ ( .A({ _11969_, _11896_ }), .Y(_12001_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36057_ ( .A({ _11970_, _11896_ }), .Y(_12002_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36058_ ( .A({ _11971_, _11896_ }), .Y(_12003_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36059_ ( .A({ _11972_, _11896_ }), .Y(_12004_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36060_ ( .A({ _11973_, _11896_ }), .Y(_12005_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36061_ ( .A({ _11974_, _11896_ }), .Y(_12006_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36062_ ( .A({ _11975_, _11896_ }), .Y(_12007_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36063_ ( .A({ _11977_, _11896_ }), .Y(_12009_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36064_ ( .A({ _11978_, _11896_ }), .Y(_12010_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36065_ ( .A({ _11979_, _11896_ }), .Y(_12011_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36066_ ( .A({ _11980_, _11896_ }), .Y(_12012_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36067_ ( .A({ _11981_, _11896_ }), .Y(_12013_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36068_ ( .A({ _11982_, _11896_ }), .Y(_12014_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36069_ ( .A({ _11983_, _11896_ }), .Y(_12015_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36070_ ( .A({ _11984_, _11896_ }), .Y(_12016_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36071_ ( .A({ _11985_, _11896_ }), .Y(_12017_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36072_ ( .A({ _11986_, _11896_ }), .Y(_12018_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36073_ ( .A({ _11988_, _11896_ }), .Y(_12020_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36074_ ( .A({ _11989_, _11896_ }), .Y(_12021_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36075_ ( .A({ _11899_, _11896_ }), .Y(_11900_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36076_ ( .A({ _11897_, _11896_ }), .Y(_11898_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36077_ ( .A({ _18556_, _05909_ }), .Y(_18557_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36078_ ( .A({ _17484_, _07122_ }), .Y(_17516_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36079_ ( .A({ _17495_, _07122_ }), .Y(_17527_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36080_ ( .A({ _17506_, _07122_ }), .Y(_17538_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36081_ ( .A({ _17509_, _07122_ }), .Y(_17541_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36082_ ( .A({ _17510_, _07122_ }), .Y(_17542_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36083_ ( .A({ _17511_, _07122_ }), .Y(_17543_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36084_ ( .A({ _17512_, _07122_ }), .Y(_17544_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36085_ ( .A({ _17513_, _07122_ }), .Y(_17545_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36086_ ( .A({ _17514_, _07122_ }), .Y(_17546_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36087_ ( .A({ _17515_, _07122_ }), .Y(_17547_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36088_ ( .A({ _17485_, _07122_ }), .Y(_17517_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36089_ ( .A({ _17486_, _07122_ }), .Y(_17518_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36090_ ( .A({ _17487_, _07122_ }), .Y(_17519_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36091_ ( .A({ _17488_, _07122_ }), .Y(_17520_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36092_ ( .A({ _17489_, _07122_ }), .Y(_17521_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36093_ ( .A({ _17490_, _07122_ }), .Y(_17522_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36094_ ( .A({ _17491_, _07122_ }), .Y(_17523_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36095_ ( .A({ _17492_, _07122_ }), .Y(_17524_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36096_ ( .A({ _17493_, _07122_ }), .Y(_17525_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36097_ ( .A({ _17494_, _07122_ }), .Y(_17526_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36098_ ( .A({ _17496_, _07122_ }), .Y(_17528_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36099_ ( .A({ _17497_, _07122_ }), .Y(_17529_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36100_ ( .A({ _17498_, _07122_ }), .Y(_17530_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36101_ ( .A({ _17499_, _07122_ }), .Y(_17531_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36102_ ( .A({ _17500_, _07122_ }), .Y(_17532_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36103_ ( .A({ _17501_, _07122_ }), .Y(_17533_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36104_ ( .A({ _17502_, _07122_ }), .Y(_17534_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36105_ ( .A({ _17503_, _07122_ }), .Y(_17535_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36106_ ( .A({ _17504_, _07122_ }), .Y(_17536_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36107_ ( .A({ _17505_, _07122_ }), .Y(_17537_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36108_ ( .A({ _17507_, _07122_ }), .Y(_17539_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36109_ ( .A({ _17508_, _07122_ }), .Y(_17540_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36110_ ( .A({ _11155_, _11146_, _11151_ }), .Y(_21880_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _36111_ ( .A({ _11150_, _11149_, _11147_ }), .Y(_11146_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36112_ ( .A({ _11148_, _04468_, _04467_, _04465_ }), .Y(_11147_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36113_ ( .A({ _04463_, _04462_, _04460_, _04457_ }), .Y(_11148_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36114_ ( .A({ _04456_, _04454_, _04453_, _04452_ }), .Y(_11149_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36115_ ( .A({ _04451_, _04450_, _04449_, _04448_ }), .Y(_11150_) );
  \$lut  #( .LUT(16'h7f00), .WIDTH(4) ) _36116_ ( .A({ _04447_, _11154_, _11153_, _11152_ }), .Y(_11151_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36117_ ( .A({ _04446_, _04445_, _04475_, _04474_ }), .Y(_11152_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36118_ ( .A({ _04473_, _04472_, _04471_, _04470_ }), .Y(_11153_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36119_ ( .A({ _04469_, _04466_, _04455_, _04444_ }), .Y(_11154_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36120_ ( .A({ _04464_, _04461_, _04459_, _04458_ }), .Y(_11155_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36121_ ( .A({ _17903_, _07122_ }), .Y(_17935_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36122_ ( .A({ _17914_, _07122_ }), .Y(_17946_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36123_ ( .A({ _17925_, _07122_ }), .Y(_17957_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36124_ ( .A({ _17928_, _07122_ }), .Y(_17960_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36125_ ( .A({ _17929_, _07122_ }), .Y(_17961_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36126_ ( .A({ _17930_, _07122_ }), .Y(_17962_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36127_ ( .A({ _17931_, _07122_ }), .Y(_17963_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36128_ ( .A({ _17932_, _07122_ }), .Y(_17964_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36129_ ( .A({ _17933_, _07122_ }), .Y(_17965_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36130_ ( .A({ _17934_, _07122_ }), .Y(_17966_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36131_ ( .A({ _17904_, _07122_ }), .Y(_17936_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36132_ ( .A({ _17905_, _07122_ }), .Y(_17937_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36133_ ( .A({ _17906_, _07122_ }), .Y(_17938_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36134_ ( .A({ _17907_, _07122_ }), .Y(_17939_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36135_ ( .A({ _17908_, _07122_ }), .Y(_17940_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36136_ ( .A({ _17909_, _07122_ }), .Y(_17941_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36137_ ( .A({ _17910_, _07122_ }), .Y(_17942_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36138_ ( .A({ _17911_, _07122_ }), .Y(_17943_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36139_ ( .A({ _17912_, _07122_ }), .Y(_17944_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36140_ ( .A({ _17913_, _07122_ }), .Y(_17945_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36141_ ( .A({ _17915_, _07122_ }), .Y(_17947_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36142_ ( .A({ _17916_, _07122_ }), .Y(_17948_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36143_ ( .A({ _17917_, _07122_ }), .Y(_17949_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36144_ ( .A({ _17918_, _07122_ }), .Y(_17950_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36145_ ( .A({ _17919_, _07122_ }), .Y(_17951_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36146_ ( .A({ _17920_, _07122_ }), .Y(_17952_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36147_ ( .A({ _17921_, _07122_ }), .Y(_17953_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36148_ ( .A({ _17922_, _07122_ }), .Y(_17954_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36149_ ( .A({ _17923_, _07122_ }), .Y(_17955_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36150_ ( .A({ _17924_, _07122_ }), .Y(_17956_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36151_ ( .A({ _17926_, _07122_ }), .Y(_17958_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36152_ ( .A({ _17927_, _07122_ }), .Y(_17959_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36153_ ( .A({ __substreamoutput_data_866[7], _11156_ }), .Y(_05261_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36154_ ( .A({ _11157_, __substreamoutput_data_866[6:4] }), .Y(_11156_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36155_ ( .A(__substreamoutput_data_866[3:0]), .Y(_11157_) );
  \$lut  #( .LUT(8'h71), .WIDTH(3) ) _36156_ ( .A({ _reducecustom_data_191[6], __variable_wdata_187[6], _11159_ }), .Y(_11158_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _36157_ ( .A({ __variable_wdata_187[5], _reducecustom_data_191[5], _11160_ }), .Y(_11159_) );
  \$lut  #( .LUT(16'hddd4), .WIDTH(4) ) _36158_ ( .A({ _11164_, _11161_, __variable_wdata_187[4], _reducecustom_data_191[4] }), .Y(_11160_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _36159_ ( .A({ _11163_, __variable_wdata_187[2], _reducecustom_data_191[2], _11162_ }), .Y(_11161_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _36160_ ( .A({ _reducecustom_data_191[0], __variable_wdata_187[0], __variable_wdata_187[1], _reducecustom_data_191[1] }), .Y(_11162_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36161_ ( .A({ _reducecustom_data_191[3], __variable_wdata_187[3] }), .Y(_11163_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36162_ ( .A({ __variable_wdata_187[3], _reducecustom_data_191[3] }), .Y(_11164_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36163_ ( .A(_reducecustom_data_191[28:25]), .Y(_11165_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36164_ ( .A({ __variable_wdata_187[7], _reducecustom_data_191[30:29], _reducecustom_data_191[24] }), .Y(_11166_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _36165_ ( .A({ __variable_wdata_187[7], _reducecustom_data_191[30:29] }), .Y(_11167_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36166_ ( .A(_reducecustom_data_191[28:25]), .Y(_11168_) );
  \$lut  #( .LUT(16'hbf00), .WIDTH(4) ) _36167_ ( .A({ _sra_data_40[39], _11169_, _11176_, _11174_ }), .Y(_05872_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36168_ ( .A({ _11173_, _11172_, _11171_, _11170_ }), .Y(_11169_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36169_ ( .A(_sra_data_40[26:23]), .Y(_11170_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36170_ ( .A(_sra_data_40[22:19]), .Y(_11171_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36171_ ( .A({ _sra_data_40[38], _sra_data_40[36:35], _sra_data_40[33] }), .Y(_11172_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36172_ ( .A(_sra_data_40[31:28]), .Y(_11173_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36173_ ( .A({ _11175_, _sra_data_40[5], _sra_data_40[3:2] }), .Y(_11174_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36174_ ( .A({ _sra_data_40[0], _sra_data_40[6], _sra_data_40[4], _sra_data_40[1] }), .Y(_11175_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36175_ ( .A({ _11180_, _11179_, _11178_, _11177_ }), .Y(_11176_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36176_ ( .A({ _sra_data_40[18:17], _sra_data_40[15:14] }), .Y(_11177_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36177_ ( .A(_sra_data_40[12:9]), .Y(_11178_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36178_ ( .A({ _sra_data_40[16], _sra_data_40[13], _sra_data_40[8:7] }), .Y(_11179_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36179_ ( .A({ _sra_data_40[37], _sra_data_40[34], _sra_data_40[32], _sra_data_40[27] }), .Y(_11180_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _36180_ ( .A({ _sra_data_40[39], _11181_, _11186_ }), .Y(_05250_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36181_ ( .A({ _11185_, _11184_, _11183_, _11182_ }), .Y(_11181_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36182_ ( .A({ _sra_data_40[18:17], _sra_data_40[15:14] }), .Y(_11182_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36183_ ( .A(_sra_data_40[12:9]), .Y(_11183_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36184_ ( .A({ _sra_data_40[16], _sra_data_40[13], _sra_data_40[8:7] }), .Y(_11184_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36185_ ( .A({ _sra_data_40[37], _sra_data_40[34], _sra_data_40[32], _sra_data_40[27] }), .Y(_11185_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36186_ ( .A({ _11190_, _11189_, _11188_, _11187_ }), .Y(_11186_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36187_ ( .A(_sra_data_40[26:23]), .Y(_11187_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36188_ ( .A(_sra_data_40[22:19]), .Y(_11188_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36189_ ( .A({ _sra_data_40[38], _sra_data_40[36:35], _sra_data_40[33] }), .Y(_11189_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36190_ ( .A(_sra_data_40[31:28]), .Y(_11190_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36191_ ( .A({ _18031_, _07122_ }), .Y(_18063_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36192_ ( .A({ _18042_, _07122_ }), .Y(_18074_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36193_ ( .A({ _18053_, _07122_ }), .Y(_18085_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36194_ ( .A({ _18056_, _07122_ }), .Y(_18088_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36195_ ( .A({ _18057_, _07122_ }), .Y(_18089_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36196_ ( .A({ _18058_, _07122_ }), .Y(_18090_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36197_ ( .A({ _18059_, _07122_ }), .Y(_18091_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36198_ ( .A({ _18060_, _07122_ }), .Y(_18092_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36199_ ( .A({ _18061_, _07122_ }), .Y(_18093_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36200_ ( .A({ _18062_, _07122_ }), .Y(_18094_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36201_ ( .A({ _18032_, _07122_ }), .Y(_18064_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36202_ ( .A({ _18033_, _07122_ }), .Y(_18065_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36203_ ( .A({ _18034_, _07122_ }), .Y(_18066_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36204_ ( .A({ _18035_, _07122_ }), .Y(_18067_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36205_ ( .A({ _18036_, _07122_ }), .Y(_18068_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36206_ ( .A({ _18037_, _07122_ }), .Y(_18069_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36207_ ( .A({ _18038_, _07122_ }), .Y(_18070_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36208_ ( .A({ _18039_, _07122_ }), .Y(_18071_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36209_ ( .A({ _18040_, _07122_ }), .Y(_18072_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36210_ ( .A({ _18041_, _07122_ }), .Y(_18073_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36211_ ( .A({ _18043_, _07122_ }), .Y(_18075_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36212_ ( .A({ _18044_, _07122_ }), .Y(_18076_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36213_ ( .A({ _18045_, _07122_ }), .Y(_18077_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36214_ ( .A({ _18046_, _07122_ }), .Y(_18078_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36215_ ( .A({ _18047_, _07122_ }), .Y(_18079_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36216_ ( .A({ _18048_, _07122_ }), .Y(_18080_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36217_ ( .A({ _18049_, _07122_ }), .Y(_18081_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36218_ ( .A({ _18050_, _07122_ }), .Y(_18082_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36219_ ( .A({ _18051_, _07122_ }), .Y(_18083_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36220_ ( .A({ _18052_, _07122_ }), .Y(_18084_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36221_ ( .A({ _18054_, _07122_ }), .Y(_18086_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36222_ ( .A({ _18055_, _07122_ }), .Y(_18087_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36223_ ( .A(matmul_15_next_out_write_size[1:0]), .Y(_21879_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36224_ ( .A(cparam_max_pool_serial_9_out_row_step[1:0]), .Y(_21878_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36225_ ( .A(cparam_max_pool_serial_9_act_offset_values_1[1:0]), .Y(_21877_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36226_ ( .A(conv2d_8_next_out_write_size[1:0]), .Y(_21876_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36227_ ( .A(cparam_conv2d_8_act_read_size[1:0]), .Y(_21875_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36228_ ( .A(cparam_conv2d_8_filter_base_step[1:0]), .Y(_21874_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36229_ ( .A({ _17646_, _07122_ }), .Y(_17678_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36230_ ( .A({ _17657_, _07122_ }), .Y(_17689_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36231_ ( .A({ _17668_, _07122_ }), .Y(_17700_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36232_ ( .A({ _17671_, _07122_ }), .Y(_17703_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36233_ ( .A({ _17672_, _07122_ }), .Y(_17704_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36234_ ( .A({ _17673_, _07122_ }), .Y(_17705_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36235_ ( .A({ _17674_, _07122_ }), .Y(_17706_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36236_ ( .A({ _17675_, _07122_ }), .Y(_17707_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36237_ ( .A({ _17676_, _07122_ }), .Y(_17708_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36238_ ( .A({ _17677_, _07122_ }), .Y(_17709_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36239_ ( .A({ _17647_, _07122_ }), .Y(_17679_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36240_ ( .A({ _17648_, _07122_ }), .Y(_17680_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36241_ ( .A({ _17649_, _07122_ }), .Y(_17681_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36242_ ( .A({ _17650_, _07122_ }), .Y(_17682_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36243_ ( .A({ _17651_, _07122_ }), .Y(_17683_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36244_ ( .A({ _17652_, _07122_ }), .Y(_17684_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36245_ ( .A({ _17653_, _07122_ }), .Y(_17685_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36246_ ( .A({ _17654_, _07122_ }), .Y(_17686_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36247_ ( .A({ _17655_, _07122_ }), .Y(_17687_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36248_ ( .A({ _17656_, _07122_ }), .Y(_17688_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36249_ ( .A({ _17658_, _07122_ }), .Y(_17690_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36250_ ( .A({ _17659_, _07122_ }), .Y(_17691_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36251_ ( .A({ _17660_, _07122_ }), .Y(_17692_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36252_ ( .A({ _17661_, _07122_ }), .Y(_17693_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36253_ ( .A({ _17662_, _07122_ }), .Y(_17694_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36254_ ( .A({ _17663_, _07122_ }), .Y(_17695_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36255_ ( .A({ _17664_, _07122_ }), .Y(_17696_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36256_ ( .A({ _17665_, _07122_ }), .Y(_17697_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36257_ ( .A({ _17666_, _07122_ }), .Y(_17698_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36258_ ( .A({ _17667_, _07122_ }), .Y(_17699_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36259_ ( .A({ _17669_, _07122_ }), .Y(_17701_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36260_ ( .A({ _17670_, _07122_ }), .Y(_17702_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36261_ ( .A({ _17711_, _07122_ }), .Y(_17743_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36262_ ( .A({ _17722_, _07122_ }), .Y(_17754_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36263_ ( .A({ _17733_, _07122_ }), .Y(_17765_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36264_ ( .A({ _17736_, _07122_ }), .Y(_17768_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36265_ ( .A({ _17737_, _07122_ }), .Y(_17769_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36266_ ( .A({ _17738_, _07122_ }), .Y(_17770_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36267_ ( .A({ _17739_, _07122_ }), .Y(_17771_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36268_ ( .A({ _17740_, _07122_ }), .Y(_17772_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36269_ ( .A({ _17741_, _07122_ }), .Y(_17773_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36270_ ( .A({ _17742_, _07122_ }), .Y(_17774_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36271_ ( .A({ _17712_, _07122_ }), .Y(_17744_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36272_ ( .A({ _17713_, _07122_ }), .Y(_17745_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36273_ ( .A({ _17714_, _07122_ }), .Y(_17746_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36274_ ( .A({ _17715_, _07122_ }), .Y(_17747_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36275_ ( .A({ _17716_, _07122_ }), .Y(_17748_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36276_ ( .A({ _17717_, _07122_ }), .Y(_17749_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36277_ ( .A({ _17718_, _07122_ }), .Y(_17750_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36278_ ( .A({ _17719_, _07122_ }), .Y(_17751_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36279_ ( .A({ _17720_, _07122_ }), .Y(_17752_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36280_ ( .A({ _17721_, _07122_ }), .Y(_17753_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36281_ ( .A({ _17723_, _07122_ }), .Y(_17755_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36282_ ( .A({ _17724_, _07122_ }), .Y(_17756_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36283_ ( .A({ _17725_, _07122_ }), .Y(_17757_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36284_ ( .A({ _17726_, _07122_ }), .Y(_17758_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36285_ ( .A({ _17727_, _07122_ }), .Y(_17759_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36286_ ( .A({ _17728_, _07122_ }), .Y(_17760_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36287_ ( .A({ _17729_, _07122_ }), .Y(_17761_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36288_ ( .A({ _17730_, _07122_ }), .Y(_17762_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36289_ ( .A({ _17731_, _07122_ }), .Y(_17763_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36290_ ( .A({ _17732_, _07122_ }), .Y(_17764_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36291_ ( .A({ _17734_, _07122_ }), .Y(_17766_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36292_ ( .A({ _17735_, _07122_ }), .Y(_17767_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36293_ ( .A({ _18163_, _07122_ }), .Y(_18195_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36294_ ( .A({ _18174_, _07122_ }), .Y(_18206_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36295_ ( .A({ _18185_, _07122_ }), .Y(_18217_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36296_ ( .A({ _18188_, _07122_ }), .Y(_18220_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36297_ ( .A({ _18189_, _07122_ }), .Y(_18221_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36298_ ( .A({ _18190_, _07122_ }), .Y(_18222_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36299_ ( .A({ _18191_, _07122_ }), .Y(_18223_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36300_ ( .A({ _18192_, _07122_ }), .Y(_18224_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36301_ ( .A({ _18193_, _07122_ }), .Y(_18225_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36302_ ( .A({ _18194_, _07122_ }), .Y(_18226_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36303_ ( .A({ _18164_, _07122_ }), .Y(_18196_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36304_ ( .A({ _18165_, _07122_ }), .Y(_18197_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36305_ ( .A({ _18166_, _07122_ }), .Y(_18198_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36306_ ( .A({ _18167_, _07122_ }), .Y(_18199_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36307_ ( .A({ _18168_, _07122_ }), .Y(_18200_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36308_ ( .A({ _18169_, _07122_ }), .Y(_18201_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36309_ ( .A({ _18170_, _07122_ }), .Y(_18202_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36310_ ( .A({ _18171_, _07122_ }), .Y(_18203_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36311_ ( .A({ _18172_, _07122_ }), .Y(_18204_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36312_ ( .A({ _18173_, _07122_ }), .Y(_18205_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36313_ ( .A({ _18175_, _07122_ }), .Y(_18207_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36314_ ( .A({ _18176_, _07122_ }), .Y(_18208_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36315_ ( .A({ _18177_, _07122_ }), .Y(_18209_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36316_ ( .A({ _18178_, _07122_ }), .Y(_18210_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36317_ ( .A({ _18179_, _07122_ }), .Y(_18211_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36318_ ( .A({ _18180_, _07122_ }), .Y(_18212_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36319_ ( .A({ _18181_, _07122_ }), .Y(_18213_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36320_ ( .A({ _18182_, _07122_ }), .Y(_18214_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36321_ ( .A({ _18183_, _07122_ }), .Y(_18215_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36322_ ( .A({ _18184_, _07122_ }), .Y(_18216_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36323_ ( .A({ _18186_, _07122_ }), .Y(_18218_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36324_ ( .A({ _18187_, _07122_ }), .Y(_18219_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36325_ ( .A({ _18095_, _07122_ }), .Y(_18127_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36326_ ( .A({ _18106_, _07122_ }), .Y(_18138_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36327_ ( .A({ _18117_, _07122_ }), .Y(_18149_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36328_ ( .A({ _18120_, _07122_ }), .Y(_18152_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36329_ ( .A({ _18121_, _07122_ }), .Y(_18153_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36330_ ( .A({ _18122_, _07122_ }), .Y(_18154_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36331_ ( .A({ _18123_, _07122_ }), .Y(_18155_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36332_ ( .A({ _18124_, _07122_ }), .Y(_18156_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36333_ ( .A({ _18125_, _07122_ }), .Y(_18157_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36334_ ( .A({ _18126_, _07122_ }), .Y(_18158_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36335_ ( .A({ _18096_, _07122_ }), .Y(_18128_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36336_ ( .A({ _18097_, _07122_ }), .Y(_18129_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36337_ ( .A({ _18098_, _07122_ }), .Y(_18130_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36338_ ( .A({ _18099_, _07122_ }), .Y(_18131_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36339_ ( .A({ _18100_, _07122_ }), .Y(_18132_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36340_ ( .A({ _18101_, _07122_ }), .Y(_18133_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36341_ ( .A({ _18102_, _07122_ }), .Y(_18134_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36342_ ( .A({ _18103_, _07122_ }), .Y(_18135_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36343_ ( .A({ _18104_, _07122_ }), .Y(_18136_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36344_ ( .A({ _18105_, _07122_ }), .Y(_18137_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36345_ ( .A({ _18107_, _07122_ }), .Y(_18139_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36346_ ( .A({ _18108_, _07122_ }), .Y(_18140_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36347_ ( .A({ _18109_, _07122_ }), .Y(_18141_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36348_ ( .A({ _18110_, _07122_ }), .Y(_18142_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36349_ ( .A({ _18111_, _07122_ }), .Y(_18143_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36350_ ( .A({ _18112_, _07122_ }), .Y(_18144_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36351_ ( .A({ _18113_, _07122_ }), .Y(_18145_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36352_ ( .A({ _18114_, _07122_ }), .Y(_18146_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36353_ ( .A({ _18115_, _07122_ }), .Y(_18147_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36354_ ( .A({ _18116_, _07122_ }), .Y(_18148_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36355_ ( .A({ _18118_, _07122_ }), .Y(_18150_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36356_ ( .A({ _18119_, _07122_ }), .Y(_18151_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36357_ ( .A({ _21388_, _04901_ }), .Y(_21387_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36358_ ( .A({ _21486_, _04902_ }), .Y(_21485_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36359_ ( .A({ _21584_, _04903_ }), .Y(_21583_) );
  \$lut  #( .LUT(16'hff80), .WIDTH(4) ) _36360_ ( .A({ _RESETN_inv_2, _saxi_register_6[0], _maxi_read_idle, _maxi_write_idle }), .Y(rst_logic) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _36361_ ( .A({ _rst_logic_2, _rst_logic_1, rst_logic }), .Y(_00000_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36362_ ( .A({ _19428_, _05909_ }), .Y(_19460_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36363_ ( .A({ _19439_, _05909_ }), .Y(_19471_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36364_ ( .A({ _19450_, _05909_ }), .Y(_19482_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36365_ ( .A({ _19453_, _05909_ }), .Y(_19485_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36366_ ( .A({ _19454_, _05909_ }), .Y(_19486_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36367_ ( .A({ _19455_, _05909_ }), .Y(_19487_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36368_ ( .A({ _19456_, _05909_ }), .Y(_19488_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36369_ ( .A({ _19457_, _05909_ }), .Y(_19489_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36370_ ( .A({ _19458_, _05909_ }), .Y(_19490_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36371_ ( .A({ _19459_, _05909_ }), .Y(_19491_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36372_ ( .A({ _19429_, _05909_ }), .Y(_19461_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36373_ ( .A({ _19430_, _05909_ }), .Y(_19462_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36374_ ( .A({ _19431_, _05909_ }), .Y(_19463_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36375_ ( .A({ _19432_, _05909_ }), .Y(_19464_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36376_ ( .A({ _19433_, _05909_ }), .Y(_19465_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36377_ ( .A({ _19434_, _05909_ }), .Y(_19466_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36378_ ( .A({ _19435_, _05909_ }), .Y(_19467_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36379_ ( .A({ _19436_, _05909_ }), .Y(_19468_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36380_ ( .A({ _19437_, _05909_ }), .Y(_19469_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36381_ ( .A({ _19438_, _05909_ }), .Y(_19470_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36382_ ( .A({ _19440_, _05909_ }), .Y(_19472_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36383_ ( .A({ _19441_, _05909_ }), .Y(_19473_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36384_ ( .A({ _19442_, _05909_ }), .Y(_19474_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36385_ ( .A({ _19443_, _05909_ }), .Y(_19475_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36386_ ( .A({ _19444_, _05909_ }), .Y(_19476_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36387_ ( .A({ _19445_, _05909_ }), .Y(_19477_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36388_ ( .A({ _19446_, _05909_ }), .Y(_19478_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36389_ ( .A({ _19447_, _05909_ }), .Y(_19479_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36390_ ( .A({ _19448_, _05909_ }), .Y(_19480_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36391_ ( .A({ _19449_, _05909_ }), .Y(_19481_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36392_ ( .A({ _19451_, _05909_ }), .Y(_19483_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36393_ ( .A({ _19452_, _05909_ }), .Y(_19484_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36394_ ( .A({ _19492_, _05909_ }), .Y(_19494_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36395_ ( .A({ _19493_, _05909_ }), .Y(_19495_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36396_ ( .A({ _19496_, _05909_ }), .Y(_19528_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36397_ ( .A({ _19507_, _05909_ }), .Y(_19539_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36398_ ( .A({ _19518_, _05909_ }), .Y(_19550_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36399_ ( .A({ _19521_, _05909_ }), .Y(_19553_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36400_ ( .A({ _19522_, _05909_ }), .Y(_19554_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36401_ ( .A({ _19523_, _05909_ }), .Y(_19555_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36402_ ( .A({ _19524_, _05909_ }), .Y(_19556_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36403_ ( .A({ _19525_, _05909_ }), .Y(_19557_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36404_ ( .A({ _19526_, _05909_ }), .Y(_19558_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36405_ ( .A({ _19527_, _05909_ }), .Y(_19559_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36406_ ( .A({ _19497_, _05909_ }), .Y(_19529_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36407_ ( .A({ _19498_, _05909_ }), .Y(_19530_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36408_ ( .A({ _19499_, _05909_ }), .Y(_19531_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36409_ ( .A({ _19500_, _05909_ }), .Y(_19532_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36410_ ( .A({ _19501_, _05909_ }), .Y(_19533_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36411_ ( .A({ _19502_, _05909_ }), .Y(_19534_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36412_ ( .A({ _19503_, _05909_ }), .Y(_19535_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36413_ ( .A({ _19504_, _05909_ }), .Y(_19536_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36414_ ( .A({ _19505_, _05909_ }), .Y(_19537_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36415_ ( .A({ _19506_, _05909_ }), .Y(_19538_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36416_ ( .A({ _19508_, _05909_ }), .Y(_19540_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36417_ ( .A({ _19509_, _05909_ }), .Y(_19541_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36418_ ( .A({ _19510_, _05909_ }), .Y(_19542_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36419_ ( .A({ _19511_, _05909_ }), .Y(_19543_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36420_ ( .A({ _19512_, _05909_ }), .Y(_19544_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36421_ ( .A({ _19513_, _05909_ }), .Y(_19545_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36422_ ( .A({ _19514_, _05909_ }), .Y(_19546_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36423_ ( .A({ _19515_, _05909_ }), .Y(_19547_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36424_ ( .A({ _19516_, _05909_ }), .Y(_19548_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36425_ ( .A({ _19517_, _05909_ }), .Y(_19549_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36426_ ( .A({ _19519_, _05909_ }), .Y(_19551_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36427_ ( .A({ _19520_, _05909_ }), .Y(_19552_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36428_ ( .A({ _19560_, _05909_ }), .Y(_19592_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36429_ ( .A({ _19571_, _05909_ }), .Y(_19603_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36430_ ( .A({ _19582_, _05909_ }), .Y(_19614_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36431_ ( .A({ _19585_, _05909_ }), .Y(_19617_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36432_ ( .A({ _19586_, _05909_ }), .Y(_19618_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36433_ ( .A({ _19587_, _05909_ }), .Y(_19619_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36434_ ( .A({ _19588_, _05909_ }), .Y(_19620_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36435_ ( .A({ _19589_, _05909_ }), .Y(_19621_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36436_ ( .A({ _19590_, _05909_ }), .Y(_19622_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36437_ ( .A({ _19591_, _05909_ }), .Y(_19623_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36438_ ( .A({ _19561_, _05909_ }), .Y(_19593_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36439_ ( .A({ _19562_, _05909_ }), .Y(_19594_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36440_ ( .A({ _19563_, _05909_ }), .Y(_19595_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36441_ ( .A({ _19564_, _05909_ }), .Y(_19596_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36442_ ( .A({ _19565_, _05909_ }), .Y(_19597_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36443_ ( .A({ _19566_, _05909_ }), .Y(_19598_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36444_ ( .A({ _19567_, _05909_ }), .Y(_19599_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36445_ ( .A({ _19568_, _05909_ }), .Y(_19600_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36446_ ( .A({ _19569_, _05909_ }), .Y(_19601_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36447_ ( .A({ _19570_, _05909_ }), .Y(_19602_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36448_ ( .A({ _19572_, _05909_ }), .Y(_19604_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36449_ ( .A({ _19573_, _05909_ }), .Y(_19605_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36450_ ( .A({ _19574_, _05909_ }), .Y(_19606_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36451_ ( .A({ _19575_, _05909_ }), .Y(_19607_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36452_ ( .A({ _19576_, _05909_ }), .Y(_19608_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36453_ ( .A({ _19577_, _05909_ }), .Y(_19609_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36454_ ( .A({ _19578_, _05909_ }), .Y(_19610_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36455_ ( .A({ _19579_, _05909_ }), .Y(_19611_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36456_ ( .A({ _19580_, _05909_ }), .Y(_19612_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36457_ ( .A({ _19581_, _05909_ }), .Y(_19613_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36458_ ( .A({ _19583_, _05909_ }), .Y(_19615_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36459_ ( .A({ _19584_, _05909_ }), .Y(_19616_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36460_ ( .A({ _19624_, _05909_ }), .Y(_19656_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36461_ ( .A({ _19635_, _05909_ }), .Y(_19667_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36462_ ( .A({ _19646_, _05909_ }), .Y(_19678_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36463_ ( .A({ _19649_, _05909_ }), .Y(_19681_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36464_ ( .A({ _19650_, _05909_ }), .Y(_19682_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36465_ ( .A({ _19651_, _05909_ }), .Y(_19683_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36466_ ( .A({ _19652_, _05909_ }), .Y(_19684_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36467_ ( .A({ _19653_, _05909_ }), .Y(_19685_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36468_ ( .A({ _19654_, _05909_ }), .Y(_19686_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36469_ ( .A({ _19655_, _05909_ }), .Y(_19687_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36470_ ( .A({ _19625_, _05909_ }), .Y(_19657_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36471_ ( .A({ _19626_, _05909_ }), .Y(_19658_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36472_ ( .A({ _19627_, _05909_ }), .Y(_19659_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36473_ ( .A({ _19628_, _05909_ }), .Y(_19660_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36474_ ( .A({ _19629_, _05909_ }), .Y(_19661_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36475_ ( .A({ _19630_, _05909_ }), .Y(_19662_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36476_ ( .A({ _19631_, _05909_ }), .Y(_19663_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36477_ ( .A({ _19632_, _05909_ }), .Y(_19664_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36478_ ( .A({ _19633_, _05909_ }), .Y(_19665_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36479_ ( .A({ _19634_, _05909_ }), .Y(_19666_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36480_ ( .A({ _19636_, _05909_ }), .Y(_19668_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36481_ ( .A({ _19637_, _05909_ }), .Y(_19669_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36482_ ( .A({ _19638_, _05909_ }), .Y(_19670_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36483_ ( .A({ _19639_, _05909_ }), .Y(_19671_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36484_ ( .A({ _19640_, _05909_ }), .Y(_19672_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36485_ ( .A({ _19641_, _05909_ }), .Y(_19673_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36486_ ( .A({ _19642_, _05909_ }), .Y(_19674_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36487_ ( .A({ _19643_, _05909_ }), .Y(_19675_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36488_ ( .A({ _19644_, _05909_ }), .Y(_19676_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36489_ ( .A({ _19645_, _05909_ }), .Y(_19677_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36490_ ( .A({ _19647_, _05909_ }), .Y(_19679_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36491_ ( .A({ _19648_, _05909_ }), .Y(_19680_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36492_ ( .A({ _03930_, _06338_ }), .Y(_19688_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36493_ ( .A({ _03941_, _06338_ }), .Y(_19699_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36494_ ( .A({ _03952_, _06338_ }), .Y(_19710_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36495_ ( .A({ _03955_, _06338_ }), .Y(_19713_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36496_ ( .A({ _03956_, _06338_ }), .Y(_19714_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36497_ ( .A({ _03957_, _06338_ }), .Y(_19715_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36498_ ( .A({ _03958_, _06338_ }), .Y(_19716_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36499_ ( .A({ _03959_, _06338_ }), .Y(_19717_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36500_ ( .A({ _03960_, _06338_ }), .Y(_19718_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36501_ ( .A({ _03961_, _06338_ }), .Y(_19719_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36502_ ( .A({ _03931_, _06338_ }), .Y(_19689_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36503_ ( .A({ _03932_, _06338_ }), .Y(_19690_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36504_ ( .A({ _03933_, _06338_ }), .Y(_19691_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36505_ ( .A({ _03934_, _06338_ }), .Y(_19692_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36506_ ( .A({ _03935_, _06338_ }), .Y(_19693_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36507_ ( .A({ _03936_, _06338_ }), .Y(_19694_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36508_ ( .A({ _03937_, _06338_ }), .Y(_19695_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36509_ ( .A({ _03938_, _06338_ }), .Y(_19696_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36510_ ( .A({ _03939_, _06338_ }), .Y(_19697_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36511_ ( .A({ _03940_, _06338_ }), .Y(_19698_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36512_ ( .A({ _03942_, _06338_ }), .Y(_19700_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36513_ ( .A({ _03943_, _06338_ }), .Y(_19701_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36514_ ( .A({ _03944_, _06338_ }), .Y(_19702_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36515_ ( .A({ _03945_, _06338_ }), .Y(_19703_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36516_ ( .A({ _03946_, _06338_ }), .Y(_19704_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36517_ ( .A({ _03947_, _06338_ }), .Y(_19705_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36518_ ( .A({ _03948_, _06338_ }), .Y(_19706_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36519_ ( .A({ _03949_, _06338_ }), .Y(_19707_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36520_ ( .A({ _03950_, _06338_ }), .Y(_19708_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36521_ ( .A({ _03951_, _06338_ }), .Y(_19709_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36522_ ( .A({ _03953_, _06338_ }), .Y(_19711_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36523_ ( .A({ _03954_, _06338_ }), .Y(_19712_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36524_ ( .A({ _19722_, _05909_ }), .Y(_19754_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36525_ ( .A({ _19733_, _05909_ }), .Y(_19765_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36526_ ( .A({ _19744_, _05909_ }), .Y(_19776_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36527_ ( .A({ _19747_, _05909_ }), .Y(_19779_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36528_ ( .A({ _19748_, _05909_ }), .Y(_19780_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36529_ ( .A({ _19749_, _05909_ }), .Y(_19781_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36530_ ( .A({ _19750_, _05909_ }), .Y(_19782_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36531_ ( .A({ _19751_, _05909_ }), .Y(_19783_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36532_ ( .A({ _19752_, _05909_ }), .Y(_19784_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36533_ ( .A({ _19753_, _05909_ }), .Y(_19785_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36534_ ( .A({ _19723_, _05909_ }), .Y(_19755_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36535_ ( .A({ _19724_, _05909_ }), .Y(_19756_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36536_ ( .A({ _19725_, _05909_ }), .Y(_19757_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36537_ ( .A({ _19726_, _05909_ }), .Y(_19758_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36538_ ( .A({ _19727_, _05909_ }), .Y(_19759_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36539_ ( .A({ _19728_, _05909_ }), .Y(_19760_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36540_ ( .A({ _19729_, _05909_ }), .Y(_19761_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36541_ ( .A({ _19730_, _05909_ }), .Y(_19762_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36542_ ( .A({ _19731_, _05909_ }), .Y(_19763_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36543_ ( .A({ _19732_, _05909_ }), .Y(_19764_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36544_ ( .A({ _19734_, _05909_ }), .Y(_19766_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36545_ ( .A({ _19735_, _05909_ }), .Y(_19767_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36546_ ( .A({ _19736_, _05909_ }), .Y(_19768_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36547_ ( .A({ _19737_, _05909_ }), .Y(_19769_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36548_ ( .A({ _19738_, _05909_ }), .Y(_19770_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36549_ ( .A({ _19739_, _05909_ }), .Y(_19771_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36550_ ( .A({ _19740_, _05909_ }), .Y(_19772_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36551_ ( .A({ _19741_, _05909_ }), .Y(_19773_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36552_ ( .A({ _19742_, _05909_ }), .Y(_19774_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36553_ ( .A({ _19743_, _05909_ }), .Y(_19775_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36554_ ( .A({ _19745_, _05909_ }), .Y(_19777_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36555_ ( .A({ _19746_, _05909_ }), .Y(_19778_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36556_ ( .A({ _18622_, _05909_ }), .Y(_18654_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36557_ ( .A({ _18633_, _05909_ }), .Y(_18665_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36558_ ( .A({ _18644_, _05909_ }), .Y(_18676_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36559_ ( .A({ _18647_, _05909_ }), .Y(_18679_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36560_ ( .A({ _18648_, _05909_ }), .Y(_18680_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36561_ ( .A({ _18649_, _05909_ }), .Y(_18681_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36562_ ( .A({ _18650_, _05909_ }), .Y(_18682_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36563_ ( .A({ _18651_, _05909_ }), .Y(_18683_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36564_ ( .A({ _18652_, _05909_ }), .Y(_18684_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36565_ ( .A({ _18653_, _05909_ }), .Y(_18685_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36566_ ( .A({ _18623_, _05909_ }), .Y(_18655_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36567_ ( .A({ _18624_, _05909_ }), .Y(_18656_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36568_ ( .A({ _18625_, _05909_ }), .Y(_18657_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36569_ ( .A({ _18626_, _05909_ }), .Y(_18658_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36570_ ( .A({ _18627_, _05909_ }), .Y(_18659_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36571_ ( .A({ _18628_, _05909_ }), .Y(_18660_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36572_ ( .A({ _18629_, _05909_ }), .Y(_18661_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36573_ ( .A({ _18630_, _05909_ }), .Y(_18662_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36574_ ( .A({ _18631_, _05909_ }), .Y(_18663_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36575_ ( .A({ _18632_, _05909_ }), .Y(_18664_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36576_ ( .A({ _18634_, _05909_ }), .Y(_18666_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36577_ ( .A({ _18635_, _05909_ }), .Y(_18667_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36578_ ( .A({ _18636_, _05909_ }), .Y(_18668_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36579_ ( .A({ _18637_, _05909_ }), .Y(_18669_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36580_ ( .A({ _18638_, _05909_ }), .Y(_18670_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36581_ ( .A({ _18639_, _05909_ }), .Y(_18671_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36582_ ( .A({ _18640_, _05909_ }), .Y(_18672_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36583_ ( .A({ _18641_, _05909_ }), .Y(_18673_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36584_ ( .A({ _18642_, _05909_ }), .Y(_18674_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36585_ ( .A({ _18643_, _05909_ }), .Y(_18675_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36586_ ( .A({ _18645_, _05909_ }), .Y(_18677_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36587_ ( .A({ _18646_, _05909_ }), .Y(_18678_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36588_ ( .A({ _19786_, _05909_ }), .Y(_19818_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36589_ ( .A({ _19797_, _05909_ }), .Y(_19829_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36590_ ( .A({ _19808_, _05909_ }), .Y(_19840_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36591_ ( .A({ _19811_, _05909_ }), .Y(_19843_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36592_ ( .A({ _19812_, _05909_ }), .Y(_19844_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36593_ ( .A({ _19813_, _05909_ }), .Y(_19845_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36594_ ( .A({ _19814_, _05909_ }), .Y(_19846_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36595_ ( .A({ _19815_, _05909_ }), .Y(_19847_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36596_ ( .A({ _19816_, _05909_ }), .Y(_19848_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36597_ ( .A({ _19817_, _05909_ }), .Y(_19849_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36598_ ( .A({ _19787_, _05909_ }), .Y(_19819_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36599_ ( .A({ _19788_, _05909_ }), .Y(_19820_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36600_ ( .A({ _19789_, _05909_ }), .Y(_19821_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36601_ ( .A({ _19790_, _05909_ }), .Y(_19822_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36602_ ( .A({ _19791_, _05909_ }), .Y(_19823_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36603_ ( .A({ _19792_, _05909_ }), .Y(_19824_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36604_ ( .A({ _19793_, _05909_ }), .Y(_19825_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36605_ ( .A({ _19794_, _05909_ }), .Y(_19826_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36606_ ( .A({ _19795_, _05909_ }), .Y(_19827_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36607_ ( .A({ _19796_, _05909_ }), .Y(_19828_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36608_ ( .A({ _19798_, _05909_ }), .Y(_19830_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36609_ ( .A({ _19799_, _05909_ }), .Y(_19831_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36610_ ( .A({ _19800_, _05909_ }), .Y(_19832_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36611_ ( .A({ _19801_, _05909_ }), .Y(_19833_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36612_ ( .A({ _19802_, _05909_ }), .Y(_19834_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36613_ ( .A({ _19803_, _05909_ }), .Y(_19835_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36614_ ( .A({ _19804_, _05909_ }), .Y(_19836_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36615_ ( .A({ _19805_, _05909_ }), .Y(_19837_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36616_ ( .A({ _19806_, _05909_ }), .Y(_19838_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36617_ ( .A({ _19807_, _05909_ }), .Y(_19839_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36618_ ( .A({ _19809_, _05909_ }), .Y(_19841_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36619_ ( .A({ _19810_, _05909_ }), .Y(_19842_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36620_ ( .A({ _19850_, _05909_ }), .Y(_19882_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36621_ ( .A({ _19861_, _05909_ }), .Y(_19893_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36622_ ( .A({ _19872_, _05909_ }), .Y(_19904_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36623_ ( .A({ _19875_, _05909_ }), .Y(_19907_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36624_ ( .A({ _19876_, _05909_ }), .Y(_19908_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36625_ ( .A({ _19877_, _05909_ }), .Y(_19909_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36626_ ( .A({ _19878_, _05909_ }), .Y(_19910_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36627_ ( .A({ _19879_, _05909_ }), .Y(_19911_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36628_ ( .A({ _19880_, _05909_ }), .Y(_19912_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36629_ ( .A({ _19881_, _05909_ }), .Y(_19913_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36630_ ( .A({ _19851_, _05909_ }), .Y(_19883_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36631_ ( .A({ _19852_, _05909_ }), .Y(_19884_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36632_ ( .A({ _19853_, _05909_ }), .Y(_19885_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36633_ ( .A({ _19854_, _05909_ }), .Y(_19886_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36634_ ( .A({ _19855_, _05909_ }), .Y(_19887_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36635_ ( .A({ _19856_, _05909_ }), .Y(_19888_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36636_ ( .A({ _19857_, _05909_ }), .Y(_19889_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36637_ ( .A({ _19858_, _05909_ }), .Y(_19890_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36638_ ( .A({ _19859_, _05909_ }), .Y(_19891_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36639_ ( .A({ _19860_, _05909_ }), .Y(_19892_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36640_ ( .A({ _19862_, _05909_ }), .Y(_19894_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36641_ ( .A({ _19863_, _05909_ }), .Y(_19895_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36642_ ( .A({ _19864_, _05909_ }), .Y(_19896_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36643_ ( .A({ _19865_, _05909_ }), .Y(_19897_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36644_ ( .A({ _19866_, _05909_ }), .Y(_19898_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36645_ ( .A({ _19867_, _05909_ }), .Y(_19899_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36646_ ( .A({ _19868_, _05909_ }), .Y(_19900_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36647_ ( .A({ _19869_, _05909_ }), .Y(_19901_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36648_ ( .A({ _19870_, _05909_ }), .Y(_19902_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36649_ ( .A({ _19871_, _05909_ }), .Y(_19903_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36650_ ( .A({ _19873_, _05909_ }), .Y(_19905_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36651_ ( .A({ _19874_, _05909_ }), .Y(_19906_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36652_ ( .A({ _18686_, _05909_ }), .Y(_18718_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36653_ ( .A({ _18697_, _05909_ }), .Y(_18729_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36654_ ( .A({ _18708_, _05909_ }), .Y(_18740_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36655_ ( .A({ _18711_, _05909_ }), .Y(_18743_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36656_ ( .A({ _18712_, _05909_ }), .Y(_18744_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36657_ ( .A({ _18713_, _05909_ }), .Y(_18745_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36658_ ( .A({ _18714_, _05909_ }), .Y(_18746_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36659_ ( .A({ _18715_, _05909_ }), .Y(_18747_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36660_ ( .A({ _18716_, _05909_ }), .Y(_18748_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36661_ ( .A({ _18717_, _05909_ }), .Y(_18749_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36662_ ( .A({ _18687_, _05909_ }), .Y(_18719_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36663_ ( .A({ _18688_, _05909_ }), .Y(_18720_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36664_ ( .A({ _18689_, _05909_ }), .Y(_18721_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36665_ ( .A({ _18690_, _05909_ }), .Y(_18722_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36666_ ( .A({ _18691_, _05909_ }), .Y(_18723_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36667_ ( .A({ _18692_, _05909_ }), .Y(_18724_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36668_ ( .A({ _18693_, _05909_ }), .Y(_18725_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36669_ ( .A({ _18694_, _05909_ }), .Y(_18726_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36670_ ( .A({ _18695_, _05909_ }), .Y(_18727_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36671_ ( .A({ _18696_, _05909_ }), .Y(_18728_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36672_ ( .A({ _18698_, _05909_ }), .Y(_18730_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36673_ ( .A({ _18699_, _05909_ }), .Y(_18731_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36674_ ( .A({ _18700_, _05909_ }), .Y(_18732_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36675_ ( .A({ _18701_, _05909_ }), .Y(_18733_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36676_ ( .A({ _18702_, _05909_ }), .Y(_18734_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36677_ ( .A({ _18703_, _05909_ }), .Y(_18735_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36678_ ( .A({ _18704_, _05909_ }), .Y(_18736_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36679_ ( .A({ _18705_, _05909_ }), .Y(_18737_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36680_ ( .A({ _18706_, _05909_ }), .Y(_18738_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36681_ ( .A({ _18707_, _05909_ }), .Y(_18739_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36682_ ( .A({ _18709_, _05909_ }), .Y(_18741_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36683_ ( .A({ _18710_, _05909_ }), .Y(_18742_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36684_ ( .A({ _18750_, _05909_ }), .Y(_18751_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36685_ ( .A({ _19914_, _05909_ }), .Y(_19946_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36686_ ( .A({ _19925_, _05909_ }), .Y(_19957_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36687_ ( .A({ _19936_, _05909_ }), .Y(_19968_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36688_ ( .A({ _19939_, _05909_ }), .Y(_19971_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36689_ ( .A({ _19940_, _05909_ }), .Y(_19972_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36690_ ( .A({ _19941_, _05909_ }), .Y(_19973_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36691_ ( .A({ _19942_, _05909_ }), .Y(_19974_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36692_ ( .A({ _19943_, _05909_ }), .Y(_19975_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36693_ ( .A({ _19944_, _05909_ }), .Y(_19976_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36694_ ( .A({ _19945_, _05909_ }), .Y(_19977_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36695_ ( .A({ _19915_, _05909_ }), .Y(_19947_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36696_ ( .A({ _19916_, _05909_ }), .Y(_19948_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36697_ ( .A({ _19917_, _05909_ }), .Y(_19949_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36698_ ( .A({ _19918_, _05909_ }), .Y(_19950_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36699_ ( .A({ _19919_, _05909_ }), .Y(_19951_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36700_ ( .A({ _19920_, _05909_ }), .Y(_19952_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36701_ ( .A({ _19921_, _05909_ }), .Y(_19953_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36702_ ( .A({ _19922_, _05909_ }), .Y(_19954_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36703_ ( .A({ _19923_, _05909_ }), .Y(_19955_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36704_ ( .A({ _19924_, _05909_ }), .Y(_19956_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36705_ ( .A({ _19926_, _05909_ }), .Y(_19958_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36706_ ( .A({ _19927_, _05909_ }), .Y(_19959_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36707_ ( .A({ _19928_, _05909_ }), .Y(_19960_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36708_ ( .A({ _19929_, _05909_ }), .Y(_19961_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36709_ ( .A({ _19930_, _05909_ }), .Y(_19962_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36710_ ( .A({ _19931_, _05909_ }), .Y(_19963_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36711_ ( .A({ _19932_, _05909_ }), .Y(_19964_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36712_ ( .A({ _19933_, _05909_ }), .Y(_19965_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36713_ ( .A({ _19934_, _05909_ }), .Y(_19966_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36714_ ( .A({ _19935_, _05909_ }), .Y(_19967_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36715_ ( .A({ _19937_, _05909_ }), .Y(_19969_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36716_ ( .A({ _19938_, _05909_ }), .Y(_19970_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36717_ ( .A({ _19978_, _05909_ }), .Y(_20010_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36718_ ( .A({ _19989_, _05909_ }), .Y(_20021_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36719_ ( .A({ _20000_, _05909_ }), .Y(_20032_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36720_ ( .A({ _20003_, _05909_ }), .Y(_20035_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36721_ ( .A({ _20004_, _05909_ }), .Y(_20036_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36722_ ( .A({ _20005_, _05909_ }), .Y(_20037_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36723_ ( .A({ _20006_, _05909_ }), .Y(_20038_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36724_ ( .A({ _20007_, _05909_ }), .Y(_20039_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36725_ ( .A({ _20008_, _05909_ }), .Y(_20040_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36726_ ( .A({ _20009_, _05909_ }), .Y(_20041_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36727_ ( .A({ _19979_, _05909_ }), .Y(_20011_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36728_ ( .A({ _19980_, _05909_ }), .Y(_20012_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36729_ ( .A({ _19981_, _05909_ }), .Y(_20013_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36730_ ( .A({ _19982_, _05909_ }), .Y(_20014_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36731_ ( .A({ _19983_, _05909_ }), .Y(_20015_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36732_ ( .A({ _19984_, _05909_ }), .Y(_20016_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36733_ ( .A({ _19985_, _05909_ }), .Y(_20017_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36734_ ( .A({ _19986_, _05909_ }), .Y(_20018_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36735_ ( .A({ _19987_, _05909_ }), .Y(_20019_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36736_ ( .A({ _19988_, _05909_ }), .Y(_20020_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36737_ ( .A({ _19990_, _05909_ }), .Y(_20022_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36738_ ( .A({ _19991_, _05909_ }), .Y(_20023_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36739_ ( .A({ _19992_, _05909_ }), .Y(_20024_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36740_ ( .A({ _19993_, _05909_ }), .Y(_20025_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36741_ ( .A({ _19994_, _05909_ }), .Y(_20026_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36742_ ( .A({ _19995_, _05909_ }), .Y(_20027_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36743_ ( .A({ _19996_, _05909_ }), .Y(_20028_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36744_ ( .A({ _19997_, _05909_ }), .Y(_20029_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36745_ ( .A({ _19998_, _05909_ }), .Y(_20030_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36746_ ( .A({ _19999_, _05909_ }), .Y(_20031_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36747_ ( .A({ _20001_, _05909_ }), .Y(_20033_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36748_ ( .A({ _20002_, _05909_ }), .Y(_20034_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36749_ ( .A({ _14441_, _06012_ }), .Y(_14473_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36750_ ( .A({ _14452_, _06012_ }), .Y(_14484_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36751_ ( .A({ _14463_, _06012_ }), .Y(_14495_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36752_ ( .A({ _14466_, _06012_ }), .Y(_14498_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36753_ ( .A({ _14467_, _06012_ }), .Y(_14499_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36754_ ( .A({ _14468_, _06012_ }), .Y(_14500_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36755_ ( .A({ _14469_, _06012_ }), .Y(_14501_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36756_ ( .A({ _14470_, _06012_ }), .Y(_14502_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36757_ ( .A({ _14471_, _06012_ }), .Y(_14503_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36758_ ( .A({ _14472_, _06012_ }), .Y(_14504_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36759_ ( .A({ _14442_, _06012_ }), .Y(_14474_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36760_ ( .A({ _14443_, _06012_ }), .Y(_14475_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36761_ ( .A({ _14444_, _06012_ }), .Y(_14476_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36762_ ( .A({ _14445_, _06012_ }), .Y(_14477_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36763_ ( .A({ _14446_, _06012_ }), .Y(_14478_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36764_ ( .A({ _14447_, _06012_ }), .Y(_14479_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36765_ ( .A({ _14448_, _06012_ }), .Y(_14480_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36766_ ( .A({ _14449_, _06012_ }), .Y(_14481_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36767_ ( .A({ _14450_, _06012_ }), .Y(_14482_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36768_ ( .A({ _14451_, _06012_ }), .Y(_14483_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36769_ ( .A({ _14453_, _06012_ }), .Y(_14485_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36770_ ( .A({ _14454_, _06012_ }), .Y(_14486_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36771_ ( .A({ _14455_, _06012_ }), .Y(_14487_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36772_ ( .A({ _14456_, _06012_ }), .Y(_14488_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36773_ ( .A({ _14457_, _06012_ }), .Y(_14489_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36774_ ( .A({ _14458_, _06012_ }), .Y(_14490_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36775_ ( .A({ _14459_, _06012_ }), .Y(_14491_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36776_ ( .A({ _14460_, _06012_ }), .Y(_14492_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36777_ ( .A({ _14461_, _06012_ }), .Y(_14493_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36778_ ( .A({ _14462_, _06012_ }), .Y(_14494_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36779_ ( .A({ _14464_, _06012_ }), .Y(_14496_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36780_ ( .A({ _14465_, _06012_ }), .Y(_14497_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36781_ ( .A({ _18752_, _05909_ }), .Y(_18784_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36782_ ( .A({ _18763_, _05909_ }), .Y(_18795_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36783_ ( .A({ _18774_, _05909_ }), .Y(_18806_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36784_ ( .A({ _18777_, _05909_ }), .Y(_18809_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36785_ ( .A({ _18778_, _05909_ }), .Y(_18810_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36786_ ( .A({ _18779_, _05909_ }), .Y(_18811_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36787_ ( .A({ _18780_, _05909_ }), .Y(_18812_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36788_ ( .A({ _18781_, _05909_ }), .Y(_18813_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36789_ ( .A({ _18782_, _05909_ }), .Y(_18814_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36790_ ( .A({ _18783_, _05909_ }), .Y(_18815_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36791_ ( .A({ _18753_, _05909_ }), .Y(_18785_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36792_ ( .A({ _18754_, _05909_ }), .Y(_18786_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36793_ ( .A({ _18755_, _05909_ }), .Y(_18787_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36794_ ( .A({ _18756_, _05909_ }), .Y(_18788_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36795_ ( .A({ _18757_, _05909_ }), .Y(_18789_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36796_ ( .A({ _18758_, _05909_ }), .Y(_18790_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36797_ ( .A({ _18759_, _05909_ }), .Y(_18791_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36798_ ( .A({ _18760_, _05909_ }), .Y(_18792_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36799_ ( .A({ _18761_, _05909_ }), .Y(_18793_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36800_ ( .A({ _18762_, _05909_ }), .Y(_18794_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36801_ ( .A({ _18764_, _05909_ }), .Y(_18796_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36802_ ( .A({ _18765_, _05909_ }), .Y(_18797_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36803_ ( .A({ _18766_, _05909_ }), .Y(_18798_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36804_ ( .A({ _18767_, _05909_ }), .Y(_18799_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36805_ ( .A({ _18768_, _05909_ }), .Y(_18800_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36806_ ( .A({ _18769_, _05909_ }), .Y(_18801_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36807_ ( .A({ _18770_, _05909_ }), .Y(_18802_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36808_ ( .A({ _18771_, _05909_ }), .Y(_18803_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36809_ ( .A({ _18772_, _05909_ }), .Y(_18804_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36810_ ( .A({ _18773_, _05909_ }), .Y(_18805_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36811_ ( .A({ _18775_, _05909_ }), .Y(_18807_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36812_ ( .A({ _18776_, _05909_ }), .Y(_18808_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36813_ ( .A({ _14505_, _06012_ }), .Y(_14537_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36814_ ( .A({ _14516_, _06012_ }), .Y(_14548_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36815_ ( .A({ _14527_, _06012_ }), .Y(_14559_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36816_ ( .A({ _14530_, _06012_ }), .Y(_14562_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36817_ ( .A({ _14531_, _06012_ }), .Y(_14563_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36818_ ( .A({ _14532_, _06012_ }), .Y(_14564_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36819_ ( .A({ _14533_, _06012_ }), .Y(_14565_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36820_ ( .A({ _14534_, _06012_ }), .Y(_14566_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36821_ ( .A({ _14535_, _06012_ }), .Y(_14567_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36822_ ( .A({ _14536_, _06012_ }), .Y(_14568_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36823_ ( .A({ _14506_, _06012_ }), .Y(_14538_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36824_ ( .A({ _14507_, _06012_ }), .Y(_14539_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36825_ ( .A({ _14508_, _06012_ }), .Y(_14540_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36826_ ( .A({ _14509_, _06012_ }), .Y(_14541_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36827_ ( .A({ _14510_, _06012_ }), .Y(_14542_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36828_ ( .A({ _14511_, _06012_ }), .Y(_14543_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36829_ ( .A({ _14512_, _06012_ }), .Y(_14544_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36830_ ( .A({ _14513_, _06012_ }), .Y(_14545_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36831_ ( .A({ _14514_, _06012_ }), .Y(_14546_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36832_ ( .A({ _14515_, _06012_ }), .Y(_14547_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36833_ ( .A({ _14517_, _06012_ }), .Y(_14549_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36834_ ( .A({ _14518_, _06012_ }), .Y(_14550_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36835_ ( .A({ _14519_, _06012_ }), .Y(_14551_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36836_ ( .A({ _14520_, _06012_ }), .Y(_14552_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36837_ ( .A({ _14521_, _06012_ }), .Y(_14553_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36838_ ( .A({ _14522_, _06012_ }), .Y(_14554_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36839_ ( .A({ _14523_, _06012_ }), .Y(_14555_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36840_ ( .A({ _14524_, _06012_ }), .Y(_14556_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36841_ ( .A({ _14525_, _06012_ }), .Y(_14557_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36842_ ( .A({ _14526_, _06012_ }), .Y(_14558_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36843_ ( .A({ _14528_, _06012_ }), .Y(_14560_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36844_ ( .A({ _14529_, _06012_ }), .Y(_14561_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36845_ ( .A({ _20042_, _05909_ }), .Y(_20074_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36846_ ( .A({ _20053_, _05909_ }), .Y(_20085_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36847_ ( .A({ _20064_, _05909_ }), .Y(_20096_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36848_ ( .A({ _20067_, _05909_ }), .Y(_20099_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36849_ ( .A({ _20068_, _05909_ }), .Y(_20100_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36850_ ( .A({ _20069_, _05909_ }), .Y(_20101_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36851_ ( .A({ _20070_, _05909_ }), .Y(_20102_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36852_ ( .A({ _20071_, _05909_ }), .Y(_20103_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36853_ ( .A({ _20072_, _05909_ }), .Y(_20104_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36854_ ( .A({ _20073_, _05909_ }), .Y(_20105_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36855_ ( .A({ _20043_, _05909_ }), .Y(_20075_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36856_ ( .A({ _20044_, _05909_ }), .Y(_20076_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36857_ ( .A({ _20045_, _05909_ }), .Y(_20077_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36858_ ( .A({ _20046_, _05909_ }), .Y(_20078_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36859_ ( .A({ _20047_, _05909_ }), .Y(_20079_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36860_ ( .A({ _20048_, _05909_ }), .Y(_20080_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36861_ ( .A({ _20049_, _05909_ }), .Y(_20081_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36862_ ( .A({ _20050_, _05909_ }), .Y(_20082_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36863_ ( .A({ _20051_, _05909_ }), .Y(_20083_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36864_ ( .A({ _20052_, _05909_ }), .Y(_20084_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36865_ ( .A({ _20054_, _05909_ }), .Y(_20086_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36866_ ( .A({ _20055_, _05909_ }), .Y(_20087_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36867_ ( .A({ _20056_, _05909_ }), .Y(_20088_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36868_ ( .A({ _20057_, _05909_ }), .Y(_20089_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36869_ ( .A({ _20058_, _05909_ }), .Y(_20090_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36870_ ( .A({ _20059_, _05909_ }), .Y(_20091_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36871_ ( .A({ _20060_, _05909_ }), .Y(_20092_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36872_ ( .A({ _20061_, _05909_ }), .Y(_20093_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36873_ ( .A({ _20062_, _05909_ }), .Y(_20094_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36874_ ( .A({ _20063_, _05909_ }), .Y(_20095_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36875_ ( .A({ _20065_, _05909_ }), .Y(_20097_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36876_ ( .A({ _20066_, _05909_ }), .Y(_20098_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36877_ ( .A({ _14313_, _06012_ }), .Y(_14345_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36878_ ( .A({ _14324_, _06012_ }), .Y(_14356_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36879_ ( .A({ _14335_, _06012_ }), .Y(_14367_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36880_ ( .A({ _14338_, _06012_ }), .Y(_14370_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36881_ ( .A({ _14339_, _06012_ }), .Y(_14371_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36882_ ( .A({ _14340_, _06012_ }), .Y(_14372_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36883_ ( .A({ _14341_, _06012_ }), .Y(_14373_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36884_ ( .A({ _14342_, _06012_ }), .Y(_14374_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36885_ ( .A({ _14343_, _06012_ }), .Y(_14375_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36886_ ( .A({ _14344_, _06012_ }), .Y(_14376_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36887_ ( .A({ _14314_, _06012_ }), .Y(_14346_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36888_ ( .A({ _14315_, _06012_ }), .Y(_14347_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36889_ ( .A({ _14316_, _06012_ }), .Y(_14348_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36890_ ( .A({ _14317_, _06012_ }), .Y(_14349_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36891_ ( .A({ _14318_, _06012_ }), .Y(_14350_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36892_ ( .A({ _14319_, _06012_ }), .Y(_14351_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36893_ ( .A({ _14320_, _06012_ }), .Y(_14352_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36894_ ( .A({ _14321_, _06012_ }), .Y(_14353_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36895_ ( .A({ _14322_, _06012_ }), .Y(_14354_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36896_ ( .A({ _14323_, _06012_ }), .Y(_14355_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36897_ ( .A({ _14325_, _06012_ }), .Y(_14357_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36898_ ( .A({ _14326_, _06012_ }), .Y(_14358_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36899_ ( .A({ _14327_, _06012_ }), .Y(_14359_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36900_ ( .A({ _14328_, _06012_ }), .Y(_14360_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36901_ ( .A({ _14329_, _06012_ }), .Y(_14361_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36902_ ( .A({ _14330_, _06012_ }), .Y(_14362_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36903_ ( .A({ _14331_, _06012_ }), .Y(_14363_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36904_ ( .A({ _14332_, _06012_ }), .Y(_14364_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36905_ ( .A({ _14333_, _06012_ }), .Y(_14365_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36906_ ( .A({ _14334_, _06012_ }), .Y(_14366_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36907_ ( .A({ _14336_, _06012_ }), .Y(_14368_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36908_ ( .A({ _14337_, _06012_ }), .Y(_14369_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36909_ ( .A({ _14377_, _06012_ }), .Y(_14409_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36910_ ( .A({ _14388_, _06012_ }), .Y(_14420_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36911_ ( .A({ _14399_, _06012_ }), .Y(_14431_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36912_ ( .A({ _14402_, _06012_ }), .Y(_14434_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36913_ ( .A({ _14403_, _06012_ }), .Y(_14435_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36914_ ( .A({ _14404_, _06012_ }), .Y(_14436_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36915_ ( .A({ _14405_, _06012_ }), .Y(_14437_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36916_ ( .A({ _14406_, _06012_ }), .Y(_14438_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36917_ ( .A({ _14407_, _06012_ }), .Y(_14439_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36918_ ( .A({ _14408_, _06012_ }), .Y(_14440_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36919_ ( .A({ _14378_, _06012_ }), .Y(_14410_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36920_ ( .A({ _14379_, _06012_ }), .Y(_14411_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36921_ ( .A({ _14380_, _06012_ }), .Y(_14412_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36922_ ( .A({ _14381_, _06012_ }), .Y(_14413_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36923_ ( .A({ _14382_, _06012_ }), .Y(_14414_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36924_ ( .A({ _14383_, _06012_ }), .Y(_14415_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36925_ ( .A({ _14384_, _06012_ }), .Y(_14416_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36926_ ( .A({ _14385_, _06012_ }), .Y(_14417_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36927_ ( .A({ _14386_, _06012_ }), .Y(_14418_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36928_ ( .A({ _14387_, _06012_ }), .Y(_14419_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36929_ ( .A({ _14389_, _06012_ }), .Y(_14421_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36930_ ( .A({ _14390_, _06012_ }), .Y(_14422_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36931_ ( .A({ _14391_, _06012_ }), .Y(_14423_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36932_ ( .A({ _14392_, _06012_ }), .Y(_14424_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36933_ ( .A({ _14393_, _06012_ }), .Y(_14425_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36934_ ( .A({ _14394_, _06012_ }), .Y(_14426_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36935_ ( .A({ _14395_, _06012_ }), .Y(_14427_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36936_ ( .A({ _14396_, _06012_ }), .Y(_14428_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36937_ ( .A({ _14397_, _06012_ }), .Y(_14429_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36938_ ( .A({ _14398_, _06012_ }), .Y(_14430_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36939_ ( .A({ _14400_, _06012_ }), .Y(_14432_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36940_ ( .A({ _14401_, _06012_ }), .Y(_14433_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36941_ ( .A({ _20106_, _05909_ }), .Y(_20138_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36942_ ( .A({ _20117_, _05909_ }), .Y(_20149_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36943_ ( .A({ _20128_, _05909_ }), .Y(_20160_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36944_ ( .A({ _20131_, _05909_ }), .Y(_20163_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36945_ ( .A({ _20132_, _05909_ }), .Y(_20164_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36946_ ( .A({ _20133_, _05909_ }), .Y(_20165_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36947_ ( .A({ _20134_, _05909_ }), .Y(_20166_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36948_ ( .A({ _20135_, _05909_ }), .Y(_20167_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36949_ ( .A({ _20136_, _05909_ }), .Y(_20168_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36950_ ( .A({ _20137_, _05909_ }), .Y(_20169_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36951_ ( .A({ _20107_, _05909_ }), .Y(_20139_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36952_ ( .A({ _20108_, _05909_ }), .Y(_20140_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36953_ ( .A({ _20109_, _05909_ }), .Y(_20141_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36954_ ( .A({ _20110_, _05909_ }), .Y(_20142_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36955_ ( .A({ _20111_, _05909_ }), .Y(_20143_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36956_ ( .A({ _20112_, _05909_ }), .Y(_20144_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36957_ ( .A({ _20113_, _05909_ }), .Y(_20145_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36958_ ( .A({ _20114_, _05909_ }), .Y(_20146_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36959_ ( .A({ _20115_, _05909_ }), .Y(_20147_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36960_ ( .A({ _20116_, _05909_ }), .Y(_20148_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36961_ ( .A({ _20118_, _05909_ }), .Y(_20150_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36962_ ( .A({ _20119_, _05909_ }), .Y(_20151_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36963_ ( .A({ _20120_, _05909_ }), .Y(_20152_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36964_ ( .A({ _20121_, _05909_ }), .Y(_20153_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36965_ ( .A({ _20122_, _05909_ }), .Y(_20154_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36966_ ( .A({ _20123_, _05909_ }), .Y(_20155_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36967_ ( .A({ _20124_, _05909_ }), .Y(_20156_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36968_ ( .A({ _20125_, _05909_ }), .Y(_20157_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36969_ ( .A({ _20126_, _05909_ }), .Y(_20158_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36970_ ( .A({ _20127_, _05909_ }), .Y(_20159_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36971_ ( .A({ _20129_, _05909_ }), .Y(_20161_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36972_ ( .A({ _20130_, _05909_ }), .Y(_20162_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36973_ ( .A({ _14249_, _06012_ }), .Y(_14281_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36974_ ( .A({ _14260_, _06012_ }), .Y(_14292_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36975_ ( .A({ _14271_, _06012_ }), .Y(_14303_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36976_ ( .A({ _14274_, _06012_ }), .Y(_14306_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36977_ ( .A({ _14275_, _06012_ }), .Y(_14307_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36978_ ( .A({ _14276_, _06012_ }), .Y(_14308_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36979_ ( .A({ _14277_, _06012_ }), .Y(_14309_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36980_ ( .A({ _14278_, _06012_ }), .Y(_14310_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36981_ ( .A({ _14279_, _06012_ }), .Y(_14311_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36982_ ( .A({ _14280_, _06012_ }), .Y(_14312_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36983_ ( .A({ _14250_, _06012_ }), .Y(_14282_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36984_ ( .A({ _14251_, _06012_ }), .Y(_14283_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36985_ ( .A({ _14252_, _06012_ }), .Y(_14284_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36986_ ( .A({ _14253_, _06012_ }), .Y(_14285_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36987_ ( .A({ _14254_, _06012_ }), .Y(_14286_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36988_ ( .A({ _14255_, _06012_ }), .Y(_14287_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36989_ ( .A({ _14256_, _06012_ }), .Y(_14288_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36990_ ( .A({ _14257_, _06012_ }), .Y(_14289_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36991_ ( .A({ _14258_, _06012_ }), .Y(_14290_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36992_ ( .A({ _14259_, _06012_ }), .Y(_14291_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36993_ ( .A({ _14261_, _06012_ }), .Y(_14293_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36994_ ( .A({ _14262_, _06012_ }), .Y(_14294_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36995_ ( .A({ _14263_, _06012_ }), .Y(_14295_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36996_ ( .A({ _14264_, _06012_ }), .Y(_14296_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36997_ ( .A({ _14265_, _06012_ }), .Y(_14297_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36998_ ( .A({ _14266_, _06012_ }), .Y(_14298_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36999_ ( .A({ _14267_, _06012_ }), .Y(_14299_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37000_ ( .A({ _14268_, _06012_ }), .Y(_14300_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37001_ ( .A({ _14269_, _06012_ }), .Y(_14301_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37002_ ( .A({ _14270_, _06012_ }), .Y(_14302_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37003_ ( .A({ _14272_, _06012_ }), .Y(_14304_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37004_ ( .A({ _14273_, _06012_ }), .Y(_14305_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37005_ ( .A({ max_pool_serial_9_row_count[0], _06012_ }), .Y(_14153_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37006_ ( .A({ max_pool_serial_9_row_count[1], _06012_ }), .Y(_14164_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37007_ ( .A({ max_pool_serial_9_row_count[2], _06012_ }), .Y(_14175_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37008_ ( .A({ max_pool_serial_9_row_count[3], _06012_ }), .Y(_14178_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37009_ ( .A({ max_pool_serial_9_row_count[4], _06012_ }), .Y(_14179_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37010_ ( .A({ max_pool_serial_9_row_count[5], _06012_ }), .Y(_14180_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37011_ ( .A({ max_pool_serial_9_row_count[6], _06012_ }), .Y(_14181_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37012_ ( .A({ max_pool_serial_9_row_count[7], _06012_ }), .Y(_14182_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37013_ ( .A({ max_pool_serial_9_row_count[8], _06012_ }), .Y(_14183_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37014_ ( .A({ max_pool_serial_9_row_count[9], _06012_ }), .Y(_14184_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37015_ ( .A({ max_pool_serial_9_row_count[10], _06012_ }), .Y(_14154_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37016_ ( .A({ max_pool_serial_9_row_count[11], _06012_ }), .Y(_14155_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37017_ ( .A({ max_pool_serial_9_row_count[12], _06012_ }), .Y(_14156_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37018_ ( .A({ max_pool_serial_9_row_count[13], _06012_ }), .Y(_14157_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37019_ ( .A({ max_pool_serial_9_row_count[14], _06012_ }), .Y(_14158_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37020_ ( .A({ max_pool_serial_9_row_count[15], _06012_ }), .Y(_14159_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37021_ ( .A({ max_pool_serial_9_row_count[16], _06012_ }), .Y(_14160_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37022_ ( .A({ max_pool_serial_9_row_count[17], _06012_ }), .Y(_14161_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37023_ ( .A({ max_pool_serial_9_row_count[18], _06012_ }), .Y(_14162_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37024_ ( .A({ max_pool_serial_9_row_count[19], _06012_ }), .Y(_14163_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37025_ ( .A({ max_pool_serial_9_row_count[20], _06012_ }), .Y(_14165_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37026_ ( .A({ max_pool_serial_9_row_count[21], _06012_ }), .Y(_14166_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37027_ ( .A({ max_pool_serial_9_row_count[22], _06012_ }), .Y(_14167_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37028_ ( .A({ max_pool_serial_9_row_count[23], _06012_ }), .Y(_14168_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37029_ ( .A({ max_pool_serial_9_row_count[24], _06012_ }), .Y(_14169_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37030_ ( .A({ max_pool_serial_9_row_count[25], _06012_ }), .Y(_14170_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37031_ ( .A({ max_pool_serial_9_row_count[26], _06012_ }), .Y(_14171_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37032_ ( .A({ max_pool_serial_9_row_count[27], _06012_ }), .Y(_14172_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37033_ ( .A({ max_pool_serial_9_row_count[28], _06012_ }), .Y(_14173_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37034_ ( .A({ max_pool_serial_9_row_count[29], _06012_ }), .Y(_14174_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37035_ ( .A({ max_pool_serial_9_row_count[30], _06012_ }), .Y(_14176_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37036_ ( .A({ max_pool_serial_9_row_count[31], _06012_ }), .Y(_14177_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37037_ ( .A({ _14185_, _06012_ }), .Y(_14217_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37038_ ( .A({ _14196_, _06012_ }), .Y(_14228_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37039_ ( .A({ _14207_, _06012_ }), .Y(_14239_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37040_ ( .A({ _14210_, _06012_ }), .Y(_14242_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37041_ ( .A({ _14211_, _06012_ }), .Y(_14243_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37042_ ( .A({ _14212_, _06012_ }), .Y(_14244_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37043_ ( .A({ _14213_, _06012_ }), .Y(_14245_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37044_ ( .A({ _14214_, _06012_ }), .Y(_14246_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37045_ ( .A({ _14215_, _06012_ }), .Y(_14247_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37046_ ( .A({ _14216_, _06012_ }), .Y(_14248_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37047_ ( .A({ _14186_, _06012_ }), .Y(_14218_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37048_ ( .A({ _14187_, _06012_ }), .Y(_14219_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37049_ ( .A({ _14188_, _06012_ }), .Y(_14220_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37050_ ( .A({ _14189_, _06012_ }), .Y(_14221_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37051_ ( .A({ _14190_, _06012_ }), .Y(_14222_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37052_ ( .A({ _14191_, _06012_ }), .Y(_14223_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37053_ ( .A({ _14192_, _06012_ }), .Y(_14224_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37054_ ( .A({ _14193_, _06012_ }), .Y(_14225_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37055_ ( .A({ _14194_, _06012_ }), .Y(_14226_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37056_ ( .A({ _14195_, _06012_ }), .Y(_14227_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37057_ ( .A({ _14197_, _06012_ }), .Y(_14229_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37058_ ( .A({ _14198_, _06012_ }), .Y(_14230_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37059_ ( .A({ _14199_, _06012_ }), .Y(_14231_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37060_ ( .A({ _14200_, _06012_ }), .Y(_14232_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37061_ ( .A({ _14201_, _06012_ }), .Y(_14233_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37062_ ( .A({ _14202_, _06012_ }), .Y(_14234_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37063_ ( .A({ _14203_, _06012_ }), .Y(_14235_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37064_ ( .A({ _14204_, _06012_ }), .Y(_14236_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37065_ ( .A({ _14205_, _06012_ }), .Y(_14237_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37066_ ( .A({ _14206_, _06012_ }), .Y(_14238_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37067_ ( .A({ _14208_, _06012_ }), .Y(_14240_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37068_ ( .A({ _14209_, _06012_ }), .Y(_14241_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37069_ ( .A({ _18816_, _05909_ }), .Y(_18848_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37070_ ( .A({ _18827_, _05909_ }), .Y(_18859_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37071_ ( .A({ _18838_, _05909_ }), .Y(_18870_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37072_ ( .A({ _18841_, _05909_ }), .Y(_18873_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37073_ ( .A({ _18842_, _05909_ }), .Y(_18874_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37074_ ( .A({ _18843_, _05909_ }), .Y(_18875_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37075_ ( .A({ _18844_, _05909_ }), .Y(_18876_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37076_ ( .A({ _18845_, _05909_ }), .Y(_18877_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37077_ ( .A({ _18846_, _05909_ }), .Y(_18878_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37078_ ( .A({ _18847_, _05909_ }), .Y(_18879_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37079_ ( .A({ _18817_, _05909_ }), .Y(_18849_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37080_ ( .A({ _18818_, _05909_ }), .Y(_18850_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37081_ ( .A({ _18819_, _05909_ }), .Y(_18851_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37082_ ( .A({ _18820_, _05909_ }), .Y(_18852_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37083_ ( .A({ _18821_, _05909_ }), .Y(_18853_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37084_ ( .A({ _18822_, _05909_ }), .Y(_18854_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37085_ ( .A({ _18823_, _05909_ }), .Y(_18855_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37086_ ( .A({ _18824_, _05909_ }), .Y(_18856_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37087_ ( .A({ _18825_, _05909_ }), .Y(_18857_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37088_ ( .A({ _18826_, _05909_ }), .Y(_18858_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37089_ ( .A({ _18828_, _05909_ }), .Y(_18860_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37090_ ( .A({ _18829_, _05909_ }), .Y(_18861_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37091_ ( .A({ _18830_, _05909_ }), .Y(_18862_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37092_ ( .A({ _18831_, _05909_ }), .Y(_18863_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37093_ ( .A({ _18832_, _05909_ }), .Y(_18864_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37094_ ( .A({ _18833_, _05909_ }), .Y(_18865_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37095_ ( .A({ _18834_, _05909_ }), .Y(_18866_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37096_ ( .A({ _18835_, _05909_ }), .Y(_18867_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37097_ ( .A({ _18836_, _05909_ }), .Y(_18868_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37098_ ( .A({ _18837_, _05909_ }), .Y(_18869_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37099_ ( .A({ _18839_, _05909_ }), .Y(_18871_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37100_ ( .A({ _18840_, _05909_ }), .Y(_18872_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37101_ ( .A({ max_pool_serial_9_bat_count[0], _06012_ }), .Y(_14121_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37102_ ( .A({ max_pool_serial_9_bat_count[1], _06012_ }), .Y(_14132_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37103_ ( .A({ max_pool_serial_9_bat_count[2], _06012_ }), .Y(_14143_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37104_ ( .A({ max_pool_serial_9_bat_count[3], _06012_ }), .Y(_14146_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37105_ ( .A({ max_pool_serial_9_bat_count[4], _06012_ }), .Y(_14147_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37106_ ( .A({ max_pool_serial_9_bat_count[5], _06012_ }), .Y(_14148_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37107_ ( .A({ max_pool_serial_9_bat_count[6], _06012_ }), .Y(_14149_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37108_ ( .A({ max_pool_serial_9_bat_count[7], _06012_ }), .Y(_14150_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37109_ ( .A({ max_pool_serial_9_bat_count[8], _06012_ }), .Y(_14151_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37110_ ( .A({ max_pool_serial_9_bat_count[9], _06012_ }), .Y(_14152_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37111_ ( .A({ max_pool_serial_9_bat_count[10], _06012_ }), .Y(_14122_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37112_ ( .A({ max_pool_serial_9_bat_count[11], _06012_ }), .Y(_14123_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37113_ ( .A({ max_pool_serial_9_bat_count[12], _06012_ }), .Y(_14124_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37114_ ( .A({ max_pool_serial_9_bat_count[13], _06012_ }), .Y(_14125_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37115_ ( .A({ max_pool_serial_9_bat_count[14], _06012_ }), .Y(_14126_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37116_ ( .A({ max_pool_serial_9_bat_count[15], _06012_ }), .Y(_14127_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37117_ ( .A({ max_pool_serial_9_bat_count[16], _06012_ }), .Y(_14128_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37118_ ( .A({ max_pool_serial_9_bat_count[17], _06012_ }), .Y(_14129_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37119_ ( .A({ max_pool_serial_9_bat_count[18], _06012_ }), .Y(_14130_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37120_ ( .A({ max_pool_serial_9_bat_count[19], _06012_ }), .Y(_14131_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37121_ ( .A({ max_pool_serial_9_bat_count[20], _06012_ }), .Y(_14133_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37122_ ( .A({ max_pool_serial_9_bat_count[21], _06012_ }), .Y(_14134_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37123_ ( .A({ max_pool_serial_9_bat_count[22], _06012_ }), .Y(_14135_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37124_ ( .A({ max_pool_serial_9_bat_count[23], _06012_ }), .Y(_14136_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37125_ ( .A({ max_pool_serial_9_bat_count[24], _06012_ }), .Y(_14137_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37126_ ( .A({ max_pool_serial_9_bat_count[25], _06012_ }), .Y(_14138_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37127_ ( .A({ max_pool_serial_9_bat_count[26], _06012_ }), .Y(_14139_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37128_ ( .A({ max_pool_serial_9_bat_count[27], _06012_ }), .Y(_14140_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37129_ ( .A({ max_pool_serial_9_bat_count[28], _06012_ }), .Y(_14141_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37130_ ( .A({ max_pool_serial_9_bat_count[29], _06012_ }), .Y(_14142_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37131_ ( .A({ max_pool_serial_9_bat_count[30], _06012_ }), .Y(_14144_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37132_ ( .A({ max_pool_serial_9_bat_count[31], _06012_ }), .Y(_14145_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _37133_ ( .A(_sra_data_40[39]), .Y(_05235_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _37134_ ( .A(maxi_rready), .Y(_05106_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _37135_ ( .A(RESETN), .Y(RESETN_inv) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _37136_ ( .A(_05269_), .Y(_05864_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _37137_ ( .A(_05273_), .Y(_05865_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _37138_ ( .A(_05385_), .Y(_05866_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _37139_ ( .A(__variable_wdata_777), .Y(_05230_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _37140_ ( .A(__variable_wdata_778), .Y(_05231_) );
  \$lut  #( .LUT(16'h035f), .WIDTH(4) ) _37141_ ( .A({ _06342_, _05951_, _06352_, _06391_ }), .Y(_11191_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37142_ ( .A({ _06448_, _06443_, _06436_, _06432_ }), .Y(_11192_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _37143_ ( .A({ _06437_, _11192_, _11191_, _06403_ }), .Y(_20213_) );
  \$lut  #( .LUT(16'h001f), .WIDTH(4) ) _37144_ ( .A({ _06403_, _05918_, _06348_, _06339_ }), .Y(_11193_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37145_ ( .A({ _06465_, _06460_, _06455_, _06454_ }), .Y(_11194_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _37146_ ( .A({ _11194_, _06453_, _11193_, _06362_ }), .Y(_20202_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _37147_ ( .A({ _05903_, _05901_, _05928_, _05918_ }), .Y(_11195_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _37148_ ( .A({ _06470_, _06341_, _05892_, _11195_ }), .Y(_11196_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _37149_ ( .A({ _06472_, _06471_, _11196_, _05944_ }), .Y(_21927_) );
  \$lut  #( .LUT(16'he0ff), .WIDTH(4) ) _37150_ ( .A({ _06566_, _06601_, _06580_, _06577_ }), .Y(_21890_) );
  \$lut  #( .LUT(16'h0ac0), .WIDTH(4) ) _37151_ ( .A({ control_matmul_15[0], control_matmul_15[1], _06591_, _06577_ }), .Y(_11197_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _37152_ ( .A({ _06598_, _13178_, _13274_, _06578_ }), .Y(_11198_) );
  \$lut  #( .LUT(16'hff80), .WIDTH(4) ) _37153_ ( .A({ _06601_, _13338_, _06583_, _06567_ }), .Y(_11199_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _37154_ ( .A({ _06644_, _06643_, _11199_, _06577_ }), .Y(_11200_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _37155_ ( .A({ _06647_, _06645_, _11200_, _11198_ }), .Y(_12858_) );
  \$lut  #( .LUT(16'h0df0), .WIDTH(4) ) _37156_ ( .A({ _06567_, _06597_, control_matmul_15[0], _06589_ }), .Y(_11201_) );
  \$lut  #( .LUT(16'h0fee), .WIDTH(4) ) _37157_ ( .A({ _06597_, _06601_, _06582_, _06593_ }), .Y(_11202_) );
  \$lut  #( .LUT(16'h5c13), .WIDTH(4) ) _37158_ ( .A({ _11201_, _11202_, _06567_, _06584_ }), .Y(_11203_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _37159_ ( .A({ _06652_, 1'h1, _06611_ }), .Y(_11204_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _37160_ ( .A({ _06659_, _06654_, _11204_, _11203_ }), .Y(_12853_) );
  \$lut  #( .LUT(16'h35ff), .WIDTH(4) ) _37161_ ( .A({ _06591_, control_matmul_15[1], _06584_, _06567_ }), .Y(_11205_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _37162_ ( .A({ _11205_, _06584_, _06630_, _06579_ }), .Y(_11206_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _37163_ ( .A({ _06664_, _05039_, _12920_, _11896_ }), .Y(_11207_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _37164_ ( .A({ _06671_, _06666_, _11207_, _11206_ }), .Y(_12856_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37165_ ( .A({ _06597_, _06587_, _06582_, _06579_ }), .Y(_11208_) );
  \$lut  #( .LUT(16'h70ff), .WIDTH(4) ) _37166_ ( .A({ _06584_, _11208_, _06591_, control_matmul_15[1] }), .Y(_11209_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _37167_ ( .A({ _11209_, _06599_, _12921_, _11896_ }), .Y(_11210_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _37168_ ( .A({ _06683_, _06678_, _06676_, _11210_ }), .Y(_12857_) );
  \$lut  #( .LUT(8'h81), .WIDTH(3) ) _37169_ ( .A({ _07430_, cparam_conv2d_8_max_col_count[3], conv2d_8_row_count[3] }), .Y(_11211_) );
  \$lut  #( .LUT(16'h2bb2), .WIDTH(4) ) _37170_ ( .A({ _11211_, conv2d_8_row_count[3], cparam_conv2d_8_max_col_count[4], conv2d_8_row_count[4] }), .Y(_11212_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _37171_ ( .A({ _07505_, _07494_, _07486_, _07462_ }), .Y(_11213_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _37172_ ( .A({ _07506_, _07500_, _11213_, _07511_ }), .Y(_05239_) );
  \$lut  #( .LUT(16'hd400), .WIDTH(4) ) _37173_ ( .A({ _07530_, _11294_, _pulse_count_193[8], _21840_ }), .Y(_05237_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _37174_ ( .A({ _07530_, _11296_, _21840_, _reducecustom_count_191[8] }), .Y(_05236_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _37175_ ( .A({ _21777_, _pulse_count_17[0], _pulse_count_17[1], _21788_ }), .Y(_11214_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _37176_ ( .A({ _07546_, _11214_, _pulse_count_17[2], _21799_ }), .Y(_11215_) );
  \$lut  #( .LUT(16'h70ff), .WIDTH(4) ) _37177_ ( .A({ _07549_, _07548_, _11215_, _07547_ }), .Y(_11216_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _37178_ ( .A({ _reduceadd_count_15[31], _21801_, _07625_, _07627_ }), .Y(_11217_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _37179_ ( .A({ _11217_, _07636_, _07624_, _07634_ }), .Y(_11218_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _37180_ ( .A({ _11218_, _21802_, _07589_, _reduceadd_count_15[32] }), .Y(_05233_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _37181_ ( .A({ _21809_, _reduceadd_count_15[9], _21808_, _reduceadd_count_15[8] }), .Y(_11219_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _37182_ ( .A({ _07601_, _11219_, _reduceadd_count_15[7], _21807_ }), .Y(_11220_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _37183_ ( .A({ _07947_, _07946_, _21349_, _07842_ }), .Y(_11221_) );
  \$lut  #( .LUT(16'h07ff), .WIDTH(4) ) _37184_ ( .A({ _07810_, _07843_, _21317_, _07838_ }), .Y(_11222_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _37185_ ( .A({ _07945_, _11222_, _07932_, _07936_ }), .Y(_11223_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _37186_ ( .A({ _07953_, _07950_, _11223_, _11221_ }), .Y(_21189_) );
  \$lut  #( .LUT(16'h001f), .WIDTH(4) ) _37187_ ( .A({ _07934_, _07922_, _07933_, _07797_ }), .Y(_11224_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _37188_ ( .A({ _07986_, _07984_, _11224_, _07833_ }), .Y(_11225_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _37189_ ( .A({ _07993_, _07990_, _07988_, _11225_ }), .Y(_21163_) );
  \$lut  #( .LUT(16'hff07), .WIDTH(4) ) _37190_ ( .A({ _maxi_write_fsm[3], _08205_, _08194_, _maxi_write_fsm[2] }), .Y(_11226_) );
  \$lut  #( .LUT(16'hfeff), .WIDTH(4) ) _37191_ ( .A({ _11226_, _08260_, _04832_, _08257_ }), .Y(_21899_) );
  \$lut  #( .LUT(16'h00bf), .WIDTH(4) ) _37192_ ( .A({ _08298_, _05875_, _08297_, control_max_pool_serial_9[2] }), .Y(_11227_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37193_ ( .A({ _05052_, _08306_, _08305_, _08304_ }), .Y(_11228_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37194_ ( .A({ _08339_, _11228_, _06012_, _05886_ }), .Y(_11229_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _37195_ ( .A({ _11229_, _11227_, _21895_ }), .Y(_21897_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _37196_ ( .A({ _05885_, _05875_, _08303_, _05886_ }), .Y(_11230_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _37197_ ( .A({ _08319_, _08316_, _08314_, _11301_ }), .Y(_14601_) );
  \$lut  #( .LUT(16'hff80), .WIDTH(4) ) _37198_ ( .A({ _08301_, _14946_, _08297_, _05886_ }), .Y(_11231_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _37199_ ( .A({ _14594_, _05052_, _11231_, _05885_ }), .Y(_11232_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37200_ ( .A({ _08327_, _08324_, _08323_, _08322_ }), .Y(_11233_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _37201_ ( .A({ _08328_, _08325_, _11233_, _11232_ }), .Y(_14626_) );
  \$lut  #( .LUT(16'h2fff), .WIDTH(4) ) _37202_ ( .A({ _08183_, _05886_, control_max_pool_serial_9[2], control_max_pool_serial_9[3] }), .Y(_11234_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37203_ ( .A({ _11234_, _05055_, _08305_, _05874_ }), .Y(_11235_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _37204_ ( .A({ _08330_, _11235_, _14708_, _08298_ }), .Y(_11236_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _37205_ ( .A({ _08333_, _08331_, _11236_ }), .Y(_14612_) );
  \$lut  #( .LUT(16'h004f), .WIDTH(4) ) _37206_ ( .A({ _08643_, _08627_, _11305_, _08631_ }), .Y(_11237_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _37207_ ( .A({ _11244_, _11241_, _11237_, _08642_ }), .Y(conv2d_8_dma_pad_mask_0) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _37208_ ( .A({ _04491_, conv2d_8_row_count[23], _04490_, conv2d_8_row_count[22] }), .Y(_11238_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _37209_ ( .A({ _08639_, _11238_, conv2d_8_row_count[16], _04483_ }), .Y(_11239_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _37210_ ( .A({ _04489_, conv2d_8_row_count[21], _04488_, conv2d_8_row_count[20] }), .Y(_11240_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37211_ ( .A({ _08640_, _08632_, _11240_, _11239_ }), .Y(_11241_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _37212_ ( .A({ _04490_, conv2d_8_row_count[22], _08653_, _08649_ }), .Y(_11242_) );
  \$lut  #( .LUT(16'h4dff), .WIDTH(4) ) _37213_ ( .A({ _08632_, conv2d_8_row_count[23], _04491_, _11242_ }), .Y(_11243_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _37214_ ( .A({ _11243_, _08644_, _07432_, _08654_ }), .Y(_11244_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37215_ ( .A({ _08788_, conv2d_8_col_count[9], _04507_ }), .Y(_11245_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _37216_ ( .A({ conv2d_8_col_count[12], _04479_, _04480_, conv2d_8_col_count[13] }), .Y(_11246_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37217_ ( .A({ _08792_, _11246_ }), .Y(_11247_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _37218_ ( .A({ _08791_, _08789_, _08790_, _08779_ }), .Y(_11248_) );
  \$lut  #( .LUT(16'h8f00), .WIDTH(4) ) _37219_ ( .A({ _11247_, _08793_, _11245_, _11248_ }), .Y(_11249_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _37220_ ( .A({ _08818_, _08807_, _08817_ }), .Y(_11250_) );
  \$lut  #( .LUT(16'hff2b), .WIDTH(4) ) _37221_ ( .A({ _08806_, _11250_, _04488_, conv2d_8_col_count[20] }), .Y(_11251_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _37222_ ( .A({ _08819_, _08820_, _11251_ }), .Y(_11252_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _37223_ ( .A({ _08809_, _11252_, _08821_ }), .Y(_11253_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _37224_ ( .A({ conv2d_8_row_count_buf[8], conv2d_8_row_count_buf[9], _04506_, _04507_ }), .Y(_11254_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _37225_ ( .A({ _08837_, _11254_, _08836_ }), .Y(_11255_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _37226_ ( .A({ _11255_, _08838_, _08840_, _08827_ }), .Y(_11256_) );
  \$lut  #( .LUT(16'h0bff), .WIDTH(4) ) _37227_ ( .A({ _08920_, _08923_, _08921_, _08886_ }), .Y(_11257_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _37228_ ( .A({ _11308_, _08904_, _11257_, _08922_ }), .Y(_11258_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _37229_ ( .A({ _04595_, _04499_, _08907_, _08939_ }), .Y(_11259_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _37230_ ( .A({ _04500_, _04596_, _11259_ }), .Y(_11260_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37231_ ( .A({ _08935_, _08933_, _08931_, _08929_ }), .Y(_11261_) );
  \$lut  #( .LUT(16'h00bf), .WIDTH(4) ) _37232_ ( .A({ _08936_, _08927_, _11261_, _04596_ }), .Y(_11262_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _37233_ ( .A({ _04484_, _04612_, _04491_, _04619_ }), .Y(_11263_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37234_ ( .A({ _08967_, _08949_, _08948_, _08946_ }), .Y(_11264_) );
  \$lut  #( .LUT(16'h9000), .WIDTH(4) ) _37235_ ( .A({ _11264_, _11263_, _04611_, _04483_ }), .Y(_11265_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _37236_ ( .A({ _11265_, _08971_, _08968_, _08950_ }), .Y(_11266_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _37237_ ( .A({ _04507_, _04699_, _04506_, _04698_ }), .Y(_11267_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37238_ ( .A({ _09075_, _11267_ }), .Y(_11268_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _37239_ ( .A({ _09076_, _11268_, _09079_, _09066_ }), .Y(_11269_) );
  \$lut  #( .LUT(16'h9000), .WIDTH(4) ) _37240_ ( .A({ _09107_, _09102_, _04675_, _04483_ }), .Y(_11270_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _37241_ ( .A({ _04484_, _04676_, _04488_, _04680_ }), .Y(_11271_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37242_ ( .A({ _09120_, _09096_, _11271_, _11270_ }), .Y(_11272_) );
  \$lut  #( .LUT(8'h81), .WIDTH(3) ) _37243_ ( .A({ _09129_, max_pool_serial_9_col_count[3], cparam_max_pool_serial_9_act_num_col[3] }), .Y(_11273_) );
  \$lut  #( .LUT(16'h4dd4), .WIDTH(4) ) _37244_ ( .A({ _11273_, cparam_max_pool_serial_9_act_num_col[3], cparam_max_pool_serial_9_act_num_col[4], max_pool_serial_9_col_count[4] }), .Y(_11274_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37245_ ( .A({ _07232_, _11274_ }), .Y(_11275_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _37246_ ( .A({ _09142_, _09132_, max_pool_serial_9_row_count_buf[4], cparam_max_pool_serial_9_act_num_col[4] }), .Y(_11276_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37247_ ( .A({ _09135_, _11276_, max_pool_serial_9_row_count_buf[7:6] }), .Y(_11277_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _37248_ ( .A({ _09146_, _09150_, _03604_, cparam_max_pool_serial_9_act_num_col[4] }), .Y(_11278_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37249_ ( .A({ _09149_, _09148_, _09145_, _09144_ }), .Y(_11279_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37250_ ( .A({ _11279_, _09143_, _11278_ }), .Y(_11280_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _37251_ ( .A({ _09163_, _09153_, _03636_, cparam_max_pool_serial_9_act_num_col[4] }), .Y(_11281_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37252_ ( .A({ _09156_, _11281_, _03639_, _03638_ }), .Y(_11282_) );
  \$lut  #( .LUT(8'h81), .WIDTH(3) ) _37253_ ( .A({ _11006_, cparam_conv2d_8_max_col_count[3], conv2d_8_prev_row_count[3] }), .Y(_11283_) );
  \$lut  #( .LUT(16'h2bb2), .WIDTH(4) ) _37254_ ( .A({ _11283_, conv2d_8_prev_row_count[3], cparam_conv2d_8_max_col_count[4], conv2d_8_prev_row_count[4] }), .Y(_11284_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _37255_ ( .A({ _11091_, _11090_, max_pool_serial_9_prev_row_count[2], cparam_max_pool_serial_9_max_col_count[2] }), .Y(_11285_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _37256_ ( .A({ _11089_, _11285_, cparam_max_pool_serial_9_max_col_count[4], max_pool_serial_9_prev_row_count[4] }), .Y(_11286_) );
  \$lut  #( .LUT(16'h007f), .WIDTH(4) ) _37257_ ( .A({ max_pool_serial_9_skip_write_out, _11081_, _11078_, _11286_ }), .Y(_05850_) );
  \$lut  #( .LUT(16'h80fe), .WIDTH(4) ) _37258_ ( .A({ _reducecustom_data_191[31], _11158_, _reducecustom_data_191[8:7] }), .Y(_11287_) );
  \$lut  #( .LUT(8'hc5), .WIDTH(3) ) _37259_ ( .A({ _11317_, _11287_, _reducecustom_data_191[31] }), .Y(_05260_) );
  \$lut  #( .LUT(16'hfff8), .WIDTH(4) ) _37260_ ( .A({ _11197_, _06595_, _13354_, _06586_ }), .Y(_11288_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _37261_ ( .A({ _12810_, _05035_, _11288_, _06567_ }), .Y(_11289_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37262_ ( .A({ _06625_, _06624_, _06623_, _06609_ }), .Y(_11290_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _37263_ ( .A({ _06613_, _11290_, _06607_, _11289_ }), .Y(_12842_) );
  \$lut  #( .LUT(8'h18), .WIDTH(3) ) _37264_ ( .A({ _07525_, _pulse_count_193[4], _21836_ }), .Y(_11291_) );
  \$lut  #( .LUT(16'hd44d), .WIDTH(4) ) _37265_ ( .A({ _21836_, _11291_, _pulse_count_193[5], _21837_ }), .Y(_11292_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _37266_ ( .A({ _21838_, _pulse_count_193[6] }), .Y(_11293_) );
  \$lut  #( .LUT(16'h008f), .WIDTH(4) ) _37267_ ( .A({ _07528_, _07529_, _11292_, _11293_ }), .Y(_11294_) );
  \$lut  #( .LUT(8'h81), .WIDTH(3) ) _37268_ ( .A({ _07538_, _21838_, _reducecustom_count_191[6] }), .Y(_11295_) );
  \$lut  #( .LUT(16'h2bb2), .WIDTH(4) ) _37269_ ( .A({ _11295_, _reducecustom_count_191[6], _21839_, _reducecustom_count_191[7] }), .Y(_11296_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _37270_ ( .A({ _21806_, _pulse_count_17[6], _pulse_count_17[7], _21807_ }), .Y(_11297_) );
  \$lut  #( .LUT(16'hf0bb), .WIDTH(4) ) _37271_ ( .A({ _11216_, _11297_, _pulse_count_17[7], _21807_ }), .Y(_11298_) );
  \$lut  #( .LUT(16'h0c0a), .WIDTH(4) ) _37272_ ( .A({ control_max_pool_serial_9[3:2], _14633_, _14761_ }), .Y(_11299_) );
  \$lut  #( .LUT(16'h07ff), .WIDTH(4) ) _37273_ ( .A({ _08297_, _11230_, _11299_, _05875_ }), .Y(_11300_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _37274_ ( .A({ _11300_, _08305_, _14697_, _08298_ }), .Y(_11301_) );
  \$lut  #( .LUT(16'h222b), .WIDTH(4) ) _37275_ ( .A({ _08622_, _08617_, _04503_, conv2d_8_row_count[5] }), .Y(_11302_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _37276_ ( .A({ _08626_, _11302_, _04504_, conv2d_8_row_count[6] }), .Y(_11303_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37277_ ( .A({ _08624_, conv2d_8_row_count[9], _04507_ }), .Y(_11304_) );
  \$lut  #( .LUT(16'h70ff), .WIDTH(4) ) _37278_ ( .A({ _11304_, _08625_, _11303_, _08623_ }), .Y(_11305_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _37279_ ( .A({ _08926_, _08924_, _04584_, _04488_ }), .Y(_11306_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _37280_ ( .A({ _08916_, _08917_, _11306_, _08915_ }), .Y(_11307_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _37281_ ( .A({ _11262_, _11260_, _11307_, _08905_ }), .Y(_11308_) );
  \$lut  #( .LUT(16'h8001), .WIDTH(4) ) _37282_ ( .A({ _reducecustom_data_191[11:9], _reducecustom_data_191[7] }), .Y(_11309_) );
  \$lut  #( .LUT(16'h8001), .WIDTH(4) ) _37283_ ( .A({ _reducecustom_data_191[16], _reducecustom_data_191[13:12], _reducecustom_data_191[7] }), .Y(_11310_) );
  \$lut  #( .LUT(16'h8001), .WIDTH(4) ) _37284_ ( .A({ _reducecustom_data_191[17], _reducecustom_data_191[15:14], _reducecustom_data_191[7] }), .Y(_11311_) );
  \$lut  #( .LUT(16'h8001), .WIDTH(4) ) _37285_ ( .A({ _reducecustom_data_191[20:18], _reducecustom_data_191[7] }), .Y(_11312_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37286_ ( .A({ _11168_, _11167_, _reducecustom_data_191[24] }), .Y(_11313_) );
  \$lut  #( .LUT(16'hf088), .WIDTH(4) ) _37287_ ( .A({ _reducecustom_data_191[7], _11313_, _11166_, _11165_ }), .Y(_11314_) );
  \$lut  #( .LUT(16'h8001), .WIDTH(4) ) _37288_ ( .A({ _reducecustom_data_191[23:21], _reducecustom_data_191[7] }), .Y(_11315_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37289_ ( .A({ _11312_, _11311_, _11310_, _11309_ }), .Y(_11316_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37290_ ( .A({ _11316_, _11315_, _11314_ }), .Y(_11317_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37291_ ( .A(max_pool_serial_9_act_base_offset_row), .B(max_pool_serial_9_act_base_offset_bat), .Y(max_pool_serial_9_act_base_offset) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37292_ ( .A(max_pool_serial_9_out_base_offset_row), .B(max_pool_serial_9_out_base_offset_bat), .Y(max_pool_serial_9_out_base_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37293_ ( .A(max_pool_serial_9_row_count), .B(1), .Y({ _03570_, _03569_, _03567_, _03566_, _03565_, _03564_, _03563_, _03562_, _03561_, _03560_, _03559_, _03558_, _03556_, _03555_, _03554_, _03553_, _03552_, _03551_, _03550_, _03549_, _03548_, _03547_, _03577_, _03576_, _03575_, _03574_, _03573_, _03572_, _03571_, _03568_, _03557_, _03546_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37294_ ( .A(max_pool_serial_9_col_count), .B(1), .Y({ _03602_, _03601_, _03599_, _03598_, _03597_, _03596_, _03595_, _03594_, _03593_, _03592_, _03591_, _03590_, _03588_, _03587_, _03586_, _03585_, _03584_, _03583_, _03582_, _03581_, _03580_, _03579_, _03609_, _03608_, _03607_, _03606_, _03605_, _03604_, _03603_, _03600_, _03589_, _03578_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37295_ ( .A(max_pool_serial_9_row_count_buf), .B(1), .Y({ _03634_, _03633_, _03631_, _03630_, _03629_, _03628_, _03627_, _03626_, _03625_, _03624_, _03623_, _03622_, _03620_, _03619_, _03618_, _03617_, _03616_, _03615_, _03614_, _03613_, _03612_, _03611_, _03641_, _03640_, _03639_, _03638_, _03637_, _03636_, _03635_, _03632_, _03621_, _03610_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37296_ ( .A(_stream_max_pool_serial_9_source_1_source_offset_buf), .B(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_0), .Y(_22041_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37297_ ( .A(_22041_), .B(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_1), .Y(_22042_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37298_ ( .A(_22042_), .B(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_2), .Y(_22043_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37299_ ( .A(_22043_), .B(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_3), .Y(_stream_max_pool_serial_9_source_1_source_pat_all_offset) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37300_ ( .A(matmul_15_act_base_offset_row), .B(matmul_15_act_base_offset_bat), .Y(matmul_15_act_base_offset) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37301_ ( .A(matmul_15_out_base_offset_val), .B(matmul_15_out_base_offset_col), .Y(_22044_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37302_ ( .A(_22044_), .B(matmul_15_out_base_offset_row), .Y(_22045_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37303_ ( .A(_22045_), .B(matmul_15_out_base_offset_bat), .Y(_22046_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37304_ ( .A(_22046_), .B(matmul_15_out_base_offset_och), .Y(matmul_15_out_base_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37305_ ( .A(matmul_15_arg_objaddr_0), .B(matmul_15_act_base_offset), .Y(_22047_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37306_ ( .A(_stream_matmul_15_source_6_source_offset_buf), .B(_source_stream_matmul_15_source_6_pat_cur_offset_0), .Y(_22048_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37307_ ( .A(_22048_), .B(_source_stream_matmul_15_source_6_pat_cur_offset_1), .Y(_22049_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37308_ ( .A(_22049_), .B(_source_stream_matmul_15_source_6_pat_cur_offset_2), .Y(_22050_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37309_ ( .A(_22050_), .B(_source_stream_matmul_15_source_6_pat_cur_offset_3), .Y(_stream_matmul_15_source_6_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37310_ ( .A(_stream_matmul_15_source_8_source_offset_buf), .B(_source_stream_matmul_15_source_8_pat_cur_offset_0), .Y(_22051_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37311_ ( .A(_22051_), .B(_source_stream_matmul_15_source_8_pat_cur_offset_1), .Y(_22052_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37312_ ( .A(_22052_), .B(_source_stream_matmul_15_source_8_pat_cur_offset_2), .Y(_22053_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37313_ ( .A(_22053_), .B(_source_stream_matmul_15_source_8_pat_cur_offset_3), .Y(_stream_matmul_15_source_8_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37314_ ( .A(_stream_matmul_15_source_19_source_offset_buf), .B(_source_stream_matmul_15_source_19_pat_cur_offset_0), .Y(_22054_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37315_ ( .A(_22054_), .B(_source_stream_matmul_15_source_19_pat_cur_offset_1), .Y(_22055_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37316_ ( .A(_22055_), .B(_source_stream_matmul_15_source_19_pat_cur_offset_2), .Y(_22056_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37317_ ( .A(_22056_), .B(_source_stream_matmul_15_source_19_pat_cur_offset_3), .Y(_stream_matmul_15_source_19_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37318_ ( .A(_stream_matmul_15_source_20_source_offset_buf), .B(_source_stream_matmul_15_source_20_pat_cur_offset_0), .Y(_22057_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37319_ ( .A(_22057_), .B(_source_stream_matmul_15_source_20_pat_cur_offset_1), .Y(_22058_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37320_ ( .A(_22058_), .B(_source_stream_matmul_15_source_20_pat_cur_offset_2), .Y(_22059_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37321_ ( .A(_22059_), .B(_source_stream_matmul_15_source_20_pat_cur_offset_3), .Y(_stream_matmul_15_source_20_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37322_ ( .A(conv2d_8_arg_objaddr_1), .B(conv2d_8_filter_base_offset), .Y(_22060_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _37323_ ( .A({ 24'h000000, cparam_conv2d_8_filter_base_step[10:2] }), .B({ 1'h0, _26478_ }), .Y(_22061_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _37324_ ( .A({ 27'h0000000, cparam_conv2d_8_act_read_size[7:2] }), .B({ 1'h0, _26479_ }), .Y(_22062_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37325_ ( .A(conv2d_8_out_laddr_offset), .B(conv2d_8_out_page_dma_offset), .Y(_22063_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37326_ ( .A(conv2d_8_objaddr), .B(conv2d_8_out_base_offset), .Y(_22064_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _37327_ ( .A({ 3'h0, conv2d_8_next_out_write_size[31:2] }), .B({ 1'h0, _26480_ }), .Y(_22065_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37328_ ( .A(max_pool_serial_9_arg_objaddr_0), .B(max_pool_serial_9_act_base_offset), .Y(_22066_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(9), .Y_WIDTH(32) ) _37329_ ( .A(max_pool_serial_9_act_page_dma_offset), .B(cparam_max_pool_serial_9_act_offset_values_1[8:0]), .Y(_22068_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37330_ ( .A(max_pool_serial_9_act_base_offset), .B(cparam_max_pool_serial_9_act_offset_values_1), .Y(_22069_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37331_ ( .A(max_pool_serial_9_arg_objaddr_0), .B(_22069_), .Y(_22070_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _37332_ ( .A({ 26'h0000000, cparam_max_pool_serial_9_act_offset_values_1[8:2] }), .B({ 1'h0, _26481_ }), .Y(_22067_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37333_ ( .A(max_pool_serial_9_objaddr), .B(max_pool_serial_9_out_base_offset), .Y(_22071_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _37334_ ( .A({ 27'h0000000, cparam_max_pool_serial_9_out_row_step[7:2] }), .B({ 1'h0, _26482_ }), .Y(_22072_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37335_ ( .A(matmul_15_arg_objaddr_1), .B(matmul_15_filter_base_offset), .Y(_22073_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37336_ ( .A(matmul_15_out_laddr_offset), .B(matmul_15_out_page_dma_offset), .Y(_22074_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37337_ ( .A(matmul_15_objaddr), .B(matmul_15_out_base_offset), .Y(_22075_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _37338_ ( .A({ 3'h0, matmul_15_next_out_write_size[31:2] }), .B({ 1'h0, _26483_ }), .Y(_22076_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37339_ ( .A(ram_w8_l4096_id0_0_1_addr), .B(_maxi_read_local_stride), .Y(_22077_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37340_ ( .A(ram_w8_l4096_id0_1_1_addr), .B(_maxi_read_local_stride), .Y(_22078_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37341_ ( .A(ram_w8_l4096_id0_2_1_addr), .B(_maxi_read_local_stride), .Y(_22079_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37342_ ( .A(ram_w8_l4096_id0_3_1_addr), .B(_maxi_read_local_stride), .Y(_22080_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37343_ ( .A(ram_w8_l2048_id0_0_1_addr), .B(_maxi_read_local_stride), .Y(_22081_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37344_ ( .A(ram_w8_l2048_id0_0_1_addr), .B(_maxi_write_local_stride), .Y(_22082_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37345_ ( .A(ram_w8_l2048_id0_1_1_addr), .B(_maxi_read_local_stride), .Y(_22083_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37346_ ( .A(ram_w8_l2048_id0_1_1_addr), .B(_maxi_write_local_stride), .Y(_22084_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37347_ ( .A(ram_w8_l2048_id0_2_1_addr), .B(_maxi_read_local_stride), .Y(_22085_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37348_ ( .A(ram_w8_l2048_id0_2_1_addr), .B(_maxi_write_local_stride), .Y(_22086_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37349_ ( .A(ram_w8_l2048_id0_3_1_addr), .B(_maxi_read_local_stride), .Y(_22087_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37350_ ( .A(ram_w8_l2048_id0_3_1_addr), .B(_maxi_write_local_stride), .Y(_22088_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37351_ ( .A(_tmp_62), .B(1), .Y(_22089_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37352_ ( .A(ram_w8_l2048_id1_0_1_addr), .B(_maxi_read_local_stride), .Y(_22090_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37353_ ( .A(ram_w8_l2048_id1_0_1_addr), .B(_maxi_write_local_stride), .Y(_22091_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37354_ ( .A(_tmp_93), .B(1), .Y(_22092_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37355_ ( .A(ram_w8_l2048_id1_1_1_addr), .B(_maxi_read_local_stride), .Y(_22093_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37356_ ( .A(ram_w8_l2048_id1_1_1_addr), .B(_maxi_write_local_stride), .Y(_22094_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37357_ ( .A(_tmp_124), .B(1), .Y(_22095_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37358_ ( .A(ram_w8_l2048_id1_2_1_addr), .B(_maxi_read_local_stride), .Y(_22096_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37359_ ( .A(ram_w8_l2048_id1_2_1_addr), .B(_maxi_write_local_stride), .Y(_22097_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37360_ ( .A(_tmp_155), .B(1), .Y(_22098_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37361_ ( .A(ram_w8_l2048_id1_3_1_addr), .B(_maxi_read_local_stride), .Y(_22099_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37362_ ( .A(ram_w8_l2048_id1_3_1_addr), .B(_maxi_write_local_stride), .Y(_22100_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37363_ ( .A(ram_w8_l2048_id2_0_1_addr), .B(_maxi_read_local_stride), .Y(_22101_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37364_ ( .A(ram_w8_l2048_id2_1_1_addr), .B(_maxi_read_local_stride), .Y(_22102_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37365_ ( .A(ram_w8_l2048_id2_2_1_addr), .B(_maxi_read_local_stride), .Y(_22103_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37366_ ( .A(ram_w8_l2048_id2_3_1_addr), .B(_maxi_read_local_stride), .Y(_22104_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37367_ ( .A(_tmp_173), .B(1), .Y(_22105_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37368_ ( .A(_tmp_186), .B(1), .Y(_22106_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37369_ ( .A(_tmp_199), .B(1), .Y(_22107_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37370_ ( .A(_tmp_212), .B(1), .Y(_22108_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37371_ ( .A(_tmp_230), .B(1), .Y(_22109_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37372_ ( .A(_tmp_243), .B(1), .Y(_22110_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37373_ ( .A(_tmp_256), .B(1), .Y(_22111_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37374_ ( .A(_tmp_269), .B(1), .Y(_22112_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37375_ ( .A(_tmp_287), .B(1), .Y(_22113_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37376_ ( .A(_tmp_300), .B(1), .Y(_22114_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37377_ ( .A(_tmp_313), .B(1), .Y(_22115_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37378_ ( .A(_tmp_326), .B(1), .Y(_22116_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37379_ ( .A(ram_w8_l2048_id19_0_1_addr), .B(_maxi_write_local_stride), .Y(_22117_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37380_ ( .A(ram_w8_l2048_id19_1_1_addr), .B(_maxi_write_local_stride), .Y(_22118_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37381_ ( .A(ram_w8_l2048_id19_2_1_addr), .B(_maxi_write_local_stride), .Y(_22119_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37382_ ( .A(ram_w8_l2048_id19_3_1_addr), .B(_maxi_write_local_stride), .Y(_22120_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(7), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37383_ ( .A(ram_w32_l128_id0_1_addr), .B(_maxi_read_local_stride), .Y(_22121_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37384_ ( .A(_reduceadd_data_15), .B(__variable_wdata_0), .Y(_22122_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _37385_ ( .A(_reduceadd_count_15), .B(1), .Y(_22123_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _37386_ ( .A(_pulse_count_17), .B(1), .Y(_22124_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37387_ ( .A(__delay_data_730), .B(_cond_data_11), .Y(_22125_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37388_ ( .A(__variable_wdata_22), .B(__variable_wdata_23), .Y(_22126_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37389_ ( .A(_22126_), .B(__variable_wdata_24), .Y(_22127_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37390_ ( .A(__variable_wdata_25), .B(__variable_wdata_26), .Y(_22128_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37391_ ( .A(_22128_), .B(__variable_wdata_27), .Y(_22129_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37392_ ( .A(__variable_wdata_28), .B(__variable_wdata_29), .Y(_22130_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37393_ ( .A(_22130_), .B(__variable_wdata_30), .Y(_22131_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37394_ ( .A(__plusn_data_32), .B(__plusn_data_33), .Y(_22132_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37395_ ( .A(_22132_), .B(__plusn_data_34), .Y(_22133_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37396_ ( .A(_reducecustom_count_191), .B(1), .Y(_22134_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37397_ ( .A(_pulse_count_193), .B(1), .Y(_22135_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(8) ) _37398_ ( .A(_cond_data_229), .B(__delay_data_916), .Y(_22136_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(8) ) _37399_ ( .A(_cond_data_236), .B(__delay_data_1229), .Y(_22137_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(4), .Y_WIDTH(8) ) _37400_ ( .A(_cond_data_243), .B(__delay_data_1300), .Y(_22138_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37401_ ( .A(__substreamoutput_data_861), .B(__delay_data_1299), .Y(_22139_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37402_ ( .A(_source_stream_conv2d_8_source_6_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_6_pat_stride_buf_0), .Y(_22140_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37403_ ( .A(_source_stream_conv2d_8_source_6_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_6_pat_stride_buf_1), .Y(_22141_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37404_ ( .A(_source_stream_conv2d_8_source_6_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_6_pat_stride_buf_2), .Y(_22142_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37405_ ( .A(_source_stream_conv2d_8_source_6_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_6_pat_stride_buf_3), .Y(_22143_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37406_ ( .A(_source_stream_conv2d_8_source_8_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_8_pat_stride_buf_0), .Y(_22144_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37407_ ( .A(_source_stream_conv2d_8_source_8_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_8_pat_stride_buf_1), .Y(_22145_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37408_ ( .A(_source_stream_conv2d_8_source_8_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_8_pat_stride_buf_2), .Y(_22146_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37409_ ( .A(_source_stream_conv2d_8_source_8_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_8_pat_stride_buf_3), .Y(_22147_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37410_ ( .A(conv2d_8_stream_act_local_0), .B(conv2d_8_act_page_comp_offset_buf_0), .Y(_22148_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37411_ ( .A(_source_stream_conv2d_8_source_19_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_19_pat_stride_buf_0), .Y(_22149_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37412_ ( .A(_source_stream_conv2d_8_source_19_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_19_pat_stride_buf_1), .Y(_22150_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37413_ ( .A(_source_stream_conv2d_8_source_19_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_19_pat_stride_buf_2), .Y(_22151_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37414_ ( .A(_source_stream_conv2d_8_source_19_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_19_pat_stride_buf_3), .Y(_22152_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37415_ ( .A(conv2d_8_stream_act_local_1), .B(conv2d_8_act_page_comp_offset_buf_0), .Y(_22153_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37416_ ( .A(_source_stream_conv2d_8_source_20_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_20_pat_stride_buf_0), .Y(_22154_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37417_ ( .A(_source_stream_conv2d_8_source_20_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_20_pat_stride_buf_1), .Y(_22155_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37418_ ( .A(_source_stream_conv2d_8_source_20_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_20_pat_stride_buf_2), .Y(_22156_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37419_ ( .A(_source_stream_conv2d_8_source_20_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_20_pat_stride_buf_3), .Y(_22157_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37420_ ( .A(conv2d_8_stream_act_local_2), .B(conv2d_8_act_page_comp_offset_buf_0), .Y(_22158_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37421_ ( .A(_source_stream_conv2d_8_source_21_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_21_pat_stride_buf_0), .Y(_22159_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37422_ ( .A(_source_stream_conv2d_8_source_21_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_21_pat_stride_buf_1), .Y(_22160_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37423_ ( .A(_source_stream_conv2d_8_source_21_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_21_pat_stride_buf_2), .Y(_22161_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37424_ ( .A(_source_stream_conv2d_8_source_21_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_21_pat_stride_buf_3), .Y(_22162_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37425_ ( .A(conv2d_8_stream_act_local_3), .B(conv2d_8_act_page_comp_offset_buf_1), .Y(_22163_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37426_ ( .A(_source_stream_conv2d_8_source_22_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_22_pat_stride_buf_0), .Y(_22164_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37427_ ( .A(_source_stream_conv2d_8_source_22_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_22_pat_stride_buf_1), .Y(_22165_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37428_ ( .A(_source_stream_conv2d_8_source_22_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_22_pat_stride_buf_2), .Y(_22166_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37429_ ( .A(_source_stream_conv2d_8_source_22_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_22_pat_stride_buf_3), .Y(_22167_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37430_ ( .A(conv2d_8_stream_act_local_4), .B(conv2d_8_act_page_comp_offset_buf_1), .Y(_22168_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37431_ ( .A(_source_stream_conv2d_8_source_23_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_23_pat_stride_buf_0), .Y(_22169_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37432_ ( .A(_source_stream_conv2d_8_source_23_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_23_pat_stride_buf_1), .Y(_22170_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37433_ ( .A(_source_stream_conv2d_8_source_23_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_23_pat_stride_buf_2), .Y(_22171_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37434_ ( .A(_source_stream_conv2d_8_source_23_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_23_pat_stride_buf_3), .Y(_22172_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37435_ ( .A(conv2d_8_stream_act_local_5), .B(conv2d_8_act_page_comp_offset_buf_1), .Y(_22173_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37436_ ( .A(_source_stream_conv2d_8_source_24_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_24_pat_stride_buf_0), .Y(_22174_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37437_ ( .A(_source_stream_conv2d_8_source_24_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_24_pat_stride_buf_1), .Y(_22175_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37438_ ( .A(_source_stream_conv2d_8_source_24_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_24_pat_stride_buf_2), .Y(_22176_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37439_ ( .A(_source_stream_conv2d_8_source_24_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_24_pat_stride_buf_3), .Y(_22177_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37440_ ( .A(conv2d_8_stream_act_local_6), .B(conv2d_8_act_page_comp_offset_buf_2), .Y(_22178_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37441_ ( .A(_source_stream_conv2d_8_source_25_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_25_pat_stride_buf_0), .Y(_22179_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37442_ ( .A(_source_stream_conv2d_8_source_25_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_25_pat_stride_buf_1), .Y(_22180_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37443_ ( .A(_source_stream_conv2d_8_source_25_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_25_pat_stride_buf_2), .Y(_22181_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37444_ ( .A(_source_stream_conv2d_8_source_25_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_25_pat_stride_buf_3), .Y(_22182_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37445_ ( .A(conv2d_8_stream_act_local_7), .B(conv2d_8_act_page_comp_offset_buf_2), .Y(_22183_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37446_ ( .A(_source_stream_conv2d_8_source_26_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_26_pat_stride_buf_0), .Y(_22184_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37447_ ( .A(_source_stream_conv2d_8_source_26_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_26_pat_stride_buf_1), .Y(_22185_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37448_ ( .A(_source_stream_conv2d_8_source_26_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_26_pat_stride_buf_2), .Y(_22186_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37449_ ( .A(_source_stream_conv2d_8_source_26_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_26_pat_stride_buf_3), .Y(_22187_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37450_ ( .A(conv2d_8_stream_act_local_8), .B(conv2d_8_act_page_comp_offset_buf_2), .Y(_22188_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37451_ ( .A(_source_stream_conv2d_8_source_27_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_27_pat_stride_buf_0), .Y(_22189_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37452_ ( .A(_source_stream_conv2d_8_source_27_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_27_pat_stride_buf_1), .Y(_22190_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37453_ ( .A(_source_stream_conv2d_8_source_27_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_27_pat_stride_buf_2), .Y(_22191_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37454_ ( .A(_source_stream_conv2d_8_source_27_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_27_pat_stride_buf_3), .Y(_22192_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37455_ ( .A(_source_stream_conv2d_8_source_28_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_28_pat_stride_buf_0), .Y(_22193_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37456_ ( .A(_source_stream_conv2d_8_source_28_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_28_pat_stride_buf_1), .Y(_22194_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37457_ ( .A(_source_stream_conv2d_8_source_28_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_28_pat_stride_buf_2), .Y(_22195_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37458_ ( .A(_source_stream_conv2d_8_source_28_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_28_pat_stride_buf_3), .Y(_22196_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37459_ ( .A(_source_stream_conv2d_8_source_29_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_29_pat_stride_buf_0), .Y(_22197_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37460_ ( .A(_source_stream_conv2d_8_source_29_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_29_pat_stride_buf_1), .Y(_22198_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37461_ ( .A(_source_stream_conv2d_8_source_29_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_29_pat_stride_buf_2), .Y(_22199_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37462_ ( .A(_source_stream_conv2d_8_source_29_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_29_pat_stride_buf_3), .Y(_22200_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37463_ ( .A(_source_stream_conv2d_8_source_30_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_30_pat_stride_buf_0), .Y(_22201_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37464_ ( .A(_source_stream_conv2d_8_source_30_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_30_pat_stride_buf_1), .Y(_22202_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37465_ ( .A(_source_stream_conv2d_8_source_30_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_30_pat_stride_buf_2), .Y(_22203_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37466_ ( .A(_source_stream_conv2d_8_source_30_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_30_pat_stride_buf_3), .Y(_22204_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37467_ ( .A(_source_stream_conv2d_8_source_31_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_31_pat_stride_buf_0), .Y(_22205_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37468_ ( .A(_source_stream_conv2d_8_source_31_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_31_pat_stride_buf_1), .Y(_22206_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37469_ ( .A(_source_stream_conv2d_8_source_31_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_31_pat_stride_buf_2), .Y(_22207_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37470_ ( .A(_source_stream_conv2d_8_source_31_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_31_pat_stride_buf_3), .Y(_22208_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37471_ ( .A(_source_stream_conv2d_8_source_32_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_32_pat_stride_buf_0), .Y(_22209_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37472_ ( .A(_source_stream_conv2d_8_source_32_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_32_pat_stride_buf_1), .Y(_22210_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37473_ ( .A(_source_stream_conv2d_8_source_32_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_32_pat_stride_buf_2), .Y(_22211_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37474_ ( .A(_source_stream_conv2d_8_source_32_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_32_pat_stride_buf_3), .Y(_22212_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37475_ ( .A(_source_stream_conv2d_8_source_33_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_33_pat_stride_buf_0), .Y(_22213_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37476_ ( .A(_source_stream_conv2d_8_source_33_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_33_pat_stride_buf_1), .Y(_22214_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37477_ ( .A(_source_stream_conv2d_8_source_33_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_33_pat_stride_buf_2), .Y(_22215_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37478_ ( .A(_source_stream_conv2d_8_source_33_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_33_pat_stride_buf_3), .Y(_22216_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37479_ ( .A(_source_stream_conv2d_8_source_34_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_34_pat_stride_buf_0), .Y(_22217_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37480_ ( .A(_source_stream_conv2d_8_source_34_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_34_pat_stride_buf_1), .Y(_22218_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37481_ ( .A(_source_stream_conv2d_8_source_34_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_34_pat_stride_buf_2), .Y(_22219_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37482_ ( .A(_source_stream_conv2d_8_source_34_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_34_pat_stride_buf_3), .Y(_22220_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37483_ ( .A(_source_stream_conv2d_8_source_35_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_35_pat_stride_buf_0), .Y(_22221_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37484_ ( .A(_source_stream_conv2d_8_source_35_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_35_pat_stride_buf_1), .Y(_22222_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37485_ ( .A(_source_stream_conv2d_8_source_35_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_35_pat_stride_buf_2), .Y(_22223_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37486_ ( .A(_source_stream_conv2d_8_source_35_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_35_pat_stride_buf_3), .Y(_22224_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37487_ ( .A(_source_stream_conv2d_8_source_36_pat_cur_offset_0), .B(_source_stream_conv2d_8_source_36_pat_stride_buf_0), .Y(_22225_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37488_ ( .A(_source_stream_conv2d_8_source_36_pat_cur_offset_1), .B(_source_stream_conv2d_8_source_36_pat_stride_buf_1), .Y(_22226_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37489_ ( .A(_source_stream_conv2d_8_source_36_pat_cur_offset_2), .B(_source_stream_conv2d_8_source_36_pat_stride_buf_2), .Y(_22227_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37490_ ( .A(_source_stream_conv2d_8_source_36_pat_cur_offset_3), .B(_source_stream_conv2d_8_source_36_pat_stride_buf_3), .Y(_22228_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37491_ ( .A(conv2d_8_stream_out_local_col), .B(conv2d_8_out_page_comp_offset_buf), .Y(_22229_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37492_ ( .A(_stream_conv2d_8_sink_37_sink_waddr), .B(_stream_conv2d_8_sink_37_sink_stride_buf), .Y(_22230_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37493_ ( .A(_counter_data_762), .B(1), .Y(_22231_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37494_ ( .A(_counter_count_762), .B(1), .Y(_22232_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37495_ ( .A(max_pool_serial_9_stream_act_local), .B(max_pool_serial_9_act_page_comp_offset_buf), .Y(_22233_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37496_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_0), .B(_source_stream_max_pool_serial_9_source_1_pat_stride_buf_0), .Y(_22234_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37497_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_1), .B(_source_stream_max_pool_serial_9_source_1_pat_stride_buf_1), .Y(_22235_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37498_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_2), .B(_source_stream_max_pool_serial_9_source_1_pat_stride_buf_2), .Y(_22236_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37499_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_3), .B(_source_stream_max_pool_serial_9_source_1_pat_stride_buf_3), .Y(_22237_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37500_ ( .A(max_pool_serial_9_stream_out_local), .B(max_pool_serial_9_out_page_comp_offset_buf), .Y(_22238_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37501_ ( .A(_stream_max_pool_serial_9_sink_3_sink_waddr), .B(_stream_max_pool_serial_9_sink_3_sink_stride_buf), .Y(_22239_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(8) ) _37502_ ( .A(_cond_data_811), .B(__delay_data_1382), .Y(_22240_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(8) ) _37503_ ( .A(_cond_data_818), .B(__delay_data_1389), .Y(_22241_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(4), .Y_WIDTH(8) ) _37504_ ( .A(_cond_data_825), .B(__delay_data_1442), .Y(_22242_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37505_ ( .A(__substreamoutput_data_861), .B(__delay_data_1441), .Y(_22243_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37506_ ( .A(_source_stream_matmul_15_source_6_pat_cur_offset_0), .B(_source_stream_matmul_15_source_6_pat_stride_buf_0), .Y(_22244_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37507_ ( .A(_source_stream_matmul_15_source_6_pat_cur_offset_1), .B(_source_stream_matmul_15_source_6_pat_stride_buf_1), .Y(_22245_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37508_ ( .A(_source_stream_matmul_15_source_6_pat_cur_offset_2), .B(_source_stream_matmul_15_source_6_pat_stride_buf_2), .Y(_22246_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37509_ ( .A(_source_stream_matmul_15_source_6_pat_cur_offset_3), .B(_source_stream_matmul_15_source_6_pat_stride_buf_3), .Y(_22247_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37510_ ( .A(_source_stream_matmul_15_source_8_pat_cur_offset_0), .B(_source_stream_matmul_15_source_8_pat_stride_buf_0), .Y(_22248_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37511_ ( .A(_source_stream_matmul_15_source_8_pat_cur_offset_1), .B(_source_stream_matmul_15_source_8_pat_stride_buf_1), .Y(_22249_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37512_ ( .A(_source_stream_matmul_15_source_8_pat_cur_offset_2), .B(_source_stream_matmul_15_source_8_pat_stride_buf_2), .Y(_22250_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37513_ ( .A(_source_stream_matmul_15_source_8_pat_cur_offset_3), .B(_source_stream_matmul_15_source_8_pat_stride_buf_3), .Y(_22251_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37514_ ( .A(matmul_15_stream_act_local_0), .B(matmul_15_act_page_comp_offset_buf_0), .Y(_22252_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37515_ ( .A(_source_stream_matmul_15_source_19_pat_cur_offset_0), .B(_source_stream_matmul_15_source_19_pat_stride_buf_0), .Y(_22253_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37516_ ( .A(_source_stream_matmul_15_source_19_pat_cur_offset_1), .B(_source_stream_matmul_15_source_19_pat_stride_buf_1), .Y(_22254_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37517_ ( .A(_source_stream_matmul_15_source_19_pat_cur_offset_2), .B(_source_stream_matmul_15_source_19_pat_stride_buf_2), .Y(_22255_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37518_ ( .A(_source_stream_matmul_15_source_19_pat_cur_offset_3), .B(_source_stream_matmul_15_source_19_pat_stride_buf_3), .Y(_22256_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37519_ ( .A(_source_stream_matmul_15_source_20_pat_cur_offset_0), .B(_source_stream_matmul_15_source_20_pat_stride_buf_0), .Y(_22257_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37520_ ( .A(_source_stream_matmul_15_source_20_pat_cur_offset_1), .B(_source_stream_matmul_15_source_20_pat_stride_buf_1), .Y(_22258_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37521_ ( .A(_source_stream_matmul_15_source_20_pat_cur_offset_2), .B(_source_stream_matmul_15_source_20_pat_stride_buf_2), .Y(_22259_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37522_ ( .A(_source_stream_matmul_15_source_20_pat_cur_offset_3), .B(_source_stream_matmul_15_source_20_pat_stride_buf_3), .Y(_22260_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37523_ ( .A(matmul_15_stream_out_local_col), .B(matmul_15_out_page_comp_offset_buf), .Y(_22261_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37524_ ( .A(_stream_matmul_15_sink_21_sink_waddr), .B(_stream_matmul_15_sink_21_sink_stride_buf), .Y(_22262_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37525_ ( .A(_saxi_register_13), .B(576), .Y({ _03666_, _03665_, _03663_, _03662_, _03661_, _03660_, _03659_, _03658_, _03657_, _03656_, _03655_, _03654_, _03652_, _03651_, _03650_, _03649_, _03648_, _03647_, _03646_, _03645_, _03644_, _03643_, _03673_, _03672_, _03671_, _03670_, _03669_, _03668_, _03667_, _03664_, _03653_, _03642_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37526_ ( .A(_saxi_register_13), .B(640), .Y({ _03698_, _03697_, _03695_, _03694_, _03693_, _03692_, _03691_, _03690_, _03689_, _03688_, _03687_, _03686_, _03684_, _03683_, _03682_, _03681_, _03680_, _03679_, _03678_, _03677_, _03676_, _03675_, _03705_, _03704_, _03703_, _03702_, _03701_, _03700_, _03699_, _03696_, _03685_, _03674_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37527_ ( .A(_saxi_register_10), .B(12544), .Y({ _03730_, _03729_, _03727_, _03726_, _03725_, _03724_, _03723_, _03722_, _03721_, _03720_, _03719_, _03718_, _03716_, _03715_, _03714_, _03713_, _03712_, _03711_, _03710_, _03709_, _03708_, _03707_, _03737_, _03736_, _03735_, _03734_, _03733_, _03732_, _03731_, _03728_, _03717_, _03706_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37528_ ( .A(_saxi_register_13), .B(704), .Y({ _03794_, _03793_, _03791_, _03790_, _03789_, _03788_, _03787_, _03786_, _03785_, _03784_, _03783_, _03782_, _03780_, _03779_, _03778_, _03777_, _03776_, _03775_, _03774_, _03773_, _03772_, _03771_, _03801_, _03800_, _03799_, _03798_, _03797_, _03796_, _03795_, _03792_, _03781_, _03770_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37529_ ( .A(_saxi_register_13), .B(1856), .Y({ _03826_, _03825_, _03823_, _03822_, _03821_, _03820_, _03819_, _03818_, _03817_, _03816_, _03815_, _03814_, _03812_, _03811_, _03810_, _03809_, _03808_, _03807_, _03806_, _03805_, _03804_, _03803_, _03833_, _03832_, _03831_, _03830_, _03829_, _03828_, _03827_, _03824_, _03813_, _03802_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37530_ ( .A(_saxi_register_13), .B(1920), .Y({ _03858_, _03857_, _03855_, _03854_, _03853_, _03852_, _03851_, _03850_, _03849_, _03848_, _03847_, _03846_, _03844_, _03843_, _03842_, _03841_, _03840_, _03839_, _03838_, _03837_, _03836_, _03835_, _03865_, _03864_, _03863_, _03862_, _03861_, _03860_, _03859_, _03856_, _03845_, _03834_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37531_ ( .A(_saxi_register_10), .B(15680), .Y({ _03762_, _03761_, _03759_, _03758_, _03757_, _03756_, _03755_, _03754_, _03753_, _03752_, _03751_, _03750_, _03748_, _03747_, _03746_, _03745_, _03744_, _03743_, _03742_, _03741_, _03740_, _03739_, _03769_, _03768_, _03767_, _03766_, _03765_, _03764_, _03763_, _03760_, _03749_, _03738_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37532_ ( .A(_saxi_register_10), .B(16832), .Y({ _03890_, _03889_, _03887_, _03886_, _03885_, _03884_, _03883_, _03882_, _03881_, _03880_, _03879_, _03878_, _03876_, _03875_, _03874_, _03873_, _03872_, _03871_, _03870_, _03869_, _03868_, _03867_, _03897_, _03896_, _03895_, _03894_, _03893_, _03892_, _03891_, _03888_, _03877_, _03866_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37533_ ( .A(_saxi_register_13), .B(1984), .Y(_22263_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37534_ ( .A(_saxi_register_13), .B(4864), .Y(_22264_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37535_ ( .A(_saxi_register_13), .B(4928), .Y(_22265_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37536_ ( .A(conv2d_8_out_laddr_offset), .B(conv2d_8_next_out_write_size), .Y(_22266_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37537_ ( .A(conv2d_8_out_ram_select), .B(1), .Y(_22267_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37538_ ( .A(conv2d_8_sync_out_count), .B(cparam_conv2d_8_inc_sync_out), .Y({ _03922_, _03921_, _03919_, _03918_, _03917_, _03916_, _03915_, _03914_, _03913_, _03912_, _03911_, _03910_, _03908_, _03907_, _03906_, _03905_, _03904_, _03903_, _03902_, _03901_, _03900_, _03899_, _03929_, _03928_, _03927_, _03926_, _03925_, _03924_, _03923_, _03920_, _03909_, _03898_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37539_ ( .A(conv2d_8_sync_out_count), .B({ 27'h0000000, cparam_conv2d_8_inc_sync_out }), .Y({ _03954_, _03953_, _03951_, _03950_, _03949_, _03948_, _03947_, _03946_, _03945_, _03944_, _03943_, _03942_, _03940_, _03939_, _03938_, _03937_, _03936_, _03935_, _03934_, _03933_, _03932_, _03931_, _03961_, _03960_, _03959_, _03958_, _03957_, _03956_, _03955_, _03952_, _03941_, _03930_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(11), .Y_WIDTH(32) ) _37540_ ( .A(conv2d_8_filter_base_offset), .B(cparam_conv2d_8_filter_base_step), .Y(_22268_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _37541_ ( .A(conv2d_8_och_count), .B(cparam_conv2d_8_och_count_step), .Y(_22269_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(8), .Y_WIDTH(32) ) _37542_ ( .A(conv2d_8_filter_page_dma_offset), .B(cparam_conv2d_8_filter_read_step), .Y(_22271_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(8), .Y_WIDTH(32) ) _37543_ ( .A(conv2d_8_filter_page_comp_offset), .B(cparam_conv2d_8_filter_read_step), .Y(_22270_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(8), .Y_WIDTH(32) ) _37544_ ( .A(_22270_), .B(cparam_conv2d_8_filter_read_step), .Y({ _03986_, _03985_, _03983_, _03982_, _03981_, _03980_, _03979_, _03978_, _03977_, _03976_, _03975_, _03974_, _03972_, _03971_, _03970_, _03969_, _03968_, _03967_, _03966_, _03965_, _03964_, _03963_, _03993_, _03992_, _03991_, _03990_, _03989_, _03988_, _03987_, _03984_, _03973_, _03962_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(8), .Y_WIDTH(32) ) _37545_ ( .A(conv2d_8_act_base_offset_row), .B(cparam_conv2d_8_act_read_size), .Y(_22272_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(32) ) _37546_ ( .A(conv2d_8_row_count), .B(1'h1), .Y(_22273_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(2) ) _37547_ ( .A(conv2d_8_row_select), .B(1'h1), .Y(_22274_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(32) ) _37548_ ( .A(conv2d_8_row_select), .B(1'h1), .Y({ _04018_, _04017_, _04015_, _04014_, _04013_, _04012_, _04011_, _04010_, _04009_, _04008_, _04007_, _04006_, _04004_, _04003_, _04002_, _04001_, _04000_, _03999_, _03998_, _03997_, _03996_, _03995_, _04025_, _04024_, _04023_, _04022_, _04021_, _04020_, _04019_, _04016_, _04005_, _03994_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _37549_ ( .A(conv2d_8_act_page_dma_offset_0), .B(cparam_conv2d_8_act_read_step), .Y(_22276_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _37550_ ( .A(conv2d_8_act_page_comp_offset_0), .B(cparam_conv2d_8_act_read_step), .Y(_22275_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _37551_ ( .A(_22275_), .B(cparam_conv2d_8_act_read_step), .Y({ _04050_, _04049_, _04047_, _04046_, _04045_, _04044_, _04043_, _04042_, _04041_, _04040_, _04039_, _04038_, _04036_, _04035_, _04034_, _04033_, _04032_, _04031_, _04030_, _04029_, _04028_, _04027_, _04057_, _04056_, _04055_, _04054_, _04053_, _04052_, _04051_, _04048_, _04037_, _04026_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _37552_ ( .A(conv2d_8_act_page_dma_offset_1), .B(cparam_conv2d_8_act_read_step), .Y(_22278_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _37553_ ( .A(conv2d_8_act_page_comp_offset_1), .B(cparam_conv2d_8_act_read_step), .Y(_22277_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _37554_ ( .A(_22277_), .B(cparam_conv2d_8_act_read_step), .Y({ _04082_, _04081_, _04079_, _04078_, _04077_, _04076_, _04075_, _04074_, _04073_, _04072_, _04071_, _04070_, _04068_, _04067_, _04066_, _04065_, _04064_, _04063_, _04062_, _04061_, _04060_, _04059_, _04089_, _04088_, _04087_, _04086_, _04085_, _04084_, _04083_, _04080_, _04069_, _04058_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _37555_ ( .A(conv2d_8_act_page_dma_offset_2), .B(cparam_conv2d_8_act_read_step), .Y(_22280_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _37556_ ( .A(conv2d_8_act_page_comp_offset_2), .B(cparam_conv2d_8_act_read_step), .Y(_22279_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _37557_ ( .A(_22279_), .B(cparam_conv2d_8_act_read_step), .Y({ _04114_, _04113_, _04111_, _04110_, _04109_, _04108_, _04107_, _04106_, _04105_, _04104_, _04103_, _04102_, _04100_, _04099_, _04098_, _04097_, _04096_, _04095_, _04094_, _04093_, _04092_, _04091_, _04121_, _04120_, _04119_, _04118_, _04117_, _04116_, _04115_, _04112_, _04101_, _04090_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37558_ ( .A(conv2d_8_out_row_count), .B(1), .Y(_22282_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37559_ ( .A(conv2d_8_out_base_offset_och), .B(cparam_conv2d_8_bias_num), .Y(_22283_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(9), .Y_WIDTH(32) ) _37560_ ( .A(conv2d_8_out_base_offset_row), .B(cparam_conv2d_8_out_row_step), .Y(_22281_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37561_ ( .A(_maxi_read_global_addr), .B(_maxi_global_base_addr), .Y(_22284_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _37562_ ( .A({ 21'h000000, _maxi_read_cur_global_addr[11:0] }), .B({ _maxi_read_rest_size[30:0], 2'h0 }), .Y({ _04147_, _04146_, _04145_, _04143_, _04142_, _04141_, _04140_, _04139_, _04138_, _04137_, _04136_, _04135_, _04134_, _04132_, _04131_, _04130_, _04129_, _04128_, _04127_, _04126_, _04125_, _04124_, _04123_, _04154_, _04153_, _04152_, _04151_, _04150_, _04149_, _04148_, _04144_, _04133_, _04122_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37563_ ( .A({ 20'h00000, _maxi_read_cur_global_addr[11:0] }), .B(1024), .Y({ _04179_, _04178_, _04176_, _04175_, _04174_, _04173_, _04172_, _04171_, _04170_, _04169_, _04168_, _04167_, _04165_, _04164_, _04163_, _04162_, _04161_, _04160_, _04159_, _04158_, _04157_, _04156_, _04186_, _04185_, _04184_, _04183_, _04182_, _04181_, _04180_, _04177_, _04166_, _04155_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _37564_ ( .A(_maxi_read_cur_global_addr), .B({ _maxi_read_cur_size[30:0], 2'h0 }), .Y(_22285_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37565_ ( .A(conv2d_8_sync_comp_count), .B(1), .Y(_22286_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37566_ ( .A(conv2d_8_stream_act_local_0), .B(cparam_conv2d_8_inc_act_laddr_large), .Y(_22287_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37567_ ( .A(conv2d_8_stream_act_local_1), .B(cparam_conv2d_8_inc_act_laddr_large), .Y(_22288_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37568_ ( .A(conv2d_8_stream_act_local_2), .B(cparam_conv2d_8_inc_act_laddr_large), .Y(_22289_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37569_ ( .A(conv2d_8_stream_act_local_3), .B(cparam_conv2d_8_inc_act_laddr_large), .Y(_22290_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37570_ ( .A(conv2d_8_stream_act_local_4), .B(cparam_conv2d_8_inc_act_laddr_large), .Y(_22291_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37571_ ( .A(conv2d_8_stream_act_local_5), .B(cparam_conv2d_8_inc_act_laddr_large), .Y(_22292_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37572_ ( .A(conv2d_8_stream_act_local_6), .B(cparam_conv2d_8_inc_act_laddr_large), .Y(_22293_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37573_ ( .A(conv2d_8_stream_act_local_7), .B(cparam_conv2d_8_inc_act_laddr_large), .Y(_22294_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37574_ ( .A(conv2d_8_stream_act_local_8), .B(cparam_conv2d_8_inc_act_laddr_large), .Y(_22295_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37575_ ( .A(conv2d_8_stream_out_local_col), .B(conv2d_8_next_stream_num_ops), .Y(_22296_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(32) ) _37576_ ( .A(conv2d_8_col_count), .B(1'h1), .Y(_22297_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(2) ) _37577_ ( .A(conv2d_8_col_select), .B(1'h1), .Y(_22298_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(32) ) _37578_ ( .A(conv2d_8_col_select), .B(1'h1), .Y({ _04211_, _04210_, _04208_, _04207_, _04206_, _04205_, _04204_, _04203_, _04202_, _04201_, _04200_, _04199_, _04197_, _04196_, _04195_, _04194_, _04193_, _04192_, _04191_, _04190_, _04189_, _04188_, _04218_, _04217_, _04216_, _04215_, _04214_, _04213_, _04212_, _04209_, _04198_, _04187_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37579_ ( .A(_maxi_write_global_addr), .B(_maxi_global_base_addr), .Y(_22299_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _37580_ ( .A({ 21'h000000, _maxi_write_cur_global_addr[11:0] }), .B({ _maxi_write_rest_size[30:0], 2'h0 }), .Y({ _04244_, _04243_, _04242_, _04240_, _04239_, _04238_, _04237_, _04236_, _04235_, _04234_, _04233_, _04232_, _04231_, _04229_, _04228_, _04227_, _04226_, _04225_, _04224_, _04223_, _04222_, _04221_, _04220_, _04251_, _04250_, _04249_, _04248_, _04247_, _04246_, _04245_, _04241_, _04230_, _04219_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37581_ ( .A({ 20'h00000, _maxi_write_cur_global_addr[11:0] }), .B(1024), .Y({ _04276_, _04275_, _04273_, _04272_, _04271_, _04270_, _04269_, _04268_, _04267_, _04266_, _04265_, _04264_, _04262_, _04261_, _04260_, _04259_, _04258_, _04257_, _04256_, _04255_, _04254_, _04253_, _04283_, _04282_, _04281_, _04280_, _04279_, _04278_, _04277_, _04274_, _04263_, _04252_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _37582_ ( .A(_maxi_write_cur_global_addr), .B({ _maxi_write_cur_size[30:0], 2'h0 }), .Y(_22300_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(8), .Y_WIDTH(32) ) _37583_ ( .A(max_pool_serial_9_out_count), .B(cparam_max_pool_serial_9_out_row_step), .Y({ _04308_, _04307_, _04305_, _04304_, _04303_, _04302_, _04301_, _04300_, _04299_, _04298_, _04297_, _04296_, _04294_, _04293_, _04292_, _04291_, _04290_, _04289_, _04288_, _04287_, _04286_, _04285_, _04315_, _04314_, _04313_, _04312_, _04311_, _04310_, _04309_, _04306_, _04295_, _04284_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(10), .Y_WIDTH(32) ) _37584_ ( .A(max_pool_serial_9_act_base_offset_row), .B(cparam_max_pool_serial_9_act_row_step), .Y(_22301_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(32) ) _37585_ ( .A(max_pool_serial_9_row_count), .B(2'h2), .Y(_22302_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(8), .Y_WIDTH(32) ) _37586_ ( .A(max_pool_serial_9_out_base_offset_row), .B(cparam_max_pool_serial_9_out_row_step), .Y(_22303_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37587_ ( .A(max_pool_serial_9_comp_count), .B(cparam_max_pool_serial_9_inc_out_laddr), .Y(_22304_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(6), .Y_WIDTH(32) ) _37588_ ( .A(max_pool_serial_9_stream_act_local), .B(cparam_max_pool_serial_9_inc_act_laddr), .Y(_22305_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _37589_ ( .A(max_pool_serial_9_stream_out_local), .B(cparam_max_pool_serial_9_inc_out_laddr), .Y(_22306_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(32) ) _37590_ ( .A(max_pool_serial_9_col_count), .B(2'h2), .Y(_22307_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37591_ ( .A(matmul_15_out_laddr_offset), .B(matmul_15_next_out_write_size), .Y(_22308_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(4), .Y_WIDTH(32) ) _37592_ ( .A(matmul_15_out_base_offset_col), .B(4'hc), .Y({ _04372_, _04371_, _04369_, _04368_, _04367_, _04366_, _04365_, _04364_, _04363_, _04362_, _04361_, _04360_, _04358_, _04357_, _04356_, _04355_, _04354_, _04353_, _04352_, _04351_, _04350_, _04349_, _04379_, _04378_, _04377_, _04376_, _04375_, _04374_, _04373_, _04370_, _04359_, _04348_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37593_ ( .A(matmul_15_out_ram_select), .B(1), .Y(_22309_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(32) ) _37594_ ( .A(matmul_15_sync_out_count), .B(1'h1), .Y({ _04340_, _04339_, _04337_, _04336_, _04335_, _04334_, _04333_, _04332_, _04331_, _04330_, _04329_, _04328_, _04326_, _04325_, _04324_, _04323_, _04322_, _04321_, _04320_, _04319_, _04318_, _04317_, _04347_, _04346_, _04345_, _04344_, _04343_, _04342_, _04341_, _04338_, _04327_, _04316_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37595_ ( .A(matmul_15_sync_out_count), .B(1), .Y({ _12503_, _12502_, _12500_, _12499_, _12498_, _12497_, _12496_, _12495_, _12494_, _12493_, _12492_, _12491_, _12489_, _12488_, _12487_, _12486_, _12485_, _12484_, _12483_, _12482_, _12481_, _12480_, _12510_, _12509_, _12508_, _12507_, _12506_, _12505_, _12504_, _12501_, _12490_, _12479_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(11), .Y_WIDTH(32) ) _37596_ ( .A(matmul_15_filter_base_offset), .B(11'h480), .Y({ _04404_, _04403_, _04401_, _04400_, _04399_, _04398_, _04397_, _04396_, _04395_, _04394_, _04393_, _04392_, _04390_, _04389_, _04388_, _04387_, _04386_, _04385_, _04384_, _04383_, _04382_, _04381_, _04411_, _04410_, _04409_, _04408_, _04407_, _04406_, _04405_, _04402_, _04391_, _04380_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(3), .Y_WIDTH(32) ) _37597_ ( .A(matmul_15_och_count), .B(3'h4), .Y({ _04436_, _04435_, _04433_, _04432_, _04431_, _04430_, _04429_, _04428_, _04427_, _04426_, _04425_, _04424_, _04422_, _04421_, _04420_, _04419_, _04418_, _04417_, _04416_, _04415_, _04414_, _04413_, _04443_, _04442_, _04441_, _04440_, _04439_, _04438_, _04437_, _04434_, _04423_, _04412_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(11), .Y_WIDTH(32) ) _37598_ ( .A(matmul_15_filter_page_dma_offset), .B(11'h480), .Y(_22311_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(11), .Y_WIDTH(32) ) _37599_ ( .A(matmul_15_filter_page_comp_offset), .B(11'h480), .Y(_22310_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(11), .Y_WIDTH(32) ) _37600_ ( .A(_22310_), .B(11'h480), .Y({ _04468_, _04467_, _04465_, _04464_, _04463_, _04462_, _04461_, _04460_, _04459_, _04458_, _04457_, _04456_, _04454_, _04453_, _04452_, _04451_, _04450_, _04449_, _04448_, _04447_, _04446_, _04445_, _04475_, _04474_, _04473_, _04472_, _04471_, _04470_, _04469_, _04466_, _04455_, _04444_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(3), .Y_WIDTH(32) ) _37601_ ( .A(matmul_15_out_base_offset_och), .B(3'h4), .Y(_22312_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37602_ ( .A(matmul_15_sync_comp_count), .B(1), .Y(_22313_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37603_ ( .A(conv2d_8_act_base_offset_row), .B(conv2d_8_act_base_offset_bat), .Y(conv2d_8_act_base_offset) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37604_ ( .A(conv2d_8_out_base_offset_val), .B(conv2d_8_out_base_offset_col), .Y(_22314_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37605_ ( .A(_22314_), .B(conv2d_8_out_base_offset_row), .Y(_22315_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37606_ ( .A(_22315_), .B(conv2d_8_out_base_offset_bat), .Y(_22316_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _37607_ ( .A(_22316_), .B(conv2d_8_out_base_offset_och), .Y(conv2d_8_out_base_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37608_ ( .A(_tmp_35), .B(_maxi_read_local_stride), .Y({ _22317_[31:9], _tmp_44 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37609_ ( .A(_tmp_36), .B(_maxi_read_local_stride), .Y({ _22318_[31:9], _tmp_45 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37610_ ( .A(_tmp_37), .B(_maxi_read_local_stride), .Y({ _22319_[31:9], _tmp_46 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37611_ ( .A(_tmp_38), .B(_maxi_read_local_stride), .Y({ _22320_[31:9], _tmp_47 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37612_ ( .A(_tmp_39), .B(_maxi_read_local_stride), .Y({ _22321_[31:9], _tmp_48 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37613_ ( .A(_tmp_40), .B(_maxi_read_local_stride), .Y({ _22322_[31:9], _tmp_49 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37614_ ( .A(_tmp_41), .B(_maxi_read_local_stride), .Y({ _22323_[31:9], _tmp_50 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37615_ ( .A(_tmp_42), .B(_maxi_read_local_stride), .Y({ _22324_[31:9], _tmp_51 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37616_ ( .A(_tmp_43), .B(_maxi_read_local_stride), .Y({ _22325_[31:9], _tmp_52 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37617_ ( .A(_tmp_66), .B(_maxi_read_local_stride), .Y({ _22326_[31:9], _tmp_75 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37618_ ( .A(_tmp_67), .B(_maxi_read_local_stride), .Y({ _22327_[31:9], _tmp_76 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37619_ ( .A(_tmp_68), .B(_maxi_read_local_stride), .Y({ _22328_[31:9], _tmp_77 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37620_ ( .A(_tmp_69), .B(_maxi_read_local_stride), .Y({ _22329_[31:9], _tmp_78 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37621_ ( .A(_tmp_70), .B(_maxi_read_local_stride), .Y({ _22330_[31:9], _tmp_79 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37622_ ( .A(_tmp_71), .B(_maxi_read_local_stride), .Y({ _22331_[31:9], _tmp_80 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37623_ ( .A(_tmp_72), .B(_maxi_read_local_stride), .Y({ _22332_[31:9], _tmp_81 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37624_ ( .A(_tmp_73), .B(_maxi_read_local_stride), .Y({ _22333_[31:9], _tmp_82 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37625_ ( .A(_tmp_74), .B(_maxi_read_local_stride), .Y({ _22334_[31:9], _tmp_83 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37626_ ( .A(_tmp_97), .B(_maxi_read_local_stride), .Y({ _22335_[31:9], _tmp_106 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37627_ ( .A(_tmp_98), .B(_maxi_read_local_stride), .Y({ _22336_[31:9], _tmp_107 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37628_ ( .A(_tmp_99), .B(_maxi_read_local_stride), .Y({ _22337_[31:9], _tmp_108 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37629_ ( .A(_tmp_100), .B(_maxi_read_local_stride), .Y({ _22338_[31:9], _tmp_109 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37630_ ( .A(_tmp_101), .B(_maxi_read_local_stride), .Y({ _22339_[31:9], _tmp_110 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37631_ ( .A(_tmp_102), .B(_maxi_read_local_stride), .Y({ _22340_[31:9], _tmp_111 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37632_ ( .A(_tmp_103), .B(_maxi_read_local_stride), .Y({ _22341_[31:9], _tmp_112 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37633_ ( .A(_tmp_104), .B(_maxi_read_local_stride), .Y({ _22342_[31:9], _tmp_113 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37634_ ( .A(_tmp_105), .B(_maxi_read_local_stride), .Y({ _22343_[31:9], _tmp_114 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37635_ ( .A(_tmp_128), .B(_maxi_read_local_stride), .Y({ _22344_[31:9], _tmp_137 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37636_ ( .A(_tmp_129), .B(_maxi_read_local_stride), .Y({ _22345_[31:9], _tmp_138 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37637_ ( .A(_tmp_130), .B(_maxi_read_local_stride), .Y({ _22346_[31:9], _tmp_139 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37638_ ( .A(_tmp_131), .B(_maxi_read_local_stride), .Y({ _22347_[31:9], _tmp_140 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37639_ ( .A(_tmp_132), .B(_maxi_read_local_stride), .Y({ _22348_[31:9], _tmp_141 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37640_ ( .A(_tmp_133), .B(_maxi_read_local_stride), .Y({ _22349_[31:9], _tmp_142 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37641_ ( .A(_tmp_134), .B(_maxi_read_local_stride), .Y({ _22350_[31:9], _tmp_143 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37642_ ( .A(_tmp_135), .B(_maxi_read_local_stride), .Y({ _22351_[31:9], _tmp_144 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37643_ ( .A(_tmp_136), .B(_maxi_read_local_stride), .Y({ _22352_[31:9], _tmp_145 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37644_ ( .A(conv2d_8_act_base_offset), .B(cparam_conv2d_8_act_offset_values_2), .Y(_22355_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37645_ ( .A(conv2d_8_arg_objaddr_0), .B(_22355_), .Y(_22356_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37646_ ( .A(conv2d_8_act_base_offset), .B(cparam_conv2d_8_act_offset_values_1), .Y(_22357_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37647_ ( .A(conv2d_8_arg_objaddr_0), .B(_22357_), .Y(_22358_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37648_ ( .A(conv2d_8_act_base_offset), .B(cparam_conv2d_8_act_offset_values_0), .Y(_22353_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37649_ ( .A(conv2d_8_arg_objaddr_0), .B(_22353_), .Y(_22354_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37650_ ( .A(conv2d_8_row_count), .B(1), .Y({ _04532_, _04531_, _04529_, _04528_, _04527_, _04526_, _04525_, _04524_, _04523_, _04522_, _04521_, _04520_, _04518_, _04517_, _04516_, _04515_, _04514_, _04513_, _04512_, _04511_, _04510_, _04509_, _04539_, _04538_, _04537_, _04536_, _04535_, _04534_, _04533_, _04530_, _04519_, _04508_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37651_ ( .A(conv2d_8_row_count), .B(2), .Y({ _04564_, _04563_, _04561_, _04560_, _04559_, _04558_, _04557_, _04556_, _04555_, _04554_, _04553_, _04552_, _04550_, _04549_, _04548_, _04547_, _04546_, _04545_, _04544_, _04543_, _04542_, _04541_, _04571_, _04570_, _04569_, _04568_, _04567_, _04566_, _04565_, _04562_, _04551_, _04540_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37652_ ( .A(_tmp_164), .B(_maxi_read_local_stride), .Y({ _22359_[31:9], _tmp_167 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37653_ ( .A(_tmp_165), .B(_maxi_read_local_stride), .Y({ _22360_[31:9], _tmp_168 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37654_ ( .A(_tmp_166), .B(_maxi_read_local_stride), .Y({ _22361_[31:9], _tmp_169 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37655_ ( .A(_tmp_177), .B(_maxi_read_local_stride), .Y({ _22362_[31:9], _tmp_180 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37656_ ( .A(_tmp_178), .B(_maxi_read_local_stride), .Y({ _22363_[31:9], _tmp_181 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37657_ ( .A(_tmp_179), .B(_maxi_read_local_stride), .Y({ _22364_[31:9], _tmp_182 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37658_ ( .A(_tmp_190), .B(_maxi_read_local_stride), .Y({ _22365_[31:9], _tmp_193 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37659_ ( .A(_tmp_191), .B(_maxi_read_local_stride), .Y({ _22366_[31:9], _tmp_194 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37660_ ( .A(_tmp_192), .B(_maxi_read_local_stride), .Y({ _22367_[31:9], _tmp_195 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37661_ ( .A(_tmp_203), .B(_maxi_read_local_stride), .Y({ _22368_[31:9], _tmp_206 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37662_ ( .A(_tmp_204), .B(_maxi_read_local_stride), .Y({ _22369_[31:9], _tmp_207 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37663_ ( .A(_tmp_205), .B(_maxi_read_local_stride), .Y({ _22370_[31:9], _tmp_208 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37664_ ( .A(_tmp_221), .B(_maxi_read_local_stride), .Y({ _22371_[31:9], _tmp_224 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37665_ ( .A(_tmp_222), .B(_maxi_read_local_stride), .Y({ _22372_[31:9], _tmp_225 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37666_ ( .A(_tmp_223), .B(_maxi_read_local_stride), .Y({ _22373_[31:9], _tmp_226 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37667_ ( .A(_tmp_234), .B(_maxi_read_local_stride), .Y({ _22374_[31:9], _tmp_237 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37668_ ( .A(_tmp_235), .B(_maxi_read_local_stride), .Y({ _22375_[31:9], _tmp_238 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37669_ ( .A(_tmp_236), .B(_maxi_read_local_stride), .Y({ _22376_[31:9], _tmp_239 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37670_ ( .A(_tmp_247), .B(_maxi_read_local_stride), .Y({ _22377_[31:9], _tmp_250 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37671_ ( .A(_tmp_248), .B(_maxi_read_local_stride), .Y({ _22378_[31:9], _tmp_251 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37672_ ( .A(_tmp_249), .B(_maxi_read_local_stride), .Y({ _22379_[31:9], _tmp_252 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37673_ ( .A(_tmp_260), .B(_maxi_read_local_stride), .Y({ _22380_[31:9], _tmp_263 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37674_ ( .A(_tmp_261), .B(_maxi_read_local_stride), .Y({ _22381_[31:9], _tmp_264 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37675_ ( .A(_tmp_262), .B(_maxi_read_local_stride), .Y({ _22382_[31:9], _tmp_265 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37676_ ( .A(_tmp_278), .B(_maxi_read_local_stride), .Y({ _22383_[31:9], _tmp_281 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37677_ ( .A(_tmp_279), .B(_maxi_read_local_stride), .Y({ _22384_[31:9], _tmp_282 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37678_ ( .A(_tmp_280), .B(_maxi_read_local_stride), .Y({ _22385_[31:9], _tmp_283 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37679_ ( .A(_tmp_291), .B(_maxi_read_local_stride), .Y({ _22386_[31:9], _tmp_294 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37680_ ( .A(_tmp_292), .B(_maxi_read_local_stride), .Y({ _22387_[31:9], _tmp_295 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37681_ ( .A(_tmp_293), .B(_maxi_read_local_stride), .Y({ _22388_[31:9], _tmp_296 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37682_ ( .A(_tmp_304), .B(_maxi_read_local_stride), .Y({ _22389_[31:9], _tmp_307 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37683_ ( .A(_tmp_305), .B(_maxi_read_local_stride), .Y({ _22390_[31:9], _tmp_308 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37684_ ( .A(_tmp_306), .B(_maxi_read_local_stride), .Y({ _22391_[31:9], _tmp_309 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37685_ ( .A(_tmp_317), .B(_maxi_read_local_stride), .Y({ _22392_[31:9], _tmp_320 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37686_ ( .A(_tmp_318), .B(_maxi_read_local_stride), .Y({ _22393_[31:9], _tmp_321 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37687_ ( .A(_tmp_319), .B(_maxi_read_local_stride), .Y({ _22394_[31:9], _tmp_322 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37688_ ( .A(conv2d_8_row_count_buf), .B(1), .Y({ _04660_, _04659_, _04657_, _04656_, _04655_, _04654_, _04653_, _04652_, _04651_, _04650_, _04649_, _04648_, _04646_, _04645_, _04644_, _04643_, _04642_, _04641_, _04640_, _04639_, _04638_, _04637_, _04667_, _04666_, _04665_, _04664_, _04663_, _04662_, _04661_, _04658_, _04647_, _04636_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37689_ ( .A(conv2d_8_col_count), .B(1), .Y({ _04596_, _04595_, _04593_, _04592_, _04591_, _04590_, _04589_, _04588_, _04587_, _04586_, _04585_, _04584_, _04582_, _04581_, _04580_, _04579_, _04578_, _04577_, _04576_, _04575_, _04574_, _04573_, _04603_, _04602_, _04601_, _04600_, _04599_, _04598_, _04597_, _04594_, _04583_, _04572_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37690_ ( .A(conv2d_8_col_count), .B(2), .Y({ _04628_, _04627_, _04625_, _04624_, _04623_, _04622_, _04621_, _04620_, _04619_, _04618_, _04617_, _04616_, _04614_, _04613_, _04612_, _04611_, _04610_, _04609_, _04608_, _04607_, _04606_, _04605_, _04635_, _04634_, _04633_, _04632_, _04631_, _04630_, _04629_, _04626_, _04615_, _04604_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37691_ ( .A(conv2d_8_row_count_buf), .B(2), .Y({ _04692_, _04691_, _04689_, _04688_, _04687_, _04686_, _04685_, _04684_, _04683_, _04682_, _04681_, _04680_, _04678_, _04677_, _04676_, _04675_, _04674_, _04673_, _04672_, _04671_, _04670_, _04669_, _04699_, _04698_, _04697_, _04696_, _04695_, _04694_, _04693_, _04690_, _04679_, _04668_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(5), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(32) ) _37692_ ( .A(cparam_conv2d_8_act_num_row), .B(cparam_conv2d_8_pad_col_left), .Y({ _04500_, _04499_, _04497_, _04496_, _04495_, _04494_, _04493_, _04492_, _04491_, _04490_, _04489_, _04488_, _04486_, _04485_, _04484_, _04483_, _04482_, _04481_, _04480_, _04479_, _04478_, _04477_, _04507_, _04506_, _04505_, _04504_, _04503_, _04502_, _04501_, _04498_, _04487_, _04476_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37693_ ( .A(_stream_conv2d_8_source_6_source_offset_buf), .B(_source_stream_conv2d_8_source_6_pat_cur_offset_0), .Y(_22395_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37694_ ( .A(_22395_), .B(_source_stream_conv2d_8_source_6_pat_cur_offset_1), .Y(_22396_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37695_ ( .A(_22396_), .B(_source_stream_conv2d_8_source_6_pat_cur_offset_2), .Y(_22397_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37696_ ( .A(_22397_), .B(_source_stream_conv2d_8_source_6_pat_cur_offset_3), .Y(_stream_conv2d_8_source_6_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37697_ ( .A(_stream_conv2d_8_source_8_source_offset_buf), .B(_source_stream_conv2d_8_source_8_pat_cur_offset_0), .Y(_22398_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37698_ ( .A(_22398_), .B(_source_stream_conv2d_8_source_8_pat_cur_offset_1), .Y(_22399_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37699_ ( .A(_22399_), .B(_source_stream_conv2d_8_source_8_pat_cur_offset_2), .Y(_22400_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37700_ ( .A(_22400_), .B(_source_stream_conv2d_8_source_8_pat_cur_offset_3), .Y(_stream_conv2d_8_source_8_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37701_ ( .A(_stream_conv2d_8_source_19_source_offset_buf), .B(_source_stream_conv2d_8_source_19_pat_cur_offset_0), .Y(_22401_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37702_ ( .A(_22401_), .B(_source_stream_conv2d_8_source_19_pat_cur_offset_1), .Y(_22402_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37703_ ( .A(_22402_), .B(_source_stream_conv2d_8_source_19_pat_cur_offset_2), .Y(_22403_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37704_ ( .A(_22403_), .B(_source_stream_conv2d_8_source_19_pat_cur_offset_3), .Y(_stream_conv2d_8_source_19_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37705_ ( .A(_stream_conv2d_8_source_20_source_offset_buf), .B(_source_stream_conv2d_8_source_20_pat_cur_offset_0), .Y(_22404_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37706_ ( .A(_22404_), .B(_source_stream_conv2d_8_source_20_pat_cur_offset_1), .Y(_22405_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37707_ ( .A(_22405_), .B(_source_stream_conv2d_8_source_20_pat_cur_offset_2), .Y(_22406_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37708_ ( .A(_22406_), .B(_source_stream_conv2d_8_source_20_pat_cur_offset_3), .Y(_stream_conv2d_8_source_20_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37709_ ( .A(_stream_conv2d_8_source_21_source_offset_buf), .B(_source_stream_conv2d_8_source_21_pat_cur_offset_0), .Y(_22407_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37710_ ( .A(_22407_), .B(_source_stream_conv2d_8_source_21_pat_cur_offset_1), .Y(_22408_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37711_ ( .A(_22408_), .B(_source_stream_conv2d_8_source_21_pat_cur_offset_2), .Y(_22409_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37712_ ( .A(_22409_), .B(_source_stream_conv2d_8_source_21_pat_cur_offset_3), .Y(_stream_conv2d_8_source_21_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37713_ ( .A(_stream_conv2d_8_source_22_source_offset_buf), .B(_source_stream_conv2d_8_source_22_pat_cur_offset_0), .Y(_22410_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37714_ ( .A(_22410_), .B(_source_stream_conv2d_8_source_22_pat_cur_offset_1), .Y(_22411_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37715_ ( .A(_22411_), .B(_source_stream_conv2d_8_source_22_pat_cur_offset_2), .Y(_22412_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37716_ ( .A(_22412_), .B(_source_stream_conv2d_8_source_22_pat_cur_offset_3), .Y(_stream_conv2d_8_source_22_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37717_ ( .A(_stream_conv2d_8_source_23_source_offset_buf), .B(_source_stream_conv2d_8_source_23_pat_cur_offset_0), .Y(_22413_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37718_ ( .A(_22413_), .B(_source_stream_conv2d_8_source_23_pat_cur_offset_1), .Y(_22414_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37719_ ( .A(_22414_), .B(_source_stream_conv2d_8_source_23_pat_cur_offset_2), .Y(_22415_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37720_ ( .A(_22415_), .B(_source_stream_conv2d_8_source_23_pat_cur_offset_3), .Y(_stream_conv2d_8_source_23_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37721_ ( .A(_stream_conv2d_8_source_24_source_offset_buf), .B(_source_stream_conv2d_8_source_24_pat_cur_offset_0), .Y(_22416_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37722_ ( .A(_22416_), .B(_source_stream_conv2d_8_source_24_pat_cur_offset_1), .Y(_22417_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37723_ ( .A(_22417_), .B(_source_stream_conv2d_8_source_24_pat_cur_offset_2), .Y(_22418_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37724_ ( .A(_22418_), .B(_source_stream_conv2d_8_source_24_pat_cur_offset_3), .Y(_stream_conv2d_8_source_24_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37725_ ( .A(_stream_conv2d_8_source_25_source_offset_buf), .B(_source_stream_conv2d_8_source_25_pat_cur_offset_0), .Y(_22419_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37726_ ( .A(_22419_), .B(_source_stream_conv2d_8_source_25_pat_cur_offset_1), .Y(_22420_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37727_ ( .A(_22420_), .B(_source_stream_conv2d_8_source_25_pat_cur_offset_2), .Y(_22421_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37728_ ( .A(_22421_), .B(_source_stream_conv2d_8_source_25_pat_cur_offset_3), .Y(_stream_conv2d_8_source_25_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37729_ ( .A(_stream_conv2d_8_source_26_source_offset_buf), .B(_source_stream_conv2d_8_source_26_pat_cur_offset_0), .Y(_22422_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37730_ ( .A(_22422_), .B(_source_stream_conv2d_8_source_26_pat_cur_offset_1), .Y(_22423_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37731_ ( .A(_22423_), .B(_source_stream_conv2d_8_source_26_pat_cur_offset_2), .Y(_22424_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37732_ ( .A(_22424_), .B(_source_stream_conv2d_8_source_26_pat_cur_offset_3), .Y(_stream_conv2d_8_source_26_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37733_ ( .A(_stream_conv2d_8_source_27_source_offset_buf), .B(_source_stream_conv2d_8_source_27_pat_cur_offset_0), .Y(_22425_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37734_ ( .A(_22425_), .B(_source_stream_conv2d_8_source_27_pat_cur_offset_1), .Y(_22426_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37735_ ( .A(_22426_), .B(_source_stream_conv2d_8_source_27_pat_cur_offset_2), .Y(_22427_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37736_ ( .A(_22427_), .B(_source_stream_conv2d_8_source_27_pat_cur_offset_3), .Y(_stream_conv2d_8_source_27_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37737_ ( .A(_stream_conv2d_8_source_28_source_offset_buf), .B(_source_stream_conv2d_8_source_28_pat_cur_offset_0), .Y(_22428_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37738_ ( .A(_22428_), .B(_source_stream_conv2d_8_source_28_pat_cur_offset_1), .Y(_22429_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37739_ ( .A(_22429_), .B(_source_stream_conv2d_8_source_28_pat_cur_offset_2), .Y(_22430_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37740_ ( .A(_22430_), .B(_source_stream_conv2d_8_source_28_pat_cur_offset_3), .Y(_stream_conv2d_8_source_28_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37741_ ( .A(_stream_conv2d_8_source_29_source_offset_buf), .B(_source_stream_conv2d_8_source_29_pat_cur_offset_0), .Y(_22431_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37742_ ( .A(_22431_), .B(_source_stream_conv2d_8_source_29_pat_cur_offset_1), .Y(_22432_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37743_ ( .A(_22432_), .B(_source_stream_conv2d_8_source_29_pat_cur_offset_2), .Y(_22433_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37744_ ( .A(_22433_), .B(_source_stream_conv2d_8_source_29_pat_cur_offset_3), .Y(_stream_conv2d_8_source_29_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37745_ ( .A(_stream_conv2d_8_source_30_source_offset_buf), .B(_source_stream_conv2d_8_source_30_pat_cur_offset_0), .Y(_22434_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37746_ ( .A(_22434_), .B(_source_stream_conv2d_8_source_30_pat_cur_offset_1), .Y(_22435_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37747_ ( .A(_22435_), .B(_source_stream_conv2d_8_source_30_pat_cur_offset_2), .Y(_22436_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37748_ ( .A(_22436_), .B(_source_stream_conv2d_8_source_30_pat_cur_offset_3), .Y(_stream_conv2d_8_source_30_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37749_ ( .A(_stream_conv2d_8_source_31_source_offset_buf), .B(_source_stream_conv2d_8_source_31_pat_cur_offset_0), .Y(_22437_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37750_ ( .A(_22437_), .B(_source_stream_conv2d_8_source_31_pat_cur_offset_1), .Y(_22438_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37751_ ( .A(_22438_), .B(_source_stream_conv2d_8_source_31_pat_cur_offset_2), .Y(_22439_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37752_ ( .A(_22439_), .B(_source_stream_conv2d_8_source_31_pat_cur_offset_3), .Y(_stream_conv2d_8_source_31_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37753_ ( .A(_stream_conv2d_8_source_32_source_offset_buf), .B(_source_stream_conv2d_8_source_32_pat_cur_offset_0), .Y(_22440_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37754_ ( .A(_22440_), .B(_source_stream_conv2d_8_source_32_pat_cur_offset_1), .Y(_22441_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37755_ ( .A(_22441_), .B(_source_stream_conv2d_8_source_32_pat_cur_offset_2), .Y(_22442_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37756_ ( .A(_22442_), .B(_source_stream_conv2d_8_source_32_pat_cur_offset_3), .Y(_stream_conv2d_8_source_32_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37757_ ( .A(_stream_conv2d_8_source_33_source_offset_buf), .B(_source_stream_conv2d_8_source_33_pat_cur_offset_0), .Y(_22443_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37758_ ( .A(_22443_), .B(_source_stream_conv2d_8_source_33_pat_cur_offset_1), .Y(_22444_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37759_ ( .A(_22444_), .B(_source_stream_conv2d_8_source_33_pat_cur_offset_2), .Y(_22445_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37760_ ( .A(_22445_), .B(_source_stream_conv2d_8_source_33_pat_cur_offset_3), .Y(_stream_conv2d_8_source_33_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37761_ ( .A(_stream_conv2d_8_source_34_source_offset_buf), .B(_source_stream_conv2d_8_source_34_pat_cur_offset_0), .Y(_22446_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37762_ ( .A(_22446_), .B(_source_stream_conv2d_8_source_34_pat_cur_offset_1), .Y(_22447_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37763_ ( .A(_22447_), .B(_source_stream_conv2d_8_source_34_pat_cur_offset_2), .Y(_22448_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37764_ ( .A(_22448_), .B(_source_stream_conv2d_8_source_34_pat_cur_offset_3), .Y(_stream_conv2d_8_source_34_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37765_ ( .A(_stream_conv2d_8_source_35_source_offset_buf), .B(_source_stream_conv2d_8_source_35_pat_cur_offset_0), .Y(_22449_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37766_ ( .A(_22449_), .B(_source_stream_conv2d_8_source_35_pat_cur_offset_1), .Y(_22450_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37767_ ( .A(_22450_), .B(_source_stream_conv2d_8_source_35_pat_cur_offset_2), .Y(_22451_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37768_ ( .A(_22451_), .B(_source_stream_conv2d_8_source_35_pat_cur_offset_3), .Y(_stream_conv2d_8_source_35_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37769_ ( .A(_stream_conv2d_8_source_36_source_offset_buf), .B(_source_stream_conv2d_8_source_36_pat_cur_offset_0), .Y(_22452_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37770_ ( .A(_22452_), .B(_source_stream_conv2d_8_source_36_pat_cur_offset_1), .Y(_22453_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37771_ ( .A(_22453_), .B(_source_stream_conv2d_8_source_36_pat_cur_offset_2), .Y(_22454_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _37772_ ( .A(_22454_), .B(_source_stream_conv2d_8_source_36_pat_cur_offset_3), .Y(_stream_conv2d_8_source_36_source_pat_all_offset) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(16), .B_SIGNED(1), .B_WIDTH(16), .Y_WIDTH(16) ) _49073_ ( .A(\__muladd_madd_110.madd._mul ), .B(\__muladd_madd_110.madd._c ), .Y(\__muladd_madd_110.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(16), .B_SIGNED(1), .B_WIDTH(16), .Y_WIDTH(16) ) _49080_ ( .A(\__muladd_madd_125.madd._mul ), .B(\__muladd_madd_125.madd._c ), .Y(\__muladd_madd_125.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(16), .B_SIGNED(1), .B_WIDTH(16), .Y_WIDTH(16) ) _49087_ ( .A(\__muladd_madd_140.madd._mul ), .B(\__muladd_madd_140.madd._c ), .Y(\__muladd_madd_140.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(16), .B_SIGNED(1), .B_WIDTH(16), .Y_WIDTH(16) ) _49094_ ( .A(\__muladd_madd_155.madd._mul ), .B(\__muladd_madd_155.madd._c ), .Y(\__muladd_madd_155.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(16), .B_SIGNED(1), .B_WIDTH(16), .Y_WIDTH(16) ) _49101_ ( .A(\__muladd_madd_170.madd._mul ), .B(\__muladd_madd_170.madd._c ), .Y(\__muladd_madd_170.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(16), .B_SIGNED(1), .B_WIDTH(16), .Y_WIDTH(16) ) _49108_ ( .A(\__muladd_madd_185.madd._mul ), .B(\__muladd_madd_185.madd._c ), .Y(\__muladd_madd_185.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(16), .B_SIGNED(1), .B_WIDTH(16), .Y_WIDTH(16) ) _49115_ ( .A(\__muladd_madd_65.madd._mul ), .B(\__muladd_madd_65.madd._c ), .Y(\__muladd_madd_65.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(16), .B_SIGNED(1), .B_WIDTH(16), .Y_WIDTH(16) ) _49122_ ( .A(\__muladd_madd_80.madd._mul ), .B(\__muladd_madd_80.madd._c ), .Y(\__muladd_madd_80.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(16), .B_SIGNED(1), .B_WIDTH(16), .Y_WIDTH(16) ) _49129_ ( .A(\__muladd_madd_95.madd._mul ), .B(\__muladd_madd_95.madd._c ), .Y(\__muladd_madd_95.madd._madd ) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48394_ ( .A(_maxi_read_cur_size), .B(1), .Y(_25935_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48395_ ( .A(_tmp_14), .B(1), .Y(_25936_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48396_ ( .A(_maxi_write_cur_size), .B(1), .Y(_25937_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48397_ ( .A(_tmp_847), .B(1), .Y(_25938_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48398_ ( .A(_tmp_964), .B(1), .Y(_25940_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48399_ ( .A(_tmp_966), .B(1), .Y(_25941_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48400_ ( .A(_tmp_968), .B(1), .Y(_25942_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48401_ ( .A(_tmp_970), .B(1), .Y(_25943_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48402_ ( .A(_tmp_19), .B(1), .Y(_25944_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48403_ ( .A(_tmp_921), .B(1), .Y(_25946_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48404_ ( .A(_tmp_21), .B(1), .Y(_25947_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48405_ ( .A(_tmp_933), .B(1), .Y(_25948_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48406_ ( .A(_tmp_23), .B(1), .Y(_25949_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48407_ ( .A(_tmp_945), .B(1), .Y(_25950_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48408_ ( .A(_tmp_25), .B(1), .Y(_25951_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48409_ ( .A(_tmp_957), .B(1), .Y(_25952_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48410_ ( .A(_tmp_32), .B(1), .Y(_25954_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48411_ ( .A(_tmp_33), .B(1), .Y(_25955_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48412_ ( .A(_tmp_853), .B(1), .Y(_25956_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48413_ ( .A(_tmp_1130), .B(1), .Y(_25957_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48414_ ( .A(_tmp_63), .B(1), .Y(_25958_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48415_ ( .A(_tmp_64), .B(1), .Y(_25959_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48416_ ( .A(_tmp_855), .B(1), .Y(_25960_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48417_ ( .A(_tmp_1142), .B(1), .Y(_25961_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48418_ ( .A(_tmp_94), .B(1), .Y(_25962_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48419_ ( .A(_tmp_95), .B(1), .Y(_25963_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48420_ ( .A(_tmp_857), .B(1), .Y(_25964_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48421_ ( .A(_tmp_1154), .B(1), .Y(_25965_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48422_ ( .A(_tmp_125), .B(1), .Y(_25966_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48423_ ( .A(_tmp_126), .B(1), .Y(_25967_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48424_ ( .A(req_block_size_27), .B(1), .Y(_25953_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48425_ ( .A(_tmp_859), .B(1), .Y(_25968_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48426_ ( .A(_tmp_1166), .B(1), .Y(_25969_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48427_ ( .A(_tmp_975), .B(1), .Y(_25970_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48428_ ( .A(_tmp_977), .B(1), .Y(_25971_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48429_ ( .A(_tmp_979), .B(1), .Y(_25972_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48430_ ( .A(_tmp_981), .B(1), .Y(_25973_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48431_ ( .A(_tmp_161), .B(1), .Y(_25975_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48432_ ( .A(_tmp_162), .B(1), .Y(_25976_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48433_ ( .A(_tmp_174), .B(1), .Y(_25977_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48434_ ( .A(_tmp_175), .B(1), .Y(_25978_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48435_ ( .A(_tmp_187), .B(1), .Y(_25979_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48436_ ( .A(_tmp_188), .B(1), .Y(_25980_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48437_ ( .A(_tmp_200), .B(1), .Y(_25981_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48438_ ( .A(_tmp_201), .B(1), .Y(_25982_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48439_ ( .A(req_block_size_156), .B(1), .Y(_25974_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48440_ ( .A(_tmp_218), .B(1), .Y(_25984_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48441_ ( .A(_tmp_219), .B(1), .Y(_25985_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48442_ ( .A(_tmp_231), .B(1), .Y(_25986_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48443_ ( .A(_tmp_232), .B(1), .Y(_25987_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48444_ ( .A(_tmp_244), .B(1), .Y(_25988_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48445_ ( .A(_tmp_245), .B(1), .Y(_25989_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48446_ ( .A(_tmp_257), .B(1), .Y(_25990_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48447_ ( .A(_tmp_258), .B(1), .Y(_25991_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48448_ ( .A(req_block_size_213), .B(1), .Y(_25983_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48449_ ( .A(_tmp_275), .B(1), .Y(_25993_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48450_ ( .A(_tmp_276), .B(1), .Y(_25994_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48451_ ( .A(_tmp_288), .B(1), .Y(_25995_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48452_ ( .A(_tmp_289), .B(1), .Y(_25996_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48453_ ( .A(_tmp_301), .B(1), .Y(_25997_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48454_ ( .A(_tmp_302), .B(1), .Y(_25998_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48455_ ( .A(_tmp_314), .B(1), .Y(_25999_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48456_ ( .A(_tmp_315), .B(1), .Y(_26000_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48457_ ( .A(req_block_size_270), .B(1), .Y(_25992_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48458_ ( .A(_tmp_810), .B(1), .Y(_26001_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48459_ ( .A(_tmp_822), .B(1), .Y(_26002_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48460_ ( .A(_tmp_834), .B(1), .Y(_26003_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48461_ ( .A(_maxi_write_size), .B(1), .Y(_25945_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48462_ ( .A(_tmp_846), .B(1), .Y(_26004_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48463_ ( .A(_maxi_read_local_addr), .B(_maxi_read_local_stride), .Y(_25939_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _48464_ ( .A(_tmp_12), .B(1), .Y(_26005_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(6), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(6) ) _48465_ ( .A(__variable_wdata_1), .B(2'h1), .Y(_26006_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48466_ ( .A(__variable_wdata_2), .B(1), .Y({ _21802_, _21801_, _21800_, _21798_, _21797_, _21796_, _21795_, _21794_, _21793_, _21792_, _21791_, _21790_, _21789_, _21787_, _21786_, _21785_, _21784_, _21783_, _21782_, _21781_, _21780_, _21779_, _21778_, _21809_, _21808_, _21807_, _21806_, _21805_, _21804_, _21803_, _21799_, _21788_, _21777_ }) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _48467_ ( .A(__variable_wdata_54), .B(2'h1), .Y(_26007_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _48468_ ( .A(__variable_wdata_69), .B(2'h1), .Y(_26008_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _48469_ ( .A(__variable_wdata_84), .B(2'h1), .Y(_26009_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _48470_ ( .A(__variable_wdata_99), .B(2'h1), .Y(_26010_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _48471_ ( .A(__variable_wdata_114), .B(2'h1), .Y(_26011_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _48472_ ( .A(__variable_wdata_129), .B(2'h1), .Y(_26012_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _48473_ ( .A(__variable_wdata_144), .B(2'h1), .Y(_26013_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _48474_ ( .A(__variable_wdata_159), .B(2'h1), .Y(_26014_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _48475_ ( .A(__variable_wdata_174), .B(2'h1), .Y(_26015_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48476_ ( .A(__variable_wdata_188), .B(1), .Y({ _21834_, _21833_, _21831_, _21830_, _21829_, _21828_, _21827_, _21826_, _21825_, _21824_, _21823_, _21822_, _21820_, _21819_, _21818_, _21817_, _21816_, _21815_, _21814_, _21813_, _21812_, _21811_, _21841_, _21840_, _21839_, _21838_, _21837_, _21836_, _21835_, _21832_, _21821_, _21810_ }) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48477_ ( .A(_source_stream_conv2d_8_source_6_pat_size_0), .B(1), .Y(_26016_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48478_ ( .A(_source_stream_conv2d_8_source_6_pat_size_1), .B(1), .Y(_26017_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48479_ ( .A(_source_stream_conv2d_8_source_6_pat_size_2), .B(1), .Y(_26018_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48480_ ( .A(_source_stream_conv2d_8_source_6_pat_size_3), .B(1), .Y(_26019_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48481_ ( .A(_source_stream_conv2d_8_source_6_pat_count_0), .B(1), .Y(_26020_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48482_ ( .A(_source_stream_conv2d_8_source_6_pat_size_buf_0), .B(1), .Y(_26021_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48483_ ( .A(_source_stream_conv2d_8_source_6_pat_count_1), .B(1), .Y(_26022_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48484_ ( .A(_source_stream_conv2d_8_source_6_pat_size_buf_1), .B(1), .Y(_26023_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48485_ ( .A(_source_stream_conv2d_8_source_6_pat_count_2), .B(1), .Y(_26024_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48486_ ( .A(_source_stream_conv2d_8_source_6_pat_size_buf_2), .B(1), .Y(_26025_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48487_ ( .A(_source_stream_conv2d_8_source_6_pat_count_3), .B(1), .Y(_26026_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48488_ ( .A(_source_stream_conv2d_8_source_6_pat_size_buf_3), .B(1), .Y(_26027_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48489_ ( .A(_source_stream_conv2d_8_source_8_pat_size_0), .B(1), .Y(_26028_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48490_ ( .A(_source_stream_conv2d_8_source_8_pat_size_1), .B(1), .Y(_26029_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48491_ ( .A(_source_stream_conv2d_8_source_8_pat_size_2), .B(1), .Y(_26030_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48492_ ( .A(_source_stream_conv2d_8_source_8_pat_size_3), .B(1), .Y(_26031_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48493_ ( .A(_source_stream_conv2d_8_source_8_pat_count_0), .B(1), .Y(_26032_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48494_ ( .A(_source_stream_conv2d_8_source_8_pat_size_buf_0), .B(1), .Y(_26033_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48495_ ( .A(_source_stream_conv2d_8_source_8_pat_count_1), .B(1), .Y(_26034_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48496_ ( .A(_source_stream_conv2d_8_source_8_pat_size_buf_1), .B(1), .Y(_26035_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48497_ ( .A(_source_stream_conv2d_8_source_8_pat_count_2), .B(1), .Y(_26036_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48498_ ( .A(_source_stream_conv2d_8_source_8_pat_size_buf_2), .B(1), .Y(_26037_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48499_ ( .A(_source_stream_conv2d_8_source_8_pat_count_3), .B(1), .Y(_26038_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48500_ ( .A(_source_stream_conv2d_8_source_8_pat_size_buf_3), .B(1), .Y(_26039_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48501_ ( .A(_source_stream_conv2d_8_source_19_pat_size_0), .B(1), .Y(_26040_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48502_ ( .A(_source_stream_conv2d_8_source_19_pat_size_1), .B(1), .Y(_26041_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48503_ ( .A(_source_stream_conv2d_8_source_19_pat_size_2), .B(1), .Y(_26042_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48504_ ( .A(_source_stream_conv2d_8_source_19_pat_size_3), .B(1), .Y(_26043_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48505_ ( .A(_source_stream_conv2d_8_source_19_pat_count_0), .B(1), .Y(_26044_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48506_ ( .A(_source_stream_conv2d_8_source_19_pat_size_buf_0), .B(1), .Y(_26045_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48507_ ( .A(_source_stream_conv2d_8_source_19_pat_count_1), .B(1), .Y(_26046_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48508_ ( .A(_source_stream_conv2d_8_source_19_pat_size_buf_1), .B(1), .Y(_26047_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48509_ ( .A(_source_stream_conv2d_8_source_19_pat_count_2), .B(1), .Y(_26048_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48510_ ( .A(_source_stream_conv2d_8_source_19_pat_size_buf_2), .B(1), .Y(_26049_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48511_ ( .A(_source_stream_conv2d_8_source_19_pat_count_3), .B(1), .Y(_26050_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48512_ ( .A(_source_stream_conv2d_8_source_19_pat_size_buf_3), .B(1), .Y(_26051_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48513_ ( .A(_source_stream_conv2d_8_source_20_pat_size_0), .B(1), .Y(_26052_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48514_ ( .A(_source_stream_conv2d_8_source_20_pat_size_1), .B(1), .Y(_26053_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48515_ ( .A(_source_stream_conv2d_8_source_20_pat_size_2), .B(1), .Y(_26054_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48516_ ( .A(_source_stream_conv2d_8_source_20_pat_size_3), .B(1), .Y(_26055_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48517_ ( .A(_source_stream_conv2d_8_source_20_pat_count_0), .B(1), .Y(_26056_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48518_ ( .A(_source_stream_conv2d_8_source_20_pat_size_buf_0), .B(1), .Y(_26057_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48519_ ( .A(_source_stream_conv2d_8_source_20_pat_count_1), .B(1), .Y(_26058_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48520_ ( .A(_source_stream_conv2d_8_source_20_pat_size_buf_1), .B(1), .Y(_26059_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48521_ ( .A(_source_stream_conv2d_8_source_20_pat_count_2), .B(1), .Y(_26060_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48522_ ( .A(_source_stream_conv2d_8_source_20_pat_size_buf_2), .B(1), .Y(_26061_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48523_ ( .A(_source_stream_conv2d_8_source_20_pat_count_3), .B(1), .Y(_26062_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48524_ ( .A(_source_stream_conv2d_8_source_20_pat_size_buf_3), .B(1), .Y(_26063_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48525_ ( .A(_source_stream_conv2d_8_source_21_pat_size_0), .B(1), .Y(_26064_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48526_ ( .A(_source_stream_conv2d_8_source_21_pat_size_1), .B(1), .Y(_26065_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48527_ ( .A(_source_stream_conv2d_8_source_21_pat_size_2), .B(1), .Y(_26066_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48528_ ( .A(_source_stream_conv2d_8_source_21_pat_size_3), .B(1), .Y(_26067_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48529_ ( .A(_source_stream_conv2d_8_source_21_pat_count_0), .B(1), .Y(_26068_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48530_ ( .A(_source_stream_conv2d_8_source_21_pat_size_buf_0), .B(1), .Y(_26069_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48531_ ( .A(_source_stream_conv2d_8_source_21_pat_count_1), .B(1), .Y(_26070_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48532_ ( .A(_source_stream_conv2d_8_source_21_pat_size_buf_1), .B(1), .Y(_26071_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48533_ ( .A(_source_stream_conv2d_8_source_21_pat_count_2), .B(1), .Y(_26072_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48534_ ( .A(_source_stream_conv2d_8_source_21_pat_size_buf_2), .B(1), .Y(_26073_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48535_ ( .A(_source_stream_conv2d_8_source_21_pat_count_3), .B(1), .Y(_26074_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48536_ ( .A(_source_stream_conv2d_8_source_21_pat_size_buf_3), .B(1), .Y(_26075_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48537_ ( .A(_source_stream_conv2d_8_source_22_pat_size_0), .B(1), .Y(_26076_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48538_ ( .A(_source_stream_conv2d_8_source_22_pat_size_1), .B(1), .Y(_26077_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48539_ ( .A(_source_stream_conv2d_8_source_22_pat_size_2), .B(1), .Y(_26078_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48540_ ( .A(_source_stream_conv2d_8_source_22_pat_size_3), .B(1), .Y(_26079_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48541_ ( .A(_source_stream_conv2d_8_source_22_pat_count_0), .B(1), .Y(_26080_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48542_ ( .A(_source_stream_conv2d_8_source_22_pat_size_buf_0), .B(1), .Y(_26081_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48543_ ( .A(_source_stream_conv2d_8_source_22_pat_count_1), .B(1), .Y(_26082_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48544_ ( .A(_source_stream_conv2d_8_source_22_pat_size_buf_1), .B(1), .Y(_26083_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48545_ ( .A(_source_stream_conv2d_8_source_22_pat_count_2), .B(1), .Y(_26084_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48546_ ( .A(_source_stream_conv2d_8_source_22_pat_size_buf_2), .B(1), .Y(_26085_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48547_ ( .A(_source_stream_conv2d_8_source_22_pat_count_3), .B(1), .Y(_26086_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48548_ ( .A(_source_stream_conv2d_8_source_22_pat_size_buf_3), .B(1), .Y(_26087_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48549_ ( .A(_source_stream_conv2d_8_source_23_pat_size_0), .B(1), .Y(_26088_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48550_ ( .A(_source_stream_conv2d_8_source_23_pat_size_1), .B(1), .Y(_26089_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48551_ ( .A(_source_stream_conv2d_8_source_23_pat_size_2), .B(1), .Y(_26090_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48552_ ( .A(_source_stream_conv2d_8_source_23_pat_size_3), .B(1), .Y(_26091_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48553_ ( .A(_source_stream_conv2d_8_source_23_pat_count_0), .B(1), .Y(_26092_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48554_ ( .A(_source_stream_conv2d_8_source_23_pat_size_buf_0), .B(1), .Y(_26093_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48555_ ( .A(_source_stream_conv2d_8_source_23_pat_count_1), .B(1), .Y(_26094_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48556_ ( .A(_source_stream_conv2d_8_source_23_pat_size_buf_1), .B(1), .Y(_26095_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48557_ ( .A(_source_stream_conv2d_8_source_23_pat_count_2), .B(1), .Y(_26096_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48558_ ( .A(_source_stream_conv2d_8_source_23_pat_size_buf_2), .B(1), .Y(_26097_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48559_ ( .A(_source_stream_conv2d_8_source_23_pat_count_3), .B(1), .Y(_26098_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48560_ ( .A(_source_stream_conv2d_8_source_23_pat_size_buf_3), .B(1), .Y(_26099_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48561_ ( .A(_source_stream_conv2d_8_source_24_pat_size_0), .B(1), .Y(_26100_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48562_ ( .A(_source_stream_conv2d_8_source_24_pat_size_1), .B(1), .Y(_26101_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48563_ ( .A(_source_stream_conv2d_8_source_24_pat_size_2), .B(1), .Y(_26102_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48564_ ( .A(_source_stream_conv2d_8_source_24_pat_size_3), .B(1), .Y(_26103_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48565_ ( .A(_source_stream_conv2d_8_source_24_pat_count_0), .B(1), .Y(_26104_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48566_ ( .A(_source_stream_conv2d_8_source_24_pat_size_buf_0), .B(1), .Y(_26105_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48567_ ( .A(_source_stream_conv2d_8_source_24_pat_count_1), .B(1), .Y(_26106_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48568_ ( .A(_source_stream_conv2d_8_source_24_pat_size_buf_1), .B(1), .Y(_26107_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48569_ ( .A(_source_stream_conv2d_8_source_24_pat_count_2), .B(1), .Y(_26108_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48570_ ( .A(_source_stream_conv2d_8_source_24_pat_size_buf_2), .B(1), .Y(_26109_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48571_ ( .A(_source_stream_conv2d_8_source_24_pat_count_3), .B(1), .Y(_26110_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48572_ ( .A(_source_stream_conv2d_8_source_24_pat_size_buf_3), .B(1), .Y(_26111_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48573_ ( .A(_source_stream_conv2d_8_source_25_pat_size_0), .B(1), .Y(_26112_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48574_ ( .A(_source_stream_conv2d_8_source_25_pat_size_1), .B(1), .Y(_26113_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48575_ ( .A(_source_stream_conv2d_8_source_25_pat_size_2), .B(1), .Y(_26114_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48576_ ( .A(_source_stream_conv2d_8_source_25_pat_size_3), .B(1), .Y(_26115_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48577_ ( .A(_source_stream_conv2d_8_source_25_pat_count_0), .B(1), .Y(_26116_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48578_ ( .A(_source_stream_conv2d_8_source_25_pat_size_buf_0), .B(1), .Y(_26117_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48579_ ( .A(_source_stream_conv2d_8_source_25_pat_count_1), .B(1), .Y(_26118_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48580_ ( .A(_source_stream_conv2d_8_source_25_pat_size_buf_1), .B(1), .Y(_26119_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48581_ ( .A(_source_stream_conv2d_8_source_25_pat_count_2), .B(1), .Y(_26120_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48582_ ( .A(_source_stream_conv2d_8_source_25_pat_size_buf_2), .B(1), .Y(_26121_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48583_ ( .A(_source_stream_conv2d_8_source_25_pat_count_3), .B(1), .Y(_26122_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48584_ ( .A(_source_stream_conv2d_8_source_25_pat_size_buf_3), .B(1), .Y(_26123_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48585_ ( .A(_source_stream_conv2d_8_source_26_pat_size_0), .B(1), .Y(_26124_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48586_ ( .A(_source_stream_conv2d_8_source_26_pat_size_1), .B(1), .Y(_26125_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48587_ ( .A(_source_stream_conv2d_8_source_26_pat_size_2), .B(1), .Y(_26126_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48588_ ( .A(_source_stream_conv2d_8_source_26_pat_size_3), .B(1), .Y(_26127_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48589_ ( .A(_source_stream_conv2d_8_source_26_pat_count_0), .B(1), .Y(_26128_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48590_ ( .A(_source_stream_conv2d_8_source_26_pat_size_buf_0), .B(1), .Y(_26129_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48591_ ( .A(_source_stream_conv2d_8_source_26_pat_count_1), .B(1), .Y(_26130_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48592_ ( .A(_source_stream_conv2d_8_source_26_pat_size_buf_1), .B(1), .Y(_26131_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48593_ ( .A(_source_stream_conv2d_8_source_26_pat_count_2), .B(1), .Y(_26132_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48594_ ( .A(_source_stream_conv2d_8_source_26_pat_size_buf_2), .B(1), .Y(_26133_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48595_ ( .A(_source_stream_conv2d_8_source_26_pat_count_3), .B(1), .Y(_26134_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48596_ ( .A(_source_stream_conv2d_8_source_26_pat_size_buf_3), .B(1), .Y(_26135_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48597_ ( .A(_source_stream_conv2d_8_source_27_pat_size_0), .B(1), .Y(_26136_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48598_ ( .A(_source_stream_conv2d_8_source_27_pat_size_1), .B(1), .Y(_26137_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48599_ ( .A(_source_stream_conv2d_8_source_27_pat_size_2), .B(1), .Y(_26138_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48600_ ( .A(_source_stream_conv2d_8_source_27_pat_size_3), .B(1), .Y(_26139_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48601_ ( .A(_source_stream_conv2d_8_source_27_pat_count_0), .B(1), .Y(_26140_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48602_ ( .A(_source_stream_conv2d_8_source_27_pat_size_buf_0), .B(1), .Y(_26141_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48603_ ( .A(_source_stream_conv2d_8_source_27_pat_count_1), .B(1), .Y(_26142_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48604_ ( .A(_source_stream_conv2d_8_source_27_pat_size_buf_1), .B(1), .Y(_26143_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48605_ ( .A(_source_stream_conv2d_8_source_27_pat_count_2), .B(1), .Y(_26144_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48606_ ( .A(_source_stream_conv2d_8_source_27_pat_size_buf_2), .B(1), .Y(_26145_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48607_ ( .A(_source_stream_conv2d_8_source_27_pat_count_3), .B(1), .Y(_26146_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48608_ ( .A(_source_stream_conv2d_8_source_27_pat_size_buf_3), .B(1), .Y(_26147_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48609_ ( .A(_source_stream_conv2d_8_source_28_pat_size_0), .B(1), .Y(_26148_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48610_ ( .A(_source_stream_conv2d_8_source_28_pat_size_1), .B(1), .Y(_26149_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48611_ ( .A(_source_stream_conv2d_8_source_28_pat_size_2), .B(1), .Y(_26150_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48612_ ( .A(_source_stream_conv2d_8_source_28_pat_size_3), .B(1), .Y(_26151_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48613_ ( .A(_source_stream_conv2d_8_source_28_pat_count_0), .B(1), .Y(_26152_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48614_ ( .A(_source_stream_conv2d_8_source_28_pat_size_buf_0), .B(1), .Y(_26153_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48615_ ( .A(_source_stream_conv2d_8_source_28_pat_count_1), .B(1), .Y(_26154_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48616_ ( .A(_source_stream_conv2d_8_source_28_pat_size_buf_1), .B(1), .Y(_26155_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48617_ ( .A(_source_stream_conv2d_8_source_28_pat_count_2), .B(1), .Y(_26156_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48618_ ( .A(_source_stream_conv2d_8_source_28_pat_size_buf_2), .B(1), .Y(_26157_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48619_ ( .A(_source_stream_conv2d_8_source_28_pat_count_3), .B(1), .Y(_26158_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48620_ ( .A(_source_stream_conv2d_8_source_28_pat_size_buf_3), .B(1), .Y(_26159_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48621_ ( .A(_source_stream_conv2d_8_source_29_pat_size_0), .B(1), .Y(_26160_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48622_ ( .A(_source_stream_conv2d_8_source_29_pat_size_1), .B(1), .Y(_26161_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48623_ ( .A(_source_stream_conv2d_8_source_29_pat_size_2), .B(1), .Y(_26162_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48624_ ( .A(_source_stream_conv2d_8_source_29_pat_size_3), .B(1), .Y(_26163_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48625_ ( .A(_source_stream_conv2d_8_source_29_pat_count_0), .B(1), .Y(_26164_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48626_ ( .A(_source_stream_conv2d_8_source_29_pat_size_buf_0), .B(1), .Y(_26165_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48627_ ( .A(_source_stream_conv2d_8_source_29_pat_count_1), .B(1), .Y(_26166_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48628_ ( .A(_source_stream_conv2d_8_source_29_pat_size_buf_1), .B(1), .Y(_26167_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48629_ ( .A(_source_stream_conv2d_8_source_29_pat_count_2), .B(1), .Y(_26168_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48630_ ( .A(_source_stream_conv2d_8_source_29_pat_size_buf_2), .B(1), .Y(_26169_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48631_ ( .A(_source_stream_conv2d_8_source_29_pat_count_3), .B(1), .Y(_26170_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48632_ ( .A(_source_stream_conv2d_8_source_29_pat_size_buf_3), .B(1), .Y(_26171_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48633_ ( .A(_source_stream_conv2d_8_source_30_pat_size_0), .B(1), .Y(_26172_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48634_ ( .A(_source_stream_conv2d_8_source_30_pat_size_1), .B(1), .Y(_26173_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48635_ ( .A(_source_stream_conv2d_8_source_30_pat_size_2), .B(1), .Y(_26174_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48636_ ( .A(_source_stream_conv2d_8_source_30_pat_size_3), .B(1), .Y(_26175_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48637_ ( .A(_source_stream_conv2d_8_source_30_pat_count_0), .B(1), .Y(_26176_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48638_ ( .A(_source_stream_conv2d_8_source_30_pat_size_buf_0), .B(1), .Y(_26177_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48639_ ( .A(_source_stream_conv2d_8_source_30_pat_count_1), .B(1), .Y(_26178_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48640_ ( .A(_source_stream_conv2d_8_source_30_pat_size_buf_1), .B(1), .Y(_26179_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48641_ ( .A(_source_stream_conv2d_8_source_30_pat_count_2), .B(1), .Y(_26180_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48642_ ( .A(_source_stream_conv2d_8_source_30_pat_size_buf_2), .B(1), .Y(_26181_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48643_ ( .A(_source_stream_conv2d_8_source_30_pat_count_3), .B(1), .Y(_26182_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48644_ ( .A(_source_stream_conv2d_8_source_30_pat_size_buf_3), .B(1), .Y(_26183_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48645_ ( .A(_source_stream_conv2d_8_source_31_pat_size_0), .B(1), .Y(_26184_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48646_ ( .A(_source_stream_conv2d_8_source_31_pat_size_1), .B(1), .Y(_26185_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48647_ ( .A(_source_stream_conv2d_8_source_31_pat_size_2), .B(1), .Y(_26186_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48648_ ( .A(_source_stream_conv2d_8_source_31_pat_size_3), .B(1), .Y(_26187_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48649_ ( .A(_source_stream_conv2d_8_source_31_pat_count_0), .B(1), .Y(_26188_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48650_ ( .A(_source_stream_conv2d_8_source_31_pat_size_buf_0), .B(1), .Y(_26189_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48651_ ( .A(_source_stream_conv2d_8_source_31_pat_count_1), .B(1), .Y(_26190_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48652_ ( .A(_source_stream_conv2d_8_source_31_pat_size_buf_1), .B(1), .Y(_26191_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48653_ ( .A(_source_stream_conv2d_8_source_31_pat_count_2), .B(1), .Y(_26192_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48654_ ( .A(_source_stream_conv2d_8_source_31_pat_size_buf_2), .B(1), .Y(_26193_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48655_ ( .A(_source_stream_conv2d_8_source_31_pat_count_3), .B(1), .Y(_26194_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48656_ ( .A(_source_stream_conv2d_8_source_31_pat_size_buf_3), .B(1), .Y(_26195_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48657_ ( .A(_source_stream_conv2d_8_source_32_pat_size_0), .B(1), .Y(_26196_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48658_ ( .A(_source_stream_conv2d_8_source_32_pat_size_1), .B(1), .Y(_26197_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48659_ ( .A(_source_stream_conv2d_8_source_32_pat_size_2), .B(1), .Y(_26198_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48660_ ( .A(_source_stream_conv2d_8_source_32_pat_size_3), .B(1), .Y(_26199_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48661_ ( .A(_source_stream_conv2d_8_source_32_pat_count_0), .B(1), .Y(_26200_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48662_ ( .A(_source_stream_conv2d_8_source_32_pat_size_buf_0), .B(1), .Y(_26201_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48663_ ( .A(_source_stream_conv2d_8_source_32_pat_count_1), .B(1), .Y(_26202_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48664_ ( .A(_source_stream_conv2d_8_source_32_pat_size_buf_1), .B(1), .Y(_26203_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48665_ ( .A(_source_stream_conv2d_8_source_32_pat_count_2), .B(1), .Y(_26204_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48666_ ( .A(_source_stream_conv2d_8_source_32_pat_size_buf_2), .B(1), .Y(_26205_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48667_ ( .A(_source_stream_conv2d_8_source_32_pat_count_3), .B(1), .Y(_26206_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48668_ ( .A(_source_stream_conv2d_8_source_32_pat_size_buf_3), .B(1), .Y(_26207_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48669_ ( .A(_source_stream_conv2d_8_source_33_pat_size_0), .B(1), .Y(_26208_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48670_ ( .A(_source_stream_conv2d_8_source_33_pat_size_1), .B(1), .Y(_26209_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48671_ ( .A(_source_stream_conv2d_8_source_33_pat_size_2), .B(1), .Y(_26210_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48672_ ( .A(_source_stream_conv2d_8_source_33_pat_size_3), .B(1), .Y(_26211_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48673_ ( .A(_source_stream_conv2d_8_source_33_pat_count_0), .B(1), .Y(_26212_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48674_ ( .A(_source_stream_conv2d_8_source_33_pat_size_buf_0), .B(1), .Y(_26213_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48675_ ( .A(_source_stream_conv2d_8_source_33_pat_count_1), .B(1), .Y(_26214_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48676_ ( .A(_source_stream_conv2d_8_source_33_pat_size_buf_1), .B(1), .Y(_26215_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48677_ ( .A(_source_stream_conv2d_8_source_33_pat_count_2), .B(1), .Y(_26216_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48678_ ( .A(_source_stream_conv2d_8_source_33_pat_size_buf_2), .B(1), .Y(_26217_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48679_ ( .A(_source_stream_conv2d_8_source_33_pat_count_3), .B(1), .Y(_26218_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48680_ ( .A(_source_stream_conv2d_8_source_33_pat_size_buf_3), .B(1), .Y(_26219_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48681_ ( .A(_source_stream_conv2d_8_source_34_pat_size_0), .B(1), .Y(_26220_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48682_ ( .A(_source_stream_conv2d_8_source_34_pat_size_1), .B(1), .Y(_26221_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48683_ ( .A(_source_stream_conv2d_8_source_34_pat_size_2), .B(1), .Y(_26222_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48684_ ( .A(_source_stream_conv2d_8_source_34_pat_size_3), .B(1), .Y(_26223_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48685_ ( .A(_source_stream_conv2d_8_source_34_pat_count_0), .B(1), .Y(_26224_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48686_ ( .A(_source_stream_conv2d_8_source_34_pat_size_buf_0), .B(1), .Y(_26225_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48687_ ( .A(_source_stream_conv2d_8_source_34_pat_count_1), .B(1), .Y(_26226_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48688_ ( .A(_source_stream_conv2d_8_source_34_pat_size_buf_1), .B(1), .Y(_26227_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48689_ ( .A(_source_stream_conv2d_8_source_34_pat_count_2), .B(1), .Y(_26228_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48690_ ( .A(_source_stream_conv2d_8_source_34_pat_size_buf_2), .B(1), .Y(_26229_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48691_ ( .A(_source_stream_conv2d_8_source_34_pat_count_3), .B(1), .Y(_26230_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48692_ ( .A(_source_stream_conv2d_8_source_34_pat_size_buf_3), .B(1), .Y(_26231_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48693_ ( .A(_source_stream_conv2d_8_source_35_pat_size_0), .B(1), .Y(_26232_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48694_ ( .A(_source_stream_conv2d_8_source_35_pat_size_1), .B(1), .Y(_26233_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48695_ ( .A(_source_stream_conv2d_8_source_35_pat_size_2), .B(1), .Y(_26234_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48696_ ( .A(_source_stream_conv2d_8_source_35_pat_size_3), .B(1), .Y(_26235_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48697_ ( .A(_source_stream_conv2d_8_source_35_pat_count_0), .B(1), .Y(_26236_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48698_ ( .A(_source_stream_conv2d_8_source_35_pat_size_buf_0), .B(1), .Y(_26237_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48699_ ( .A(_source_stream_conv2d_8_source_35_pat_count_1), .B(1), .Y(_26238_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48700_ ( .A(_source_stream_conv2d_8_source_35_pat_size_buf_1), .B(1), .Y(_26239_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48701_ ( .A(_source_stream_conv2d_8_source_35_pat_count_2), .B(1), .Y(_26240_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48702_ ( .A(_source_stream_conv2d_8_source_35_pat_size_buf_2), .B(1), .Y(_26241_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48703_ ( .A(_source_stream_conv2d_8_source_35_pat_count_3), .B(1), .Y(_26242_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48704_ ( .A(_source_stream_conv2d_8_source_35_pat_size_buf_3), .B(1), .Y(_26243_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48705_ ( .A(_source_stream_conv2d_8_source_36_pat_size_0), .B(1), .Y(_26244_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48706_ ( .A(_source_stream_conv2d_8_source_36_pat_size_1), .B(1), .Y(_26245_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48707_ ( .A(_source_stream_conv2d_8_source_36_pat_size_2), .B(1), .Y(_26246_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48708_ ( .A(_source_stream_conv2d_8_source_36_pat_size_3), .B(1), .Y(_26247_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48709_ ( .A(_source_stream_conv2d_8_source_36_pat_count_0), .B(1), .Y(_26248_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48710_ ( .A(_source_stream_conv2d_8_source_36_pat_size_buf_0), .B(1), .Y(_26249_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48711_ ( .A(_source_stream_conv2d_8_source_36_pat_count_1), .B(1), .Y(_26250_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48712_ ( .A(_source_stream_conv2d_8_source_36_pat_size_buf_1), .B(1), .Y(_26251_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48713_ ( .A(_source_stream_conv2d_8_source_36_pat_count_2), .B(1), .Y(_26252_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48714_ ( .A(_source_stream_conv2d_8_source_36_pat_size_buf_2), .B(1), .Y(_26253_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48715_ ( .A(_source_stream_conv2d_8_source_36_pat_count_3), .B(1), .Y(_26254_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48716_ ( .A(_source_stream_conv2d_8_source_36_pat_size_buf_3), .B(1), .Y(_26255_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48717_ ( .A(_stream_conv2d_8_sink_37_sink_offset), .B(_stream_conv2d_8_sink_37_sink_stride), .Y(_26256_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48718_ ( .A(_stream_conv2d_8_sink_37_sink_count), .B(1), .Y(_26257_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(3), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48719_ ( .A(__variable_wdata_757), .B(1), .Y({ _21866_, _21865_, _21863_, _21862_, _21861_, _21860_, _21859_, _21858_, _21857_, _21856_, _21855_, _21854_, _21852_, _21851_, _21850_, _21849_, _21848_, _21847_, _21846_, _21845_, _21844_, _21843_, _21873_, _21872_, _21871_, _21870_, _21869_, _21868_, _21867_, _21864_, _21853_, _21842_ }) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48720_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_0), .B(1), .Y(_26258_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48721_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_1), .B(1), .Y(_26259_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48722_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_2), .B(1), .Y(_26260_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48723_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_3), .B(1), .Y(_26261_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48724_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_0), .B(1), .Y(_26262_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48725_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_buf_0), .B(1), .Y(_26263_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48726_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_1), .B(1), .Y(_26264_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48727_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_buf_1), .B(1), .Y(_26265_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48728_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_2), .B(1), .Y(_26266_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48729_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_buf_2), .B(1), .Y(_26267_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48730_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_3), .B(1), .Y(_26268_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48731_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_buf_3), .B(1), .Y(_26269_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48732_ ( .A(_stream_max_pool_serial_9_sink_3_sink_offset), .B(_stream_max_pool_serial_9_sink_3_sink_stride), .Y(_26270_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48733_ ( .A(_stream_max_pool_serial_9_sink_3_sink_count), .B(1), .Y(_26271_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48734_ ( .A(_source_stream_matmul_15_source_6_pat_size_0), .B(1), .Y(_26272_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48735_ ( .A(_source_stream_matmul_15_source_6_pat_size_1), .B(1), .Y(_26273_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48736_ ( .A(_source_stream_matmul_15_source_6_pat_size_2), .B(1), .Y(_26274_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48737_ ( .A(_source_stream_matmul_15_source_6_pat_size_3), .B(1), .Y(_26275_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48738_ ( .A(_source_stream_matmul_15_source_6_pat_count_0), .B(1), .Y(_26276_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48739_ ( .A(_source_stream_matmul_15_source_6_pat_size_buf_0), .B(1), .Y(_26277_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48740_ ( .A(_source_stream_matmul_15_source_6_pat_count_1), .B(1), .Y(_26278_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48741_ ( .A(_source_stream_matmul_15_source_6_pat_size_buf_1), .B(1), .Y(_26279_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48742_ ( .A(_source_stream_matmul_15_source_6_pat_count_2), .B(1), .Y(_26280_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48743_ ( .A(_source_stream_matmul_15_source_6_pat_size_buf_2), .B(1), .Y(_26281_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48744_ ( .A(_source_stream_matmul_15_source_6_pat_count_3), .B(1), .Y(_26282_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48745_ ( .A(_source_stream_matmul_15_source_6_pat_size_buf_3), .B(1), .Y(_26283_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48746_ ( .A(_source_stream_matmul_15_source_8_pat_size_0), .B(1), .Y(_26284_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48747_ ( .A(_source_stream_matmul_15_source_8_pat_size_1), .B(1), .Y(_26285_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48748_ ( .A(_source_stream_matmul_15_source_8_pat_size_2), .B(1), .Y(_26286_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48749_ ( .A(_source_stream_matmul_15_source_8_pat_size_3), .B(1), .Y(_26287_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48750_ ( .A(_source_stream_matmul_15_source_8_pat_count_0), .B(1), .Y(_26288_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48751_ ( .A(_source_stream_matmul_15_source_8_pat_size_buf_0), .B(1), .Y(_26289_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48752_ ( .A(_source_stream_matmul_15_source_8_pat_count_1), .B(1), .Y(_26290_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48753_ ( .A(_source_stream_matmul_15_source_8_pat_size_buf_1), .B(1), .Y(_26291_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48754_ ( .A(_source_stream_matmul_15_source_8_pat_count_2), .B(1), .Y(_26292_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48755_ ( .A(_source_stream_matmul_15_source_8_pat_size_buf_2), .B(1), .Y(_26293_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48756_ ( .A(_source_stream_matmul_15_source_8_pat_count_3), .B(1), .Y(_26294_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48757_ ( .A(_source_stream_matmul_15_source_8_pat_size_buf_3), .B(1), .Y(_26295_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48758_ ( .A(_source_stream_matmul_15_source_19_pat_size_0), .B(1), .Y(_26296_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48759_ ( .A(_source_stream_matmul_15_source_19_pat_size_1), .B(1), .Y(_26297_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48760_ ( .A(_source_stream_matmul_15_source_19_pat_size_2), .B(1), .Y(_26298_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48761_ ( .A(_source_stream_matmul_15_source_19_pat_size_3), .B(1), .Y(_26299_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48762_ ( .A(_source_stream_matmul_15_source_19_pat_count_0), .B(1), .Y(_26300_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48763_ ( .A(_source_stream_matmul_15_source_19_pat_size_buf_0), .B(1), .Y(_26301_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48764_ ( .A(_source_stream_matmul_15_source_19_pat_count_1), .B(1), .Y(_26302_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48765_ ( .A(_source_stream_matmul_15_source_19_pat_size_buf_1), .B(1), .Y(_26303_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48766_ ( .A(_source_stream_matmul_15_source_19_pat_count_2), .B(1), .Y(_26304_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48767_ ( .A(_source_stream_matmul_15_source_19_pat_size_buf_2), .B(1), .Y(_26305_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48768_ ( .A(_source_stream_matmul_15_source_19_pat_count_3), .B(1), .Y(_26306_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48769_ ( .A(_source_stream_matmul_15_source_19_pat_size_buf_3), .B(1), .Y(_26307_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48770_ ( .A(_source_stream_matmul_15_source_20_pat_size_0), .B(1), .Y(_26308_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48771_ ( .A(_source_stream_matmul_15_source_20_pat_size_1), .B(1), .Y(_26309_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48772_ ( .A(_source_stream_matmul_15_source_20_pat_size_2), .B(1), .Y(_26310_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48773_ ( .A(_source_stream_matmul_15_source_20_pat_size_3), .B(1), .Y(_26311_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48774_ ( .A(_source_stream_matmul_15_source_20_pat_count_0), .B(1), .Y(_26312_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48775_ ( .A(_source_stream_matmul_15_source_20_pat_size_buf_0), .B(1), .Y(_26313_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48776_ ( .A(_source_stream_matmul_15_source_20_pat_count_1), .B(1), .Y(_26314_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48777_ ( .A(_source_stream_matmul_15_source_20_pat_size_buf_1), .B(1), .Y(_26315_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48778_ ( .A(_source_stream_matmul_15_source_20_pat_count_2), .B(1), .Y(_26316_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48779_ ( .A(_source_stream_matmul_15_source_20_pat_size_buf_2), .B(1), .Y(_26317_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48780_ ( .A(_source_stream_matmul_15_source_20_pat_count_3), .B(1), .Y(_26318_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48781_ ( .A(_source_stream_matmul_15_source_20_pat_size_buf_3), .B(1), .Y(_26319_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48782_ ( .A(_stream_matmul_15_sink_21_sink_offset), .B(_stream_matmul_15_sink_21_sink_stride), .Y(_26320_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48783_ ( .A(_stream_matmul_15_sink_21_sink_count), .B(1), .Y(_26321_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _48784_ ( .A(conv2d_8_row_select), .B(2), .Y(_26322_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _48785_ ( .A(4096), .B({ 21'h000000, _maxi_read_cur_global_addr[11:0] }), .Y({ _25922_[30:0], _26323_[1:0] }) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _48786_ ( .A(_maxi_read_rest_size), .B({ 2'h0, _25922_[30:0] }), .Y(_26324_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48787_ ( .A(_maxi_read_rest_size), .B(256), .Y(_26325_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(2) ) _48788_ ( .A(conv2d_8_col_select), .B(2'h2), .Y(_26326_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _48789_ ( .A(4096), .B({ 21'h000000, _maxi_write_cur_global_addr[11:0] }), .Y({ _25923_[30:0], _26327_[1:0] }) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _48790_ ( .A(_maxi_write_rest_size), .B({ 2'h0, _25923_[30:0] }), .Y(_26328_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _48791_ ( .A(_maxi_write_rest_size), .B(256), .Y(_26329_) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(16) ) _49074_ ( .A(\__muladd_madd_110.madd._a ), .B(\__muladd_madd_110.madd._b ), .Y(\__muladd_madd_110.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(16) ) _49081_ ( .A(\__muladd_madd_125.madd._a ), .B(\__muladd_madd_125.madd._b ), .Y(\__muladd_madd_125.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(16) ) _49088_ ( .A(\__muladd_madd_140.madd._a ), .B(\__muladd_madd_140.madd._b ), .Y(\__muladd_madd_140.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(16) ) _49095_ ( .A(\__muladd_madd_155.madd._a ), .B(\__muladd_madd_155.madd._b ), .Y(\__muladd_madd_155.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(16) ) _49102_ ( .A(\__muladd_madd_170.madd._a ), .B(\__muladd_madd_170.madd._b ), .Y(\__muladd_madd_170.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(16) ) _49109_ ( .A(\__muladd_madd_185.madd._a ), .B(\__muladd_madd_185.madd._b ), .Y(\__muladd_madd_185.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(16) ) _49116_ ( .A(\__muladd_madd_65.madd._a ), .B(\__muladd_madd_65.madd._b ), .Y(\__muladd_madd_65.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(16) ) _49123_ ( .A(\__muladd_madd_80.madd._a ), .B(\__muladd_madd_80.madd._b ), .Y(\__muladd_madd_80.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(16) ) _49130_ ( .A(\__muladd_madd_95.madd._a ), .B(\__muladd_madd_95.madd._b ), .Y(\__muladd_madd_95.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(40) ) _49136_ ( .A(\_times_mul_39.mult._a ), .B(\_times_mul_39.mult._b ), .Y(\_times_mul_39.mult._mul ) );
  \$mux  #( .WIDTH(32) ) _41323_ ( .A(_stream_matmul_15_sink_21_sink_fsm_4), .B(0), .S(_05862_), .Y(_22455_) );
  \$mux  #( .WIDTH(32) ) _41324_ ( .A(_22455_), .B(0), .S(_stream_matmul_15_term_sink), .Y({ _11342_, _11341_, _11339_, _11338_, _11337_, _11336_, _11335_, _11334_, _11333_, _11332_, _11331_, _11330_, _11328_, _11327_, _11326_, _11325_, _11324_, _11323_, _11322_, _11321_, _11320_, _11319_, _11349_, _11348_, _11347_, _11346_, _11345_, _11344_, _11343_, _11340_, _11329_, _11318_ }) );
  \$mux  #( .WIDTH(32) ) _41325_ ( .A(_stream_matmul_15_sink_21_sink_fsm_4), .B(1), .S(_05803_), .Y({ _11406_, _11405_, _11403_, _11402_, _11401_, _11400_, _11399_, _11398_, _11397_, _11396_, _11395_, _11394_, _11392_, _11391_, _11390_, _11389_, _11388_, _11387_, _11386_, _11385_, _11384_, _11383_, _11413_, _11412_, _11411_, _11410_, _11409_, _11408_, _11407_, _11404_, _11393_, _11382_ }) );
  \$mux  #( .WIDTH(32) ) _41327_ ( .A(_stream_matmul_15_source_20_source_pat_fsm_3), .B(2), .S(_05861_), .Y({ _11470_, _11469_, _11467_, _11466_, _11465_, _11464_, _11463_, _11462_, _11461_, _11460_, _11459_, _11458_, _11456_, _11455_, _11454_, _11453_, _11452_, _11451_, _11450_, _11449_, _11448_, _11447_, _11477_, _11476_, _11475_, _11474_, _11473_, _11472_, _11471_, _11468_, _11457_, _11446_ }) );
  \$mux  #( .WIDTH(32) ) _41328_ ( .A(_stream_matmul_15_source_20_source_pat_fsm_3), .B(1), .S(_05798_), .Y({ _11502_, _11501_, _11499_, _11498_, _11497_, _11496_, _11495_, _11494_, _11493_, _11492_, _11491_, _11490_, _11488_, _11487_, _11486_, _11485_, _11484_, _11483_, _11482_, _11481_, _11480_, _11479_, _11509_, _11508_, _11507_, _11506_, _11505_, _11504_, _11503_, _11500_, _11489_, _11478_ }) );
  \$mux  #( .WIDTH(32) ) _41332_ ( .A(_stream_matmul_15_source_19_source_pat_fsm_2), .B(2), .S(_05860_), .Y({ _11566_, _11565_, _11563_, _11562_, _11561_, _11560_, _11559_, _11558_, _11557_, _11556_, _11555_, _11554_, _11552_, _11551_, _11550_, _11549_, _11548_, _11547_, _11546_, _11545_, _11544_, _11543_, _11573_, _11572_, _11571_, _11570_, _11569_, _11568_, _11567_, _11564_, _11553_, _11542_ }) );
  \$mux  #( .WIDTH(32) ) _41333_ ( .A(_stream_matmul_15_source_19_source_pat_fsm_2), .B(1), .S(_05793_), .Y({ _11598_, _11597_, _11595_, _11594_, _11593_, _11592_, _11591_, _11590_, _11589_, _11588_, _11587_, _11586_, _11584_, _11583_, _11582_, _11581_, _11580_, _11579_, _11578_, _11577_, _11576_, _11575_, _11605_, _11604_, _11603_, _11602_, _11601_, _11600_, _11599_, _11596_, _11585_, _11574_ }) );
  \$mux  #( .WIDTH(32) ) _41335_ ( .A(_stream_matmul_15_source_8_source_pat_fsm_1), .B(2), .S(_05859_), .Y({ _11662_, _11661_, _11659_, _11658_, _11657_, _11656_, _11655_, _11654_, _11653_, _11652_, _11651_, _11650_, _11648_, _11647_, _11646_, _11645_, _11644_, _11643_, _11642_, _11641_, _11640_, _11639_, _11669_, _11668_, _11667_, _11666_, _11665_, _11664_, _11663_, _11660_, _11649_, _11638_ }) );
  \$mux  #( .WIDTH(32) ) _41336_ ( .A(_stream_matmul_15_source_8_source_pat_fsm_1), .B(1), .S(_05788_), .Y({ _11694_, _11693_, _11691_, _11690_, _11689_, _11688_, _11687_, _11686_, _11685_, _11684_, _11683_, _11682_, _11680_, _11679_, _11678_, _11677_, _11676_, _11675_, _11674_, _11673_, _11672_, _11671_, _11701_, _11700_, _11699_, _11698_, _11697_, _11696_, _11695_, _11692_, _11681_, _11670_ }) );
  \$mux  #( .WIDTH(32) ) _41338_ ( .A(_stream_matmul_15_source_6_source_pat_fsm_0), .B(2), .S(_05858_), .Y({ _11758_, _11757_, _11755_, _11754_, _11753_, _11752_, _11751_, _11750_, _11749_, _11748_, _11747_, _11746_, _11744_, _11743_, _11742_, _11741_, _11740_, _11739_, _11738_, _11737_, _11736_, _11735_, _11765_, _11764_, _11763_, _11762_, _11761_, _11760_, _11759_, _11756_, _11745_, _11734_ }) );
  \$mux  #( .WIDTH(32) ) _41339_ ( .A(_stream_matmul_15_source_6_source_pat_fsm_0), .B(1), .S(_05783_), .Y({ _11790_, _11789_, _11787_, _11786_, _11785_, _11784_, _11783_, _11782_, _11781_, _11780_, _11779_, _11778_, _11776_, _11775_, _11774_, _11773_, _11772_, _11771_, _11770_, _11769_, _11768_, _11767_, _11797_, _11796_, _11795_, _11794_, _11793_, _11792_, _11791_, _11788_, _11777_, _11766_ }) );
  \$mux  #( .WIDTH(1) ) _41341_ ( .A(matmul_15_stream_pad_mask_0_0), .B(matmul_15_stream_pad_masks), .S(_05028_), .Y(_22461_) );
  \$mux  #( .WIDTH(32) ) _41343_ ( .A(matmul_15_och_count), .B(matmul_15_och_count_buf), .S(_05030_), .Y(_22462_) );
  \$mux  #( .WIDTH(1) ) _41345_ ( .A(matmul_15_row_select), .B(matmul_15_row_select_buf), .S(_05030_), .Y(_22463_) );
  \$mux  #( .WIDTH(32) ) _41347_ ( .A(matmul_15_row_count), .B(matmul_15_row_count_buf), .S(_05030_), .Y(_22464_) );
  \$mux  #( .WIDTH(32) ) _41349_ ( .A(matmul_15_out_page_comp_offset), .B(matmul_15_out_page_comp_offset_buf), .S(_05030_), .Y(_22465_) );
  \$mux  #( .WIDTH(32) ) _41351_ ( .A(matmul_15_act_page_comp_offset_0), .B(matmul_15_act_page_comp_offset_buf_0), .S(_05030_), .Y(_22466_) );
  \$mux  #( .WIDTH(32) ) _41353_ ( .A(matmul_15_filter_page_comp_offset), .B(matmul_15_filter_page_comp_offset_buf), .S(_05030_), .Y(_22467_) );
  \$mux  #( .WIDTH(32) ) _41355_ ( .A(5), .B(matmul_15_comp_fsm), .S(_stream_matmul_15_source_busy), .Y({ _11854_, _11853_, _11851_, _11850_, _11849_, _11848_, _11847_, _11846_, _11845_, _11844_, _11843_, _11842_, _11840_, _11839_, _11838_, _11837_, _11836_, _11835_, _11834_, _11833_, _11832_, _11831_, _11861_, _11860_, _11859_, _11858_, _11857_, _11856_, _11855_, _11852_, _11841_, _11830_ }) );
  \$mux  #( .WIDTH(32) ) _41356_ ( .A(matmul_15_comp_fsm), .B(1), .S(_05857_), .Y({ _11886_, _11885_, _11883_, _11882_, _11881_, _11880_, _11879_, _11878_, _11877_, _11876_, _11875_, _11874_, _11872_, _11871_, _11870_, _11869_, _11868_, _11867_, _11866_, _11865_, _11864_, _11863_, _11893_, _11892_, _11891_, _11890_, _11889_, _11888_, _11887_, _11884_, _11873_, _11862_ }) );
  \$mux  #( .WIDTH(32) ) _41362_ ( .A(matmul_15_sync_comp_count), .B(_22313_), .S(_stream_matmul_15_end_flag), .Y(_22473_) );
  \$mux  #( .WIDTH(32) ) _41363_ ( .A(0), .B(_22473_), .S(_05038_), .Y(_22474_) );
  \$mux  #( .WIDTH(32) ) _41365_ ( .A(4), .B(matmul_15_next_stream_num_ops), .S(_05030_), .Y(_22475_) );
  \$mux  #( .WIDTH(1) ) _41367_ ( .A(1'h1), .B(_control_matmul_15_cond_32_4_1), .S(_05036_), .Y(_22476_) );
  \$mux  #( .WIDTH(1) ) _41369_ ( .A(axim_flag_1118), .B(1'h0), .S(_control_matmul_15_cond_32_4_1), .Y(_22477_) );
  \$mux  #( .WIDTH(1) ) _41370_ ( .A(_22477_), .B(axim_flag_1118), .S(_05029_), .Y(_22478_) );
  \$mux  #( .WIDTH(1) ) _41371_ ( .A(1'h1), .B(_22478_), .S(_05036_), .Y(_22479_) );
  \$mux  #( .WIDTH(1) ) _41373_ ( .A(1'h1), .B(_control_matmul_15_cond_22_3_1), .S(_05037_), .Y(_22480_) );
  \$mux  #( .WIDTH(1) ) _41375_ ( .A(axim_flag_972), .B(1'h0), .S(_control_matmul_15_cond_22_3_1), .Y(_22481_) );
  \$mux  #( .WIDTH(1) ) _41376_ ( .A(_22481_), .B(axim_flag_972), .S(_05031_), .Y(_22482_) );
  \$mux  #( .WIDTH(1) ) _41377_ ( .A(1'h1), .B(_22482_), .S(_05037_), .Y(_22483_) );
  \$mux  #( .WIDTH(1) ) _41379_ ( .A(1'h1), .B(_control_matmul_15_cond_14_2_1), .S(_05039_), .Y(_22484_) );
  \$mux  #( .WIDTH(1) ) _41381_ ( .A(axim_flag_961), .B(1'h0), .S(_control_matmul_15_cond_14_2_1), .Y(_22485_) );
  \$mux  #( .WIDTH(1) ) _41382_ ( .A(_22485_), .B(axim_flag_961), .S(_05032_), .Y(_22486_) );
  \$mux  #( .WIDTH(1) ) _41383_ ( .A(1'h1), .B(_22486_), .S(_05039_), .Y(_22487_) );
  \$mux  #( .WIDTH(1) ) _41385_ ( .A(1'h1), .B(_control_matmul_15_cond_8_1_1), .S(_05040_), .Y(_22488_) );
  \$mux  #( .WIDTH(1) ) _41387_ ( .A(axim_flag_960), .B(1'h0), .S(_control_matmul_15_cond_8_1_1), .Y(_22489_) );
  \$mux  #( .WIDTH(1) ) _41388_ ( .A(_22489_), .B(axim_flag_960), .S(_05033_), .Y(_22490_) );
  \$mux  #( .WIDTH(1) ) _41389_ ( .A(1'h1), .B(_22490_), .S(_05040_), .Y(_22491_) );
  \$mux  #( .WIDTH(1) ) _41391_ ( .A(1'h1), .B(_control_matmul_15_cond_3_0_1), .S(_05041_), .Y(_22492_) );
  \$mux  #( .WIDTH(1) ) _41394_ ( .A(axim_flag_959), .B(1'h0), .S(_control_matmul_15_cond_3_0_1), .Y(_22493_) );
  \$mux  #( .WIDTH(1) ) _41395_ ( .A(_22493_), .B(axim_flag_959), .S(_05034_), .Y(_22494_) );
  \$mux  #( .WIDTH(1) ) _41396_ ( .A(1'h1), .B(_22494_), .S(_05041_), .Y(_22495_) );
  \$mux  #( .WIDTH(1) ) _41398_ ( .A(matmul_15_skip_write_out), .B(1'h0), .S(_05855_), .Y(_11894_) );
  \$mux  #( .WIDTH(1) ) _41399_ ( .A(_22496_), .B(1'h1), .S(RST), .Y(_03133_) );
  \$mux  #( .WIDTH(1) ) _41400_ ( .A(matmul_15_skip_comp), .B(1'h1), .S(_05232_), .Y(_11897_) );
  \$mux  #( .WIDTH(1) ) _41403_ ( .A(matmul_15_skip_read_filter), .B(1'h1), .S(_05232_), .Y(_11899_) );
  \$mux  #( .WIDTH(32) ) _41405_ ( .A(0), .B(matmul_15_out_laddr_offset), .S(matmul_15_skip_write_out), .Y({ _11925_, _11924_, _11922_, _11921_, _11920_, _11919_, _11918_, _11917_, _11916_, _11915_, _11914_, _11913_, _11911_, _11910_, _11909_, _11908_, _11907_, _11906_, _11905_, _11904_, _11903_, _11902_, _11932_, _11931_, _11930_, _11929_, _11928_, _11927_, _11926_, _11923_, _11912_, _11901_ }) );
  \$mux  #( .WIDTH(32) ) _41406_ ( .A(_22308_), .B(matmul_15_out_laddr_offset), .S(_04896_), .Y({ _11957_, _11956_, _11954_, _11953_, _11952_, _11951_, _11950_, _11949_, _11948_, _11947_, _11946_, _11945_, _11943_, _11942_, _11941_, _11940_, _11939_, _11938_, _11937_, _11936_, _11935_, _11934_, _11964_, _11963_, _11962_, _11961_, _11960_, _11959_, _11958_, _11955_, _11944_, _11933_ }) );
  \$mux  #( .WIDTH(32) ) _41408_ ( .A(0), .B(1024), .S(matmul_15_out_page), .Y({ _11989_, _11988_, _11986_, _11985_, _11984_, _11983_, _11982_, _11981_, _11980_, _11979_, _11978_, _11977_, _11975_, _11974_, _11973_, _11972_, _11971_, _11970_, _11969_, _11968_, _11967_, _11966_, _11996_, _11995_, _11994_, _11993_, _11992_, _11991_, _11990_, _11987_, _11976_, _11965_ }) );
  \$mux  #( .WIDTH(32) ) _41410_ ( .A(1024), .B(0), .S(matmul_15_out_page), .Y({ _12053_, _12052_, _12050_, _12049_, _12048_, _12047_, _12046_, _12045_, _12044_, _12043_, _12042_, _12041_, _12039_, _12038_, _12037_, _12036_, _12035_, _12034_, _12033_, _12032_, _12031_, _12030_, _12060_, _12059_, _12058_, _12057_, _12056_, _12055_, _12054_, _12051_, _12040_, _12029_ }) );
  \$mux  #( .WIDTH(1) ) _41412_ ( .A(1'h1), .B(1'h0), .S(matmul_15_out_page), .Y(_12093_) );
  \$mux  #( .WIDTH(32) ) _41414_ ( .A(0), .B(_22311_), .S(_21880_), .Y({ _12119_, _12118_, _12116_, _12115_, _12114_, _12113_, _12112_, _12111_, _12110_, _12109_, _12108_, _12107_, _12105_, _12104_, _12103_, _12102_, _12101_, _12100_, _12099_, _12098_, _12097_, _12096_, _12126_, _12125_, _12124_, _12123_, _12122_, _12121_, _12120_, _12117_, _12106_, _12095_ }) );
  \$mux  #( .WIDTH(32) ) _41416_ ( .A(0), .B(_22310_), .S(_21880_), .Y({ _12183_, _12182_, _12180_, _12179_, _12178_, _12177_, _12176_, _12175_, _12174_, _12173_, _12172_, _12171_, _12169_, _12168_, _12167_, _12166_, _12165_, _12164_, _12163_, _12162_, _12161_, _12160_, _12190_, _12189_, _12188_, _12187_, _12186_, _12185_, _12184_, _12181_, _12170_, _12159_ }) );
  \$mux  #( .WIDTH(1) ) _41420_ ( .A(matmul_15_prev_row_select), .B(1'h0), .S(_04701_), .Y(_22508_) );
  \$mux  #( .WIDTH(32) ) _41425_ ( .A(0), .B(matmul_15_out_ram_select), .S(matmul_15_skip_write_out), .Y({ _12343_, _12342_, _12340_, _12339_, _12338_, _12337_, _12336_, _12335_, _12334_, _12333_, _12332_, _12331_, _12329_, _12328_, _12327_, _12326_, _12325_, _12324_, _12323_, _12322_, _12321_, _12320_, _12350_, _12349_, _12348_, _12347_, _12346_, _12345_, _12344_, _12341_, _12330_, _12319_ }) );
  \$mux  #( .WIDTH(32) ) _41426_ ( .A(0), .B(_22309_), .S(_04896_), .Y({ _12375_, _12374_, _12372_, _12371_, _12370_, _12369_, _12368_, _12367_, _12366_, _12365_, _12364_, _12363_, _12361_, _12360_, _12359_, _12358_, _12357_, _12356_, _12355_, _12354_, _12353_, _12352_, _12382_, _12381_, _12380_, _12379_, _12378_, _12377_, _12376_, _12373_, _12362_, _12351_ }) );
  \$mux  #( .WIDTH(32) ) _41428_ ( .A(0), .B(matmul_15_out_row_count), .S(matmul_15_skip_write_out), .Y({ _12407_, _12406_, _12404_, _12403_, _12402_, _12401_, _12400_, _12399_, _12398_, _12397_, _12396_, _12395_, _12393_, _12392_, _12391_, _12390_, _12389_, _12388_, _12387_, _12386_, _12385_, _12384_, _12414_, _12413_, _12412_, _12411_, _12410_, _12409_, _12408_, _12405_, _12394_, _12383_ }) );
  \$mux  #( .WIDTH(1) ) _41430_ ( .A(matmul_15_row_select), .B(1'h0), .S(_04701_), .Y(_22514_) );
  \$mux  #( .WIDTH(32) ) _41435_ ( .A(matmul_15_next_out_write_size), .B(4), .S(_04701_), .Y(_22518_) );
  \$mux  #( .WIDTH(1) ) _41438_ ( .A(matmul_15_dma_flag_0), .B(1'h1), .S(_04701_), .Y(_22520_) );
  \$mux  #( .WIDTH(32) ) _41440_ ( .A(_22312_), .B(matmul_15_out_base_offset_och), .S(matmul_15_skip_write_out), .Y({ _12567_, _12566_, _12564_, _12563_, _12562_, _12561_, _12560_, _12559_, _12558_, _12557_, _12556_, _12555_, _12553_, _12552_, _12551_, _12550_, _12549_, _12548_, _12547_, _12546_, _12545_, _12544_, _12574_, _12573_, _12572_, _12571_, _12570_, _12569_, _12568_, _12565_, _12554_, _12543_ }) );
  \$mux  #( .WIDTH(32) ) _41442_ ( .A(0), .B(matmul_15_out_base_offset_bat), .S(matmul_15_skip_write_out), .Y({ _12631_, _12630_, _12628_, _12627_, _12626_, _12625_, _12624_, _12623_, _12622_, _12621_, _12620_, _12619_, _12617_, _12616_, _12615_, _12614_, _12613_, _12612_, _12611_, _12610_, _12609_, _12608_, _12638_, _12637_, _12636_, _12635_, _12634_, _12633_, _12632_, _12629_, _12618_, _12607_ }) );
  \$mux  #( .WIDTH(32) ) _41444_ ( .A(0), .B(matmul_15_out_base_offset_row), .S(matmul_15_skip_write_out), .Y({ _12695_, _12694_, _12692_, _12691_, _12690_, _12689_, _12688_, _12687_, _12686_, _12685_, _12684_, _12683_, _12681_, _12680_, _12679_, _12678_, _12677_, _12676_, _12675_, _12674_, _12673_, _12672_, _12702_, _12701_, _12700_, _12699_, _12698_, _12697_, _12696_, _12693_, _12682_, _12671_ }) );
  \$mux  #( .WIDTH(32) ) _41446_ ( .A(0), .B(matmul_15_out_base_offset_col), .S(matmul_15_skip_write_out), .Y({ _12759_, _12758_, _12756_, _12755_, _12754_, _12753_, _12752_, _12751_, _12750_, _12749_, _12748_, _12747_, _12745_, _12744_, _12743_, _12742_, _12741_, _12740_, _12739_, _12738_, _12737_, _12736_, _12766_, _12765_, _12764_, _12763_, _12762_, _12761_, _12760_, _12757_, _12746_, _12735_ }) );
  \$mux  #( .WIDTH(32) ) _41448_ ( .A(0), .B(matmul_15_out_base_offset_val), .S(_05042_), .Y(_22525_) );
  \$mux  #( .WIDTH(32) ) _41453_ ( .A(0), .B(control_matmul_15), .S(_05134_), .Y({ _12823_, _12822_, _12820_, _12819_, _12818_, _12817_, _12816_, _12815_, _12814_, _12813_, _12812_, _12811_, _12809_, _12808_, _12807_, _12806_, _12805_, _12804_, _12803_, _12802_, _12801_, _12800_, _12830_, _12829_, _12828_, _12827_, _12826_, _12825_, _12824_, _12821_, _12810_, _12799_ }) );
  \$mux  #( .WIDTH(32) ) _41454_ ( .A(control_matmul_15), .B(39), .S(_maxi_write_idle), .Y({ _12887_, _12886_, _12884_, _12883_, _12882_, _12881_, _12880_, _12879_, _12878_, _12877_, _12876_, _12875_, _12873_, _12872_, _12871_, _12870_, _12869_, _12868_, _12867_, _12866_, _12865_, _12864_, _12894_, _12893_, _12892_, _12891_, _12890_, _12889_, _12888_, _12885_, _12874_, _12863_ }) );
  \$mux  #( .WIDTH(32) ) _41455_ ( .A(13), .B(38), .S(_05856_), .Y({ _12919_, _12918_, _12916_, _12915_, _12914_, _12913_, _12912_, _12911_, _12910_, _12909_, _12908_, _12907_, _12905_, _12904_, _12903_, _12902_, _12901_, _12900_, _12899_, _12898_, _12897_, _12896_, _12926_, _12925_, _12924_, _12923_, _12922_, _12921_, _12920_, _12917_, _12906_, _12895_ }) );
  \$mux  #( .WIDTH(32) ) _41456_ ( .A(control_matmul_15), .B(32), .S(_maxi_write_idle), .Y({ _12951_, _12950_, _12948_, _12947_, _12946_, _12945_, _12944_, _12943_, _12942_, _12941_, _12940_, _12939_, _12937_, _12936_, _12935_, _12934_, _12933_, _12932_, _12931_, _12930_, _12929_, _12928_, _12958_, _12957_, _12956_, _12955_, _12954_, _12953_, _12952_, _12949_, _12938_, _12927_ }) );
  \$mux  #( .WIDTH(32) ) _41457_ ( .A(31), .B(35), .S(matmul_15_dma_out_mask_0), .Y({ _12983_, _12982_, _12980_, _12979_, _12978_, _12977_, _12976_, _12975_, _12974_, _12973_, _12972_, _12971_, _12969_, _12968_, _12967_, _12966_, _12965_, _12964_, _12963_, _12962_, _12961_, _12960_, _12990_, _12989_, _12988_, _12987_, _12986_, _12985_, _12984_, _12981_, _12970_, _12959_ }) );
  \$mux  #( .WIDTH(32) ) _41458_ ( .A(control_matmul_15), .B(30), .S(_05248_), .Y(_22530_) );
  \$mux  #( .WIDTH(32) ) _41459_ ( .A(_22530_), .B(37), .S(matmul_15_skip_write_out), .Y({ _13015_, _13014_, _13012_, _13011_, _13010_, _13009_, _13008_, _13007_, _13006_, _13005_, _13004_, _13003_, _13001_, _13000_, _12999_, _12998_, _12997_, _12996_, _12995_, _12994_, _12993_, _12992_, _13022_, _13021_, _13020_, _13019_, _13018_, _13017_, _13016_, _13013_, _13002_, _12991_ }) );
  \$mux  #( .WIDTH(32) ) _41460_ ( .A(29), .B(control_matmul_15), .S(_04897_), .Y({ _13047_, _13046_, _13044_, _13043_, _13042_, _13041_, _13040_, _13039_, _13038_, _13037_, _13036_, _13035_, _13033_, _13032_, _13031_, _13030_, _13029_, _13028_, _13027_, _13026_, _13025_, _13024_, _13054_, _13053_, _13052_, _13051_, _13050_, _13049_, _13048_, _13045_, _13034_, _13023_ }) );
  \$mux  #( .WIDTH(32) ) _41461_ ( .A(control_matmul_15), .B(26), .S(_maxi_read_idle), .Y({ _13079_, _13078_, _13076_, _13075_, _13074_, _13073_, _13072_, _13071_, _13070_, _13069_, _13068_, _13067_, _13065_, _13064_, _13063_, _13062_, _13061_, _13060_, _13059_, _13058_, _13057_, _13056_, _13086_, _13085_, _13084_, _13083_, _13082_, _13081_, _13080_, _13077_, _13066_, _13055_ }) );
  \$mux  #( .WIDTH(32) ) _41462_ ( .A(control_matmul_15), .B(22), .S(_maxi_read_idle), .Y({ _13111_, _13110_, _13108_, _13107_, _13106_, _13105_, _13104_, _13103_, _13102_, _13101_, _13100_, _13099_, _13097_, _13096_, _13095_, _13094_, _13093_, _13092_, _13091_, _13090_, _13089_, _13088_, _13118_, _13117_, _13116_, _13115_, _13114_, _13113_, _13112_, _13109_, _13098_, _13087_ }) );
  \$mux  #( .WIDTH(32) ) _41463_ ( .A(21), .B(26), .S(_05871_), .Y(_22531_) );
  \$mux  #( .WIDTH(32) ) _41464_ ( .A(_22531_), .B(27), .S(matmul_15_skip_read_act), .Y({ _13143_, _13142_, _13140_, _13139_, _13138_, _13137_, _13136_, _13135_, _13134_, _13133_, _13132_, _13131_, _13129_, _13128_, _13127_, _13126_, _13125_, _13124_, _13123_, _13122_, _13121_, _13120_, _13150_, _13149_, _13148_, _13147_, _13146_, _13145_, _13144_, _13141_, _13130_, _13119_ }) );
  \$mux  #( .WIDTH(32) ) _41465_ ( .A(control_matmul_15), .B(18), .S(_maxi_read_idle), .Y({ _13175_, _13174_, _13172_, _13171_, _13170_, _13169_, _13168_, _13167_, _13166_, _13165_, _13164_, _13163_, _13161_, _13160_, _13159_, _13158_, _13157_, _13156_, _13155_, _13154_, _13153_, _13152_, _13182_, _13181_, _13180_, _13179_, _13178_, _13177_, _13176_, _13173_, _13162_, _13151_ }) );
  \$mux  #( .WIDTH(32) ) _41466_ ( .A(control_matmul_15), .B(14), .S(_maxi_read_idle), .Y(_22532_) );
  \$mux  #( .WIDTH(32) ) _41467_ ( .A(_22532_), .B(19), .S(matmul_15_skip_read_filter), .Y({ _13207_, _13206_, _13204_, _13203_, _13202_, _13201_, _13200_, _13199_, _13198_, _13197_, _13196_, _13195_, _13193_, _13192_, _13191_, _13190_, _13189_, _13188_, _13187_, _13186_, _13185_, _13184_, _13214_, _13213_, _13212_, _13211_, _13210_, _13209_, _13208_, _13205_, _13194_, _13183_ }) );
  \$mux  #( .WIDTH(32) ) _41468_ ( .A(control_matmul_15), .B(12), .S(_maxi_read_idle), .Y({ _13239_, _13238_, _13236_, _13235_, _13234_, _13233_, _13232_, _13231_, _13230_, _13229_, _13228_, _13227_, _13225_, _13224_, _13223_, _13222_, _13221_, _13220_, _13219_, _13218_, _13217_, _13216_, _13246_, _13245_, _13244_, _13243_, _13242_, _13241_, _13240_, _13237_, _13226_, _13215_ }) );
  \$mux  #( .WIDTH(32) ) _41469_ ( .A(control_matmul_15), .B(8), .S(_maxi_read_idle), .Y({ _13271_, _13270_, _13268_, _13267_, _13266_, _13265_, _13264_, _13263_, _13262_, _13261_, _13260_, _13259_, _13257_, _13256_, _13255_, _13254_, _13253_, _13252_, _13251_, _13250_, _13249_, _13248_, _13278_, _13277_, _13276_, _13275_, _13274_, _13273_, _13272_, _13269_, _13258_, _13247_ }) );
  \$mux  #( .WIDTH(32) ) _41470_ ( .A(control_matmul_15), .B(7), .S(_maxi_read_idle), .Y({ _13303_, _13302_, _13300_, _13299_, _13298_, _13297_, _13296_, _13295_, _13294_, _13293_, _13292_, _13291_, _13289_, _13288_, _13287_, _13286_, _13285_, _13284_, _13283_, _13282_, _13281_, _13280_, _13310_, _13309_, _13308_, _13307_, _13306_, _13305_, _13304_, _13301_, _13290_, _13279_ }) );
  \$mux  #( .WIDTH(32) ) _41471_ ( .A(control_matmul_15), .B(3), .S(_maxi_read_idle), .Y({ _13335_, _13334_, _13332_, _13331_, _13330_, _13329_, _13328_, _13327_, _13326_, _13325_, _13324_, _13323_, _13321_, _13320_, _13319_, _13318_, _13317_, _13316_, _13315_, _13314_, _13313_, _13312_, _13342_, _13341_, _13340_, _13339_, _13338_, _13337_, _13336_, _13333_, _13322_, _13311_ }) );
  \$mux  #( .WIDTH(32) ) _41472_ ( .A(1), .B(control_matmul_15), .S(_05135_), .Y({ _13367_, _13366_, _13364_, _13363_, _13362_, _13361_, _13360_, _13359_, _13358_, _13357_, _13356_, _13355_, _13353_, _13352_, _13351_, _13350_, _13349_, _13348_, _13347_, _13346_, _13345_, _13344_, _13374_, _13373_, _13372_, _13371_, _13370_, _13369_, _13368_, _13365_, _13354_, _13343_ }) );
  \$mux  #( .WIDTH(32) ) _41474_ ( .A(_stream_max_pool_serial_9_sink_3_sink_fsm_1), .B(0), .S(_05854_), .Y(_22533_) );
  \$mux  #( .WIDTH(32) ) _41475_ ( .A(_22533_), .B(0), .S(_stream_max_pool_serial_9_term_sink), .Y({ _13399_, _13398_, _13396_, _13395_, _13394_, _13393_, _13392_, _13391_, _13390_, _13389_, _13388_, _13387_, _13385_, _13384_, _13383_, _13382_, _13381_, _13380_, _13379_, _13378_, _13377_, _13376_, _13406_, _13405_, _13404_, _13403_, _13402_, _13401_, _13400_, _13397_, _13386_, _13375_ }) );
  \$mux  #( .WIDTH(32) ) _41476_ ( .A(_stream_max_pool_serial_9_sink_3_sink_fsm_1), .B(1), .S(_05781_), .Y({ _13463_, _13462_, _13460_, _13459_, _13458_, _13457_, _13456_, _13455_, _13454_, _13453_, _13452_, _13451_, _13449_, _13448_, _13447_, _13446_, _13445_, _13444_, _13443_, _13442_, _13441_, _13440_, _13470_, _13469_, _13468_, _13467_, _13466_, _13465_, _13464_, _13461_, _13450_, _13439_ }) );
  \$mux  #( .WIDTH(32) ) _41478_ ( .A(_stream_max_pool_serial_9_source_1_source_pat_fsm_0), .B(2), .S(_05853_), .Y({ _13527_, _13526_, _13524_, _13523_, _13522_, _13521_, _13520_, _13519_, _13518_, _13517_, _13516_, _13515_, _13513_, _13512_, _13511_, _13510_, _13509_, _13508_, _13507_, _13506_, _13505_, _13504_, _13534_, _13533_, _13532_, _13531_, _13530_, _13529_, _13528_, _13525_, _13514_, _13503_ }) );
  \$mux  #( .WIDTH(32) ) _41479_ ( .A(_stream_max_pool_serial_9_source_1_source_pat_fsm_0), .B(1), .S(_05776_), .Y({ _13559_, _13558_, _13556_, _13555_, _13554_, _13553_, _13552_, _13551_, _13550_, _13549_, _13548_, _13547_, _13545_, _13544_, _13543_, _13542_, _13541_, _13540_, _13539_, _13538_, _13537_, _13536_, _13566_, _13565_, _13564_, _13563_, _13562_, _13561_, _13560_, _13557_, _13546_, _13535_ }) );
  \$mux  #( .WIDTH(4) ) _41481_ ( .A({ max_pool_serial_9_stream_pad_mask_1_1, max_pool_serial_9_stream_pad_mask_1_0, max_pool_serial_9_stream_pad_mask_0_1, max_pool_serial_9_stream_pad_mask_0_0 }), .B(max_pool_serial_9_stream_pad_masks), .S(_05047_), .Y(_22536_) );
  \$mux  #( .WIDTH(32) ) _41483_ ( .A(max_pool_serial_9_row_count), .B(max_pool_serial_9_row_count_buf), .S(_05048_), .Y(_22537_) );
  \$mux  #( .WIDTH(32) ) _41485_ ( .A(max_pool_serial_9_out_page_comp_offset), .B(max_pool_serial_9_out_page_comp_offset_buf), .S(_05048_), .Y(_22538_) );
  \$mux  #( .WIDTH(32) ) _41487_ ( .A(max_pool_serial_9_act_page_comp_offset), .B(max_pool_serial_9_act_page_comp_offset_buf), .S(_05048_), .Y(_22539_) );
  \$mux  #( .WIDTH(32) ) _41489_ ( .A(2), .B(0), .S(_05247_), .Y({ _13591_, _13590_, _13588_, _13587_, _13586_, _13585_, _13584_, _13583_, _13582_, _13581_, _13580_, _13579_, _13577_, _13576_, _13575_, _13574_, _13573_, _13572_, _13571_, _13570_, _13569_, _13568_, _13598_, _13597_, _13596_, _13595_, _13594_, _13593_, _13592_, _13589_, _13578_, _13567_ }) );
  \$mux  #( .WIDTH(32) ) _41490_ ( .A(4), .B(max_pool_serial_9_comp_fsm), .S(_stream_max_pool_serial_9_source_busy), .Y({ _13655_, _13654_, _13652_, _13651_, _13650_, _13649_, _13648_, _13647_, _13646_, _13645_, _13644_, _13643_, _13641_, _13640_, _13639_, _13638_, _13637_, _13636_, _13635_, _13634_, _13633_, _13632_, _13662_, _13661_, _13660_, _13659_, _13658_, _13657_, _13656_, _13653_, _13642_, _13631_ }) );
  \$mux  #( .WIDTH(32) ) _41491_ ( .A(max_pool_serial_9_comp_fsm), .B(1), .S(_05852_), .Y({ _13687_, _13686_, _13684_, _13683_, _13682_, _13681_, _13680_, _13679_, _13678_, _13677_, _13676_, _13675_, _13673_, _13672_, _13671_, _13670_, _13669_, _13668_, _13667_, _13666_, _13665_, _13664_, _13694_, _13693_, _13692_, _13691_, _13690_, _13689_, _13688_, _13685_, _13674_, _13663_ }) );
  \$mux  #( .WIDTH(32) ) _41493_ ( .A(0), .B(max_pool_serial_9_comp_count), .S(_05055_), .Y(_22541_) );
  \$mux  #( .WIDTH(32) ) _41494_ ( .A(_22541_), .B(_22304_), .S(_stream_max_pool_serial_9_end_flag), .Y(_22542_) );
  \$mux  #( .WIDTH(32) ) _41496_ ( .A(_22306_), .B(0), .S(_05247_), .Y({ _13719_, _13718_, _13716_, _13715_, _13714_, _13713_, _13712_, _13711_, _13710_, _13709_, _13708_, _13707_, _13705_, _13704_, _13703_, _13702_, _13701_, _13700_, _13699_, _13698_, _13697_, _13696_, _13726_, _13725_, _13724_, _13723_, _13722_, _13721_, _13720_, _13717_, _13706_, _13695_ }) );
  \$mux  #( .WIDTH(32) ) _41498_ ( .A(_22305_), .B(0), .S(_05247_), .Y({ _13783_, _13782_, _13780_, _13779_, _13778_, _13777_, _13776_, _13775_, _13774_, _13773_, _13772_, _13771_, _13769_, _13768_, _13767_, _13766_, _13765_, _13764_, _13763_, _13762_, _13761_, _13760_, _13790_, _13789_, _13788_, _13787_, _13786_, _13785_, _13784_, _13781_, _13770_, _13759_ }) );
  \$mux  #( .WIDTH(32) ) _41500_ ( .A(_22307_), .B(0), .S(_05247_), .Y({ _13847_, _13846_, _13844_, _13843_, _13842_, _13841_, _13840_, _13839_, _13838_, _13837_, _13836_, _13835_, _13833_, _13832_, _13831_, _13830_, _13829_, _13828_, _13827_, _13826_, _13825_, _13824_, _13854_, _13853_, _13852_, _13851_, _13850_, _13849_, _13848_, _13845_, _13834_, _13823_ }) );
  \$mux  #( .WIDTH(1) ) _41502_ ( .A(1'h1), .B(_control_max_pool_serial_9_cond_19_2_1), .S(_05053_), .Y(_22546_) );
  \$mux  #( .WIDTH(1) ) _41504_ ( .A(axim_flag_909), .B(1'h0), .S(_control_max_pool_serial_9_cond_19_2_1), .Y(_22547_) );
  \$mux  #( .WIDTH(1) ) _41505_ ( .A(_22547_), .B(axim_flag_909), .S(_05049_), .Y(_22548_) );
  \$mux  #( .WIDTH(1) ) _41506_ ( .A(1'h1), .B(_22548_), .S(_05053_), .Y(_22549_) );
  \$mux  #( .WIDTH(1) ) _41508_ ( .A(1'h1), .B(_control_max_pool_serial_9_cond_11_1_1), .S(_05054_), .Y(_22550_) );
  \$mux  #( .WIDTH(1) ) _41510_ ( .A(axim_flag_861), .B(1'h0), .S(_control_max_pool_serial_9_cond_11_1_1), .Y(_22551_) );
  \$mux  #( .WIDTH(1) ) _41511_ ( .A(_22551_), .B(axim_flag_861), .S(_05050_), .Y(_22552_) );
  \$mux  #( .WIDTH(1) ) _41512_ ( .A(1'h1), .B(_22552_), .S(_05054_), .Y(_22553_) );
  \$mux  #( .WIDTH(1) ) _41514_ ( .A(1'h1), .B(_control_max_pool_serial_9_cond_5_0_1), .S(_05056_), .Y(_22554_) );
  \$mux  #( .WIDTH(1) ) _41517_ ( .A(axim_flag_850), .B(1'h0), .S(_control_max_pool_serial_9_cond_5_0_1), .Y(_22555_) );
  \$mux  #( .WIDTH(1) ) _41518_ ( .A(_22555_), .B(axim_flag_850), .S(_05051_), .Y(_22556_) );
  \$mux  #( .WIDTH(1) ) _41519_ ( .A(1'h1), .B(_22556_), .S(_05056_), .Y(_22557_) );
  \$mux  #( .WIDTH(1) ) _41522_ ( .A(max_pool_serial_9_skip_write_out), .B(1'h0), .S(_05851_), .Y(_13919_) );
  \$mux  #( .WIDTH(1) ) _41524_ ( .A(max_pool_serial_9_skip_comp), .B(1'h1), .S(_05246_), .Y(_13921_) );
  \$mux  #( .WIDTH(1) ) _41526_ ( .A(max_pool_serial_9_skip_read_act), .B(1'h1), .S(_05246_), .Y(_13923_) );
  \$mux  #( .WIDTH(32) ) _41528_ ( .A(0), .B(1024), .S(max_pool_serial_9_out_page), .Y({ _13949_, _13948_, _13946_, _13945_, _13944_, _13943_, _13942_, _13941_, _13940_, _13939_, _13938_, _13937_, _13935_, _13934_, _13933_, _13932_, _13931_, _13930_, _13929_, _13928_, _13927_, _13926_, _13956_, _13955_, _13954_, _13953_, _13952_, _13951_, _13950_, _13947_, _13936_, _13925_ }) );
  \$mux  #( .WIDTH(32) ) _41530_ ( .A(1024), .B(0), .S(max_pool_serial_9_out_page), .Y({ _14013_, _14012_, _14010_, _14009_, _14008_, _14007_, _14006_, _14005_, _14004_, _14003_, _14002_, _14001_, _13999_, _13998_, _13997_, _13996_, _13995_, _13994_, _13993_, _13992_, _13991_, _13990_, _14020_, _14019_, _14018_, _14017_, _14016_, _14015_, _14014_, _14011_, _14000_, _13989_ }) );
  \$mux  #( .WIDTH(1) ) _41532_ ( .A(1'h1), .B(1'h0), .S(max_pool_serial_9_out_page), .Y(_14053_) );
  \$mux  #( .WIDTH(32) ) _41535_ ( .A(1024), .B(0), .S(max_pool_serial_9_act_page), .Y({ _14079_, _14078_, _14076_, _14075_, _14074_, _14073_, _14072_, _14071_, _14070_, _14069_, _14068_, _14067_, _14065_, _14064_, _14063_, _14062_, _14061_, _14060_, _14059_, _14058_, _14057_, _14056_, _14086_, _14085_, _14084_, _14083_, _14082_, _14081_, _14080_, _14077_, _14066_, _14055_ }) );
  \$mux  #( .WIDTH(1) ) _41537_ ( .A(1'h1), .B(1'h0), .S(max_pool_serial_9_act_page), .Y(_14119_) );
  \$mux  #( .WIDTH(32) ) _41541_ ( .A(max_pool_serial_9_bat_count), .B(0), .S(_05246_), .Y({ _14209_, _14208_, _14206_, _14205_, _14204_, _14203_, _14202_, _14201_, _14200_, _14199_, _14198_, _14197_, _14195_, _14194_, _14193_, _14192_, _14191_, _14190_, _14189_, _14188_, _14187_, _14186_, _14216_, _14215_, _14214_, _14213_, _14212_, _14211_, _14210_, _14207_, _14196_, _14185_ }) );
  \$mux  #( .WIDTH(32) ) _41543_ ( .A(_22302_), .B(0), .S(_05246_), .Y({ _14273_, _14272_, _14270_, _14269_, _14268_, _14267_, _14266_, _14265_, _14264_, _14263_, _14262_, _14261_, _14259_, _14258_, _14257_, _14256_, _14255_, _14254_, _14253_, _14252_, _14251_, _14250_, _14280_, _14279_, _14278_, _14277_, _14276_, _14275_, _14274_, _14271_, _14260_, _14249_ }) );
  \$mux  #( .WIDTH(32) ) _41545_ ( .A(max_pool_serial_9_out_base_offset_bat), .B(0), .S(_05850_), .Y({ _14337_, _14336_, _14334_, _14333_, _14332_, _14331_, _14330_, _14329_, _14328_, _14327_, _14326_, _14325_, _14323_, _14322_, _14321_, _14320_, _14319_, _14318_, _14317_, _14316_, _14315_, _14314_, _14344_, _14343_, _14342_, _14341_, _14340_, _14339_, _14338_, _14335_, _14324_, _14313_ }) );
  \$mux  #( .WIDTH(32) ) _41547_ ( .A(_22303_), .B(max_pool_serial_9_out_base_offset_row), .S(max_pool_serial_9_skip_write_out), .Y(_22573_) );
  \$mux  #( .WIDTH(32) ) _41548_ ( .A(_22573_), .B(0), .S(_05850_), .Y({ _14401_, _14400_, _14398_, _14397_, _14396_, _14395_, _14394_, _14393_, _14392_, _14391_, _14390_, _14389_, _14387_, _14386_, _14385_, _14384_, _14383_, _14382_, _14381_, _14380_, _14379_, _14378_, _14408_, _14407_, _14406_, _14405_, _14404_, _14403_, _14402_, _14399_, _14388_, _14377_ }) );
  \$mux  #( .WIDTH(32) ) _41550_ ( .A(max_pool_serial_9_act_base_offset_bat), .B(0), .S(_05246_), .Y({ _14465_, _14464_, _14462_, _14461_, _14460_, _14459_, _14458_, _14457_, _14456_, _14455_, _14454_, _14453_, _14451_, _14450_, _14449_, _14448_, _14447_, _14446_, _14445_, _14444_, _14443_, _14442_, _14472_, _14471_, _14470_, _14469_, _14468_, _14467_, _14466_, _14463_, _14452_, _14441_ }) );
  \$mux  #( .WIDTH(32) ) _41552_ ( .A(_22301_), .B(0), .S(_05246_), .Y({ _14529_, _14528_, _14526_, _14525_, _14524_, _14523_, _14522_, _14521_, _14520_, _14519_, _14518_, _14517_, _14515_, _14514_, _14513_, _14512_, _14511_, _14510_, _14509_, _14508_, _14507_, _14506_, _14536_, _14535_, _14534_, _14533_, _14532_, _14531_, _14530_, _14527_, _14516_, _14505_ }) );
  \$mux  #( .WIDTH(32) ) _41554_ ( .A(0), .B(control_max_pool_serial_9), .S(_05145_), .Y(_22577_) );
  \$mux  #( .WIDTH(32) ) _41555_ ( .A(0), .B(_22577_), .S(_05141_), .Y({ _14593_, _14592_, _14590_, _14589_, _14588_, _14587_, _14586_, _14585_, _14584_, _14583_, _14582_, _14581_, _14579_, _14578_, _14577_, _14576_, _14575_, _14574_, _14573_, _14572_, _14571_, _14570_, _14600_, _14599_, _14598_, _14597_, _14596_, _14595_, _14594_, _14591_, _14580_, _14569_ }) );
  \$mux  #( .WIDTH(32) ) _41556_ ( .A(control_max_pool_serial_9), .B(25), .S(_maxi_write_idle), .Y({ _14657_, _14656_, _14654_, _14653_, _14652_, _14651_, _14650_, _14649_, _14648_, _14647_, _14646_, _14645_, _14643_, _14642_, _14641_, _14640_, _14639_, _14638_, _14637_, _14636_, _14635_, _14634_, _14664_, _14663_, _14662_, _14661_, _14660_, _14659_, _14658_, _14655_, _14644_, _14633_ }) );
  \$mux  #( .WIDTH(32) ) _41557_ ( .A(3), .B(24), .S(_05850_), .Y({ _14689_, _14688_, _14686_, _14685_, _14684_, _14683_, _14682_, _14681_, _14680_, _14679_, _14678_, _14677_, _14675_, _14674_, _14673_, _14672_, _14671_, _14670_, _14669_, _14668_, _14667_, _14666_, _14696_, _14695_, _14694_, _14693_, _14692_, _14691_, _14690_, _14687_, _14676_, _14665_ }) );
  \$mux  #( .WIDTH(32) ) _41558_ ( .A(control_max_pool_serial_9), .B(19), .S(_maxi_write_idle), .Y({ _14721_, _14720_, _14718_, _14717_, _14716_, _14715_, _14714_, _14713_, _14712_, _14711_, _14710_, _14709_, _14707_, _14706_, _14705_, _14704_, _14703_, _14702_, _14701_, _14700_, _14699_, _14698_, _14728_, _14727_, _14726_, _14725_, _14724_, _14723_, _14722_, _14719_, _14708_, _14697_ }) );
  \$mux  #( .WIDTH(32) ) _41559_ ( .A(control_max_pool_serial_9), .B(18), .S(_05245_), .Y(_22579_) );
  \$mux  #( .WIDTH(32) ) _41560_ ( .A(_22579_), .B(23), .S(max_pool_serial_9_skip_write_out), .Y({ _14753_, _14752_, _14750_, _14749_, _14748_, _14747_, _14746_, _14745_, _14744_, _14743_, _14742_, _14741_, _14739_, _14738_, _14737_, _14736_, _14735_, _14734_, _14733_, _14732_, _14731_, _14730_, _14760_, _14759_, _14758_, _14757_, _14756_, _14755_, _14754_, _14751_, _14740_, _14729_ }) );
  \$mux  #( .WIDTH(32) ) _41561_ ( .A(17), .B(control_max_pool_serial_9), .S(_04898_), .Y({ _14785_, _14784_, _14782_, _14781_, _14780_, _14779_, _14778_, _14777_, _14776_, _14775_, _14774_, _14773_, _14771_, _14770_, _14769_, _14768_, _14767_, _14766_, _14765_, _14764_, _14763_, _14762_, _14792_, _14791_, _14790_, _14789_, _14788_, _14787_, _14786_, _14783_, _14772_, _14761_ }) );
  \$mux  #( .WIDTH(32) ) _41562_ ( .A(control_max_pool_serial_9), .B(15), .S(_maxi_read_idle), .Y({ _14817_, _14816_, _14814_, _14813_, _14812_, _14811_, _14810_, _14809_, _14808_, _14807_, _14806_, _14805_, _14803_, _14802_, _14801_, _14800_, _14799_, _14798_, _14797_, _14796_, _14795_, _14794_, _14824_, _14823_, _14822_, _14821_, _14820_, _14819_, _14818_, _14815_, _14804_, _14793_ }) );
  \$mux  #( .WIDTH(32) ) _41563_ ( .A(control_max_pool_serial_9), .B(11), .S(_maxi_read_idle), .Y({ _14849_, _14848_, _14846_, _14845_, _14844_, _14843_, _14842_, _14841_, _14840_, _14839_, _14838_, _14837_, _14835_, _14834_, _14833_, _14832_, _14831_, _14830_, _14829_, _14828_, _14827_, _14826_, _14856_, _14855_, _14854_, _14853_, _14852_, _14851_, _14850_, _14847_, _14836_, _14825_ }) );
  \$mux  #( .WIDTH(32) ) _41564_ ( .A(10), .B(15), .S(max_pool_serial_9_dma_pad_mask_1), .Y({ _14881_, _14880_, _14878_, _14877_, _14876_, _14875_, _14874_, _14873_, _14872_, _14871_, _14870_, _14869_, _14867_, _14866_, _14865_, _14864_, _14863_, _14862_, _14861_, _14860_, _14859_, _14858_, _14888_, _14887_, _14886_, _14885_, _14884_, _14883_, _14882_, _14879_, _14868_, _14857_ }) );
  \$mux  #( .WIDTH(32) ) _41565_ ( .A(control_max_pool_serial_9), .B(9), .S(_maxi_read_idle), .Y({ _14913_, _14912_, _14910_, _14909_, _14908_, _14907_, _14906_, _14905_, _14904_, _14903_, _14902_, _14901_, _14899_, _14898_, _14897_, _14896_, _14895_, _14894_, _14893_, _14892_, _14891_, _14890_, _14920_, _14919_, _14918_, _14917_, _14916_, _14915_, _14914_, _14911_, _14900_, _14889_ }) );
  \$mux  #( .WIDTH(32) ) _41566_ ( .A(control_max_pool_serial_9), .B(5), .S(_maxi_read_idle), .Y({ _14945_, _14944_, _14942_, _14941_, _14940_, _14939_, _14938_, _14937_, _14936_, _14935_, _14934_, _14933_, _14931_, _14930_, _14929_, _14928_, _14927_, _14926_, _14925_, _14924_, _14923_, _14922_, _14952_, _14951_, _14950_, _14949_, _14948_, _14947_, _14946_, _14943_, _14932_, _14921_ }) );
  \$mux  #( .WIDTH(32) ) _41567_ ( .A(4), .B(9), .S(max_pool_serial_9_dma_pad_mask_0), .Y(_22580_) );
  \$mux  #( .WIDTH(32) ) _41568_ ( .A(_22580_), .B(16), .S(max_pool_serial_9_skip_read_act), .Y({ _14977_, _14976_, _14974_, _14973_, _14972_, _14971_, _14970_, _14969_, _14968_, _14967_, _14966_, _14965_, _14963_, _14962_, _14961_, _14960_, _14959_, _14958_, _14957_, _14956_, _14955_, _14954_, _14984_, _14983_, _14982_, _14981_, _14980_, _14979_, _14978_, _14975_, _14964_, _14953_ }) );
  \$mux  #( .WIDTH(32) ) _41569_ ( .A(1), .B(control_max_pool_serial_9), .S(_05146_), .Y(_22581_) );
  \$mux  #( .WIDTH(32) ) _41570_ ( .A(1), .B(_22581_), .S(_05142_), .Y({ _15009_, _15008_, _15006_, _15005_, _15004_, _15003_, _15002_, _15001_, _15000_, _14999_, _14998_, _14997_, _14995_, _14994_, _14993_, _14992_, _14991_, _14990_, _14989_, _14988_, _14987_, _14986_, _15016_, _15015_, _15014_, _15013_, _15012_, _15011_, _15010_, _15007_, _14996_, _14985_ }) );
  \$mux  #( .WIDTH(1) ) _41572_ ( .A(1'h1), .B(__maxi_write_fsm_cond_4_0_1), .S(_05058_), .Y(_22582_) );
  \$mux  #( .WIDTH(1) ) _41575_ ( .A(axim_flag_849), .B(1'h0), .S(__maxi_write_fsm_cond_4_0_1), .Y(_22583_) );
  \$mux  #( .WIDTH(1) ) _41576_ ( .A(_22583_), .B(axim_flag_849), .S(_05057_), .Y(_22584_) );
  \$mux  #( .WIDTH(1) ) _41577_ ( .A(1'h1), .B(_22584_), .S(_05058_), .Y(_22585_) );
  \$mux  #( .WIDTH(33) ) _41579_ ( .A(_26329_), .B(_26328_), .S(_05244_), .Y(_22586_) );
  \$mux  #( .WIDTH(33) ) _41580_ ( .A(_22586_), .B(33'h000000000), .S(_05263_), .Y(_22587_) );
  \$mux  #( .WIDTH(33) ) _41581_ ( .A(_22587_), .B(_26328_), .S(_05847_), .Y({ _15042_, _15041_, _15040_, _15038_, _15037_, _15036_, _15035_, _15034_, _15033_, _15032_, _15031_, _15030_, _15029_, _15027_, _15026_, _15025_, _15024_, _15023_, _15022_, _15021_, _15020_, _15019_, _15018_, _15049_, _15048_, _15047_, _15046_, _15045_, _15044_, _15043_, _15039_, _15028_, _15017_ }) );
  \$mux  #( .WIDTH(33) ) _41582_ ( .A(_maxi_write_rest_size), .B(_maxi_write_size), .S(_maxi_write_start), .Y({ _15108_, _15107_, _15106_, _15104_, _15103_, _15102_, _15101_, _15100_, _15099_, _15098_, _15097_, _15096_, _15095_, _15093_, _15092_, _15091_, _15090_, _15089_, _15088_, _15087_, _15086_, _15085_, _15084_, _15115_, _15114_, _15113_, _15112_, _15111_, _15110_, _15109_, _15105_, _15094_, _15083_ }) );
  \$mux  #( .WIDTH(33) ) _41584_ ( .A(33'h000000100), .B({ 2'h0, _25923_[30:0] }), .S(_05244_), .Y(_22589_) );
  \$mux  #( .WIDTH(33) ) _41585_ ( .A(_22589_), .B(_maxi_write_rest_size), .S(_05263_), .Y(_22590_) );
  \$mux  #( .WIDTH(33) ) _41586_ ( .A(_22590_), .B({ 2'h0, _25923_[30:0] }), .S(_05847_), .Y(_22591_) );
  \$mux  #( .WIDTH(33) ) _41587_ ( .A(_22591_), .B(_maxi_write_cur_size), .S(_05059_), .Y(_22592_) );
  \$mux  #( .WIDTH(32) ) _41589_ ( .A(_maxi_write_cur_global_addr), .B(_22300_[31:0]), .S(_maxi_write_data_done), .Y({ _15140_, _15139_, _15137_, _15136_, _15135_, _15134_, _15133_, _15132_, _15131_, _15130_, _15129_, _15128_, _15126_, _15125_, _15124_, _15123_, _15122_, _15121_, _15120_, _15119_, _15118_, _15117_, _15147_, _15146_, _15145_, _15144_, _15143_, _15142_, _15141_, _15138_, _15127_, _15116_ }) );
  \$mux  #( .WIDTH(32) ) _41590_ ( .A(_maxi_write_cur_global_addr), .B({ _22299_[31:2], 2'h0 }), .S(_maxi_write_start), .Y({ _15204_, _15203_, _15201_, _15200_, _15199_, _15198_, _15197_, _15196_, _15195_, _15194_, _15193_, _15192_, _15190_, _15189_, _15188_, _15187_, _15186_, _15185_, _15184_, _15183_, _15182_, _15181_, _15211_, _15210_, _15209_, _15208_, _15207_, _15206_, _15205_, _15202_, _15191_, _15180_ }) );
  \$mux  #( .WIDTH(32) ) _41592_ ( .A(_maxi_write_fsm), .B(1), .S(_05848_), .Y(_22595_) );
  \$mux  #( .WIDTH(32) ) _41593_ ( .A(_22595_), .B(4), .S(_05849_), .Y({ _15268_, _15267_, _15265_, _15264_, _15263_, _15262_, _15261_, _15260_, _15259_, _15258_, _15257_, _15256_, _15254_, _15253_, _15252_, _15251_, _15250_, _15249_, _15248_, _15247_, _15246_, _15245_, _15275_, _15274_, _15273_, _15272_, _15271_, _15270_, _15269_, _15266_, _15255_, _15244_ }) );
  \$mux  #( .WIDTH(32) ) _41594_ ( .A(_maxi_write_fsm), .B(3), .S(_05865_), .Y({ _15300_, _15299_, _15297_, _15296_, _15295_, _15294_, _15293_, _15292_, _15291_, _15290_, _15289_, _15288_, _15286_, _15285_, _15284_, _15283_, _15282_, _15281_, _15280_, _15279_, _15278_, _15277_, _15307_, _15306_, _15305_, _15304_, _15303_, _15302_, _15301_, _15298_, _15287_, _15276_ }) );
  \$mux  #( .WIDTH(32) ) _41595_ ( .A(_maxi_write_fsm), .B(1), .S(_05647_), .Y(_22596_) );
  \$mux  #( .WIDTH(32) ) _41596_ ( .A(_22596_), .B(1), .S(_05429_), .Y(_22597_) );
  \$mux  #( .WIDTH(32) ) _41597_ ( .A(_22597_), .B(1), .S(_05479_), .Y({ _15332_, _15331_, _15329_, _15328_, _15327_, _15326_, _15325_, _15324_, _15323_, _15322_, _15321_, _15320_, _15318_, _15317_, _15316_, _15315_, _15314_, _15313_, _15312_, _15311_, _15310_, _15309_, _15339_, _15338_, _15337_, _15336_, _15335_, _15334_, _15333_, _15330_, _15319_, _15308_ }) );
  \$mux  #( .WIDTH(32) ) _41599_ ( .A(_stream_conv2d_8_sink_37_sink_fsm_20), .B(0), .S(_05846_), .Y(_22598_) );
  \$mux  #( .WIDTH(32) ) _41600_ ( .A(_22598_), .B(0), .S(_stream_conv2d_8_term_sink), .Y({ _15364_, _15363_, _15361_, _15360_, _15359_, _15358_, _15357_, _15356_, _15355_, _15354_, _15353_, _15352_, _15350_, _15349_, _15348_, _15347_, _15346_, _15345_, _15344_, _15343_, _15342_, _15341_, _15371_, _15370_, _15369_, _15368_, _15367_, _15366_, _15365_, _15362_, _15351_, _15340_ }) );
  \$mux  #( .WIDTH(32) ) _41601_ ( .A(_stream_conv2d_8_sink_37_sink_fsm_20), .B(1), .S(_05774_), .Y({ _15428_, _15427_, _15425_, _15424_, _15423_, _15422_, _15421_, _15420_, _15419_, _15418_, _15417_, _15416_, _15414_, _15413_, _15412_, _15411_, _15410_, _15409_, _15408_, _15407_, _15406_, _15405_, _15435_, _15434_, _15433_, _15432_, _15431_, _15430_, _15429_, _15426_, _15415_, _15404_ }) );
  \$mux  #( .WIDTH(32) ) _41603_ ( .A(_stream_conv2d_8_source_36_source_pat_fsm_19), .B(2), .S(_05845_), .Y({ _15492_, _15491_, _15489_, _15488_, _15487_, _15486_, _15485_, _15484_, _15483_, _15482_, _15481_, _15480_, _15478_, _15477_, _15476_, _15475_, _15474_, _15473_, _15472_, _15471_, _15470_, _15469_, _15499_, _15498_, _15497_, _15496_, _15495_, _15494_, _15493_, _15490_, _15479_, _15468_ }) );
  \$mux  #( .WIDTH(32) ) _41604_ ( .A(_stream_conv2d_8_source_36_source_pat_fsm_19), .B(1), .S(_05769_), .Y({ _15524_, _15523_, _15521_, _15520_, _15519_, _15518_, _15517_, _15516_, _15515_, _15514_, _15513_, _15512_, _15510_, _15509_, _15508_, _15507_, _15506_, _15505_, _15504_, _15503_, _15502_, _15501_, _15531_, _15530_, _15529_, _15528_, _15527_, _15526_, _15525_, _15522_, _15511_, _15500_ }) );
  \$mux  #( .WIDTH(32) ) _41608_ ( .A(_stream_conv2d_8_source_35_source_pat_fsm_18), .B(2), .S(_05844_), .Y({ _15588_, _15587_, _15585_, _15584_, _15583_, _15582_, _15581_, _15580_, _15579_, _15578_, _15577_, _15576_, _15574_, _15573_, _15572_, _15571_, _15570_, _15569_, _15568_, _15567_, _15566_, _15565_, _15595_, _15594_, _15593_, _15592_, _15591_, _15590_, _15589_, _15586_, _15575_, _15564_ }) );
  \$mux  #( .WIDTH(32) ) _41609_ ( .A(_stream_conv2d_8_source_35_source_pat_fsm_18), .B(1), .S(_05764_), .Y({ _15620_, _15619_, _15617_, _15616_, _15615_, _15614_, _15613_, _15612_, _15611_, _15610_, _15609_, _15608_, _15606_, _15605_, _15604_, _15603_, _15602_, _15601_, _15600_, _15599_, _15598_, _15597_, _15627_, _15626_, _15625_, _15624_, _15623_, _15622_, _15621_, _15618_, _15607_, _15596_ }) );
  \$mux  #( .WIDTH(32) ) _41613_ ( .A(_stream_conv2d_8_source_34_source_pat_fsm_17), .B(2), .S(_05843_), .Y({ _15684_, _15683_, _15681_, _15680_, _15679_, _15678_, _15677_, _15676_, _15675_, _15674_, _15673_, _15672_, _15670_, _15669_, _15668_, _15667_, _15666_, _15665_, _15664_, _15663_, _15662_, _15661_, _15691_, _15690_, _15689_, _15688_, _15687_, _15686_, _15685_, _15682_, _15671_, _15660_ }) );
  \$mux  #( .WIDTH(32) ) _41614_ ( .A(_stream_conv2d_8_source_34_source_pat_fsm_17), .B(1), .S(_05759_), .Y({ _15716_, _15715_, _15713_, _15712_, _15711_, _15710_, _15709_, _15708_, _15707_, _15706_, _15705_, _15704_, _15702_, _15701_, _15700_, _15699_, _15698_, _15697_, _15696_, _15695_, _15694_, _15693_, _15723_, _15722_, _15721_, _15720_, _15719_, _15718_, _15717_, _15714_, _15703_, _15692_ }) );
  \$mux  #( .WIDTH(32) ) _41618_ ( .A(_stream_conv2d_8_source_33_source_pat_fsm_16), .B(2), .S(_05842_), .Y({ _15780_, _15779_, _15777_, _15776_, _15775_, _15774_, _15773_, _15772_, _15771_, _15770_, _15769_, _15768_, _15766_, _15765_, _15764_, _15763_, _15762_, _15761_, _15760_, _15759_, _15758_, _15757_, _15787_, _15786_, _15785_, _15784_, _15783_, _15782_, _15781_, _15778_, _15767_, _15756_ }) );
  \$mux  #( .WIDTH(32) ) _41619_ ( .A(_stream_conv2d_8_source_33_source_pat_fsm_16), .B(1), .S(_05754_), .Y({ _15812_, _15811_, _15809_, _15808_, _15807_, _15806_, _15805_, _15804_, _15803_, _15802_, _15801_, _15800_, _15798_, _15797_, _15796_, _15795_, _15794_, _15793_, _15792_, _15791_, _15790_, _15789_, _15819_, _15818_, _15817_, _15816_, _15815_, _15814_, _15813_, _15810_, _15799_, _15788_ }) );
  \$mux  #( .WIDTH(32) ) _41623_ ( .A(_stream_conv2d_8_source_32_source_pat_fsm_15), .B(2), .S(_05841_), .Y({ _15876_, _15875_, _15873_, _15872_, _15871_, _15870_, _15869_, _15868_, _15867_, _15866_, _15865_, _15864_, _15862_, _15861_, _15860_, _15859_, _15858_, _15857_, _15856_, _15855_, _15854_, _15853_, _15883_, _15882_, _15881_, _15880_, _15879_, _15878_, _15877_, _15874_, _15863_, _15852_ }) );
  \$mux  #( .WIDTH(32) ) _41624_ ( .A(_stream_conv2d_8_source_32_source_pat_fsm_15), .B(1), .S(_05749_), .Y({ _15908_, _15907_, _15905_, _15904_, _15903_, _15902_, _15901_, _15900_, _15899_, _15898_, _15897_, _15896_, _15894_, _15893_, _15892_, _15891_, _15890_, _15889_, _15888_, _15887_, _15886_, _15885_, _15915_, _15914_, _15913_, _15912_, _15911_, _15910_, _15909_, _15906_, _15895_, _15884_ }) );
  \$mux  #( .WIDTH(32) ) _41628_ ( .A(_stream_conv2d_8_source_31_source_pat_fsm_14), .B(2), .S(_05840_), .Y({ _15972_, _15971_, _15969_, _15968_, _15967_, _15966_, _15965_, _15964_, _15963_, _15962_, _15961_, _15960_, _15958_, _15957_, _15956_, _15955_, _15954_, _15953_, _15952_, _15951_, _15950_, _15949_, _15979_, _15978_, _15977_, _15976_, _15975_, _15974_, _15973_, _15970_, _15959_, _15948_ }) );
  \$mux  #( .WIDTH(32) ) _41629_ ( .A(_stream_conv2d_8_source_31_source_pat_fsm_14), .B(1), .S(_05744_), .Y({ _16004_, _16003_, _16001_, _16000_, _15999_, _15998_, _15997_, _15996_, _15995_, _15994_, _15993_, _15992_, _15990_, _15989_, _15988_, _15987_, _15986_, _15985_, _15984_, _15983_, _15982_, _15981_, _16011_, _16010_, _16009_, _16008_, _16007_, _16006_, _16005_, _16002_, _15991_, _15980_ }) );
  \$mux  #( .WIDTH(32) ) _41633_ ( .A(_stream_conv2d_8_source_30_source_pat_fsm_13), .B(2), .S(_05839_), .Y({ _16068_, _16067_, _16065_, _16064_, _16063_, _16062_, _16061_, _16060_, _16059_, _16058_, _16057_, _16056_, _16054_, _16053_, _16052_, _16051_, _16050_, _16049_, _16048_, _16047_, _16046_, _16045_, _16075_, _16074_, _16073_, _16072_, _16071_, _16070_, _16069_, _16066_, _16055_, _16044_ }) );
  \$mux  #( .WIDTH(32) ) _41634_ ( .A(_stream_conv2d_8_source_30_source_pat_fsm_13), .B(1), .S(_05739_), .Y({ _16100_, _16099_, _16097_, _16096_, _16095_, _16094_, _16093_, _16092_, _16091_, _16090_, _16089_, _16088_, _16086_, _16085_, _16084_, _16083_, _16082_, _16081_, _16080_, _16079_, _16078_, _16077_, _16107_, _16106_, _16105_, _16104_, _16103_, _16102_, _16101_, _16098_, _16087_, _16076_ }) );
  \$mux  #( .WIDTH(32) ) _41638_ ( .A(_stream_conv2d_8_source_29_source_pat_fsm_12), .B(2), .S(_05838_), .Y({ _16164_, _16163_, _16161_, _16160_, _16159_, _16158_, _16157_, _16156_, _16155_, _16154_, _16153_, _16152_, _16150_, _16149_, _16148_, _16147_, _16146_, _16145_, _16144_, _16143_, _16142_, _16141_, _16171_, _16170_, _16169_, _16168_, _16167_, _16166_, _16165_, _16162_, _16151_, _16140_ }) );
  \$mux  #( .WIDTH(32) ) _41639_ ( .A(_stream_conv2d_8_source_29_source_pat_fsm_12), .B(1), .S(_05734_), .Y({ _16196_, _16195_, _16193_, _16192_, _16191_, _16190_, _16189_, _16188_, _16187_, _16186_, _16185_, _16184_, _16182_, _16181_, _16180_, _16179_, _16178_, _16177_, _16176_, _16175_, _16174_, _16173_, _16203_, _16202_, _16201_, _16200_, _16199_, _16198_, _16197_, _16194_, _16183_, _16172_ }) );
  \$mux  #( .WIDTH(32) ) _41645_ ( .A(_stream_conv2d_8_source_28_source_pat_fsm_11), .B(2), .S(_05837_), .Y({ _16260_, _16259_, _16257_, _16256_, _16255_, _16254_, _16253_, _16252_, _16251_, _16250_, _16249_, _16248_, _16246_, _16245_, _16244_, _16243_, _16242_, _16241_, _16240_, _16239_, _16238_, _16237_, _16267_, _16266_, _16265_, _16264_, _16263_, _16262_, _16261_, _16258_, _16247_, _16236_ }) );
  \$mux  #( .WIDTH(32) ) _41646_ ( .A(_stream_conv2d_8_source_28_source_pat_fsm_11), .B(1), .S(_05729_), .Y({ _16292_, _16291_, _16289_, _16288_, _16287_, _16286_, _16285_, _16284_, _16283_, _16282_, _16281_, _16280_, _16278_, _16277_, _16276_, _16275_, _16274_, _16273_, _16272_, _16271_, _16270_, _16269_, _16299_, _16298_, _16297_, _16296_, _16295_, _16294_, _16293_, _16290_, _16279_, _16268_ }) );
  \$mux  #( .WIDTH(32) ) _41652_ ( .A(_stream_conv2d_8_source_27_source_pat_fsm_10), .B(2), .S(_05836_), .Y({ _16356_, _16355_, _16353_, _16352_, _16351_, _16350_, _16349_, _16348_, _16347_, _16346_, _16345_, _16344_, _16342_, _16341_, _16340_, _16339_, _16338_, _16337_, _16336_, _16335_, _16334_, _16333_, _16363_, _16362_, _16361_, _16360_, _16359_, _16358_, _16357_, _16354_, _16343_, _16332_ }) );
  \$mux  #( .WIDTH(32) ) _41653_ ( .A(_stream_conv2d_8_source_27_source_pat_fsm_10), .B(1), .S(_05724_), .Y({ _16388_, _16387_, _16385_, _16384_, _16383_, _16382_, _16381_, _16380_, _16379_, _16378_, _16377_, _16376_, _16374_, _16373_, _16372_, _16371_, _16370_, _16369_, _16368_, _16367_, _16366_, _16365_, _16395_, _16394_, _16393_, _16392_, _16391_, _16390_, _16389_, _16386_, _16375_, _16364_ }) );
  \$mux  #( .WIDTH(32) ) _41657_ ( .A(_stream_conv2d_8_source_26_source_pat_fsm_9), .B(2), .S(_05835_), .Y({ _16452_, _16451_, _16449_, _16448_, _16447_, _16446_, _16445_, _16444_, _16443_, _16442_, _16441_, _16440_, _16438_, _16437_, _16436_, _16435_, _16434_, _16433_, _16432_, _16431_, _16430_, _16429_, _16459_, _16458_, _16457_, _16456_, _16455_, _16454_, _16453_, _16450_, _16439_, _16428_ }) );
  \$mux  #( .WIDTH(32) ) _41658_ ( .A(_stream_conv2d_8_source_26_source_pat_fsm_9), .B(1), .S(_05719_), .Y({ _16484_, _16483_, _16481_, _16480_, _16479_, _16478_, _16477_, _16476_, _16475_, _16474_, _16473_, _16472_, _16470_, _16469_, _16468_, _16467_, _16466_, _16465_, _16464_, _16463_, _16462_, _16461_, _16491_, _16490_, _16489_, _16488_, _16487_, _16486_, _16485_, _16482_, _16471_, _16460_ }) );
  \$mux  #( .WIDTH(32) ) _41662_ ( .A(_stream_conv2d_8_source_25_source_pat_fsm_8), .B(2), .S(_05834_), .Y({ _16548_, _16547_, _16545_, _16544_, _16543_, _16542_, _16541_, _16540_, _16539_, _16538_, _16537_, _16536_, _16534_, _16533_, _16532_, _16531_, _16530_, _16529_, _16528_, _16527_, _16526_, _16525_, _16555_, _16554_, _16553_, _16552_, _16551_, _16550_, _16549_, _16546_, _16535_, _16524_ }) );
  \$mux  #( .WIDTH(32) ) _41663_ ( .A(_stream_conv2d_8_source_25_source_pat_fsm_8), .B(1), .S(_05714_), .Y({ _16580_, _16579_, _16577_, _16576_, _16575_, _16574_, _16573_, _16572_, _16571_, _16570_, _16569_, _16568_, _16566_, _16565_, _16564_, _16563_, _16562_, _16561_, _16560_, _16559_, _16558_, _16557_, _16587_, _16586_, _16585_, _16584_, _16583_, _16582_, _16581_, _16578_, _16567_, _16556_ }) );
  \$mux  #( .WIDTH(32) ) _41667_ ( .A(_stream_conv2d_8_source_24_source_pat_fsm_7), .B(2), .S(_05833_), .Y({ _16644_, _16643_, _16641_, _16640_, _16639_, _16638_, _16637_, _16636_, _16635_, _16634_, _16633_, _16632_, _16630_, _16629_, _16628_, _16627_, _16626_, _16625_, _16624_, _16623_, _16622_, _16621_, _16651_, _16650_, _16649_, _16648_, _16647_, _16646_, _16645_, _16642_, _16631_, _16620_ }) );
  \$mux  #( .WIDTH(32) ) _41668_ ( .A(_stream_conv2d_8_source_24_source_pat_fsm_7), .B(1), .S(_05709_), .Y({ _16676_, _16675_, _16673_, _16672_, _16671_, _16670_, _16669_, _16668_, _16667_, _16666_, _16665_, _16664_, _16662_, _16661_, _16660_, _16659_, _16658_, _16657_, _16656_, _16655_, _16654_, _16653_, _16683_, _16682_, _16681_, _16680_, _16679_, _16678_, _16677_, _16674_, _16663_, _16652_ }) );
  \$mux  #( .WIDTH(32) ) _41672_ ( .A(_stream_conv2d_8_source_23_source_pat_fsm_6), .B(2), .S(_05832_), .Y({ _16740_, _16739_, _16737_, _16736_, _16735_, _16734_, _16733_, _16732_, _16731_, _16730_, _16729_, _16728_, _16726_, _16725_, _16724_, _16723_, _16722_, _16721_, _16720_, _16719_, _16718_, _16717_, _16747_, _16746_, _16745_, _16744_, _16743_, _16742_, _16741_, _16738_, _16727_, _16716_ }) );
  \$mux  #( .WIDTH(32) ) _41673_ ( .A(_stream_conv2d_8_source_23_source_pat_fsm_6), .B(1), .S(_05704_), .Y({ _16772_, _16771_, _16769_, _16768_, _16767_, _16766_, _16765_, _16764_, _16763_, _16762_, _16761_, _16760_, _16758_, _16757_, _16756_, _16755_, _16754_, _16753_, _16752_, _16751_, _16750_, _16749_, _16779_, _16778_, _16777_, _16776_, _16775_, _16774_, _16773_, _16770_, _16759_, _16748_ }) );
  \$mux  #( .WIDTH(32) ) _41677_ ( .A(_stream_conv2d_8_source_22_source_pat_fsm_5), .B(2), .S(_05831_), .Y({ _16836_, _16835_, _16833_, _16832_, _16831_, _16830_, _16829_, _16828_, _16827_, _16826_, _16825_, _16824_, _16822_, _16821_, _16820_, _16819_, _16818_, _16817_, _16816_, _16815_, _16814_, _16813_, _16843_, _16842_, _16841_, _16840_, _16839_, _16838_, _16837_, _16834_, _16823_, _16812_ }) );
  \$mux  #( .WIDTH(32) ) _41678_ ( .A(_stream_conv2d_8_source_22_source_pat_fsm_5), .B(1), .S(_05699_), .Y({ _16868_, _16867_, _16865_, _16864_, _16863_, _16862_, _16861_, _16860_, _16859_, _16858_, _16857_, _16856_, _16854_, _16853_, _16852_, _16851_, _16850_, _16849_, _16848_, _16847_, _16846_, _16845_, _16875_, _16874_, _16873_, _16872_, _16871_, _16870_, _16869_, _16866_, _16855_, _16844_ }) );
  \$mux  #( .WIDTH(32) ) _41682_ ( .A(_stream_conv2d_8_source_21_source_pat_fsm_4), .B(2), .S(_05830_), .Y({ _16932_, _16931_, _16929_, _16928_, _16927_, _16926_, _16925_, _16924_, _16923_, _16922_, _16921_, _16920_, _16918_, _16917_, _16916_, _16915_, _16914_, _16913_, _16912_, _16911_, _16910_, _16909_, _16939_, _16938_, _16937_, _16936_, _16935_, _16934_, _16933_, _16930_, _16919_, _16908_ }) );
  \$mux  #( .WIDTH(32) ) _41683_ ( .A(_stream_conv2d_8_source_21_source_pat_fsm_4), .B(1), .S(_05694_), .Y({ _16964_, _16963_, _16961_, _16960_, _16959_, _16958_, _16957_, _16956_, _16955_, _16954_, _16953_, _16952_, _16950_, _16949_, _16948_, _16947_, _16946_, _16945_, _16944_, _16943_, _16942_, _16941_, _16971_, _16970_, _16969_, _16968_, _16967_, _16966_, _16965_, _16962_, _16951_, _16940_ }) );
  \$mux  #( .WIDTH(32) ) _41687_ ( .A(_stream_conv2d_8_source_20_source_pat_fsm_3), .B(2), .S(_05829_), .Y({ _17028_, _17027_, _17025_, _17024_, _17023_, _17022_, _17021_, _17020_, _17019_, _17018_, _17017_, _17016_, _17014_, _17013_, _17012_, _17011_, _17010_, _17009_, _17008_, _17007_, _17006_, _17005_, _17035_, _17034_, _17033_, _17032_, _17031_, _17030_, _17029_, _17026_, _17015_, _17004_ }) );
  \$mux  #( .WIDTH(32) ) _41688_ ( .A(_stream_conv2d_8_source_20_source_pat_fsm_3), .B(1), .S(_05689_), .Y({ _17060_, _17059_, _17057_, _17056_, _17055_, _17054_, _17053_, _17052_, _17051_, _17050_, _17049_, _17048_, _17046_, _17045_, _17044_, _17043_, _17042_, _17041_, _17040_, _17039_, _17038_, _17037_, _17067_, _17066_, _17065_, _17064_, _17063_, _17062_, _17061_, _17058_, _17047_, _17036_ }) );
  \$mux  #( .WIDTH(32) ) _41692_ ( .A(_stream_conv2d_8_source_19_source_pat_fsm_2), .B(2), .S(_05828_), .Y({ _17124_, _17123_, _17121_, _17120_, _17119_, _17118_, _17117_, _17116_, _17115_, _17114_, _17113_, _17112_, _17110_, _17109_, _17108_, _17107_, _17106_, _17105_, _17104_, _17103_, _17102_, _17101_, _17131_, _17130_, _17129_, _17128_, _17127_, _17126_, _17125_, _17122_, _17111_, _17100_ }) );
  \$mux  #( .WIDTH(32) ) _41693_ ( .A(_stream_conv2d_8_source_19_source_pat_fsm_2), .B(1), .S(_05684_), .Y({ _17156_, _17155_, _17153_, _17152_, _17151_, _17150_, _17149_, _17148_, _17147_, _17146_, _17145_, _17144_, _17142_, _17141_, _17140_, _17139_, _17138_, _17137_, _17136_, _17135_, _17134_, _17133_, _17163_, _17162_, _17161_, _17160_, _17159_, _17158_, _17157_, _17154_, _17143_, _17132_ }) );
  \$mux  #( .WIDTH(32) ) _41697_ ( .A(_stream_conv2d_8_source_8_source_pat_fsm_1), .B(2), .S(_05827_), .Y({ _17220_, _17219_, _17217_, _17216_, _17215_, _17214_, _17213_, _17212_, _17211_, _17210_, _17209_, _17208_, _17206_, _17205_, _17204_, _17203_, _17202_, _17201_, _17200_, _17199_, _17198_, _17197_, _17227_, _17226_, _17225_, _17224_, _17223_, _17222_, _17221_, _17218_, _17207_, _17196_ }) );
  \$mux  #( .WIDTH(32) ) _41698_ ( .A(_stream_conv2d_8_source_8_source_pat_fsm_1), .B(1), .S(_05679_), .Y({ _17252_, _17251_, _17249_, _17248_, _17247_, _17246_, _17245_, _17244_, _17243_, _17242_, _17241_, _17240_, _17238_, _17237_, _17236_, _17235_, _17234_, _17233_, _17232_, _17231_, _17230_, _17229_, _17259_, _17258_, _17257_, _17256_, _17255_, _17254_, _17253_, _17250_, _17239_, _17228_ }) );
  \$mux  #( .WIDTH(32) ) _41704_ ( .A(_stream_conv2d_8_source_6_source_pat_fsm_0), .B(2), .S(_05826_), .Y({ _17316_, _17315_, _17313_, _17312_, _17311_, _17310_, _17309_, _17308_, _17307_, _17306_, _17305_, _17304_, _17302_, _17301_, _17300_, _17299_, _17298_, _17297_, _17296_, _17295_, _17294_, _17293_, _17323_, _17322_, _17321_, _17320_, _17319_, _17318_, _17317_, _17314_, _17303_, _17292_ }) );
  \$mux  #( .WIDTH(32) ) _41705_ ( .A(_stream_conv2d_8_source_6_source_pat_fsm_0), .B(1), .S(_05674_), .Y({ _17348_, _17347_, _17345_, _17344_, _17343_, _17342_, _17341_, _17340_, _17339_, _17338_, _17337_, _17336_, _17334_, _17333_, _17332_, _17331_, _17330_, _17329_, _17328_, _17327_, _17326_, _17325_, _17355_, _17354_, _17353_, _17352_, _17351_, _17350_, _17349_, _17346_, _17335_, _17324_ }) );
  \$mux  #( .WIDTH(9) ) _41707_ ( .A({ conv2d_8_stream_pad_mask_2_2, conv2d_8_stream_pad_mask_2_1, conv2d_8_stream_pad_mask_2_0, conv2d_8_stream_pad_mask_1_2, conv2d_8_stream_pad_mask_1_1, conv2d_8_stream_pad_mask_1_0, conv2d_8_stream_pad_mask_0_2, conv2d_8_stream_pad_mask_0_1, conv2d_8_stream_pad_mask_0_0 }), .B(conv2d_8_stream_pad_masks), .S(_05100_), .Y(_22620_) );
  \$mux  #( .WIDTH(32) ) _41709_ ( .A(conv2d_8_och_count), .B(conv2d_8_och_count_buf), .S(_05102_), .Y(_22621_) );
  \$mux  #( .WIDTH(2) ) _41711_ ( .A(conv2d_8_row_select), .B(conv2d_8_row_select_buf), .S(_05102_), .Y(_22622_) );
  \$mux  #( .WIDTH(32) ) _41713_ ( .A(conv2d_8_row_count), .B(conv2d_8_row_count_buf), .S(_05102_), .Y(_22623_) );
  \$mux  #( .WIDTH(32) ) _41715_ ( .A(conv2d_8_out_page_comp_offset), .B(conv2d_8_out_page_comp_offset_buf), .S(_05102_), .Y(_22624_) );
  \$mux  #( .WIDTH(32) ) _41717_ ( .A(conv2d_8_act_page_comp_offset_2), .B(conv2d_8_act_page_comp_offset_buf_2), .S(_05102_), .Y(_22625_) );
  \$mux  #( .WIDTH(32) ) _41719_ ( .A(conv2d_8_act_page_comp_offset_1), .B(conv2d_8_act_page_comp_offset_buf_1), .S(_05102_), .Y(_22626_) );
  \$mux  #( .WIDTH(32) ) _41721_ ( .A(conv2d_8_act_page_comp_offset_0), .B(conv2d_8_act_page_comp_offset_buf_0), .S(_05102_), .Y(_22627_) );
  \$mux  #( .WIDTH(32) ) _41723_ ( .A(conv2d_8_filter_page_comp_offset), .B(conv2d_8_filter_page_comp_offset_buf), .S(_05102_), .Y(_22628_) );
  \$mux  #( .WIDTH(32) ) _41725_ ( .A(2), .B(0), .S(_05242_), .Y({ _17380_, _17379_, _17377_, _17376_, _17375_, _17374_, _17373_, _17372_, _17371_, _17370_, _17369_, _17368_, _17366_, _17365_, _17364_, _17363_, _17362_, _17361_, _17360_, _17359_, _17358_, _17357_, _17387_, _17386_, _17385_, _17384_, _17383_, _17382_, _17381_, _17378_, _17367_, _17356_ }) );
  \$mux  #( .WIDTH(32) ) _41726_ ( .A(5), .B(conv2d_8_comp_fsm), .S(_stream_conv2d_8_source_busy), .Y({ _17444_, _17443_, _17441_, _17440_, _17439_, _17438_, _17437_, _17436_, _17435_, _17434_, _17433_, _17432_, _17430_, _17429_, _17428_, _17427_, _17426_, _17425_, _17424_, _17423_, _17422_, _17421_, _17451_, _17450_, _17449_, _17448_, _17447_, _17446_, _17445_, _17442_, _17431_, _17420_ }) );
  \$mux  #( .WIDTH(32) ) _41727_ ( .A(conv2d_8_comp_fsm), .B(1), .S(_05824_), .Y({ _17476_, _17475_, _17473_, _17472_, _17471_, _17470_, _17469_, _17468_, _17467_, _17466_, _17465_, _17464_, _17462_, _17461_, _17460_, _17459_, _17458_, _17457_, _17456_, _17455_, _17454_, _17453_, _17483_, _17482_, _17481_, _17480_, _17479_, _17478_, _17477_, _17474_, _17463_, _17452_ }) );
  \$mux  #( .WIDTH(32) ) _41729_ ( .A(_22296_), .B(0), .S(_05242_), .Y({ _17508_, _17507_, _17505_, _17504_, _17503_, _17502_, _17501_, _17500_, _17499_, _17498_, _17497_, _17496_, _17494_, _17493_, _17492_, _17491_, _17490_, _17489_, _17488_, _17487_, _17486_, _17485_, _17515_, _17514_, _17513_, _17512_, _17511_, _17510_, _17509_, _17506_, _17495_, _17484_ }) );
  \$mux  #( .WIDTH(32) ) _41731_ ( .A(conv2d_8_stream_act_local_8), .B(_22295_), .S(_17548_), .Y(_22631_) );
  \$mux  #( .WIDTH(32) ) _41732_ ( .A(_22631_), .B(0), .S(_05242_), .Y(_22632_) );
  \$mux  #( .WIDTH(32) ) _41733_ ( .A(_22632_), .B({ cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset }), .S(_05825_), .Y({ _17573_, _17572_, _17570_, _17569_, _17568_, _17567_, _17566_, _17565_, _17564_, _17563_, _17562_, _17561_, _17559_, _17558_, _17557_, _17556_, _17555_, _17554_, _17553_, _17552_, _17551_, _17550_, _17580_, _17579_, _17578_, _17577_, _17576_, _17575_, _17574_, _17571_, _17560_, _17549_ }) );
  \$mux  #( .WIDTH(32) ) _41735_ ( .A(conv2d_8_stream_act_local_7), .B(_22294_), .S(_17645_), .Y(_22634_) );
  \$mux  #( .WIDTH(32) ) _41736_ ( .A(_22634_), .B(0), .S(_05242_), .Y({ _17670_, _17669_, _17667_, _17666_, _17665_, _17664_, _17663_, _17662_, _17661_, _17660_, _17659_, _17658_, _17656_, _17655_, _17654_, _17653_, _17652_, _17651_, _17650_, _17649_, _17648_, _17647_, _17677_, _17676_, _17675_, _17674_, _17673_, _17672_, _17671_, _17668_, _17657_, _17646_ }) );
  \$mux  #( .WIDTH(32) ) _41738_ ( .A(conv2d_8_stream_act_local_6), .B(_22293_), .S(_17710_), .Y(_22636_) );
  \$mux  #( .WIDTH(32) ) _41739_ ( .A(_22636_), .B(0), .S(_05242_), .Y({ _17735_, _17734_, _17732_, _17731_, _17730_, _17729_, _17728_, _17727_, _17726_, _17725_, _17724_, _17723_, _17721_, _17720_, _17719_, _17718_, _17717_, _17716_, _17715_, _17714_, _17713_, _17712_, _17742_, _17741_, _17740_, _17739_, _17738_, _17737_, _17736_, _17733_, _17722_, _17711_ }) );
  \$mux  #( .WIDTH(32) ) _41741_ ( .A(conv2d_8_stream_act_local_5), .B(_22292_), .S(_17548_), .Y(_22638_) );
  \$mux  #( .WIDTH(32) ) _41742_ ( .A(_22638_), .B(0), .S(_05242_), .Y(_22639_) );
  \$mux  #( .WIDTH(32) ) _41743_ ( .A(_22639_), .B({ cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset }), .S(_05825_), .Y({ _17799_, _17798_, _17796_, _17795_, _17794_, _17793_, _17792_, _17791_, _17790_, _17789_, _17788_, _17787_, _17785_, _17784_, _17783_, _17782_, _17781_, _17780_, _17779_, _17778_, _17777_, _17776_, _17806_, _17805_, _17804_, _17803_, _17802_, _17801_, _17800_, _17797_, _17786_, _17775_ }) );
  \$mux  #( .WIDTH(32) ) _41745_ ( .A(conv2d_8_stream_act_local_4), .B(_22291_), .S(_17645_), .Y(_22641_) );
  \$mux  #( .WIDTH(32) ) _41746_ ( .A(_22641_), .B(0), .S(_05242_), .Y({ _17863_, _17862_, _17860_, _17859_, _17858_, _17857_, _17856_, _17855_, _17854_, _17853_, _17852_, _17851_, _17849_, _17848_, _17847_, _17846_, _17845_, _17844_, _17843_, _17842_, _17841_, _17840_, _17870_, _17869_, _17868_, _17867_, _17866_, _17865_, _17864_, _17861_, _17850_, _17839_ }) );
  \$mux  #( .WIDTH(32) ) _41748_ ( .A(conv2d_8_stream_act_local_3), .B(_22290_), .S(_17710_), .Y(_22643_) );
  \$mux  #( .WIDTH(32) ) _41749_ ( .A(_22643_), .B(0), .S(_05242_), .Y({ _17927_, _17926_, _17924_, _17923_, _17922_, _17921_, _17920_, _17919_, _17918_, _17917_, _17916_, _17915_, _17913_, _17912_, _17911_, _17910_, _17909_, _17908_, _17907_, _17906_, _17905_, _17904_, _17934_, _17933_, _17932_, _17931_, _17930_, _17929_, _17928_, _17925_, _17914_, _17903_ }) );
  \$mux  #( .WIDTH(32) ) _41751_ ( .A(conv2d_8_stream_act_local_2), .B(_22289_), .S(_17548_), .Y(_22645_) );
  \$mux  #( .WIDTH(32) ) _41752_ ( .A(_22645_), .B(0), .S(_05242_), .Y(_22646_) );
  \$mux  #( .WIDTH(32) ) _41753_ ( .A(_22646_), .B({ cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset }), .S(_05825_), .Y({ _17991_, _17990_, _17988_, _17987_, _17986_, _17985_, _17984_, _17983_, _17982_, _17981_, _17980_, _17979_, _17977_, _17976_, _17975_, _17974_, _17973_, _17972_, _17971_, _17970_, _17969_, _17968_, _17998_, _17997_, _17996_, _17995_, _17994_, _17993_, _17992_, _17989_, _17978_, _17967_ }) );
  \$mux  #( .WIDTH(32) ) _41754_ ( .A(0), .B({ cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset[3], cparam_conv2d_8_stream_act_local_large_offset }), .S(cparam_conv2d_8_pad_col_left), .Y({ _17637_, _17636_, _17634_, _17633_, _17632_, _17631_, _17630_, _17629_, _17628_, _17627_, _17626_, _17625_, _17623_, _17622_, _17621_, _17620_, _17619_, _17618_, _17617_, _17616_, _17615_, _17614_, _17644_, _17643_, _17642_, _17641_, _17640_, _17639_, _17638_, _17635_, _17624_, _17613_ }) );
  \$mux  #( .WIDTH(32) ) _41756_ ( .A(conv2d_8_stream_act_local_1), .B(_22288_), .S(_17645_), .Y(_22648_) );
  \$mux  #( .WIDTH(32) ) _41757_ ( .A(_22648_), .B(0), .S(_05242_), .Y({ _18055_, _18054_, _18052_, _18051_, _18050_, _18049_, _18048_, _18047_, _18046_, _18045_, _18044_, _18043_, _18041_, _18040_, _18039_, _18038_, _18037_, _18036_, _18035_, _18034_, _18033_, _18032_, _18062_, _18061_, _18060_, _18059_, _18058_, _18057_, _18056_, _18053_, _18042_, _18031_ }) );
  \$mux  #( .WIDTH(32) ) _41759_ ( .A(conv2d_8_stream_act_local_0), .B(_22287_), .S(_17710_), .Y(_22650_) );
  \$mux  #( .WIDTH(32) ) _41760_ ( .A(_22650_), .B(0), .S(_05242_), .Y({ _18119_, _18118_, _18116_, _18115_, _18114_, _18113_, _18112_, _18111_, _18110_, _18109_, _18108_, _18107_, _18105_, _18104_, _18103_, _18102_, _18101_, _18100_, _18099_, _18098_, _18097_, _18096_, _18126_, _18125_, _18124_, _18123_, _18122_, _18121_, _18120_, _18117_, _18106_, _18095_ }) );
  \$mux  #( .WIDTH(2) ) _41762_ ( .A(_22298_), .B(_26326_), .S(_05243_), .Y(_22652_) );
  \$mux  #( .WIDTH(2) ) _41763_ ( .A(_22652_), .B(cparam_conv2d_8_col_select_initval), .S(_05242_), .Y({ _18160_, _18159_ }) );
  \$mux  #( .WIDTH(32) ) _41765_ ( .A(_22297_), .B(0), .S(_05242_), .Y({ _18187_, _18186_, _18184_, _18183_, _18182_, _18181_, _18180_, _18179_, _18178_, _18177_, _18176_, _18175_, _18173_, _18172_, _18171_, _18170_, _18169_, _18168_, _18167_, _18166_, _18165_, _18164_, _18194_, _18193_, _18192_, _18191_, _18190_, _18189_, _18188_, _18185_, _18174_, _18163_ }) );
  \$mux  #( .WIDTH(32) ) _41767_ ( .A(conv2d_8_sync_comp_count), .B(_22286_), .S(_stream_conv2d_8_end_flag), .Y(_22655_) );
  \$mux  #( .WIDTH(32) ) _41768_ ( .A(0), .B(_22655_), .S(_05129_), .Y(_22656_) );
  \$mux  #( .WIDTH(32) ) _41770_ ( .A({ 27'h0000000, cparam_conv2d_8_bias_num }), .B(conv2d_8_next_stream_num_ops), .S(_05102_), .Y(_22657_) );
  \$mux  #( .WIDTH(9) ) _41772_ ( .A(req_block_size_270), .B({ 6'h00, cparam_conv2d_8_inc_act_laddr_large[4:2] }), .S(set_req_271), .Y(_22658_) );
  \$mux  #( .WIDTH(9) ) _41774_ ( .A(req_block_size_213), .B({ 6'h00, cparam_conv2d_8_inc_act_laddr_large[4:2] }), .S(set_req_214), .Y(_22659_) );
  \$mux  #( .WIDTH(9) ) _41776_ ( .A(req_block_size_156), .B({ 6'h00, cparam_conv2d_8_inc_act_laddr_large[4:2] }), .S(set_req_157), .Y(_22660_) );
  \$mux  #( .WIDTH(9) ) _41778_ ( .A(req_block_size_27), .B({ 6'h00, cparam_conv2d_8_inc_act_laddr_large[4:2] }), .S(set_req_28), .Y(_22661_) );
  \$mux  #( .WIDTH(1) ) _41780_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_9_1), .S(_05106_), .Y(_22662_) );
  \$mux  #( .WIDTH(1) ) _41782_ ( .A(_wvalid_974), .B(1'h0), .S(__maxi_read_fsm_cond_3_9_1), .Y(_22663_) );
  \$mux  #( .WIDTH(1) ) _41783_ ( .A(_22663_), .B(_wvalid_974), .S(_05104_), .Y(_22664_) );
  \$mux  #( .WIDTH(1) ) _41784_ ( .A(_22664_), .B(1'h1), .S(_05821_), .Y(_22665_) );
  \$mux  #( .WIDTH(1) ) _41785_ ( .A(_22665_), .B(_22664_), .S(_05106_), .Y(_22666_) );
  \$mux  #( .WIDTH(32) ) _41787_ ( .A(_wdata_973), .B(maxi_rdata), .S(_05821_), .Y(_22667_) );
  \$mux  #( .WIDTH(32) ) _41788_ ( .A(_22667_), .B(_wdata_973), .S(_05106_), .Y(_22668_) );
  \$mux  #( .WIDTH(1) ) _41790_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_8_1), .S(_05106_), .Y(_22669_) );
  \$mux  #( .WIDTH(1) ) _41792_ ( .A(_wvalid_963), .B(1'h0), .S(__maxi_read_fsm_cond_3_8_1), .Y(_22670_) );
  \$mux  #( .WIDTH(1) ) _41793_ ( .A(_22670_), .B(_wvalid_963), .S(_05104_), .Y(_22671_) );
  \$mux  #( .WIDTH(1) ) _41794_ ( .A(_22671_), .B(1'h1), .S(_05820_), .Y(_22672_) );
  \$mux  #( .WIDTH(1) ) _41795_ ( .A(_22672_), .B(_22671_), .S(_05106_), .Y(_22673_) );
  \$mux  #( .WIDTH(32) ) _41797_ ( .A(_wdata_962), .B(maxi_rdata), .S(_05820_), .Y(_22674_) );
  \$mux  #( .WIDTH(32) ) _41798_ ( .A(_22674_), .B(_wdata_962), .S(_05106_), .Y(_22675_) );
  \$mux  #( .WIDTH(1) ) _41800_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_7_1), .S(_05106_), .Y(_22676_) );
  \$mux  #( .WIDTH(1) ) _41802_ ( .A(_wvalid_852), .B(1'h0), .S(__maxi_read_fsm_cond_3_7_1), .Y(_22677_) );
  \$mux  #( .WIDTH(1) ) _41803_ ( .A(_22677_), .B(_wvalid_852), .S(_05104_), .Y(_22678_) );
  \$mux  #( .WIDTH(1) ) _41804_ ( .A(_22678_), .B(1'h1), .S(_05819_), .Y(_22679_) );
  \$mux  #( .WIDTH(1) ) _41805_ ( .A(_22679_), .B(_22678_), .S(_05106_), .Y(_22680_) );
  \$mux  #( .WIDTH(32) ) _41807_ ( .A(_wdata_851), .B(maxi_rdata), .S(_05819_), .Y(_22681_) );
  \$mux  #( .WIDTH(32) ) _41808_ ( .A(_22681_), .B(_wdata_851), .S(_05106_), .Y(_22682_) );
  \$mux  #( .WIDTH(1) ) _41810_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_6_1), .S(_05106_), .Y(_22683_) );
  \$mux  #( .WIDTH(1) ) _41812_ ( .A(_wvalid_274), .B(1'h0), .S(__maxi_read_fsm_cond_3_6_1), .Y(_22684_) );
  \$mux  #( .WIDTH(1) ) _41813_ ( .A(_22684_), .B(_wvalid_274), .S(_05104_), .Y(_22685_) );
  \$mux  #( .WIDTH(1) ) _41814_ ( .A(_22685_), .B(1'h1), .S(_05818_), .Y(_22686_) );
  \$mux  #( .WIDTH(1) ) _41815_ ( .A(_22686_), .B(_22685_), .S(_05106_), .Y(_22687_) );
  \$mux  #( .WIDTH(32) ) _41817_ ( .A(_wdata_273), .B(maxi_rdata), .S(_05818_), .Y(_22688_) );
  \$mux  #( .WIDTH(32) ) _41818_ ( .A(_22688_), .B(_wdata_273), .S(_05106_), .Y(_22689_) );
  \$mux  #( .WIDTH(1) ) _41820_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_5_1), .S(_05106_), .Y(_22690_) );
  \$mux  #( .WIDTH(1) ) _41822_ ( .A(_wvalid_217), .B(1'h0), .S(__maxi_read_fsm_cond_3_5_1), .Y(_22691_) );
  \$mux  #( .WIDTH(1) ) _41823_ ( .A(_22691_), .B(_wvalid_217), .S(_05104_), .Y(_22692_) );
  \$mux  #( .WIDTH(1) ) _41824_ ( .A(_22692_), .B(1'h1), .S(_05817_), .Y(_22693_) );
  \$mux  #( .WIDTH(1) ) _41825_ ( .A(_22693_), .B(_22692_), .S(_05106_), .Y(_22694_) );
  \$mux  #( .WIDTH(32) ) _41827_ ( .A(_wdata_216), .B(maxi_rdata), .S(_05817_), .Y(_22695_) );
  \$mux  #( .WIDTH(32) ) _41828_ ( .A(_22695_), .B(_wdata_216), .S(_05106_), .Y(_22696_) );
  \$mux  #( .WIDTH(1) ) _41830_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_4_1), .S(_05106_), .Y(_22697_) );
  \$mux  #( .WIDTH(1) ) _41832_ ( .A(_wvalid_160), .B(1'h0), .S(__maxi_read_fsm_cond_3_4_1), .Y(_22698_) );
  \$mux  #( .WIDTH(1) ) _41833_ ( .A(_22698_), .B(_wvalid_160), .S(_05104_), .Y(_22699_) );
  \$mux  #( .WIDTH(1) ) _41834_ ( .A(_22699_), .B(1'h1), .S(_05816_), .Y(_22700_) );
  \$mux  #( .WIDTH(1) ) _41835_ ( .A(_22700_), .B(_22699_), .S(_05106_), .Y(_22701_) );
  \$mux  #( .WIDTH(32) ) _41837_ ( .A(_wdata_159), .B(maxi_rdata), .S(_05816_), .Y(_22702_) );
  \$mux  #( .WIDTH(32) ) _41838_ ( .A(_22702_), .B(_wdata_159), .S(_05106_), .Y(_22703_) );
  \$mux  #( .WIDTH(1) ) _41840_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_3_1), .S(_05106_), .Y(_22704_) );
  \$mux  #( .WIDTH(1) ) _41842_ ( .A(_wvalid_31), .B(1'h0), .S(__maxi_read_fsm_cond_3_3_1), .Y(_22705_) );
  \$mux  #( .WIDTH(1) ) _41843_ ( .A(_22705_), .B(_wvalid_31), .S(_05104_), .Y(_22706_) );
  \$mux  #( .WIDTH(1) ) _41844_ ( .A(_22706_), .B(1'h1), .S(_05815_), .Y(_22707_) );
  \$mux  #( .WIDTH(1) ) _41845_ ( .A(_22707_), .B(_22706_), .S(_05106_), .Y(_22708_) );
  \$mux  #( .WIDTH(32) ) _41847_ ( .A(_wdata_30), .B(maxi_rdata), .S(_05815_), .Y(_22709_) );
  \$mux  #( .WIDTH(32) ) _41848_ ( .A(_22709_), .B(_wdata_30), .S(_05106_), .Y(_22710_) );
  \$mux  #( .WIDTH(1) ) _41850_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_2_1), .S(_05106_), .Y(_22711_) );
  \$mux  #( .WIDTH(1) ) _41852_ ( .A(_wvalid_18), .B(1'h0), .S(__maxi_read_fsm_cond_3_2_1), .Y(_22712_) );
  \$mux  #( .WIDTH(1) ) _41853_ ( .A(_22712_), .B(_wvalid_18), .S(_05104_), .Y(_22713_) );
  \$mux  #( .WIDTH(1) ) _41854_ ( .A(_22713_), .B(1'h1), .S(_05814_), .Y(_22714_) );
  \$mux  #( .WIDTH(1) ) _41855_ ( .A(_22714_), .B(_22713_), .S(_05106_), .Y(_22715_) );
  \$mux  #( .WIDTH(32) ) _41857_ ( .A(_wdata_17), .B(maxi_rdata), .S(_05814_), .Y(_22716_) );
  \$mux  #( .WIDTH(32) ) _41858_ ( .A(_22716_), .B(_wdata_17), .S(_05106_), .Y(_22717_) );
  \$mux  #( .WIDTH(1) ) _41860_ ( .A(1'h1), .B(__maxi_read_fsm_cond_4_1_1), .S(_05105_), .Y(_22718_) );
  \$mux  #( .WIDTH(1) ) _41862_ ( .A(axim_flag_15), .B(1'h0), .S(__maxi_read_fsm_cond_4_1_1), .Y(_22719_) );
  \$mux  #( .WIDTH(1) ) _41863_ ( .A(_22719_), .B(axim_flag_15), .S(_05103_), .Y(_22720_) );
  \$mux  #( .WIDTH(1) ) _41864_ ( .A(1'h1), .B(_22720_), .S(_05105_), .Y(_22721_) );
  \$mux  #( .WIDTH(1) ) _41866_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_0_1), .S(_05106_), .Y(_22722_) );
  \$mux  #( .WIDTH(1) ) _41869_ ( .A(_wvalid_11), .B(1'h0), .S(__maxi_read_fsm_cond_3_0_1), .Y(_22723_) );
  \$mux  #( .WIDTH(1) ) _41870_ ( .A(_22723_), .B(_wvalid_11), .S(_05104_), .Y(_22724_) );
  \$mux  #( .WIDTH(1) ) _41871_ ( .A(_22724_), .B(1'h1), .S(_05812_), .Y(_22725_) );
  \$mux  #( .WIDTH(1) ) _41872_ ( .A(_22725_), .B(_22724_), .S(_05106_), .Y(_22726_) );
  \$mux  #( .WIDTH(32) ) _41874_ ( .A(_wdata_10), .B(maxi_rdata), .S(_05812_), .Y(_22727_) );
  \$mux  #( .WIDTH(32) ) _41875_ ( .A(_22727_), .B(_wdata_10), .S(_05106_), .Y(_22728_) );
  \$mux  #( .WIDTH(33) ) _41877_ ( .A(_26325_), .B(_26324_), .S(_05241_), .Y(_22729_) );
  \$mux  #( .WIDTH(33) ) _41878_ ( .A(_22729_), .B(33'h000000000), .S(_05262_), .Y(_22730_) );
  \$mux  #( .WIDTH(33) ) _41879_ ( .A(_22730_), .B(_26324_), .S(_05811_), .Y({ _18252_, _18251_, _18250_, _18248_, _18247_, _18246_, _18245_, _18244_, _18243_, _18242_, _18241_, _18240_, _18239_, _18237_, _18236_, _18235_, _18234_, _18233_, _18232_, _18231_, _18230_, _18229_, _18228_, _18259_, _18258_, _18257_, _18256_, _18255_, _18254_, _18253_, _18249_, _18238_, _18227_ }) );
  \$mux  #( .WIDTH(33) ) _41880_ ( .A(_maxi_read_rest_size), .B(_maxi_read_size), .S(_maxi_read_start), .Y({ _18318_, _18317_, _18316_, _18314_, _18313_, _18312_, _18311_, _18310_, _18309_, _18308_, _18307_, _18306_, _18305_, _18303_, _18302_, _18301_, _18300_, _18299_, _18298_, _18297_, _18296_, _18295_, _18294_, _18325_, _18324_, _18323_, _18322_, _18321_, _18320_, _18319_, _18315_, _18304_, _18293_ }) );
  \$mux  #( .WIDTH(33) ) _41882_ ( .A(33'h000000100), .B({ 2'h0, _25922_[30:0] }), .S(_05241_), .Y(_22732_) );
  \$mux  #( .WIDTH(33) ) _41883_ ( .A(_22732_), .B(_maxi_read_rest_size), .S(_05262_), .Y(_22733_) );
  \$mux  #( .WIDTH(33) ) _41884_ ( .A(_22733_), .B({ 2'h0, _25922_[30:0] }), .S(_05811_), .Y(_22734_) );
  \$mux  #( .WIDTH(33) ) _41885_ ( .A(_22734_), .B(_maxi_read_cur_size), .S(_05107_), .Y(_22735_) );
  \$mux  #( .WIDTH(32) ) _41887_ ( .A(_maxi_read_cur_global_addr), .B(_22285_[31:0]), .S(_05813_), .Y({ _18350_, _18349_, _18347_, _18346_, _18345_, _18344_, _18343_, _18342_, _18341_, _18340_, _18339_, _18338_, _18336_, _18335_, _18334_, _18333_, _18332_, _18331_, _18330_, _18329_, _18328_, _18327_, _18357_, _18356_, _18355_, _18354_, _18353_, _18352_, _18351_, _18348_, _18337_, _18326_ }) );
  \$mux  #( .WIDTH(32) ) _41888_ ( .A(_maxi_read_cur_global_addr), .B({ _22284_[31:2], 2'h0 }), .S(_maxi_read_start), .Y({ _18414_, _18413_, _18411_, _18410_, _18409_, _18408_, _18407_, _18406_, _18405_, _18404_, _18403_, _18402_, _18400_, _18399_, _18398_, _18397_, _18396_, _18395_, _18394_, _18393_, _18392_, _18391_, _18421_, _18420_, _18419_, _18418_, _18417_, _18416_, _18415_, _18412_, _18401_, _18390_ }) );
  \$mux  #( .WIDTH(32) ) _41890_ ( .A(_maxi_read_fsm), .B(1), .S(_05822_), .Y(_22738_) );
  \$mux  #( .WIDTH(32) ) _41891_ ( .A(_22738_), .B(4), .S(_05823_), .Y({ _18478_, _18477_, _18475_, _18474_, _18473_, _18472_, _18471_, _18470_, _18469_, _18468_, _18467_, _18466_, _18464_, _18463_, _18462_, _18461_, _18460_, _18459_, _18458_, _18457_, _18456_, _18455_, _18485_, _18484_, _18483_, _18482_, _18481_, _18480_, _18479_, _18476_, _18465_, _18454_ }) );
  \$mux  #( .WIDTH(32) ) _41892_ ( .A(_maxi_read_fsm), .B(3), .S(_05864_), .Y({ _18510_, _18509_, _18507_, _18506_, _18505_, _18504_, _18503_, _18502_, _18501_, _18500_, _18499_, _18498_, _18496_, _18495_, _18494_, _18493_, _18492_, _18491_, _18490_, _18489_, _18488_, _18487_, _18517_, _18516_, _18515_, _18514_, _18513_, _18512_, _18511_, _18508_, _18497_, _18486_ }) );
  \$mux  #( .WIDTH(32) ) _41893_ ( .A(_maxi_read_fsm), .B(1), .S(_05671_), .Y(_22739_) );
  \$mux  #( .WIDTH(32) ) _41894_ ( .A(_22739_), .B(1), .S(_05423_), .Y(_22740_) );
  \$mux  #( .WIDTH(32) ) _41895_ ( .A(_22740_), .B(1), .S(_05459_), .Y(_22741_) );
  \$mux  #( .WIDTH(32) ) _41896_ ( .A(_22741_), .B(1), .S(_05557_), .Y(_22742_) );
  \$mux  #( .WIDTH(32) ) _41897_ ( .A(_22742_), .B(1), .S(_05586_), .Y(_22743_) );
  \$mux  #( .WIDTH(32) ) _41898_ ( .A(_22743_), .B(1), .S(_05615_), .Y(_22744_) );
  \$mux  #( .WIDTH(32) ) _41899_ ( .A(_22744_), .B(1), .S(_05473_), .Y(_22745_) );
  \$mux  #( .WIDTH(32) ) _41900_ ( .A(_22745_), .B(1), .S(_05414_), .Y(_22746_) );
  \$mux  #( .WIDTH(32) ) _41901_ ( .A(_22746_), .B(1), .S(_05548_), .Y({ _18542_, _18541_, _18539_, _18538_, _18537_, _18536_, _18535_, _18534_, _18533_, _18532_, _18531_, _18530_, _18528_, _18527_, _18526_, _18525_, _18524_, _18523_, _18522_, _18521_, _18520_, _18519_, _18549_, _18548_, _18547_, _18546_, _18545_, _18544_, _18543_, _18540_, _18529_, _18518_ }) );
  \$mux  #( .WIDTH(1) ) _41903_ ( .A(1'h1), .B(_control_conv2d_8_cond_48_10_1), .S(_05120_), .Y(_22747_) );
  \$mux  #( .WIDTH(1) ) _41905_ ( .A(axim_flag_798), .B(1'h0), .S(_control_conv2d_8_cond_48_10_1), .Y(_22748_) );
  \$mux  #( .WIDTH(1) ) _41906_ ( .A(_22748_), .B(axim_flag_798), .S(_05108_), .Y(_22749_) );
  \$mux  #( .WIDTH(1) ) _41907_ ( .A(1'h1), .B(_22749_), .S(_05120_), .Y(_22750_) );
  \$mux  #( .WIDTH(1) ) _41909_ ( .A(1'h1), .B(_control_conv2d_8_cond_38_9_1), .S(_05121_), .Y(_22751_) );
  \$mux  #( .WIDTH(1) ) _41911_ ( .A(axim_flag_272), .B(1'h0), .S(_control_conv2d_8_cond_38_9_1), .Y(_22752_) );
  \$mux  #( .WIDTH(1) ) _41912_ ( .A(_22752_), .B(axim_flag_272), .S(_05109_), .Y(_22753_) );
  \$mux  #( .WIDTH(1) ) _41913_ ( .A(1'h1), .B(_22753_), .S(_05121_), .Y(_22754_) );
  \$mux  #( .WIDTH(1) ) _41915_ ( .A(1'h1), .B(_control_conv2d_8_cond_37_8_1), .S(_05122_), .Y(_22755_) );
  \$mux  #( .WIDTH(1) ) _41917_ ( .A(set_req_271), .B(1'h0), .S(_control_conv2d_8_cond_37_8_1), .Y(_22756_) );
  \$mux  #( .WIDTH(1) ) _41918_ ( .A(_22756_), .B(set_req_271), .S(_05110_), .Y(_22757_) );
  \$mux  #( .WIDTH(1) ) _41919_ ( .A(1'h1), .B(_22757_), .S(_05122_), .Y(_22758_) );
  \$mux  #( .WIDTH(1) ) _41921_ ( .A(1'h1), .B(_control_conv2d_8_cond_31_7_1), .S(_05123_), .Y(_22759_) );
  \$mux  #( .WIDTH(1) ) _41923_ ( .A(axim_flag_215), .B(1'h0), .S(_control_conv2d_8_cond_31_7_1), .Y(_22760_) );
  \$mux  #( .WIDTH(1) ) _41924_ ( .A(_22760_), .B(axim_flag_215), .S(_05111_), .Y(_22761_) );
  \$mux  #( .WIDTH(1) ) _41925_ ( .A(1'h1), .B(_22761_), .S(_05123_), .Y(_22762_) );
  \$mux  #( .WIDTH(1) ) _41927_ ( .A(1'h1), .B(_control_conv2d_8_cond_30_6_1), .S(_05124_), .Y(_22763_) );
  \$mux  #( .WIDTH(1) ) _41929_ ( .A(set_req_214), .B(1'h0), .S(_control_conv2d_8_cond_30_6_1), .Y(_22764_) );
  \$mux  #( .WIDTH(1) ) _41930_ ( .A(_22764_), .B(set_req_214), .S(_05112_), .Y(_22765_) );
  \$mux  #( .WIDTH(1) ) _41931_ ( .A(1'h1), .B(_22765_), .S(_05124_), .Y(_22766_) );
  \$mux  #( .WIDTH(1) ) _41933_ ( .A(1'h1), .B(_control_conv2d_8_cond_24_5_1), .S(_05125_), .Y(_22767_) );
  \$mux  #( .WIDTH(1) ) _41935_ ( .A(axim_flag_158), .B(1'h0), .S(_control_conv2d_8_cond_24_5_1), .Y(_22768_) );
  \$mux  #( .WIDTH(1) ) _41936_ ( .A(_22768_), .B(axim_flag_158), .S(_05113_), .Y(_22769_) );
  \$mux  #( .WIDTH(1) ) _41937_ ( .A(1'h1), .B(_22769_), .S(_05125_), .Y(_22770_) );
  \$mux  #( .WIDTH(1) ) _41939_ ( .A(1'h1), .B(_control_conv2d_8_cond_23_4_1), .S(_05126_), .Y(_22771_) );
  \$mux  #( .WIDTH(1) ) _41941_ ( .A(set_req_157), .B(1'h0), .S(_control_conv2d_8_cond_23_4_1), .Y(_22772_) );
  \$mux  #( .WIDTH(1) ) _41942_ ( .A(_22772_), .B(set_req_157), .S(_05114_), .Y(_22773_) );
  \$mux  #( .WIDTH(1) ) _41943_ ( .A(1'h1), .B(_22773_), .S(_05126_), .Y(_22774_) );
  \$mux  #( .WIDTH(1) ) _41945_ ( .A(1'h1), .B(_control_conv2d_8_cond_15_3_1), .S(_05127_), .Y(_22775_) );
  \$mux  #( .WIDTH(1) ) _41947_ ( .A(axim_flag_29), .B(1'h0), .S(_control_conv2d_8_cond_15_3_1), .Y(_22776_) );
  \$mux  #( .WIDTH(1) ) _41948_ ( .A(_22776_), .B(axim_flag_29), .S(_05115_), .Y(_22777_) );
  \$mux  #( .WIDTH(1) ) _41949_ ( .A(1'h1), .B(_22777_), .S(_05127_), .Y(_22778_) );
  \$mux  #( .WIDTH(1) ) _41951_ ( .A(1'h1), .B(_control_conv2d_8_cond_14_2_1), .S(_05128_), .Y(_22779_) );
  \$mux  #( .WIDTH(1) ) _41953_ ( .A(set_req_28), .B(1'h0), .S(_control_conv2d_8_cond_14_2_1), .Y(_22780_) );
  \$mux  #( .WIDTH(1) ) _41954_ ( .A(_22780_), .B(set_req_28), .S(_05116_), .Y(_22781_) );
  \$mux  #( .WIDTH(1) ) _41955_ ( .A(1'h1), .B(_22781_), .S(_05128_), .Y(_22782_) );
  \$mux  #( .WIDTH(1) ) _41957_ ( .A(1'h1), .B(_control_conv2d_8_cond_8_1_1), .S(_05130_), .Y(_22783_) );
  \$mux  #( .WIDTH(1) ) _41959_ ( .A(axim_flag_16), .B(1'h0), .S(_control_conv2d_8_cond_8_1_1), .Y(_22784_) );
  \$mux  #( .WIDTH(1) ) _41960_ ( .A(_22784_), .B(axim_flag_16), .S(_05117_), .Y(_22785_) );
  \$mux  #( .WIDTH(1) ) _41961_ ( .A(1'h1), .B(_22785_), .S(_05130_), .Y(_22786_) );
  \$mux  #( .WIDTH(1) ) _41963_ ( .A(1'h1), .B(_control_conv2d_8_cond_3_0_1), .S(_05131_), .Y(_22787_) );
  \$mux  #( .WIDTH(1) ) _41966_ ( .A(axim_flag_9), .B(1'h0), .S(_control_conv2d_8_cond_3_0_1), .Y(_22788_) );
  \$mux  #( .WIDTH(1) ) _41967_ ( .A(_22788_), .B(axim_flag_9), .S(_05118_), .Y(_22789_) );
  \$mux  #( .WIDTH(1) ) _41968_ ( .A(1'h1), .B(_22789_), .S(_05131_), .Y(_22790_) );
  \$mux  #( .WIDTH(1) ) _41970_ ( .A(conv2d_8_skip_write_out), .B(1'h0), .S(_05810_), .Y(_18550_) );
  \$mux  #( .WIDTH(1) ) _41971_ ( .A(_22791_), .B(1'h1), .S(RST), .Y(_03072_) );
  \$mux  #( .WIDTH(1) ) _41972_ ( .A(conv2d_8_skip_comp), .B(1'h1), .S(conv2d_8_update_filter), .Y(_18552_) );
  \$mux  #( .WIDTH(1) ) _41974_ ( .A(conv2d_8_skip_read_act), .B(1'h1), .S(conv2d_8_update_filter), .Y(_18554_) );
  \$mux  #( .WIDTH(1) ) _41976_ ( .A(conv2d_8_skip_read_filter), .B(1'h1), .S(conv2d_8_update_filter), .Y(_18556_) );
  \$mux  #( .WIDTH(32) ) _41978_ ( .A(0), .B(conv2d_8_out_laddr_offset), .S(conv2d_8_skip_write_out), .Y({ _18582_, _18581_, _18579_, _18578_, _18577_, _18576_, _18575_, _18574_, _18573_, _18572_, _18571_, _18570_, _18568_, _18567_, _18566_, _18565_, _18564_, _18563_, _18562_, _18561_, _18560_, _18559_, _18589_, _18588_, _18587_, _18586_, _18585_, _18584_, _18583_, _18580_, _18569_, _18558_ }) );
  \$mux  #( .WIDTH(32) ) _41979_ ( .A(_22266_), .B(conv2d_8_out_laddr_offset), .S(_04894_), .Y({ _18614_, _18613_, _18611_, _18610_, _18609_, _18608_, _18607_, _18606_, _18605_, _18604_, _18603_, _18602_, _18600_, _18599_, _18598_, _18597_, _18596_, _18595_, _18594_, _18593_, _18592_, _18591_, _18621_, _18620_, _18619_, _18618_, _18617_, _18616_, _18615_, _18612_, _18601_, _18590_ }) );
  \$mux  #( .WIDTH(32) ) _41981_ ( .A(0), .B(1024), .S(conv2d_8_out_page), .Y({ _18646_, _18645_, _18643_, _18642_, _18641_, _18640_, _18639_, _18638_, _18637_, _18636_, _18635_, _18634_, _18632_, _18631_, _18630_, _18629_, _18628_, _18627_, _18626_, _18625_, _18624_, _18623_, _18653_, _18652_, _18651_, _18650_, _18649_, _18648_, _18647_, _18644_, _18633_, _18622_ }) );
  \$mux  #( .WIDTH(32) ) _41983_ ( .A(1024), .B(0), .S(conv2d_8_out_page), .Y({ _18710_, _18709_, _18707_, _18706_, _18705_, _18704_, _18703_, _18702_, _18701_, _18700_, _18699_, _18698_, _18696_, _18695_, _18694_, _18693_, _18692_, _18691_, _18690_, _18689_, _18688_, _18687_, _18717_, _18716_, _18715_, _18714_, _18713_, _18712_, _18711_, _18708_, _18697_, _18686_ }) );
  \$mux  #( .WIDTH(1) ) _41985_ ( .A(1'h1), .B(1'h0), .S(conv2d_8_out_page), .Y(_18750_) );
  \$mux  #( .WIDTH(32) ) _41987_ ( .A(conv2d_8_filter_page_dma_offset), .B(_22271_), .S(conv2d_8_update_filter), .Y(_22799_) );
  \$mux  #( .WIDTH(32) ) _41988_ ( .A(_22799_), .B(0), .S(_05805_), .Y({ _18776_, _18775_, _18773_, _18772_, _18771_, _18770_, _18769_, _18768_, _18767_, _18766_, _18765_, _18764_, _18762_, _18761_, _18760_, _18759_, _18758_, _18757_, _18756_, _18755_, _18754_, _18753_, _18783_, _18782_, _18781_, _18780_, _18779_, _18778_, _18777_, _18774_, _18763_, _18752_ }) );
  \$mux  #( .WIDTH(32) ) _41990_ ( .A(conv2d_8_filter_page_comp_offset), .B(_22270_), .S(conv2d_8_update_filter), .Y(_22801_) );
  \$mux  #( .WIDTH(32) ) _41991_ ( .A(_22801_), .B(0), .S(_05805_), .Y({ _18840_, _18839_, _18837_, _18836_, _18835_, _18834_, _18833_, _18832_, _18831_, _18830_, _18829_, _18828_, _18826_, _18825_, _18824_, _18823_, _18822_, _18821_, _18820_, _18819_, _18818_, _18817_, _18847_, _18846_, _18845_, _18844_, _18843_, _18842_, _18841_, _18838_, _18827_, _18816_ }) );
  \$mux  #( .WIDTH(32) ) _41993_ ( .A(conv2d_8_act_page_dma_offset_2), .B(_22280_), .S(conv2d_8_mux_next_dma_flag_2), .Y(_22803_) );
  \$mux  #( .WIDTH(32) ) _41994_ ( .A(_22803_), .B(0), .S(_05808_), .Y(_22804_) );
  \$mux  #( .WIDTH(32) ) _41995_ ( .A(_22804_), .B(0), .S(conv2d_8_update_filter), .Y({ _18904_, _18903_, _18901_, _18900_, _18899_, _18898_, _18897_, _18896_, _18895_, _18894_, _18893_, _18892_, _18890_, _18889_, _18888_, _18887_, _18886_, _18885_, _18884_, _18883_, _18882_, _18881_, _18911_, _18910_, _18909_, _18908_, _18907_, _18906_, _18905_, _18902_, _18891_, _18880_ }) );
  \$mux  #( .WIDTH(32) ) _41997_ ( .A(conv2d_8_act_page_dma_offset_1), .B(_22278_), .S(conv2d_8_mux_next_dma_flag_1), .Y(_22806_) );
  \$mux  #( .WIDTH(32) ) _41998_ ( .A(_22806_), .B(0), .S(_05807_), .Y(_22807_) );
  \$mux  #( .WIDTH(32) ) _41999_ ( .A(_22807_), .B(0), .S(conv2d_8_update_filter), .Y({ _18968_, _18967_, _18965_, _18964_, _18963_, _18962_, _18961_, _18960_, _18959_, _18958_, _18957_, _18956_, _18954_, _18953_, _18952_, _18951_, _18950_, _18949_, _18948_, _18947_, _18946_, _18945_, _18975_, _18974_, _18973_, _18972_, _18971_, _18970_, _18969_, _18966_, _18955_, _18944_ }) );
  \$mux  #( .WIDTH(32) ) _42001_ ( .A(conv2d_8_act_page_dma_offset_0), .B(_22276_), .S(conv2d_8_mux_next_dma_flag_0), .Y(_22809_) );
  \$mux  #( .WIDTH(32) ) _42002_ ( .A(_22809_), .B(0), .S(_05806_), .Y(_22810_) );
  \$mux  #( .WIDTH(32) ) _42003_ ( .A(_22810_), .B(0), .S(conv2d_8_update_filter), .Y({ _19032_, _19031_, _19029_, _19028_, _19027_, _19026_, _19025_, _19024_, _19023_, _19022_, _19021_, _19020_, _19018_, _19017_, _19016_, _19015_, _19014_, _19013_, _19012_, _19011_, _19010_, _19009_, _19039_, _19038_, _19037_, _19036_, _19035_, _19034_, _19033_, _19030_, _19019_, _19008_ }) );
  \$mux  #( .WIDTH(32) ) _42005_ ( .A(conv2d_8_act_page_comp_offset_2), .B(_22279_), .S(conv2d_8_mux_next_dma_flag_2), .Y(_22812_) );
  \$mux  #( .WIDTH(32) ) _42006_ ( .A(_22812_), .B(0), .S(_05808_), .Y(_22813_) );
  \$mux  #( .WIDTH(32) ) _42007_ ( .A(_22813_), .B(0), .S(conv2d_8_update_filter), .Y({ _19096_, _19095_, _19093_, _19092_, _19091_, _19090_, _19089_, _19088_, _19087_, _19086_, _19085_, _19084_, _19082_, _19081_, _19080_, _19079_, _19078_, _19077_, _19076_, _19075_, _19074_, _19073_, _19103_, _19102_, _19101_, _19100_, _19099_, _19098_, _19097_, _19094_, _19083_, _19072_ }) );
  \$mux  #( .WIDTH(32) ) _42009_ ( .A(conv2d_8_act_page_comp_offset_1), .B(_22277_), .S(conv2d_8_mux_next_dma_flag_1), .Y(_22815_) );
  \$mux  #( .WIDTH(32) ) _42010_ ( .A(_22815_), .B(0), .S(_05807_), .Y(_22816_) );
  \$mux  #( .WIDTH(32) ) _42011_ ( .A(_22816_), .B(0), .S(conv2d_8_update_filter), .Y({ _19160_, _19159_, _19157_, _19156_, _19155_, _19154_, _19153_, _19152_, _19151_, _19150_, _19149_, _19148_, _19146_, _19145_, _19144_, _19143_, _19142_, _19141_, _19140_, _19139_, _19138_, _19137_, _19167_, _19166_, _19165_, _19164_, _19163_, _19162_, _19161_, _19158_, _19147_, _19136_ }) );
  \$mux  #( .WIDTH(32) ) _42013_ ( .A(conv2d_8_act_page_comp_offset_0), .B(_22275_), .S(conv2d_8_mux_next_dma_flag_0), .Y(_22818_) );
  \$mux  #( .WIDTH(32) ) _42014_ ( .A(_22818_), .B(0), .S(_05806_), .Y(_22819_) );
  \$mux  #( .WIDTH(32) ) _42015_ ( .A(_22819_), .B(0), .S(conv2d_8_update_filter), .Y({ _19224_, _19223_, _19221_, _19220_, _19219_, _19218_, _19217_, _19216_, _19215_, _19214_, _19213_, _19212_, _19210_, _19209_, _19208_, _19207_, _19206_, _19205_, _19204_, _19203_, _19202_, _19201_, _19231_, _19230_, _19229_, _19228_, _19227_, _19226_, _19225_, _19222_, _19211_, _19200_ }) );
  \$mux  #( .WIDTH(2) ) _42017_ ( .A(conv2d_8_row_select), .B(2'h0), .S(conv2d_8_update_filter), .Y({ _19265_, _19264_ }) );
  \$mux  #( .WIDTH(32) ) _42022_ ( .A(0), .B(conv2d_8_out_ram_select), .S(conv2d_8_skip_write_out), .Y({ _19388_, _19387_, _19385_, _19384_, _19383_, _19382_, _19381_, _19380_, _19379_, _19378_, _19377_, _19376_, _19374_, _19373_, _19372_, _19371_, _19370_, _19369_, _19368_, _19367_, _19366_, _19365_, _19395_, _19394_, _19393_, _19392_, _19391_, _19390_, _19389_, _19386_, _19375_, _19364_ }) );
  \$mux  #( .WIDTH(32) ) _42023_ ( .A(0), .B(_22267_), .S(_04894_), .Y({ _19420_, _19419_, _19417_, _19416_, _19415_, _19414_, _19413_, _19412_, _19411_, _19410_, _19409_, _19408_, _19406_, _19405_, _19404_, _19403_, _19402_, _19401_, _19400_, _19399_, _19398_, _19397_, _19427_, _19426_, _19425_, _19424_, _19423_, _19422_, _19421_, _19418_, _19407_, _19396_ }) );
  \$mux  #( .WIDTH(32) ) _42025_ ( .A(_22282_), .B(conv2d_8_out_row_count), .S(conv2d_8_skip_write_out), .Y(_22826_) );
  \$mux  #( .WIDTH(32) ) _42026_ ( .A(_22826_), .B(0), .S(_05809_), .Y({ _19452_, _19451_, _19449_, _19448_, _19447_, _19446_, _19445_, _19444_, _19443_, _19442_, _19441_, _19440_, _19438_, _19437_, _19436_, _19435_, _19434_, _19433_, _19432_, _19431_, _19430_, _19429_, _19459_, _19458_, _19457_, _19456_, _19455_, _19454_, _19453_, _19450_, _19439_, _19428_ }) );
  \$mux  #( .WIDTH(2) ) _42028_ ( .A(_22274_), .B(_26322_[1:0]), .S(_05240_), .Y(_22828_) );
  \$mux  #( .WIDTH(2) ) _42029_ ( .A(_22828_), .B(2'h0), .S(conv2d_8_update_filter), .Y({ _19493_, _19492_ }) );
  \$mux  #( .WIDTH(32) ) _42031_ ( .A(conv2d_8_och_count), .B(_22269_), .S(conv2d_8_update_filter), .Y({ _19520_, _19519_, _19517_, _19516_, _19515_, _19514_, _19513_, _19512_, _19511_, _19510_, _19509_, _19508_, _19506_, _19505_, _19504_, _19503_, _19502_, _19501_, _19500_, _19499_, _19498_, _19497_, _19527_, _19526_, _19525_, _19524_, _19523_, _19522_, _19521_, _19518_, _19507_, _19496_ }) );
  \$mux  #( .WIDTH(32) ) _42033_ ( .A(conv2d_8_bat_count), .B(0), .S(conv2d_8_update_filter), .Y({ _19584_, _19583_, _19581_, _19580_, _19579_, _19578_, _19577_, _19576_, _19575_, _19574_, _19573_, _19572_, _19570_, _19569_, _19568_, _19567_, _19566_, _19565_, _19564_, _19563_, _19562_, _19561_, _19591_, _19590_, _19589_, _19588_, _19587_, _19586_, _19585_, _19582_, _19571_, _19560_ }) );
  \$mux  #( .WIDTH(32) ) _42035_ ( .A(_22273_), .B(0), .S(conv2d_8_update_filter), .Y({ _19648_, _19647_, _19645_, _19644_, _19643_, _19642_, _19641_, _19640_, _19639_, _19638_, _19637_, _19636_, _19634_, _19633_, _19632_, _19631_, _19630_, _19629_, _19628_, _19627_, _19626_, _19625_, _19655_, _19654_, _19653_, _19652_, _19651_, _19650_, _19649_, _19646_, _19635_, _19624_ }) );
  \$mux  #( .WIDTH(32) ) _42037_ ( .A(conv2d_8_next_out_write_size), .B({ 23'h000000, cparam_conv2d_8_out_row_step }), .S(_04700_), .Y(_22833_) );
  \$mux  #( .WIDTH(1) ) _42041_ ( .A(1'h0), .B(1'h1), .S(conv2d_8_update_filter), .Y(_19720_) );
  \$mux  #( .WIDTH(1) ) _42043_ ( .A(conv2d_8_dma_flag_0), .B(1'h1), .S(_04700_), .Y(_22837_) );
  \$mux  #( .WIDTH(32) ) _42045_ ( .A(conv2d_8_out_base_offset_och), .B(_22283_), .S(_05809_), .Y({ _19746_, _19745_, _19743_, _19742_, _19741_, _19740_, _19739_, _19738_, _19737_, _19736_, _19735_, _19734_, _19732_, _19731_, _19730_, _19729_, _19728_, _19727_, _19726_, _19725_, _19724_, _19723_, _19753_, _19752_, _19751_, _19750_, _19749_, _19748_, _19747_, _19744_, _19733_, _19722_ }) );
  \$mux  #( .WIDTH(32) ) _42047_ ( .A(conv2d_8_out_base_offset_bat), .B(0), .S(_05809_), .Y({ _19810_, _19809_, _19807_, _19806_, _19805_, _19804_, _19803_, _19802_, _19801_, _19800_, _19799_, _19798_, _19796_, _19795_, _19794_, _19793_, _19792_, _19791_, _19790_, _19789_, _19788_, _19787_, _19817_, _19816_, _19815_, _19814_, _19813_, _19812_, _19811_, _19808_, _19797_, _19786_ }) );
  \$mux  #( .WIDTH(32) ) _42049_ ( .A(_22281_), .B(conv2d_8_out_base_offset_row), .S(conv2d_8_skip_write_out), .Y(_22840_) );
  \$mux  #( .WIDTH(32) ) _42050_ ( .A(_22840_), .B(0), .S(_05809_), .Y({ _19874_, _19873_, _19871_, _19870_, _19869_, _19868_, _19867_, _19866_, _19865_, _19864_, _19863_, _19862_, _19860_, _19859_, _19858_, _19857_, _19856_, _19855_, _19854_, _19853_, _19852_, _19851_, _19881_, _19880_, _19879_, _19878_, _19877_, _19876_, _19875_, _19872_, _19861_, _19850_ }) );
  \$mux  #( .WIDTH(32) ) _42052_ ( .A(0), .B(conv2d_8_out_base_offset_col), .S(conv2d_8_skip_write_out), .Y({ _19938_, _19937_, _19935_, _19934_, _19933_, _19932_, _19931_, _19930_, _19929_, _19928_, _19927_, _19926_, _19924_, _19923_, _19922_, _19921_, _19920_, _19919_, _19918_, _19917_, _19916_, _19915_, _19945_, _19944_, _19943_, _19942_, _19941_, _19940_, _19939_, _19936_, _19925_, _19914_ }) );
  \$mux  #( .WIDTH(32) ) _42054_ ( .A(0), .B(conv2d_8_out_base_offset_val), .S(_05132_), .Y(_22843_) );
  \$mux  #( .WIDTH(32) ) _42056_ ( .A(conv2d_8_filter_base_offset), .B(_22268_), .S(conv2d_8_update_filter), .Y({ _20002_, _20001_, _19999_, _19998_, _19997_, _19996_, _19995_, _19994_, _19993_, _19992_, _19991_, _19990_, _19988_, _19987_, _19986_, _19985_, _19984_, _19983_, _19982_, _19981_, _19980_, _19979_, _20009_, _20008_, _20007_, _20006_, _20005_, _20004_, _20003_, _20000_, _19989_, _19978_ }) );
  \$mux  #( .WIDTH(32) ) _42058_ ( .A(conv2d_8_act_base_offset_bat), .B(0), .S(conv2d_8_update_filter), .Y({ _20066_, _20065_, _20063_, _20062_, _20061_, _20060_, _20059_, _20058_, _20057_, _20056_, _20055_, _20054_, _20052_, _20051_, _20050_, _20049_, _20048_, _20047_, _20046_, _20045_, _20044_, _20043_, _20073_, _20072_, _20071_, _20070_, _20069_, _20068_, _20067_, _20064_, _20053_, _20042_ }) );
  \$mux  #( .WIDTH(32) ) _42060_ ( .A(_22272_), .B(0), .S(conv2d_8_update_filter), .Y({ _20130_, _20129_, _20127_, _20126_, _20125_, _20124_, _20123_, _20122_, _20121_, _20120_, _20119_, _20118_, _20116_, _20115_, _20114_, _20113_, _20112_, _20111_, _20110_, _20109_, _20108_, _20107_, _20137_, _20136_, _20135_, _20134_, _20133_, _20132_, _20131_, _20128_, _20117_, _20106_ }) );
  \$mux  #( .WIDTH(32) ) _42062_ ( .A(0), .B(control_conv2d_8), .S(_05147_), .Y(_22847_) );
  \$mux  #( .WIDTH(32) ) _42063_ ( .A(0), .B(_22847_), .S(_05143_), .Y({ _20194_, _20193_, _20191_, _20190_, _20189_, _20188_, _20187_, _20186_, _20185_, _20184_, _20183_, _20182_, _20180_, _20179_, _20178_, _20177_, _20176_, _20175_, _20174_, _20173_, _20172_, _20171_, _20201_, _20200_, _20199_, _20198_, _20197_, _20196_, _20195_, _20192_, _20181_, _20170_ }) );
  \$mux  #( .WIDTH(32) ) _42064_ ( .A(control_conv2d_8), .B(55), .S(_maxi_write_idle), .Y({ _20258_, _20257_, _20255_, _20254_, _20253_, _20252_, _20251_, _20250_, _20249_, _20248_, _20247_, _20246_, _20244_, _20243_, _20242_, _20241_, _20240_, _20239_, _20238_, _20237_, _20236_, _20235_, _20265_, _20264_, _20263_, _20262_, _20261_, _20260_, _20259_, _20256_, _20245_, _20234_ }) );
  \$mux  #( .WIDTH(32) ) _42065_ ( .A(21), .B(13), .S(conv2d_8_update_filter), .Y(_22849_) );
  \$mux  #( .WIDTH(32) ) _42066_ ( .A(_22849_), .B(54), .S(_05809_), .Y({ _20290_, _20289_, _20287_, _20286_, _20285_, _20284_, _20283_, _20282_, _20281_, _20280_, _20279_, _20278_, _20276_, _20275_, _20274_, _20273_, _20272_, _20271_, _20270_, _20269_, _20268_, _20267_, _20297_, _20296_, _20295_, _20294_, _20293_, _20292_, _20291_, _20288_, _20277_, _20266_ }) );
  \$mux  #( .WIDTH(32) ) _42067_ ( .A(control_conv2d_8), .B(48), .S(_maxi_write_idle), .Y({ _20322_, _20321_, _20319_, _20318_, _20317_, _20316_, _20315_, _20314_, _20313_, _20312_, _20311_, _20310_, _20308_, _20307_, _20306_, _20305_, _20304_, _20303_, _20302_, _20301_, _20300_, _20299_, _20329_, _20328_, _20327_, _20326_, _20325_, _20324_, _20323_, _20320_, _20309_, _20298_ }) );
  \$mux  #( .WIDTH(32) ) _42068_ ( .A(47), .B(51), .S(conv2d_8_dma_out_mask_0), .Y({ _20354_, _20353_, _20351_, _20350_, _20349_, _20348_, _20347_, _20346_, _20345_, _20344_, _20343_, _20342_, _20340_, _20339_, _20338_, _20337_, _20336_, _20335_, _20334_, _20333_, _20332_, _20331_, _20361_, _20360_, _20359_, _20358_, _20357_, _20356_, _20355_, _20352_, _20341_, _20330_ }) );
  \$mux  #( .WIDTH(32) ) _42069_ ( .A(control_conv2d_8), .B(46), .S(_05239_), .Y(_22850_) );
  \$mux  #( .WIDTH(32) ) _42070_ ( .A(_22850_), .B(53), .S(conv2d_8_skip_write_out), .Y({ _20386_, _20385_, _20383_, _20382_, _20381_, _20380_, _20379_, _20378_, _20377_, _20376_, _20375_, _20374_, _20372_, _20371_, _20370_, _20369_, _20368_, _20367_, _20366_, _20365_, _20364_, _20363_, _20393_, _20392_, _20391_, _20390_, _20389_, _20388_, _20387_, _20384_, _20373_, _20362_ }) );
  \$mux  #( .WIDTH(32) ) _42071_ ( .A(45), .B(control_conv2d_8), .S(_04899_), .Y({ _20418_, _20417_, _20415_, _20414_, _20413_, _20412_, _20411_, _20410_, _20409_, _20408_, _20407_, _20406_, _20404_, _20403_, _20402_, _20401_, _20400_, _20399_, _20398_, _20397_, _20396_, _20395_, _20425_, _20424_, _20423_, _20422_, _20421_, _20420_, _20419_, _20416_, _20405_, _20394_ }) );
  \$mux  #( .WIDTH(32) ) _42072_ ( .A(control_conv2d_8), .B(42), .S(_maxi_read_idle), .Y({ _20450_, _20449_, _20447_, _20446_, _20445_, _20444_, _20443_, _20442_, _20441_, _20440_, _20439_, _20438_, _20436_, _20435_, _20434_, _20433_, _20432_, _20431_, _20430_, _20429_, _20428_, _20427_, _20457_, _20456_, _20455_, _20454_, _20453_, _20452_, _20451_, _20448_, _20437_, _20426_ }) );
  \$mux  #( .WIDTH(32) ) _42073_ ( .A(control_conv2d_8), .B(37), .S(_maxi_read_idle), .Y({ _20482_, _20481_, _20479_, _20478_, _20477_, _20476_, _20475_, _20474_, _20473_, _20472_, _20471_, _20470_, _20468_, _20467_, _20466_, _20465_, _20464_, _20463_, _20462_, _20461_, _20460_, _20459_, _20489_, _20488_, _20487_, _20486_, _20485_, _20484_, _20483_, _20480_, _20469_, _20458_ }) );
  \$mux  #( .WIDTH(32) ) _42074_ ( .A(36), .B(42), .S(_05870_), .Y({ _20514_, _20513_, _20511_, _20510_, _20509_, _20508_, _20507_, _20506_, _20505_, _20504_, _20503_, _20502_, _20500_, _20499_, _20498_, _20497_, _20496_, _20495_, _20494_, _20493_, _20492_, _20491_, _20521_, _20520_, _20519_, _20518_, _20517_, _20516_, _20515_, _20512_, _20501_, _20490_ }) );
  \$mux  #( .WIDTH(32) ) _42075_ ( .A(control_conv2d_8), .B(35), .S(_maxi_read_idle), .Y({ _20546_, _20545_, _20543_, _20542_, _20541_, _20540_, _20539_, _20538_, _20537_, _20536_, _20535_, _20534_, _20532_, _20531_, _20530_, _20529_, _20528_, _20527_, _20526_, _20525_, _20524_, _20523_, _20553_, _20552_, _20551_, _20550_, _20549_, _20548_, _20547_, _20544_, _20533_, _20522_ }) );
  \$mux  #( .WIDTH(32) ) _42076_ ( .A(control_conv2d_8), .B(30), .S(_maxi_read_idle), .Y({ _20578_, _20577_, _20575_, _20574_, _20573_, _20572_, _20571_, _20570_, _20569_, _20568_, _20567_, _20566_, _20564_, _20563_, _20562_, _20561_, _20560_, _20559_, _20558_, _20557_, _20556_, _20555_, _20585_, _20584_, _20583_, _20582_, _20581_, _20580_, _20579_, _20576_, _20565_, _20554_ }) );
  \$mux  #( .WIDTH(32) ) _42077_ ( .A(29), .B(35), .S(_05869_), .Y({ _20610_, _20609_, _20607_, _20606_, _20605_, _20604_, _20603_, _20602_, _20601_, _20600_, _20599_, _20598_, _20596_, _20595_, _20594_, _20593_, _20592_, _20591_, _20590_, _20589_, _20588_, _20587_, _20617_, _20616_, _20615_, _20614_, _20613_, _20612_, _20611_, _20608_, _20597_, _20586_ }) );
  \$mux  #( .WIDTH(32) ) _42078_ ( .A(control_conv2d_8), .B(28), .S(_maxi_read_idle), .Y({ _20642_, _20641_, _20639_, _20638_, _20637_, _20636_, _20635_, _20634_, _20633_, _20632_, _20631_, _20630_, _20628_, _20627_, _20626_, _20625_, _20624_, _20623_, _20622_, _20621_, _20620_, _20619_, _20649_, _20648_, _20647_, _20646_, _20645_, _20644_, _20643_, _20640_, _20629_, _20618_ }) );
  \$mux  #( .WIDTH(32) ) _42079_ ( .A(control_conv2d_8), .B(23), .S(_maxi_read_idle), .Y({ _20674_, _20673_, _20671_, _20670_, _20669_, _20668_, _20667_, _20666_, _20665_, _20664_, _20663_, _20662_, _20660_, _20659_, _20658_, _20657_, _20656_, _20655_, _20654_, _20653_, _20652_, _20651_, _20681_, _20680_, _20679_, _20678_, _20677_, _20676_, _20675_, _20672_, _20661_, _20650_ }) );
  \$mux  #( .WIDTH(32) ) _42080_ ( .A(22), .B(28), .S(_05868_), .Y(_22851_) );
  \$mux  #( .WIDTH(32) ) _42081_ ( .A(_22851_), .B(43), .S(conv2d_8_skip_read_act), .Y({ _20706_, _20705_, _20703_, _20702_, _20701_, _20700_, _20699_, _20698_, _20697_, _20696_, _20695_, _20694_, _20692_, _20691_, _20690_, _20689_, _20688_, _20687_, _20686_, _20685_, _20684_, _20683_, _20713_, _20712_, _20711_, _20710_, _20709_, _20708_, _20707_, _20704_, _20693_, _20682_ }) );
  \$mux  #( .WIDTH(32) ) _42082_ ( .A(control_conv2d_8), .B(19), .S(_maxi_read_idle), .Y({ _20738_, _20737_, _20735_, _20734_, _20733_, _20732_, _20731_, _20730_, _20729_, _20728_, _20727_, _20726_, _20724_, _20723_, _20722_, _20721_, _20720_, _20719_, _20718_, _20717_, _20716_, _20715_, _20745_, _20744_, _20743_, _20742_, _20741_, _20740_, _20739_, _20736_, _20725_, _20714_ }) );
  \$mux  #( .WIDTH(32) ) _42083_ ( .A(control_conv2d_8), .B(14), .S(_maxi_read_idle), .Y(_22852_) );
  \$mux  #( .WIDTH(32) ) _42084_ ( .A(_22852_), .B(20), .S(conv2d_8_skip_read_filter), .Y({ _20770_, _20769_, _20767_, _20766_, _20765_, _20764_, _20763_, _20762_, _20761_, _20760_, _20759_, _20758_, _20756_, _20755_, _20754_, _20753_, _20752_, _20751_, _20750_, _20749_, _20748_, _20747_, _20777_, _20776_, _20775_, _20774_, _20773_, _20772_, _20771_, _20768_, _20757_, _20746_ }) );
  \$mux  #( .WIDTH(32) ) _42085_ ( .A(control_conv2d_8), .B(12), .S(_maxi_read_idle), .Y({ _20802_, _20801_, _20799_, _20798_, _20797_, _20796_, _20795_, _20794_, _20793_, _20792_, _20791_, _20790_, _20788_, _20787_, _20786_, _20785_, _20784_, _20783_, _20782_, _20781_, _20780_, _20779_, _20809_, _20808_, _20807_, _20806_, _20805_, _20804_, _20803_, _20800_, _20789_, _20778_ }) );
  \$mux  #( .WIDTH(32) ) _42086_ ( .A(control_conv2d_8), .B(8), .S(_maxi_read_idle), .Y({ _20834_, _20833_, _20831_, _20830_, _20829_, _20828_, _20827_, _20826_, _20825_, _20824_, _20823_, _20822_, _20820_, _20819_, _20818_, _20817_, _20816_, _20815_, _20814_, _20813_, _20812_, _20811_, _20841_, _20840_, _20839_, _20838_, _20837_, _20836_, _20835_, _20832_, _20821_, _20810_ }) );
  \$mux  #( .WIDTH(32) ) _42087_ ( .A(control_conv2d_8), .B(7), .S(_maxi_read_idle), .Y({ _20866_, _20865_, _20863_, _20862_, _20861_, _20860_, _20859_, _20858_, _20857_, _20856_, _20855_, _20854_, _20852_, _20851_, _20850_, _20849_, _20848_, _20847_, _20846_, _20845_, _20844_, _20843_, _20873_, _20872_, _20871_, _20870_, _20869_, _20868_, _20867_, _20864_, _20853_, _20842_ }) );
  \$mux  #( .WIDTH(32) ) _42088_ ( .A(control_conv2d_8), .B(3), .S(_maxi_read_idle), .Y({ _20898_, _20897_, _20895_, _20894_, _20893_, _20892_, _20891_, _20890_, _20889_, _20888_, _20887_, _20886_, _20884_, _20883_, _20882_, _20881_, _20880_, _20879_, _20878_, _20877_, _20876_, _20875_, _20905_, _20904_, _20903_, _20902_, _20901_, _20900_, _20899_, _20896_, _20885_, _20874_ }) );
  \$mux  #( .WIDTH(32) ) _42089_ ( .A(1), .B(control_conv2d_8), .S(_05148_), .Y(_22853_) );
  \$mux  #( .WIDTH(32) ) _42090_ ( .A(1), .B(_22853_), .S(_05144_), .Y({ _20930_, _20929_, _20927_, _20926_, _20925_, _20924_, _20923_, _20922_, _20921_, _20920_, _20919_, _20918_, _20916_, _20915_, _20914_, _20913_, _20912_, _20911_, _20910_, _20909_, _20908_, _20907_, _20937_, _20936_, _20935_, _20934_, _20933_, _20932_, _20931_, _20928_, _20917_, _20906_ }) );
  \$mux  #( .WIDTH(32) ) _42092_ ( .A(_22265_), .B(matmul_15_arg_objaddr_3), .S(_05136_), .Y(_22854_) );
  \$mux  #( .WIDTH(32) ) _42094_ ( .A(_22264_), .B(matmul_15_arg_objaddr_2), .S(_05137_), .Y(_22855_) );
  \$mux  #( .WIDTH(32) ) _42096_ ( .A(_22263_), .B(matmul_15_arg_objaddr_1), .S(_05138_), .Y(_22856_) );
  \$mux  #( .WIDTH(32) ) _42098_ ( .A({ _03890_, _03889_, _03887_, _03886_, _03885_, _03884_, _03883_, _03882_, _03881_, _03880_, _03879_, _03878_, _03876_, _03875_, _03874_, _03873_, _03872_, _03871_, _03870_, _03869_, _03868_, _03867_, _03897_, _03896_, _03895_, _03894_, _03893_, _03892_, _03891_, _03888_, _03877_, _03866_ }), .B(matmul_15_arg_objaddr_0), .S(_05139_), .Y(_22857_) );
  \$mux  #( .WIDTH(32) ) _42100_ ( .A(_saxi_register_11), .B(matmul_15_objaddr), .S(_05140_), .Y(_22858_) );
  \$mux  #( .WIDTH(32) ) _42109_ ( .A(49), .B(main_fsm), .S(_05035_), .Y({ _21219_, _21218_, _21216_, _21215_, _21214_, _21213_, _21212_, _21211_, _21210_, _21209_, _21208_, _21207_, _21205_, _21204_, _21203_, _21202_, _21201_, _21200_, _21199_, _21198_, _21197_, _21196_, _21226_, _21225_, _21224_, _21223_, _21222_, _21221_, _21220_, _21217_, _21206_, _21195_ }) );
  \$mux  #( .WIDTH(32) ) _42110_ ( .A(38), .B(main_fsm), .S(_05052_), .Y({ _21251_, _21250_, _21248_, _21247_, _21246_, _21245_, _21244_, _21243_, _21242_, _21241_, _21240_, _21239_, _21237_, _21236_, _21235_, _21234_, _21233_, _21232_, _21231_, _21230_, _21229_, _21228_, _21258_, _21257_, _21256_, _21255_, _21254_, _21253_, _21252_, _21249_, _21238_, _21227_ }) );
  \$mux  #( .WIDTH(32) ) _42111_ ( .A(31), .B(main_fsm), .S(_05119_), .Y({ _21283_, _21282_, _21280_, _21279_, _21278_, _21277_, _21276_, _21275_, _21274_, _21273_, _21272_, _21271_, _21269_, _21268_, _21267_, _21266_, _21265_, _21264_, _21263_, _21262_, _21261_, _21260_, _21290_, _21289_, _21288_, _21287_, _21286_, _21285_, _21284_, _21281_, _21270_, _21259_ }) );
  \$mux  #( .WIDTH(32) ) _42112_ ( .A(21), .B(main_fsm), .S(_05052_), .Y({ _21315_, _21314_, _21312_, _21311_, _21310_, _21309_, _21308_, _21307_, _21306_, _21305_, _21304_, _21303_, _21301_, _21300_, _21299_, _21298_, _21297_, _21296_, _21295_, _21294_, _21293_, _21292_, _21322_, _21321_, _21320_, _21319_, _21318_, _21317_, _21316_, _21313_, _21302_, _21291_ }) );
  \$mux  #( .WIDTH(32) ) _42113_ ( .A(14), .B(main_fsm), .S(_05119_), .Y({ _21347_, _21346_, _21344_, _21343_, _21342_, _21341_, _21340_, _21339_, _21338_, _21337_, _21336_, _21335_, _21333_, _21332_, _21331_, _21330_, _21329_, _21328_, _21327_, _21326_, _21325_, _21324_, _21354_, _21353_, _21352_, _21351_, _21350_, _21349_, _21348_, _21345_, _21334_, _21323_ }) );
  \$mux  #( .WIDTH(32) ) _42114_ ( .A(main_fsm), .B(1), .S(_05873_), .Y({ _21379_, _21378_, _21376_, _21375_, _21374_, _21373_, _21372_, _21371_, _21370_, _21369_, _21368_, _21367_, _21365_, _21364_, _21363_, _21362_, _21361_, _21360_, _21359_, _21358_, _21357_, _21356_, _21386_, _21385_, _21384_, _21383_, _21382_, _21381_, _21380_, _21377_, _21366_, _21355_ }) );
  \$mux  #( .WIDTH(1) ) _42118_ ( .A(_stream_matmul_15_source_busy), .B(1'h1), .S(_stream_matmul_15_start_flag), .Y(_21388_) );
  \$mux  #( .WIDTH(1) ) _42120_ ( .A(1'h0), .B(1'h1), .S(__tmp_1117_34), .Y(_22870_) );
  \$mux  #( .WIDTH(1) ) _42122_ ( .A(1'h0), .B(1'h1), .S(__tmp_1115_38), .Y(_22871_) );
  \$mux  #( .WIDTH(1) ) _42124_ ( .A(1'h0), .B(1'h1), .S(_stream_matmul_15_start_flag), .Y(_22872_) );
  \$mux  #( .WIDTH(1) ) _42125_ ( .A(_22872_), .B(1'h0), .S(_04901_), .Y(_22873_) );
  \$mux  #( .WIDTH(32) ) _42127_ ( .A(_stream_matmul_15_fsm), .B(3), .S(_stream_matmul_15_done), .Y({ _21445_, _21444_, _21442_, _21441_, _21440_, _21439_, _21438_, _21437_, _21436_, _21435_, _21434_, _21433_, _21431_, _21430_, _21429_, _21428_, _21427_, _21426_, _21425_, _21424_, _21423_, _21422_, _21452_, _21451_, _21450_, _21449_, _21448_, _21447_, _21446_, _21443_, _21432_, _21421_ }) );
  \$mux  #( .WIDTH(32) ) _42128_ ( .A(_stream_matmul_15_fsm), .B(1), .S(_stream_matmul_15_start_flag), .Y({ _21477_, _21476_, _21474_, _21473_, _21472_, _21471_, _21470_, _21469_, _21468_, _21467_, _21466_, _21465_, _21463_, _21462_, _21461_, _21460_, _21459_, _21458_, _21457_, _21456_, _21455_, _21454_, _21484_, _21483_, _21482_, _21481_, _21480_, _21479_, _21478_, _21475_, _21464_, _21453_ }) );
  \$mux  #( .WIDTH(8) ) _42333_ ( .A(__variable_wdata_844), .B(_stream_matmul_15_source_20_source_ram_rdata), .S(_stream_matmul_15_source_20_source_ram_rvalid), .Y(_22876_) );
  \$mux  #( .WIDTH(32) ) _42335_ ( .A(_source_stream_matmul_15_source_20_pat_stride_buf_3), .B(_source_stream_matmul_15_source_20_pat_stride_3), .S(_05798_), .Y(_22877_) );
  \$mux  #( .WIDTH(32) ) _42337_ ( .A(_source_stream_matmul_15_source_20_pat_stride_buf_2), .B(_source_stream_matmul_15_source_20_pat_stride_2), .S(_05798_), .Y(_22878_) );
  \$mux  #( .WIDTH(32) ) _42339_ ( .A(_source_stream_matmul_15_source_20_pat_stride_buf_1), .B(_source_stream_matmul_15_source_20_pat_stride_1), .S(_05798_), .Y(_22879_) );
  \$mux  #( .WIDTH(32) ) _42341_ ( .A(_source_stream_matmul_15_source_20_pat_stride_buf_0), .B(_source_stream_matmul_15_source_20_pat_stride_0), .S(_05798_), .Y(_22880_) );
  \$mux  #( .WIDTH(33) ) _42343_ ( .A(_source_stream_matmul_15_source_20_pat_size_buf_3), .B(_source_stream_matmul_15_source_20_pat_size_3), .S(_05798_), .Y(_22881_) );
  \$mux  #( .WIDTH(33) ) _42345_ ( .A(_source_stream_matmul_15_source_20_pat_size_buf_2), .B(_source_stream_matmul_15_source_20_pat_size_2), .S(_05798_), .Y(_22882_) );
  \$mux  #( .WIDTH(33) ) _42347_ ( .A(_source_stream_matmul_15_source_20_pat_size_buf_1), .B(_source_stream_matmul_15_source_20_pat_size_1), .S(_05798_), .Y(_22883_) );
  \$mux  #( .WIDTH(33) ) _42349_ ( .A(_source_stream_matmul_15_source_20_pat_size_buf_0), .B(_source_stream_matmul_15_source_20_pat_size_0), .S(_05798_), .Y(_22884_) );
  \$mux  #( .WIDTH(33) ) _42351_ ( .A(_source_stream_matmul_15_source_20_pat_count_3), .B(_26311_), .S(_05798_), .Y(_22885_) );
  \$mux  #( .WIDTH(33) ) _42352_ ( .A(_22885_), .B(_26318_), .S(_05801_), .Y(_22886_) );
  \$mux  #( .WIDTH(33) ) _42353_ ( .A(_22886_), .B(_26319_), .S(_05802_), .Y(_22887_) );
  \$mux  #( .WIDTH(33) ) _42355_ ( .A(_source_stream_matmul_15_source_20_pat_count_2), .B(_26310_), .S(_05798_), .Y(_22888_) );
  \$mux  #( .WIDTH(33) ) _42356_ ( .A(_22888_), .B(_26316_), .S(_05800_), .Y(_22889_) );
  \$mux  #( .WIDTH(33) ) _42357_ ( .A(_22889_), .B(_26317_), .S(_05801_), .Y(_22890_) );
  \$mux  #( .WIDTH(33) ) _42359_ ( .A(_source_stream_matmul_15_source_20_pat_count_1), .B(_26309_), .S(_05798_), .Y(_22891_) );
  \$mux  #( .WIDTH(33) ) _42360_ ( .A(_22891_), .B(_26314_), .S(_05799_), .Y(_22892_) );
  \$mux  #( .WIDTH(33) ) _42361_ ( .A(_22892_), .B(_26315_), .S(_05800_), .Y(_22893_) );
  \$mux  #( .WIDTH(33) ) _42363_ ( .A(_source_stream_matmul_15_source_20_pat_count_0), .B(_26308_), .S(_05798_), .Y(_22894_) );
  \$mux  #( .WIDTH(33) ) _42364_ ( .A(_26312_), .B(_22894_), .S(_05020_), .Y(_22895_) );
  \$mux  #( .WIDTH(33) ) _42365_ ( .A(_22895_), .B(_26313_), .S(_05799_), .Y(_22896_) );
  \$mux  #( .WIDTH(32) ) _42367_ ( .A(_source_stream_matmul_15_source_20_pat_stride_3), .B(0), .S(_set_flag_1034), .Y(_22897_) );
  \$mux  #( .WIDTH(32) ) _42369_ ( .A(_source_stream_matmul_15_source_20_pat_stride_2), .B(0), .S(_set_flag_1034), .Y(_22898_) );
  \$mux  #( .WIDTH(32) ) _42371_ ( .A(_source_stream_matmul_15_source_20_pat_stride_1), .B(288), .S(_set_flag_1034), .Y(_22899_) );
  \$mux  #( .WIDTH(32) ) _42373_ ( .A(_source_stream_matmul_15_source_20_pat_stride_0), .B(1), .S(_set_flag_1034), .Y(_22900_) );
  \$mux  #( .WIDTH(33) ) _42375_ ( .A(_source_stream_matmul_15_source_20_pat_size_3), .B(33'h000000001), .S(_set_flag_1034), .Y(_22901_) );
  \$mux  #( .WIDTH(33) ) _42377_ ( .A(_source_stream_matmul_15_source_20_pat_size_2), .B(33'h000000001), .S(_set_flag_1034), .Y(_22902_) );
  \$mux  #( .WIDTH(33) ) _42379_ ( .A(_source_stream_matmul_15_source_20_pat_size_1), .B({ 1'h0, matmul_15_next_stream_num_ops }), .S(_set_flag_1034), .Y(_22903_) );
  \$mux  #( .WIDTH(33) ) _42381_ ( .A(_source_stream_matmul_15_source_20_pat_size_0), .B(33'h000000120), .S(_set_flag_1034), .Y(_22904_) );
  \$mux  #( .WIDTH(32) ) _42383_ ( .A(_source_stream_matmul_15_source_20_pat_cur_offset_3), .B(0), .S(_05798_), .Y(_22905_) );
  \$mux  #( .WIDTH(32) ) _42384_ ( .A(_22905_), .B(_22260_), .S(_05801_), .Y(_22906_) );
  \$mux  #( .WIDTH(32) ) _42385_ ( .A(_22906_), .B(0), .S(_05802_), .Y(_22907_) );
  \$mux  #( .WIDTH(32) ) _42387_ ( .A(_source_stream_matmul_15_source_20_pat_cur_offset_2), .B(0), .S(_05798_), .Y(_22908_) );
  \$mux  #( .WIDTH(32) ) _42388_ ( .A(_22908_), .B(_22259_), .S(_05800_), .Y(_22909_) );
  \$mux  #( .WIDTH(32) ) _42389_ ( .A(_22909_), .B(0), .S(_05801_), .Y(_22910_) );
  \$mux  #( .WIDTH(32) ) _42391_ ( .A(_source_stream_matmul_15_source_20_pat_cur_offset_1), .B(0), .S(_05798_), .Y(_22911_) );
  \$mux  #( .WIDTH(32) ) _42392_ ( .A(_22911_), .B(_22258_), .S(_05799_), .Y(_22912_) );
  \$mux  #( .WIDTH(32) ) _42393_ ( .A(_22912_), .B(0), .S(_05800_), .Y(_22913_) );
  \$mux  #( .WIDTH(32) ) _42395_ ( .A(_source_stream_matmul_15_source_20_pat_cur_offset_0), .B(0), .S(_05798_), .Y(_22914_) );
  \$mux  #( .WIDTH(32) ) _42396_ ( .A(_22257_), .B(_22914_), .S(_05020_), .Y(_22915_) );
  \$mux  #( .WIDTH(32) ) _42397_ ( .A(_22915_), .B(0), .S(_05799_), .Y(_22916_) );
  \$mux  #( .WIDTH(8) ) _42399_ ( .A(__variable_wdata_830), .B(_stream_matmul_15_source_19_source_ram_rdata), .S(_stream_matmul_15_source_19_source_ram_rvalid), .Y(_22917_) );
  \$mux  #( .WIDTH(32) ) _42401_ ( .A(_source_stream_matmul_15_source_19_pat_stride_buf_3), .B(_source_stream_matmul_15_source_19_pat_stride_3), .S(_05793_), .Y(_22918_) );
  \$mux  #( .WIDTH(32) ) _42403_ ( .A(_source_stream_matmul_15_source_19_pat_stride_buf_2), .B(_source_stream_matmul_15_source_19_pat_stride_2), .S(_05793_), .Y(_22919_) );
  \$mux  #( .WIDTH(32) ) _42405_ ( .A(_source_stream_matmul_15_source_19_pat_stride_buf_1), .B(_source_stream_matmul_15_source_19_pat_stride_1), .S(_05793_), .Y(_22920_) );
  \$mux  #( .WIDTH(32) ) _42407_ ( .A(_source_stream_matmul_15_source_19_pat_stride_buf_0), .B(_source_stream_matmul_15_source_19_pat_stride_0), .S(_05793_), .Y(_22921_) );
  \$mux  #( .WIDTH(33) ) _42409_ ( .A(_source_stream_matmul_15_source_19_pat_size_buf_3), .B(_source_stream_matmul_15_source_19_pat_size_3), .S(_05793_), .Y(_22922_) );
  \$mux  #( .WIDTH(33) ) _42411_ ( .A(_source_stream_matmul_15_source_19_pat_size_buf_2), .B(_source_stream_matmul_15_source_19_pat_size_2), .S(_05793_), .Y(_22923_) );
  \$mux  #( .WIDTH(33) ) _42413_ ( .A(_source_stream_matmul_15_source_19_pat_size_buf_1), .B(_source_stream_matmul_15_source_19_pat_size_1), .S(_05793_), .Y(_22924_) );
  \$mux  #( .WIDTH(33) ) _42415_ ( .A(_source_stream_matmul_15_source_19_pat_size_buf_0), .B(_source_stream_matmul_15_source_19_pat_size_0), .S(_05793_), .Y(_22925_) );
  \$mux  #( .WIDTH(33) ) _42417_ ( .A(_source_stream_matmul_15_source_19_pat_count_3), .B(_26299_), .S(_05793_), .Y(_22926_) );
  \$mux  #( .WIDTH(33) ) _42418_ ( .A(_22926_), .B(_26306_), .S(_05796_), .Y(_22927_) );
  \$mux  #( .WIDTH(33) ) _42419_ ( .A(_22927_), .B(_26307_), .S(_05797_), .Y(_22928_) );
  \$mux  #( .WIDTH(33) ) _42421_ ( .A(_source_stream_matmul_15_source_19_pat_count_2), .B(_26298_), .S(_05793_), .Y(_22929_) );
  \$mux  #( .WIDTH(33) ) _42422_ ( .A(_22929_), .B(_26304_), .S(_05795_), .Y(_22930_) );
  \$mux  #( .WIDTH(33) ) _42423_ ( .A(_22930_), .B(_26305_), .S(_05796_), .Y(_22931_) );
  \$mux  #( .WIDTH(33) ) _42425_ ( .A(_source_stream_matmul_15_source_19_pat_count_1), .B(_26297_), .S(_05793_), .Y(_22932_) );
  \$mux  #( .WIDTH(33) ) _42426_ ( .A(_22932_), .B(_26302_), .S(_05794_), .Y(_22933_) );
  \$mux  #( .WIDTH(33) ) _42427_ ( .A(_22933_), .B(_26303_), .S(_05795_), .Y(_22934_) );
  \$mux  #( .WIDTH(33) ) _42429_ ( .A(_source_stream_matmul_15_source_19_pat_count_0), .B(_26296_), .S(_05793_), .Y(_22935_) );
  \$mux  #( .WIDTH(33) ) _42430_ ( .A(_26300_), .B(_22935_), .S(_05021_), .Y(_22936_) );
  \$mux  #( .WIDTH(33) ) _42431_ ( .A(_22936_), .B(_26301_), .S(_05794_), .Y(_22937_) );
  \$mux  #( .WIDTH(32) ) _42433_ ( .A(_source_stream_matmul_15_source_19_pat_stride_3), .B(0), .S(_set_flag_1034), .Y(_22938_) );
  \$mux  #( .WIDTH(32) ) _42435_ ( .A(_source_stream_matmul_15_source_19_pat_stride_2), .B(0), .S(_set_flag_1034), .Y(_22939_) );
  \$mux  #( .WIDTH(32) ) _42437_ ( .A(_source_stream_matmul_15_source_19_pat_stride_1), .B(0), .S(_set_flag_1034), .Y(_22940_) );
  \$mux  #( .WIDTH(32) ) _42439_ ( .A(_source_stream_matmul_15_source_19_pat_stride_0), .B(1), .S(_set_flag_1034), .Y(_22941_) );
  \$mux  #( .WIDTH(33) ) _42441_ ( .A(_source_stream_matmul_15_source_19_pat_size_3), .B(33'h000000001), .S(_set_flag_1034), .Y(_22942_) );
  \$mux  #( .WIDTH(33) ) _42443_ ( .A(_source_stream_matmul_15_source_19_pat_size_2), .B(33'h000000001), .S(_set_flag_1034), .Y(_22943_) );
  \$mux  #( .WIDTH(33) ) _42445_ ( .A(_source_stream_matmul_15_source_19_pat_size_1), .B({ 1'h0, matmul_15_next_stream_num_ops }), .S(_set_flag_1034), .Y(_22944_) );
  \$mux  #( .WIDTH(33) ) _42447_ ( .A(_source_stream_matmul_15_source_19_pat_size_0), .B(33'h000000120), .S(_set_flag_1034), .Y(_22945_) );
  \$mux  #( .WIDTH(32) ) _42449_ ( .A(_source_stream_matmul_15_source_19_pat_cur_offset_3), .B(0), .S(_05793_), .Y(_22946_) );
  \$mux  #( .WIDTH(32) ) _42450_ ( .A(_22946_), .B(_22256_), .S(_05796_), .Y(_22947_) );
  \$mux  #( .WIDTH(32) ) _42451_ ( .A(_22947_), .B(0), .S(_05797_), .Y(_22948_) );
  \$mux  #( .WIDTH(32) ) _42453_ ( .A(_source_stream_matmul_15_source_19_pat_cur_offset_2), .B(0), .S(_05793_), .Y(_22949_) );
  \$mux  #( .WIDTH(32) ) _42454_ ( .A(_22949_), .B(_22255_), .S(_05795_), .Y(_22950_) );
  \$mux  #( .WIDTH(32) ) _42455_ ( .A(_22950_), .B(0), .S(_05796_), .Y(_22951_) );
  \$mux  #( .WIDTH(32) ) _42457_ ( .A(_source_stream_matmul_15_source_19_pat_cur_offset_1), .B(0), .S(_05793_), .Y(_22952_) );
  \$mux  #( .WIDTH(32) ) _42458_ ( .A(_22952_), .B(_22254_), .S(_05794_), .Y(_22953_) );
  \$mux  #( .WIDTH(32) ) _42459_ ( .A(_22953_), .B(0), .S(_05795_), .Y(_22954_) );
  \$mux  #( .WIDTH(32) ) _42461_ ( .A(_source_stream_matmul_15_source_19_pat_cur_offset_0), .B(0), .S(_05793_), .Y(_22955_) );
  \$mux  #( .WIDTH(32) ) _42462_ ( .A(_22253_), .B(_22955_), .S(_05021_), .Y(_22956_) );
  \$mux  #( .WIDTH(32) ) _42463_ ( .A(_22956_), .B(0), .S(_05794_), .Y(_22957_) );
  \$mux  #( .WIDTH(4) ) _42465_ ( .A(__variable_wdata_828), .B(_stream_matmul_15_constant_17_next_constant_data), .S(_stream_matmul_15_start), .Y(_22958_) );
  \$mux  #( .WIDTH(1) ) _42467_ ( .A(__variable_wdata_827), .B(_stream_matmul_15_constant_16_next_constant_data), .S(_stream_matmul_15_start), .Y(_22959_) );
  \$mux  #( .WIDTH(1) ) _42469_ ( .A(__variable_wdata_826), .B(_stream_matmul_15_constant_15_next_constant_data), .S(_stream_matmul_15_start), .Y(_22960_) );
  \$mux  #( .WIDTH(8) ) _42471_ ( .A(__variable_wdata_820), .B(_stream_matmul_15_source_14_source_empty_data), .S(_stream_matmul_15_start), .Y(_22961_) );
  \$mux  #( .WIDTH(8) ) _42473_ ( .A(__variable_wdata_813), .B(_stream_matmul_15_source_12_source_empty_data), .S(_stream_matmul_15_start), .Y(_22962_) );
  \$mux  #( .WIDTH(8) ) _42475_ ( .A(__variable_wdata_806), .B(_stream_matmul_15_source_10_source_empty_data), .S(_stream_matmul_15_start), .Y(_22963_) );
  \$mux  #( .WIDTH(8) ) _42477_ ( .A(__variable_wdata_799), .B(_stream_matmul_15_source_8_source_ram_rdata), .S(_stream_matmul_15_source_8_source_ram_rvalid), .Y(_22964_) );
  \$mux  #( .WIDTH(32) ) _42479_ ( .A(_source_stream_matmul_15_source_8_pat_stride_buf_3), .B(_source_stream_matmul_15_source_8_pat_stride_3), .S(_05788_), .Y(_22965_) );
  \$mux  #( .WIDTH(32) ) _42481_ ( .A(_source_stream_matmul_15_source_8_pat_stride_buf_2), .B(_source_stream_matmul_15_source_8_pat_stride_2), .S(_05788_), .Y(_22966_) );
  \$mux  #( .WIDTH(32) ) _42483_ ( .A(_source_stream_matmul_15_source_8_pat_stride_buf_1), .B(_source_stream_matmul_15_source_8_pat_stride_1), .S(_05788_), .Y(_22967_) );
  \$mux  #( .WIDTH(32) ) _42485_ ( .A(_source_stream_matmul_15_source_8_pat_stride_buf_0), .B(_source_stream_matmul_15_source_8_pat_stride_0), .S(_05788_), .Y(_22968_) );
  \$mux  #( .WIDTH(33) ) _42487_ ( .A(_source_stream_matmul_15_source_8_pat_size_buf_3), .B(_source_stream_matmul_15_source_8_pat_size_3), .S(_05788_), .Y(_22969_) );
  \$mux  #( .WIDTH(33) ) _42489_ ( .A(_source_stream_matmul_15_source_8_pat_size_buf_2), .B(_source_stream_matmul_15_source_8_pat_size_2), .S(_05788_), .Y(_22970_) );
  \$mux  #( .WIDTH(33) ) _42491_ ( .A(_source_stream_matmul_15_source_8_pat_size_buf_1), .B(_source_stream_matmul_15_source_8_pat_size_1), .S(_05788_), .Y(_22971_) );
  \$mux  #( .WIDTH(33) ) _42493_ ( .A(_source_stream_matmul_15_source_8_pat_size_buf_0), .B(_source_stream_matmul_15_source_8_pat_size_0), .S(_05788_), .Y(_22972_) );
  \$mux  #( .WIDTH(33) ) _42495_ ( .A(_source_stream_matmul_15_source_8_pat_count_3), .B(_26287_), .S(_05788_), .Y(_22973_) );
  \$mux  #( .WIDTH(33) ) _42496_ ( .A(_22973_), .B(_26294_), .S(_05791_), .Y(_22974_) );
  \$mux  #( .WIDTH(33) ) _42497_ ( .A(_22974_), .B(_26295_), .S(_05792_), .Y(_22975_) );
  \$mux  #( .WIDTH(33) ) _42499_ ( .A(_source_stream_matmul_15_source_8_pat_count_2), .B(_26286_), .S(_05788_), .Y(_22976_) );
  \$mux  #( .WIDTH(33) ) _42500_ ( .A(_22976_), .B(_26292_), .S(_05790_), .Y(_22977_) );
  \$mux  #( .WIDTH(33) ) _42501_ ( .A(_22977_), .B(_26293_), .S(_05791_), .Y(_22978_) );
  \$mux  #( .WIDTH(33) ) _42503_ ( .A(_source_stream_matmul_15_source_8_pat_count_1), .B(_26285_), .S(_05788_), .Y(_22979_) );
  \$mux  #( .WIDTH(33) ) _42504_ ( .A(_22979_), .B(_26290_), .S(_05789_), .Y(_22980_) );
  \$mux  #( .WIDTH(33) ) _42505_ ( .A(_22980_), .B(_26291_), .S(_05790_), .Y(_22981_) );
  \$mux  #( .WIDTH(33) ) _42507_ ( .A(_source_stream_matmul_15_source_8_pat_count_0), .B(_26284_), .S(_05788_), .Y(_22982_) );
  \$mux  #( .WIDTH(33) ) _42508_ ( .A(_26288_), .B(_22982_), .S(_05025_), .Y(_22983_) );
  \$mux  #( .WIDTH(33) ) _42509_ ( .A(_22983_), .B(_26289_), .S(_05789_), .Y(_22984_) );
  \$mux  #( .WIDTH(32) ) _42511_ ( .A(_source_stream_matmul_15_source_8_pat_stride_3), .B(0), .S(_set_flag_1034), .Y(_22985_) );
  \$mux  #( .WIDTH(32) ) _42513_ ( .A(_source_stream_matmul_15_source_8_pat_stride_2), .B(0), .S(_set_flag_1034), .Y(_22986_) );
  \$mux  #( .WIDTH(32) ) _42515_ ( .A(_source_stream_matmul_15_source_8_pat_stride_1), .B(0), .S(_set_flag_1034), .Y(_22987_) );
  \$mux  #( .WIDTH(32) ) _42517_ ( .A(_source_stream_matmul_15_source_8_pat_stride_0), .B(0), .S(_set_flag_1034), .Y(_22988_) );
  \$mux  #( .WIDTH(33) ) _42519_ ( .A(_source_stream_matmul_15_source_8_pat_size_3), .B(33'h000000001), .S(_set_flag_1034), .Y(_22989_) );
  \$mux  #( .WIDTH(33) ) _42521_ ( .A(_source_stream_matmul_15_source_8_pat_size_2), .B(33'h000000001), .S(_set_flag_1034), .Y(_22990_) );
  \$mux  #( .WIDTH(33) ) _42523_ ( .A(_source_stream_matmul_15_source_8_pat_size_1), .B({ 1'h0, matmul_15_next_stream_num_ops }), .S(_set_flag_1034), .Y(_22991_) );
  \$mux  #( .WIDTH(33) ) _42525_ ( .A(_source_stream_matmul_15_source_8_pat_size_0), .B(33'h000000120), .S(_set_flag_1034), .Y(_22992_) );
  \$mux  #( .WIDTH(32) ) _42527_ ( .A(_source_stream_matmul_15_source_8_pat_cur_offset_3), .B(0), .S(_05788_), .Y(_22993_) );
  \$mux  #( .WIDTH(32) ) _42528_ ( .A(_22993_), .B(_22251_), .S(_05791_), .Y(_22994_) );
  \$mux  #( .WIDTH(32) ) _42529_ ( .A(_22994_), .B(0), .S(_05792_), .Y(_22995_) );
  \$mux  #( .WIDTH(32) ) _42531_ ( .A(_source_stream_matmul_15_source_8_pat_cur_offset_2), .B(0), .S(_05788_), .Y(_22996_) );
  \$mux  #( .WIDTH(32) ) _42532_ ( .A(_22996_), .B(_22250_), .S(_05790_), .Y(_22997_) );
  \$mux  #( .WIDTH(32) ) _42533_ ( .A(_22997_), .B(0), .S(_05791_), .Y(_22998_) );
  \$mux  #( .WIDTH(32) ) _42535_ ( .A(_source_stream_matmul_15_source_8_pat_cur_offset_1), .B(0), .S(_05788_), .Y(_22999_) );
  \$mux  #( .WIDTH(32) ) _42536_ ( .A(_22999_), .B(_22249_), .S(_05789_), .Y(_23000_) );
  \$mux  #( .WIDTH(32) ) _42537_ ( .A(_23000_), .B(0), .S(_05790_), .Y(_23001_) );
  \$mux  #( .WIDTH(32) ) _42539_ ( .A(_source_stream_matmul_15_source_8_pat_cur_offset_0), .B(0), .S(_05788_), .Y(_23002_) );
  \$mux  #( .WIDTH(32) ) _42540_ ( .A(_22248_), .B(_23002_), .S(_05025_), .Y(_23003_) );
  \$mux  #( .WIDTH(32) ) _42541_ ( .A(_23003_), .B(0), .S(_05789_), .Y(_23004_) );
  \$mux  #( .WIDTH(32) ) _42543_ ( .A(__variable_wdata_792), .B(_stream_matmul_15_source_6_source_ram_rdata), .S(_stream_matmul_15_source_6_source_ram_rvalid), .Y(_23005_) );
  \$mux  #( .WIDTH(32) ) _42545_ ( .A(_source_stream_matmul_15_source_6_pat_stride_buf_3), .B(_source_stream_matmul_15_source_6_pat_stride_3), .S(_05783_), .Y(_23006_) );
  \$mux  #( .WIDTH(32) ) _42547_ ( .A(_source_stream_matmul_15_source_6_pat_stride_buf_2), .B(_source_stream_matmul_15_source_6_pat_stride_2), .S(_05783_), .Y(_23007_) );
  \$mux  #( .WIDTH(32) ) _42549_ ( .A(_source_stream_matmul_15_source_6_pat_stride_buf_1), .B(_source_stream_matmul_15_source_6_pat_stride_1), .S(_05783_), .Y(_23008_) );
  \$mux  #( .WIDTH(32) ) _42551_ ( .A(_source_stream_matmul_15_source_6_pat_stride_buf_0), .B(_source_stream_matmul_15_source_6_pat_stride_0), .S(_05783_), .Y(_23009_) );
  \$mux  #( .WIDTH(33) ) _42553_ ( .A(_source_stream_matmul_15_source_6_pat_size_buf_3), .B(_source_stream_matmul_15_source_6_pat_size_3), .S(_05783_), .Y(_23010_) );
  \$mux  #( .WIDTH(33) ) _42555_ ( .A(_source_stream_matmul_15_source_6_pat_size_buf_2), .B(_source_stream_matmul_15_source_6_pat_size_2), .S(_05783_), .Y(_23011_) );
  \$mux  #( .WIDTH(33) ) _42557_ ( .A(_source_stream_matmul_15_source_6_pat_size_buf_1), .B(_source_stream_matmul_15_source_6_pat_size_1), .S(_05783_), .Y(_23012_) );
  \$mux  #( .WIDTH(33) ) _42559_ ( .A(_source_stream_matmul_15_source_6_pat_size_buf_0), .B(_source_stream_matmul_15_source_6_pat_size_0), .S(_05783_), .Y(_23013_) );
  \$mux  #( .WIDTH(33) ) _42561_ ( .A(_source_stream_matmul_15_source_6_pat_count_3), .B(_26275_), .S(_05783_), .Y(_23014_) );
  \$mux  #( .WIDTH(33) ) _42562_ ( .A(_23014_), .B(_26282_), .S(_05786_), .Y(_23015_) );
  \$mux  #( .WIDTH(33) ) _42563_ ( .A(_23015_), .B(_26283_), .S(_05787_), .Y(_23016_) );
  \$mux  #( .WIDTH(33) ) _42565_ ( .A(_source_stream_matmul_15_source_6_pat_count_2), .B(_26274_), .S(_05783_), .Y(_23017_) );
  \$mux  #( .WIDTH(33) ) _42566_ ( .A(_23017_), .B(_26280_), .S(_05785_), .Y(_23018_) );
  \$mux  #( .WIDTH(33) ) _42567_ ( .A(_23018_), .B(_26281_), .S(_05786_), .Y(_23019_) );
  \$mux  #( .WIDTH(33) ) _42569_ ( .A(_source_stream_matmul_15_source_6_pat_count_1), .B(_26273_), .S(_05783_), .Y(_23020_) );
  \$mux  #( .WIDTH(33) ) _42570_ ( .A(_23020_), .B(_26278_), .S(_05784_), .Y(_23021_) );
  \$mux  #( .WIDTH(33) ) _42571_ ( .A(_23021_), .B(_26279_), .S(_05785_), .Y(_23022_) );
  \$mux  #( .WIDTH(33) ) _42573_ ( .A(_source_stream_matmul_15_source_6_pat_count_0), .B(_26272_), .S(_05783_), .Y(_23023_) );
  \$mux  #( .WIDTH(33) ) _42574_ ( .A(_26276_), .B(_23023_), .S(_05023_), .Y(_23024_) );
  \$mux  #( .WIDTH(33) ) _42575_ ( .A(_23024_), .B(_26277_), .S(_05784_), .Y(_23025_) );
  \$mux  #( .WIDTH(32) ) _42577_ ( .A(_source_stream_matmul_15_source_6_pat_stride_3), .B(0), .S(_set_flag_1034), .Y(_23026_) );
  \$mux  #( .WIDTH(32) ) _42579_ ( .A(_source_stream_matmul_15_source_6_pat_stride_2), .B(0), .S(_set_flag_1034), .Y(_23027_) );
  \$mux  #( .WIDTH(32) ) _42581_ ( .A(_source_stream_matmul_15_source_6_pat_stride_1), .B(1), .S(_set_flag_1034), .Y(_23028_) );
  \$mux  #( .WIDTH(32) ) _42583_ ( .A(_source_stream_matmul_15_source_6_pat_stride_0), .B(0), .S(_set_flag_1034), .Y(_23029_) );
  \$mux  #( .WIDTH(33) ) _42585_ ( .A(_source_stream_matmul_15_source_6_pat_size_3), .B(33'h000000001), .S(_set_flag_1034), .Y(_23030_) );
  \$mux  #( .WIDTH(33) ) _42587_ ( .A(_source_stream_matmul_15_source_6_pat_size_2), .B(33'h000000001), .S(_set_flag_1034), .Y(_23031_) );
  \$mux  #( .WIDTH(33) ) _42589_ ( .A(_source_stream_matmul_15_source_6_pat_size_1), .B({ 1'h0, matmul_15_next_stream_num_ops }), .S(_set_flag_1034), .Y(_23032_) );
  \$mux  #( .WIDTH(33) ) _42591_ ( .A(_source_stream_matmul_15_source_6_pat_size_0), .B(33'h000000120), .S(_set_flag_1034), .Y(_23033_) );
  \$mux  #( .WIDTH(32) ) _42593_ ( .A(_source_stream_matmul_15_source_6_pat_cur_offset_3), .B(0), .S(_05783_), .Y(_23034_) );
  \$mux  #( .WIDTH(32) ) _42594_ ( .A(_23034_), .B(_22247_), .S(_05786_), .Y(_23035_) );
  \$mux  #( .WIDTH(32) ) _42595_ ( .A(_23035_), .B(0), .S(_05787_), .Y(_23036_) );
  \$mux  #( .WIDTH(32) ) _42597_ ( .A(_source_stream_matmul_15_source_6_pat_cur_offset_2), .B(0), .S(_05783_), .Y(_23037_) );
  \$mux  #( .WIDTH(32) ) _42598_ ( .A(_23037_), .B(_22246_), .S(_05785_), .Y(_23038_) );
  \$mux  #( .WIDTH(32) ) _42599_ ( .A(_23038_), .B(0), .S(_05786_), .Y(_23039_) );
  \$mux  #( .WIDTH(32) ) _42601_ ( .A(_source_stream_matmul_15_source_6_pat_cur_offset_1), .B(0), .S(_05783_), .Y(_23040_) );
  \$mux  #( .WIDTH(32) ) _42602_ ( .A(_23040_), .B(_22245_), .S(_05784_), .Y(_23041_) );
  \$mux  #( .WIDTH(32) ) _42603_ ( .A(_23041_), .B(0), .S(_05785_), .Y(_23042_) );
  \$mux  #( .WIDTH(32) ) _42605_ ( .A(_source_stream_matmul_15_source_6_pat_cur_offset_0), .B(0), .S(_05783_), .Y(_23043_) );
  \$mux  #( .WIDTH(32) ) _42606_ ( .A(_22244_), .B(_23043_), .S(_05023_), .Y(_23044_) );
  \$mux  #( .WIDTH(32) ) _42607_ ( .A(_23044_), .B(0), .S(_05784_), .Y(_23045_) );
  \$mux  #( .WIDTH(1) ) _42609_ ( .A(__variable_wdata_779), .B(_stream_matmul_15_constant_3_next_constant_data), .S(_stream_matmul_15_start), .Y(_23046_) );
  \$mux  #( .WIDTH(1) ) _42611_ ( .A(__variable_wdata_778), .B(_stream_matmul_15_constant_2_next_constant_data), .S(_stream_matmul_15_start), .Y(_23047_) );
  \$mux  #( .WIDTH(1) ) _42613_ ( .A(__variable_wdata_777), .B(_stream_matmul_15_constant_1_next_constant_data), .S(_stream_matmul_15_start), .Y(_23048_) );
  \$mux  #( .WIDTH(9) ) _42615_ ( .A(__variable_wdata_776), .B(_stream_matmul_15_constant_0_next_constant_data), .S(_stream_matmul_15_start), .Y(_23049_) );
  \$mux  #( .WIDTH(1) ) _42617_ ( .A(1'h1), .B(1'h0), .S(_05027_), .Y(_22875_) );
  \$mux  #( .WIDTH(8) ) _42746_ ( .A(_stream_matmul_15_sink_21_sink_wdata), .B(__substreamoutput_data_866), .S(_05804_), .Y(_23050_) );
  \$mux  #( .WIDTH(1) ) _42748_ ( .A(1'h0), .B(1'h1), .S(_05804_), .Y(_23051_) );
  \$mux  #( .WIDTH(32) ) _42750_ ( .A(_stream_matmul_15_sink_21_sink_waddr), .B(_26320_), .S(_05803_), .Y(_23052_) );
  \$mux  #( .WIDTH(32) ) _42751_ ( .A(_23052_), .B(_22262_), .S(_05804_), .Y(_23053_) );
  \$mux  #( .WIDTH(8) ) _42753_ ( .A(_stream_matmul_15_sink_21_sink_ram_sel), .B(8'h05), .S(__set_flag_1034_37), .Y(_23054_) );
  \$mux  #( .WIDTH(32) ) _42755_ ( .A(_stream_matmul_15_sink_21_sink_stride_buf), .B(_stream_matmul_15_sink_21_sink_stride), .S(_05803_), .Y(_23055_) );
  \$mux  #( .WIDTH(33) ) _42757_ ( .A(_stream_matmul_15_sink_21_sink_count), .B(_stream_matmul_15_sink_21_sink_size), .S(_05803_), .Y(_23056_) );
  \$mux  #( .WIDTH(33) ) _42758_ ( .A(_23056_), .B(_26321_), .S(_05804_), .Y(_23057_) );
  \$mux  #( .WIDTH(32) ) _42760_ ( .A(_stream_matmul_15_sink_21_sink_stride), .B(1), .S(__set_flag_1034_37), .Y(_23058_) );
  \$mux  #( .WIDTH(33) ) _42762_ ( .A(_stream_matmul_15_sink_21_sink_size), .B(__stream_matmul_15_sink_21_sink_size_1_37), .S(__set_flag_1034_37), .Y(_23059_) );
  \$mux  #( .WIDTH(32) ) _42764_ ( .A(_stream_matmul_15_sink_21_sink_offset), .B(__stream_matmul_15_sink_21_sink_offset_0_37), .S(__set_flag_1034_37), .Y(_23060_) );
  \$mux  #( .WIDTH(3) ) _42766_ ( .A(_stream_matmul_15_sink_21_sink_mode), .B(3'h1), .S(__set_flag_1034_37), .Y(_23061_) );
  \$mux  #( .WIDTH(1) ) _42768_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l4096_id0_3_cond_1_1), .Y(_23062_) );
  \$mux  #( .WIDTH(1) ) _42770_ ( .A(1'h1), .B(_stream_matmul_15_source_20_source_ram_renable), .S(_05020_), .Y(_23063_) );
  \$mux  #( .WIDTH(1) ) _42771_ ( .A(1'h0), .B(_23063_), .S(_05019_), .Y(_23064_) );
  \$mux  #( .WIDTH(32) ) _42773_ ( .A(_stream_matmul_15_source_20_source_pat_all_offset), .B(_stream_matmul_15_source_20_source_ram_raddr), .S(_05020_), .Y(_23065_) );
  \$mux  #( .WIDTH(8) ) _42775_ ( .A(_stream_matmul_15_source_20_source_ram_sel), .B(8'h04), .S(_set_flag_1034), .Y(_23066_) );
  \$mux  #( .WIDTH(32) ) _42777_ ( .A(_stream_matmul_15_source_20_source_offset_buf), .B(_stream_matmul_15_source_20_source_offset), .S(_05798_), .Y(_23067_) );
  \$mux  #( .WIDTH(32) ) _42779_ ( .A(_stream_matmul_15_source_20_source_offset), .B(matmul_15_filter_page_comp_offset_buf), .S(_set_flag_1034), .Y(_23068_) );
  \$mux  #( .WIDTH(3) ) _42781_ ( .A(_stream_matmul_15_source_20_source_mode), .B(3'h2), .S(_set_flag_1034), .Y(_23069_) );
  \$mux  #( .WIDTH(1) ) _42783_ ( .A(_stream_matmul_15_source_20_idle), .B(1'h0), .S(_05798_), .Y(_23070_) );
  \$mux  #( .WIDTH(1) ) _42784_ ( .A(1'h1), .B(_23070_), .S(_05019_), .Y(_23071_) );
  \$mux  #( .WIDTH(1) ) _42785_ ( .A(_23071_), .B(1'h1), .S(RST), .Y(_02613_) );
  \$mux  #( .WIDTH(1) ) _42786_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id2_3_cond_4_1), .Y(_23072_) );
  \$mux  #( .WIDTH(1) ) _42788_ ( .A(1'h1), .B(_stream_matmul_15_source_19_source_ram_renable), .S(_05021_), .Y(_23073_) );
  \$mux  #( .WIDTH(1) ) _42789_ ( .A(1'h0), .B(_23073_), .S(_05022_), .Y(_23074_) );
  \$mux  #( .WIDTH(32) ) _42791_ ( .A(_stream_matmul_15_source_19_source_pat_all_offset), .B(_stream_matmul_15_source_19_source_ram_raddr), .S(_05021_), .Y(_23075_) );
  \$mux  #( .WIDTH(8) ) _42793_ ( .A(_stream_matmul_15_source_19_source_ram_sel), .B(8'h03), .S(_set_flag_1034), .Y(_23076_) );
  \$mux  #( .WIDTH(32) ) _42795_ ( .A(_stream_matmul_15_source_19_source_offset_buf), .B(_stream_matmul_15_source_19_source_offset), .S(_05793_), .Y(_23077_) );
  \$mux  #( .WIDTH(32) ) _42797_ ( .A(_stream_matmul_15_source_19_source_offset), .B(_22252_), .S(_set_flag_1034), .Y(_23078_) );
  \$mux  #( .WIDTH(3) ) _42799_ ( .A(_stream_matmul_15_source_19_source_mode), .B(3'h2), .S(_set_flag_1034), .Y(_23079_) );
  \$mux  #( .WIDTH(1) ) _42801_ ( .A(_stream_matmul_15_source_19_idle), .B(1'h0), .S(_05793_), .Y(_23080_) );
  \$mux  #( .WIDTH(1) ) _42802_ ( .A(1'h1), .B(_23080_), .S(_05022_), .Y(_23081_) );
  \$mux  #( .WIDTH(1) ) _42803_ ( .A(_23081_), .B(1'h1), .S(RST), .Y(_02604_) );
  \$mux  #( .WIDTH(4) ) _42804_ ( .A(_stream_matmul_15_constant_17_next_constant_data), .B(4'h8), .S(_set_flag_1034), .Y(_23082_) );
  \$mux  #( .WIDTH(1) ) _42806_ ( .A(_stream_matmul_15_constant_16_next_constant_data), .B(1'h0), .S(_set_flag_1034), .Y(_23083_) );
  \$mux  #( .WIDTH(1) ) _42808_ ( .A(_stream_matmul_15_constant_15_next_constant_data), .B(1'h0), .S(_set_flag_1034), .Y(_23084_) );
  \$mux  #( .WIDTH(8) ) _42810_ ( .A(_stream_matmul_15_source_14_source_empty_data), .B(8'h00), .S(_set_flag_1034), .Y(_23085_) );
  \$mux  #( .WIDTH(1) ) _42812_ ( .A(_stream_matmul_15_source_14_idle), .B(1'h1), .S(_stream_matmul_15_start), .Y(_23086_) );
  \$mux  #( .WIDTH(1) ) _42813_ ( .A(_23086_), .B(1'h1), .S(RST), .Y(_02602_) );
  \$mux  #( .WIDTH(8) ) _42814_ ( .A(_stream_matmul_15_source_12_source_empty_data), .B(8'h00), .S(_set_flag_1034), .Y(_23087_) );
  \$mux  #( .WIDTH(1) ) _42816_ ( .A(_stream_matmul_15_source_12_idle), .B(1'h1), .S(_stream_matmul_15_start), .Y(_23088_) );
  \$mux  #( .WIDTH(1) ) _42817_ ( .A(_23088_), .B(1'h1), .S(RST), .Y(_02600_) );
  \$mux  #( .WIDTH(8) ) _42818_ ( .A(_stream_matmul_15_source_10_source_empty_data), .B(8'h00), .S(_set_flag_1034), .Y(_23089_) );
  \$mux  #( .WIDTH(1) ) _42820_ ( .A(_stream_matmul_15_source_10_idle), .B(1'h1), .S(_stream_matmul_15_start), .Y(_23090_) );
  \$mux  #( .WIDTH(1) ) _42821_ ( .A(_23090_), .B(1'h1), .S(RST), .Y(_02598_) );
  \$mux  #( .WIDTH(1) ) _42822_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id0_3_cond_4_1), .Y(_23091_) );
  \$mux  #( .WIDTH(1) ) _42824_ ( .A(1'h1), .B(_stream_matmul_15_source_8_source_ram_renable), .S(_05025_), .Y(_23092_) );
  \$mux  #( .WIDTH(1) ) _42825_ ( .A(1'h0), .B(_23092_), .S(_05024_), .Y(_23093_) );
  \$mux  #( .WIDTH(32) ) _42827_ ( .A(_stream_matmul_15_source_8_source_pat_all_offset), .B(_stream_matmul_15_source_8_source_ram_raddr), .S(_05025_), .Y(_23094_) );
  \$mux  #( .WIDTH(8) ) _42829_ ( .A(_stream_matmul_15_source_8_source_ram_sel), .B(8'h02), .S(_set_flag_1034), .Y(_23095_) );
  \$mux  #( .WIDTH(32) ) _42831_ ( .A(_stream_matmul_15_source_8_source_offset_buf), .B(_stream_matmul_15_source_8_source_offset), .S(_05788_), .Y(_23096_) );
  \$mux  #( .WIDTH(32) ) _42833_ ( .A(_stream_matmul_15_source_8_source_offset), .B(0), .S(_set_flag_1034), .Y(_23097_) );
  \$mux  #( .WIDTH(3) ) _42835_ ( .A(_stream_matmul_15_source_8_source_mode), .B(3'h2), .S(_set_flag_1034), .Y(_23098_) );
  \$mux  #( .WIDTH(1) ) _42837_ ( .A(_stream_matmul_15_source_8_idle), .B(1'h0), .S(_05788_), .Y(_23099_) );
  \$mux  #( .WIDTH(1) ) _42838_ ( .A(1'h1), .B(_23099_), .S(_05024_), .Y(_23100_) );
  \$mux  #( .WIDTH(1) ) _42839_ ( .A(_23100_), .B(1'h1), .S(RST), .Y(_02631_) );
  \$mux  #( .WIDTH(1) ) _42840_ ( .A(1'h0), .B(1'h1), .S(_ram_w32_l128_id0_cond_4_1), .Y(_23101_) );
  \$mux  #( .WIDTH(1) ) _42842_ ( .A(1'h1), .B(_stream_matmul_15_source_6_source_ram_renable), .S(_05023_), .Y(_23102_) );
  \$mux  #( .WIDTH(1) ) _42843_ ( .A(1'h0), .B(_23102_), .S(_05026_), .Y(_23103_) );
  \$mux  #( .WIDTH(32) ) _42845_ ( .A(_stream_matmul_15_source_6_source_pat_all_offset), .B(_stream_matmul_15_source_6_source_ram_raddr), .S(_05023_), .Y(_23104_) );
  \$mux  #( .WIDTH(8) ) _42847_ ( .A(_stream_matmul_15_source_6_source_ram_sel), .B(8'h01), .S(_set_flag_1034), .Y(_23105_) );
  \$mux  #( .WIDTH(32) ) _42849_ ( .A(_stream_matmul_15_source_6_source_offset_buf), .B(_stream_matmul_15_source_6_source_offset), .S(_05783_), .Y(_23106_) );
  \$mux  #( .WIDTH(32) ) _42851_ ( .A(_stream_matmul_15_source_6_source_offset), .B(matmul_15_och_count_buf), .S(_set_flag_1034), .Y(_23107_) );
  \$mux  #( .WIDTH(3) ) _42853_ ( .A(_stream_matmul_15_source_6_source_mode), .B(3'h2), .S(_set_flag_1034), .Y(_23108_) );
  \$mux  #( .WIDTH(1) ) _42855_ ( .A(_stream_matmul_15_source_6_idle), .B(1'h0), .S(_05783_), .Y(_23109_) );
  \$mux  #( .WIDTH(1) ) _42856_ ( .A(1'h1), .B(_23109_), .S(_05026_), .Y(_23110_) );
  \$mux  #( .WIDTH(1) ) _42857_ ( .A(_23110_), .B(1'h1), .S(RST), .Y(_02622_) );
  \$mux  #( .WIDTH(1) ) _42858_ ( .A(_stream_matmul_15_constant_3_next_constant_data), .B(matmul_15_stream_pad_masks), .S(_set_flag_1034), .Y(_23111_) );
  \$mux  #( .WIDTH(1) ) _42860_ ( .A(_stream_matmul_15_constant_2_next_constant_data), .B(matmul_15_row_select_buf), .S(_set_flag_1034), .Y(_23112_) );
  \$mux  #( .WIDTH(1) ) _42862_ ( .A(_stream_matmul_15_constant_1_next_constant_data), .B(matmul_15_col_select), .S(_set_flag_1034), .Y(_23113_) );
  \$mux  #( .WIDTH(9) ) _42864_ ( .A(_stream_matmul_15_constant_0_next_constant_data), .B(9'h120), .S(_set_flag_1034), .Y(_23114_) );
  \$mux  #( .WIDTH(1) ) _42866_ ( .A(_stream_max_pool_serial_9_reduce_reset), .B(1'h0), .S(__tmp_884_5), .Y(_23115_) );
  \$mux  #( .WIDTH(1) ) _42867_ ( .A(_23115_), .B(1'h1), .S(__tmp_908_1), .Y(_23116_) );
  \$mux  #( .WIDTH(1) ) _42868_ ( .A(_23116_), .B(1'h1), .S(RST), .Y(_02647_) );
  \$mux  #( .WIDTH(1) ) _42869_ ( .A(_stream_max_pool_serial_9_source_busy), .B(1'h1), .S(_stream_max_pool_serial_9_start_flag), .Y(_21486_) );
  \$mux  #( .WIDTH(1) ) _42871_ ( .A(1'h0), .B(1'h1), .S(__tmp_908_6), .Y(_23118_) );
  \$mux  #( .WIDTH(1) ) _42873_ ( .A(1'h0), .B(1'h1), .S(__tmp_906_10), .Y(_23119_) );
  \$mux  #( .WIDTH(1) ) _42875_ ( .A(1'h0), .B(1'h1), .S(_stream_max_pool_serial_9_start_flag), .Y(_23120_) );
  \$mux  #( .WIDTH(1) ) _42876_ ( .A(_23120_), .B(1'h0), .S(_04902_), .Y(_23121_) );
  \$mux  #( .WIDTH(32) ) _42878_ ( .A(_stream_max_pool_serial_9_fsm), .B(3), .S(_stream_max_pool_serial_9_source_1_idle), .Y({ _21543_, _21542_, _21540_, _21539_, _21538_, _21537_, _21536_, _21535_, _21534_, _21533_, _21532_, _21531_, _21529_, _21528_, _21527_, _21526_, _21525_, _21524_, _21523_, _21522_, _21521_, _21520_, _21550_, _21549_, _21548_, _21547_, _21546_, _21545_, _21544_, _21541_, _21530_, _21519_ }) );
  \$mux  #( .WIDTH(32) ) _42879_ ( .A(_stream_max_pool_serial_9_fsm), .B(1), .S(_stream_max_pool_serial_9_start_flag), .Y({ _21575_, _21574_, _21572_, _21571_, _21570_, _21569_, _21568_, _21567_, _21566_, _21565_, _21564_, _21563_, _21561_, _21560_, _21559_, _21558_, _21557_, _21556_, _21555_, _21554_, _21553_, _21552_, _21582_, _21581_, _21580_, _21579_, _21578_, _21577_, _21576_, _21573_, _21562_, _21551_ }) );
  \$mux  #( .WIDTH(1) ) _42895_ ( .A(1'h1), .B(1'h0), .S(_05046_), .Y(_23123_) );
  \$mux  #( .WIDTH(8) ) _42934_ ( .A(__variable_wdata_758), .B(_stream_max_pool_serial_9_source_1_source_ram_rdata), .S(_stream_max_pool_serial_9_source_1_source_ram_rvalid), .Y(_23125_) );
  \$mux  #( .WIDTH(32) ) _42936_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_stride_buf_3), .B(_source_stream_max_pool_serial_9_source_1_pat_stride_3), .S(_05776_), .Y(_23126_) );
  \$mux  #( .WIDTH(32) ) _42938_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_stride_buf_2), .B(_source_stream_max_pool_serial_9_source_1_pat_stride_2), .S(_05776_), .Y(_23127_) );
  \$mux  #( .WIDTH(32) ) _42940_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_stride_buf_1), .B(_source_stream_max_pool_serial_9_source_1_pat_stride_1), .S(_05776_), .Y(_23128_) );
  \$mux  #( .WIDTH(32) ) _42942_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_stride_buf_0), .B(_source_stream_max_pool_serial_9_source_1_pat_stride_0), .S(_05776_), .Y(_23129_) );
  \$mux  #( .WIDTH(33) ) _42944_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_buf_3), .B(_source_stream_max_pool_serial_9_source_1_pat_size_3), .S(_05776_), .Y(_23130_) );
  \$mux  #( .WIDTH(33) ) _42946_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_buf_2), .B(_source_stream_max_pool_serial_9_source_1_pat_size_2), .S(_05776_), .Y(_23131_) );
  \$mux  #( .WIDTH(33) ) _42948_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_buf_1), .B(_source_stream_max_pool_serial_9_source_1_pat_size_1), .S(_05776_), .Y(_23132_) );
  \$mux  #( .WIDTH(33) ) _42950_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_buf_0), .B(_source_stream_max_pool_serial_9_source_1_pat_size_0), .S(_05776_), .Y(_23133_) );
  \$mux  #( .WIDTH(33) ) _42952_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_3), .B(_26261_), .S(_05776_), .Y(_23134_) );
  \$mux  #( .WIDTH(33) ) _42953_ ( .A(_23134_), .B(_26268_), .S(_05779_), .Y(_23135_) );
  \$mux  #( .WIDTH(33) ) _42954_ ( .A(_23135_), .B(_26269_), .S(_05780_), .Y(_23136_) );
  \$mux  #( .WIDTH(33) ) _42956_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_2), .B(_26260_), .S(_05776_), .Y(_23137_) );
  \$mux  #( .WIDTH(33) ) _42957_ ( .A(_23137_), .B(_26266_), .S(_05778_), .Y(_23138_) );
  \$mux  #( .WIDTH(33) ) _42958_ ( .A(_23138_), .B(_26267_), .S(_05779_), .Y(_23139_) );
  \$mux  #( .WIDTH(33) ) _42960_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_1), .B(_26259_), .S(_05776_), .Y(_23140_) );
  \$mux  #( .WIDTH(33) ) _42961_ ( .A(_23140_), .B(_26264_), .S(_05777_), .Y(_23141_) );
  \$mux  #( .WIDTH(33) ) _42962_ ( .A(_23141_), .B(_26265_), .S(_05778_), .Y(_23142_) );
  \$mux  #( .WIDTH(33) ) _42964_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_count_0), .B(_26258_), .S(_05776_), .Y(_23143_) );
  \$mux  #( .WIDTH(33) ) _42965_ ( .A(_26262_), .B(_23143_), .S(_05043_), .Y(_23144_) );
  \$mux  #( .WIDTH(33) ) _42966_ ( .A(_23144_), .B(_26263_), .S(_05777_), .Y(_23145_) );
  \$mux  #( .WIDTH(32) ) _42968_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_stride_3), .B(0), .S(_set_flag_874), .Y(_23146_) );
  \$mux  #( .WIDTH(32) ) _42970_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_stride_2), .B(1), .S(_set_flag_874), .Y(_23147_) );
  \$mux  #( .WIDTH(32) ) _42972_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_stride_1), .B({ 23'h000000, cparam_max_pool_serial_9_act_offset_values_1[8:0] }), .S(_set_flag_874), .Y(_23148_) );
  \$mux  #( .WIDTH(32) ) _42974_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_stride_0), .B({ 27'h0000000, cparam_max_pool_serial_9_inc_out_laddr }), .S(_set_flag_874), .Y(_23149_) );
  \$mux  #( .WIDTH(33) ) _42976_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_3), .B(33'h000000001), .S(_set_flag_874), .Y(_23150_) );
  \$mux  #( .WIDTH(33) ) _42978_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_2), .B({ 28'h0000000, cparam_max_pool_serial_9_inc_out_laddr }), .S(_set_flag_874), .Y(_23151_) );
  \$mux  #( .WIDTH(33) ) _42980_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_1), .B(33'h000000002), .S(_set_flag_874), .Y(_23152_) );
  \$mux  #( .WIDTH(33) ) _42982_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_size_0), .B(33'h000000002), .S(_set_flag_874), .Y(_23153_) );
  \$mux  #( .WIDTH(32) ) _42984_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_3), .B(0), .S(_05776_), .Y(_23154_) );
  \$mux  #( .WIDTH(32) ) _42985_ ( .A(_23154_), .B(_22237_), .S(_05779_), .Y(_23155_) );
  \$mux  #( .WIDTH(32) ) _42986_ ( .A(_23155_), .B(0), .S(_05780_), .Y(_23156_) );
  \$mux  #( .WIDTH(32) ) _42988_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_2), .B(0), .S(_05776_), .Y(_23157_) );
  \$mux  #( .WIDTH(32) ) _42989_ ( .A(_23157_), .B(_22236_), .S(_05778_), .Y(_23158_) );
  \$mux  #( .WIDTH(32) ) _42990_ ( .A(_23158_), .B(0), .S(_05779_), .Y(_23159_) );
  \$mux  #( .WIDTH(32) ) _42992_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_1), .B(0), .S(_05776_), .Y(_23160_) );
  \$mux  #( .WIDTH(32) ) _42993_ ( .A(_23160_), .B(_22235_), .S(_05777_), .Y(_23161_) );
  \$mux  #( .WIDTH(32) ) _42994_ ( .A(_23161_), .B(0), .S(_05778_), .Y(_23162_) );
  \$mux  #( .WIDTH(32) ) _42996_ ( .A(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_0), .B(0), .S(_05776_), .Y(_23163_) );
  \$mux  #( .WIDTH(32) ) _42997_ ( .A(_22234_), .B(_23163_), .S(_05043_), .Y(_23164_) );
  \$mux  #( .WIDTH(32) ) _42998_ ( .A(_23164_), .B(0), .S(_05777_), .Y(_23165_) );
  \$mux  #( .WIDTH(4) ) _43000_ ( .A(__variable_wdata_759), .B(_stream_max_pool_serial_9_constant_2_next_constant_data), .S(_stream_max_pool_serial_9_start), .Y(_23166_) );
  \$mux  #( .WIDTH(3) ) _43002_ ( .A(__variable_wdata_757), .B(_stream_max_pool_serial_9_constant_0_next_constant_data), .S(_stream_max_pool_serial_9_start), .Y(_23167_) );
  \$mux  #( .WIDTH(1) ) _43004_ ( .A(1'h1), .B(1'h0), .S(_05045_), .Y(_23124_) );
  \$mux  #( .WIDTH(4) ) _43016_ ( .A(_26630_[3:0]), .B(4'h0), .S(_stream_max_pool_serial_9_reduce_reset), .Y(_23168_) );
  \$mux  #( .WIDTH(32) ) _43018_ ( .A(_22231_), .B(0), .S(_stream_max_pool_serial_9_reduce_reset), .Y(_23169_) );
  \$mux  #( .WIDTH(32) ) _43019_ ( .A(0), .B(_23169_), .S(_04893_), .Y(_23170_) );
  \$mux  #( .WIDTH(32) ) _43020_ ( .A(_23170_), .B(-1), .S(RST), .Y(_01468_) );
  \$mux  #( .WIDTH(8) ) _43021_ ( .A(_stream_max_pool_serial_9_sink_3_sink_wdata), .B(__substreamoutput_data_773[7:0]), .S(_05782_), .Y(_23171_) );
  \$mux  #( .WIDTH(1) ) _43023_ ( .A(1'h0), .B(1'h1), .S(_05782_), .Y(_23172_) );
  \$mux  #( .WIDTH(32) ) _43025_ ( .A(_stream_max_pool_serial_9_sink_3_sink_waddr), .B(_26270_), .S(_05781_), .Y(_23173_) );
  \$mux  #( .WIDTH(32) ) _43026_ ( .A(_23173_), .B(_22239_), .S(_05782_), .Y(_23174_) );
  \$mux  #( .WIDTH(8) ) _43028_ ( .A(_stream_max_pool_serial_9_sink_3_sink_ram_sel), .B(8'h02), .S(__set_flag_874_9), .Y(_23175_) );
  \$mux  #( .WIDTH(32) ) _43030_ ( .A(_stream_max_pool_serial_9_sink_3_sink_stride_buf), .B(_stream_max_pool_serial_9_sink_3_sink_stride), .S(_05781_), .Y(_23176_) );
  \$mux  #( .WIDTH(33) ) _43032_ ( .A(_stream_max_pool_serial_9_sink_3_sink_count), .B(_stream_max_pool_serial_9_sink_3_sink_size), .S(_05781_), .Y(_23177_) );
  \$mux  #( .WIDTH(33) ) _43033_ ( .A(_23177_), .B(_26271_), .S(_05782_), .Y(_23178_) );
  \$mux  #( .WIDTH(32) ) _43035_ ( .A(_stream_max_pool_serial_9_sink_3_sink_stride), .B(1), .S(__set_flag_874_9), .Y(_23179_) );
  \$mux  #( .WIDTH(33) ) _43037_ ( .A(_stream_max_pool_serial_9_sink_3_sink_size), .B(__stream_max_pool_serial_9_sink_3_sink_size_1_9), .S(__set_flag_874_9), .Y(_23180_) );
  \$mux  #( .WIDTH(32) ) _43039_ ( .A(_stream_max_pool_serial_9_sink_3_sink_offset), .B(__stream_max_pool_serial_9_sink_3_sink_offset_0_9), .S(__set_flag_874_9), .Y(_23181_) );
  \$mux  #( .WIDTH(3) ) _43041_ ( .A(_stream_max_pool_serial_9_sink_3_sink_mode), .B(3'h1), .S(__set_flag_874_9), .Y(_23182_) );
  \$mux  #( .WIDTH(4) ) _43043_ ( .A(_stream_max_pool_serial_9_constant_2_next_constant_data), .B(max_pool_serial_9_stream_pad_masks), .S(_set_flag_874), .Y(_23183_) );
  \$mux  #( .WIDTH(1) ) _43045_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id1_3_cond_5_1), .Y(_23184_) );
  \$mux  #( .WIDTH(1) ) _43047_ ( .A(1'h1), .B(_stream_max_pool_serial_9_source_1_source_ram_renable), .S(_05043_), .Y(_23185_) );
  \$mux  #( .WIDTH(1) ) _43048_ ( .A(1'h0), .B(_23185_), .S(_05044_), .Y(_23186_) );
  \$mux  #( .WIDTH(32) ) _43050_ ( .A(_stream_max_pool_serial_9_source_1_source_pat_all_offset), .B(_stream_max_pool_serial_9_source_1_source_ram_raddr), .S(_05043_), .Y(_23187_) );
  \$mux  #( .WIDTH(8) ) _43052_ ( .A(_stream_max_pool_serial_9_source_1_source_ram_sel), .B(8'h01), .S(_set_flag_874), .Y(_23188_) );
  \$mux  #( .WIDTH(32) ) _43054_ ( .A(_stream_max_pool_serial_9_source_1_source_offset_buf), .B(_stream_max_pool_serial_9_source_1_source_offset), .S(_05776_), .Y(_23189_) );
  \$mux  #( .WIDTH(32) ) _43056_ ( .A(_stream_max_pool_serial_9_source_1_source_offset), .B(_22233_), .S(_set_flag_874), .Y(_23190_) );
  \$mux  #( .WIDTH(3) ) _43058_ ( .A(_stream_max_pool_serial_9_source_1_source_mode), .B(3'h2), .S(_set_flag_874), .Y(_23191_) );
  \$mux  #( .WIDTH(1) ) _43060_ ( .A(_stream_max_pool_serial_9_source_1_idle), .B(1'h0), .S(_05776_), .Y(_23192_) );
  \$mux  #( .WIDTH(1) ) _43061_ ( .A(1'h1), .B(_23192_), .S(_05044_), .Y(_23193_) );
  \$mux  #( .WIDTH(1) ) _43062_ ( .A(_23193_), .B(1'h1), .S(RST), .Y(_02659_) );
  \$mux  #( .WIDTH(3) ) _43063_ ( .A(_stream_max_pool_serial_9_constant_0_next_constant_data), .B(3'h4), .S(_set_flag_874), .Y(_23194_) );
  \$mux  #( .WIDTH(1) ) _43065_ ( .A(_stream_conv2d_8_source_busy), .B(1'h1), .S(_stream_conv2d_8_start_flag), .Y(_21584_) );
  \$mux  #( .WIDTH(1) ) _43067_ ( .A(1'h0), .B(1'h1), .S(__tmp_797_42), .Y(_23196_) );
  \$mux  #( .WIDTH(1) ) _43069_ ( .A(1'h0), .B(1'h1), .S(__tmp_795_46), .Y(_23197_) );
  \$mux  #( .WIDTH(1) ) _43071_ ( .A(1'h0), .B(1'h1), .S(_stream_conv2d_8_start_flag), .Y(_23198_) );
  \$mux  #( .WIDTH(1) ) _43072_ ( .A(_23198_), .B(1'h0), .S(_04903_), .Y(_23199_) );
  \$mux  #( .WIDTH(32) ) _43074_ ( .A(_stream_conv2d_8_fsm), .B(3), .S(_stream_conv2d_8_done), .Y({ _21641_, _21640_, _21638_, _21637_, _21636_, _21635_, _21634_, _21633_, _21632_, _21631_, _21630_, _21629_, _21627_, _21626_, _21625_, _21624_, _21623_, _21622_, _21621_, _21620_, _21619_, _21618_, _21648_, _21647_, _21646_, _21645_, _21644_, _21643_, _21642_, _21639_, _21628_, _21617_ }) );
  \$mux  #( .WIDTH(32) ) _43075_ ( .A(_stream_conv2d_8_fsm), .B(1), .S(_stream_conv2d_8_start_flag), .Y({ _21673_, _21672_, _21670_, _21669_, _21668_, _21667_, _21666_, _21665_, _21664_, _21663_, _21662_, _21661_, _21659_, _21658_, _21657_, _21656_, _21655_, _21654_, _21653_, _21652_, _21651_, _21650_, _21680_, _21679_, _21678_, _21677_, _21676_, _21675_, _21674_, _21671_, _21660_, _21649_ }) );
  \$mux  #( .WIDTH(8) ) _43326_ ( .A(__variable_wdata_490), .B(_stream_conv2d_8_source_36_source_ram_rdata), .S(_stream_conv2d_8_source_36_source_ram_rvalid), .Y(_23202_) );
  \$mux  #( .WIDTH(32) ) _43328_ ( .A(_source_stream_conv2d_8_source_36_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_36_pat_stride_3), .S(_05769_), .Y(_23203_) );
  \$mux  #( .WIDTH(32) ) _43330_ ( .A(_source_stream_conv2d_8_source_36_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_36_pat_stride_2), .S(_05769_), .Y(_23204_) );
  \$mux  #( .WIDTH(32) ) _43332_ ( .A(_source_stream_conv2d_8_source_36_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_36_pat_stride_1), .S(_05769_), .Y(_23205_) );
  \$mux  #( .WIDTH(32) ) _43334_ ( .A(_source_stream_conv2d_8_source_36_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_36_pat_stride_0), .S(_05769_), .Y(_23206_) );
  \$mux  #( .WIDTH(33) ) _43336_ ( .A(_source_stream_conv2d_8_source_36_pat_size_buf_3), .B(_source_stream_conv2d_8_source_36_pat_size_3), .S(_05769_), .Y(_23207_) );
  \$mux  #( .WIDTH(33) ) _43338_ ( .A(_source_stream_conv2d_8_source_36_pat_size_buf_2), .B(_source_stream_conv2d_8_source_36_pat_size_2), .S(_05769_), .Y(_23208_) );
  \$mux  #( .WIDTH(33) ) _43340_ ( .A(_source_stream_conv2d_8_source_36_pat_size_buf_1), .B(_source_stream_conv2d_8_source_36_pat_size_1), .S(_05769_), .Y(_23209_) );
  \$mux  #( .WIDTH(33) ) _43342_ ( .A(_source_stream_conv2d_8_source_36_pat_size_buf_0), .B(_source_stream_conv2d_8_source_36_pat_size_0), .S(_05769_), .Y(_23210_) );
  \$mux  #( .WIDTH(33) ) _43344_ ( .A(_source_stream_conv2d_8_source_36_pat_count_3), .B(_26247_), .S(_05769_), .Y(_23211_) );
  \$mux  #( .WIDTH(33) ) _43345_ ( .A(_23211_), .B(_26254_), .S(_05772_), .Y(_23212_) );
  \$mux  #( .WIDTH(33) ) _43346_ ( .A(_23212_), .B(_26255_), .S(_05773_), .Y(_23213_) );
  \$mux  #( .WIDTH(33) ) _43348_ ( .A(_source_stream_conv2d_8_source_36_pat_count_2), .B(_26246_), .S(_05769_), .Y(_23214_) );
  \$mux  #( .WIDTH(33) ) _43349_ ( .A(_23214_), .B(_26252_), .S(_05771_), .Y(_23215_) );
  \$mux  #( .WIDTH(33) ) _43350_ ( .A(_23215_), .B(_26253_), .S(_05772_), .Y(_23216_) );
  \$mux  #( .WIDTH(33) ) _43352_ ( .A(_source_stream_conv2d_8_source_36_pat_count_1), .B(_26245_), .S(_05769_), .Y(_23217_) );
  \$mux  #( .WIDTH(33) ) _43353_ ( .A(_23217_), .B(_26250_), .S(_05770_), .Y(_23218_) );
  \$mux  #( .WIDTH(33) ) _43354_ ( .A(_23218_), .B(_26251_), .S(_05771_), .Y(_23219_) );
  \$mux  #( .WIDTH(33) ) _43356_ ( .A(_source_stream_conv2d_8_source_36_pat_count_0), .B(_26244_), .S(_05769_), .Y(_23220_) );
  \$mux  #( .WIDTH(33) ) _43357_ ( .A(_26248_), .B(_23220_), .S(_05061_), .Y(_23221_) );
  \$mux  #( .WIDTH(33) ) _43358_ ( .A(_23221_), .B(_26249_), .S(_05770_), .Y(_23222_) );
  \$mux  #( .WIDTH(32) ) _43360_ ( .A(_source_stream_conv2d_8_source_36_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23223_) );
  \$mux  #( .WIDTH(32) ) _43362_ ( .A(_source_stream_conv2d_8_source_36_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23224_) );
  \$mux  #( .WIDTH(32) ) _43364_ ( .A(_source_stream_conv2d_8_source_36_pat_stride_1), .B({ 27'h0000000, cparam_conv2d_8_inc_act_laddr_large }), .S(_set_flag_538), .Y(_23225_) );
  \$mux  #( .WIDTH(32) ) _43366_ ( .A(_source_stream_conv2d_8_source_36_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23226_) );
  \$mux  #( .WIDTH(33) ) _43368_ ( .A(_source_stream_conv2d_8_source_36_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23227_) );
  \$mux  #( .WIDTH(33) ) _43370_ ( .A(_source_stream_conv2d_8_source_36_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23228_) );
  \$mux  #( .WIDTH(33) ) _43372_ ( .A(_source_stream_conv2d_8_source_36_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23229_) );
  \$mux  #( .WIDTH(33) ) _43374_ ( .A(_source_stream_conv2d_8_source_36_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23230_) );
  \$mux  #( .WIDTH(32) ) _43376_ ( .A(_source_stream_conv2d_8_source_36_pat_cur_offset_3), .B(0), .S(_05769_), .Y(_23231_) );
  \$mux  #( .WIDTH(32) ) _43377_ ( .A(_23231_), .B(_22228_), .S(_05772_), .Y(_23232_) );
  \$mux  #( .WIDTH(32) ) _43378_ ( .A(_23232_), .B(0), .S(_05773_), .Y(_23233_) );
  \$mux  #( .WIDTH(32) ) _43380_ ( .A(_source_stream_conv2d_8_source_36_pat_cur_offset_2), .B(0), .S(_05769_), .Y(_23234_) );
  \$mux  #( .WIDTH(32) ) _43381_ ( .A(_23234_), .B(_22227_), .S(_05771_), .Y(_23235_) );
  \$mux  #( .WIDTH(32) ) _43382_ ( .A(_23235_), .B(0), .S(_05772_), .Y(_23236_) );
  \$mux  #( .WIDTH(32) ) _43384_ ( .A(_source_stream_conv2d_8_source_36_pat_cur_offset_1), .B(0), .S(_05769_), .Y(_23237_) );
  \$mux  #( .WIDTH(32) ) _43385_ ( .A(_23237_), .B(_22226_), .S(_05770_), .Y(_23238_) );
  \$mux  #( .WIDTH(32) ) _43386_ ( .A(_23238_), .B(0), .S(_05771_), .Y(_23239_) );
  \$mux  #( .WIDTH(32) ) _43388_ ( .A(_source_stream_conv2d_8_source_36_pat_cur_offset_0), .B(0), .S(_05769_), .Y(_23240_) );
  \$mux  #( .WIDTH(32) ) _43389_ ( .A(_22225_), .B(_23240_), .S(_05061_), .Y(_23241_) );
  \$mux  #( .WIDTH(32) ) _43390_ ( .A(_23241_), .B(0), .S(_05770_), .Y(_23242_) );
  \$mux  #( .WIDTH(8) ) _43392_ ( .A(__variable_wdata_489), .B(_stream_conv2d_8_source_35_source_ram_rdata), .S(_stream_conv2d_8_source_35_source_ram_rvalid), .Y(_23243_) );
  \$mux  #( .WIDTH(32) ) _43394_ ( .A(_source_stream_conv2d_8_source_35_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_35_pat_stride_3), .S(_05764_), .Y(_23244_) );
  \$mux  #( .WIDTH(32) ) _43396_ ( .A(_source_stream_conv2d_8_source_35_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_35_pat_stride_2), .S(_05764_), .Y(_23245_) );
  \$mux  #( .WIDTH(32) ) _43398_ ( .A(_source_stream_conv2d_8_source_35_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_35_pat_stride_1), .S(_05764_), .Y(_23246_) );
  \$mux  #( .WIDTH(32) ) _43400_ ( .A(_source_stream_conv2d_8_source_35_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_35_pat_stride_0), .S(_05764_), .Y(_23247_) );
  \$mux  #( .WIDTH(33) ) _43402_ ( .A(_source_stream_conv2d_8_source_35_pat_size_buf_3), .B(_source_stream_conv2d_8_source_35_pat_size_3), .S(_05764_), .Y(_23248_) );
  \$mux  #( .WIDTH(33) ) _43404_ ( .A(_source_stream_conv2d_8_source_35_pat_size_buf_2), .B(_source_stream_conv2d_8_source_35_pat_size_2), .S(_05764_), .Y(_23249_) );
  \$mux  #( .WIDTH(33) ) _43406_ ( .A(_source_stream_conv2d_8_source_35_pat_size_buf_1), .B(_source_stream_conv2d_8_source_35_pat_size_1), .S(_05764_), .Y(_23250_) );
  \$mux  #( .WIDTH(33) ) _43408_ ( .A(_source_stream_conv2d_8_source_35_pat_size_buf_0), .B(_source_stream_conv2d_8_source_35_pat_size_0), .S(_05764_), .Y(_23251_) );
  \$mux  #( .WIDTH(33) ) _43410_ ( .A(_source_stream_conv2d_8_source_35_pat_count_3), .B(_26235_), .S(_05764_), .Y(_23252_) );
  \$mux  #( .WIDTH(33) ) _43411_ ( .A(_23252_), .B(_26242_), .S(_05767_), .Y(_23253_) );
  \$mux  #( .WIDTH(33) ) _43412_ ( .A(_23253_), .B(_26243_), .S(_05768_), .Y(_23254_) );
  \$mux  #( .WIDTH(33) ) _43414_ ( .A(_source_stream_conv2d_8_source_35_pat_count_2), .B(_26234_), .S(_05764_), .Y(_23255_) );
  \$mux  #( .WIDTH(33) ) _43415_ ( .A(_23255_), .B(_26240_), .S(_05766_), .Y(_23256_) );
  \$mux  #( .WIDTH(33) ) _43416_ ( .A(_23256_), .B(_26241_), .S(_05767_), .Y(_23257_) );
  \$mux  #( .WIDTH(33) ) _43418_ ( .A(_source_stream_conv2d_8_source_35_pat_count_1), .B(_26233_), .S(_05764_), .Y(_23258_) );
  \$mux  #( .WIDTH(33) ) _43419_ ( .A(_23258_), .B(_26238_), .S(_05765_), .Y(_23259_) );
  \$mux  #( .WIDTH(33) ) _43420_ ( .A(_23259_), .B(_26239_), .S(_05766_), .Y(_23260_) );
  \$mux  #( .WIDTH(33) ) _43422_ ( .A(_source_stream_conv2d_8_source_35_pat_count_0), .B(_26232_), .S(_05764_), .Y(_23261_) );
  \$mux  #( .WIDTH(33) ) _43423_ ( .A(_26236_), .B(_23261_), .S(_05064_), .Y(_23262_) );
  \$mux  #( .WIDTH(33) ) _43424_ ( .A(_23262_), .B(_26237_), .S(_05765_), .Y(_23263_) );
  \$mux  #( .WIDTH(32) ) _43426_ ( .A(_source_stream_conv2d_8_source_35_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23264_) );
  \$mux  #( .WIDTH(32) ) _43428_ ( .A(_source_stream_conv2d_8_source_35_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23265_) );
  \$mux  #( .WIDTH(32) ) _43430_ ( .A(_source_stream_conv2d_8_source_35_pat_stride_1), .B({ 27'h0000000, cparam_conv2d_8_inc_act_laddr_large }), .S(_set_flag_538), .Y(_23266_) );
  \$mux  #( .WIDTH(32) ) _43432_ ( .A(_source_stream_conv2d_8_source_35_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23267_) );
  \$mux  #( .WIDTH(33) ) _43434_ ( .A(_source_stream_conv2d_8_source_35_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23268_) );
  \$mux  #( .WIDTH(33) ) _43436_ ( .A(_source_stream_conv2d_8_source_35_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23269_) );
  \$mux  #( .WIDTH(33) ) _43438_ ( .A(_source_stream_conv2d_8_source_35_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23270_) );
  \$mux  #( .WIDTH(33) ) _43440_ ( .A(_source_stream_conv2d_8_source_35_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23271_) );
  \$mux  #( .WIDTH(32) ) _43442_ ( .A(_source_stream_conv2d_8_source_35_pat_cur_offset_3), .B(0), .S(_05764_), .Y(_23272_) );
  \$mux  #( .WIDTH(32) ) _43443_ ( .A(_23272_), .B(_22224_), .S(_05767_), .Y(_23273_) );
  \$mux  #( .WIDTH(32) ) _43444_ ( .A(_23273_), .B(0), .S(_05768_), .Y(_23274_) );
  \$mux  #( .WIDTH(32) ) _43446_ ( .A(_source_stream_conv2d_8_source_35_pat_cur_offset_2), .B(0), .S(_05764_), .Y(_23275_) );
  \$mux  #( .WIDTH(32) ) _43447_ ( .A(_23275_), .B(_22223_), .S(_05766_), .Y(_23276_) );
  \$mux  #( .WIDTH(32) ) _43448_ ( .A(_23276_), .B(0), .S(_05767_), .Y(_23277_) );
  \$mux  #( .WIDTH(32) ) _43450_ ( .A(_source_stream_conv2d_8_source_35_pat_cur_offset_1), .B(0), .S(_05764_), .Y(_23278_) );
  \$mux  #( .WIDTH(32) ) _43451_ ( .A(_23278_), .B(_22222_), .S(_05765_), .Y(_23279_) );
  \$mux  #( .WIDTH(32) ) _43452_ ( .A(_23279_), .B(0), .S(_05766_), .Y(_23280_) );
  \$mux  #( .WIDTH(32) ) _43454_ ( .A(_source_stream_conv2d_8_source_35_pat_cur_offset_0), .B(0), .S(_05764_), .Y(_23281_) );
  \$mux  #( .WIDTH(32) ) _43455_ ( .A(_22221_), .B(_23281_), .S(_05064_), .Y(_23282_) );
  \$mux  #( .WIDTH(32) ) _43456_ ( .A(_23282_), .B(0), .S(_05765_), .Y(_23283_) );
  \$mux  #( .WIDTH(8) ) _43458_ ( .A(__variable_wdata_488), .B(_stream_conv2d_8_source_34_source_ram_rdata), .S(_stream_conv2d_8_source_34_source_ram_rvalid), .Y(_23284_) );
  \$mux  #( .WIDTH(32) ) _43460_ ( .A(_source_stream_conv2d_8_source_34_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_34_pat_stride_3), .S(_05759_), .Y(_23285_) );
  \$mux  #( .WIDTH(32) ) _43462_ ( .A(_source_stream_conv2d_8_source_34_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_34_pat_stride_2), .S(_05759_), .Y(_23286_) );
  \$mux  #( .WIDTH(32) ) _43464_ ( .A(_source_stream_conv2d_8_source_34_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_34_pat_stride_1), .S(_05759_), .Y(_23287_) );
  \$mux  #( .WIDTH(32) ) _43466_ ( .A(_source_stream_conv2d_8_source_34_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_34_pat_stride_0), .S(_05759_), .Y(_23288_) );
  \$mux  #( .WIDTH(33) ) _43468_ ( .A(_source_stream_conv2d_8_source_34_pat_size_buf_3), .B(_source_stream_conv2d_8_source_34_pat_size_3), .S(_05759_), .Y(_23289_) );
  \$mux  #( .WIDTH(33) ) _43470_ ( .A(_source_stream_conv2d_8_source_34_pat_size_buf_2), .B(_source_stream_conv2d_8_source_34_pat_size_2), .S(_05759_), .Y(_23290_) );
  \$mux  #( .WIDTH(33) ) _43472_ ( .A(_source_stream_conv2d_8_source_34_pat_size_buf_1), .B(_source_stream_conv2d_8_source_34_pat_size_1), .S(_05759_), .Y(_23291_) );
  \$mux  #( .WIDTH(33) ) _43474_ ( .A(_source_stream_conv2d_8_source_34_pat_size_buf_0), .B(_source_stream_conv2d_8_source_34_pat_size_0), .S(_05759_), .Y(_23292_) );
  \$mux  #( .WIDTH(33) ) _43476_ ( .A(_source_stream_conv2d_8_source_34_pat_count_3), .B(_26223_), .S(_05759_), .Y(_23293_) );
  \$mux  #( .WIDTH(33) ) _43477_ ( .A(_23293_), .B(_26230_), .S(_05762_), .Y(_23294_) );
  \$mux  #( .WIDTH(33) ) _43478_ ( .A(_23294_), .B(_26231_), .S(_05763_), .Y(_23295_) );
  \$mux  #( .WIDTH(33) ) _43480_ ( .A(_source_stream_conv2d_8_source_34_pat_count_2), .B(_26222_), .S(_05759_), .Y(_23296_) );
  \$mux  #( .WIDTH(33) ) _43481_ ( .A(_23296_), .B(_26228_), .S(_05761_), .Y(_23297_) );
  \$mux  #( .WIDTH(33) ) _43482_ ( .A(_23297_), .B(_26229_), .S(_05762_), .Y(_23298_) );
  \$mux  #( .WIDTH(33) ) _43484_ ( .A(_source_stream_conv2d_8_source_34_pat_count_1), .B(_26221_), .S(_05759_), .Y(_23299_) );
  \$mux  #( .WIDTH(33) ) _43485_ ( .A(_23299_), .B(_26226_), .S(_05760_), .Y(_23300_) );
  \$mux  #( .WIDTH(33) ) _43486_ ( .A(_23300_), .B(_26227_), .S(_05761_), .Y(_23301_) );
  \$mux  #( .WIDTH(33) ) _43488_ ( .A(_source_stream_conv2d_8_source_34_pat_count_0), .B(_26220_), .S(_05759_), .Y(_23302_) );
  \$mux  #( .WIDTH(33) ) _43489_ ( .A(_26224_), .B(_23302_), .S(_05066_), .Y(_23303_) );
  \$mux  #( .WIDTH(33) ) _43490_ ( .A(_23303_), .B(_26225_), .S(_05760_), .Y(_23304_) );
  \$mux  #( .WIDTH(32) ) _43492_ ( .A(_source_stream_conv2d_8_source_34_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23305_) );
  \$mux  #( .WIDTH(32) ) _43494_ ( .A(_source_stream_conv2d_8_source_34_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23306_) );
  \$mux  #( .WIDTH(32) ) _43496_ ( .A(_source_stream_conv2d_8_source_34_pat_stride_1), .B({ 27'h0000000, cparam_conv2d_8_inc_act_laddr_large }), .S(_set_flag_538), .Y(_23307_) );
  \$mux  #( .WIDTH(32) ) _43498_ ( .A(_source_stream_conv2d_8_source_34_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23308_) );
  \$mux  #( .WIDTH(33) ) _43500_ ( .A(_source_stream_conv2d_8_source_34_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23309_) );
  \$mux  #( .WIDTH(33) ) _43502_ ( .A(_source_stream_conv2d_8_source_34_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23310_) );
  \$mux  #( .WIDTH(33) ) _43504_ ( .A(_source_stream_conv2d_8_source_34_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23311_) );
  \$mux  #( .WIDTH(33) ) _43506_ ( .A(_source_stream_conv2d_8_source_34_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23312_) );
  \$mux  #( .WIDTH(32) ) _43508_ ( .A(_source_stream_conv2d_8_source_34_pat_cur_offset_3), .B(0), .S(_05759_), .Y(_23313_) );
  \$mux  #( .WIDTH(32) ) _43509_ ( .A(_23313_), .B(_22220_), .S(_05762_), .Y(_23314_) );
  \$mux  #( .WIDTH(32) ) _43510_ ( .A(_23314_), .B(0), .S(_05763_), .Y(_23315_) );
  \$mux  #( .WIDTH(32) ) _43512_ ( .A(_source_stream_conv2d_8_source_34_pat_cur_offset_2), .B(0), .S(_05759_), .Y(_23316_) );
  \$mux  #( .WIDTH(32) ) _43513_ ( .A(_23316_), .B(_22219_), .S(_05761_), .Y(_23317_) );
  \$mux  #( .WIDTH(32) ) _43514_ ( .A(_23317_), .B(0), .S(_05762_), .Y(_23318_) );
  \$mux  #( .WIDTH(32) ) _43516_ ( .A(_source_stream_conv2d_8_source_34_pat_cur_offset_1), .B(0), .S(_05759_), .Y(_23319_) );
  \$mux  #( .WIDTH(32) ) _43517_ ( .A(_23319_), .B(_22218_), .S(_05760_), .Y(_23320_) );
  \$mux  #( .WIDTH(32) ) _43518_ ( .A(_23320_), .B(0), .S(_05761_), .Y(_23321_) );
  \$mux  #( .WIDTH(32) ) _43520_ ( .A(_source_stream_conv2d_8_source_34_pat_cur_offset_0), .B(0), .S(_05759_), .Y(_23322_) );
  \$mux  #( .WIDTH(32) ) _43521_ ( .A(_22217_), .B(_23322_), .S(_05066_), .Y(_23323_) );
  \$mux  #( .WIDTH(32) ) _43522_ ( .A(_23323_), .B(0), .S(_05760_), .Y(_23324_) );
  \$mux  #( .WIDTH(8) ) _43524_ ( .A(__variable_wdata_487), .B(_stream_conv2d_8_source_33_source_ram_rdata), .S(_stream_conv2d_8_source_33_source_ram_rvalid), .Y(_23325_) );
  \$mux  #( .WIDTH(32) ) _43526_ ( .A(_source_stream_conv2d_8_source_33_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_33_pat_stride_3), .S(_05754_), .Y(_23326_) );
  \$mux  #( .WIDTH(32) ) _43528_ ( .A(_source_stream_conv2d_8_source_33_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_33_pat_stride_2), .S(_05754_), .Y(_23327_) );
  \$mux  #( .WIDTH(32) ) _43530_ ( .A(_source_stream_conv2d_8_source_33_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_33_pat_stride_1), .S(_05754_), .Y(_23328_) );
  \$mux  #( .WIDTH(32) ) _43532_ ( .A(_source_stream_conv2d_8_source_33_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_33_pat_stride_0), .S(_05754_), .Y(_23329_) );
  \$mux  #( .WIDTH(33) ) _43534_ ( .A(_source_stream_conv2d_8_source_33_pat_size_buf_3), .B(_source_stream_conv2d_8_source_33_pat_size_3), .S(_05754_), .Y(_23330_) );
  \$mux  #( .WIDTH(33) ) _43536_ ( .A(_source_stream_conv2d_8_source_33_pat_size_buf_2), .B(_source_stream_conv2d_8_source_33_pat_size_2), .S(_05754_), .Y(_23331_) );
  \$mux  #( .WIDTH(33) ) _43538_ ( .A(_source_stream_conv2d_8_source_33_pat_size_buf_1), .B(_source_stream_conv2d_8_source_33_pat_size_1), .S(_05754_), .Y(_23332_) );
  \$mux  #( .WIDTH(33) ) _43540_ ( .A(_source_stream_conv2d_8_source_33_pat_size_buf_0), .B(_source_stream_conv2d_8_source_33_pat_size_0), .S(_05754_), .Y(_23333_) );
  \$mux  #( .WIDTH(33) ) _43542_ ( .A(_source_stream_conv2d_8_source_33_pat_count_3), .B(_26211_), .S(_05754_), .Y(_23334_) );
  \$mux  #( .WIDTH(33) ) _43543_ ( .A(_23334_), .B(_26218_), .S(_05757_), .Y(_23335_) );
  \$mux  #( .WIDTH(33) ) _43544_ ( .A(_23335_), .B(_26219_), .S(_05758_), .Y(_23336_) );
  \$mux  #( .WIDTH(33) ) _43546_ ( .A(_source_stream_conv2d_8_source_33_pat_count_2), .B(_26210_), .S(_05754_), .Y(_23337_) );
  \$mux  #( .WIDTH(33) ) _43547_ ( .A(_23337_), .B(_26216_), .S(_05756_), .Y(_23338_) );
  \$mux  #( .WIDTH(33) ) _43548_ ( .A(_23338_), .B(_26217_), .S(_05757_), .Y(_23339_) );
  \$mux  #( .WIDTH(33) ) _43550_ ( .A(_source_stream_conv2d_8_source_33_pat_count_1), .B(_26209_), .S(_05754_), .Y(_23340_) );
  \$mux  #( .WIDTH(33) ) _43551_ ( .A(_23340_), .B(_26214_), .S(_05755_), .Y(_23341_) );
  \$mux  #( .WIDTH(33) ) _43552_ ( .A(_23341_), .B(_26215_), .S(_05756_), .Y(_23342_) );
  \$mux  #( .WIDTH(33) ) _43554_ ( .A(_source_stream_conv2d_8_source_33_pat_count_0), .B(_26208_), .S(_05754_), .Y(_23343_) );
  \$mux  #( .WIDTH(33) ) _43555_ ( .A(_26212_), .B(_23343_), .S(_05067_), .Y(_23344_) );
  \$mux  #( .WIDTH(33) ) _43556_ ( .A(_23344_), .B(_26213_), .S(_05755_), .Y(_23345_) );
  \$mux  #( .WIDTH(32) ) _43558_ ( .A(_source_stream_conv2d_8_source_33_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23346_) );
  \$mux  #( .WIDTH(32) ) _43560_ ( .A(_source_stream_conv2d_8_source_33_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23347_) );
  \$mux  #( .WIDTH(32) ) _43562_ ( .A(_source_stream_conv2d_8_source_33_pat_stride_1), .B({ 27'h0000000, cparam_conv2d_8_inc_act_laddr_large }), .S(_set_flag_538), .Y(_23348_) );
  \$mux  #( .WIDTH(32) ) _43564_ ( .A(_source_stream_conv2d_8_source_33_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23349_) );
  \$mux  #( .WIDTH(33) ) _43566_ ( .A(_source_stream_conv2d_8_source_33_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23350_) );
  \$mux  #( .WIDTH(33) ) _43568_ ( .A(_source_stream_conv2d_8_source_33_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23351_) );
  \$mux  #( .WIDTH(33) ) _43570_ ( .A(_source_stream_conv2d_8_source_33_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23352_) );
  \$mux  #( .WIDTH(33) ) _43572_ ( .A(_source_stream_conv2d_8_source_33_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23353_) );
  \$mux  #( .WIDTH(32) ) _43574_ ( .A(_source_stream_conv2d_8_source_33_pat_cur_offset_3), .B(0), .S(_05754_), .Y(_23354_) );
  \$mux  #( .WIDTH(32) ) _43575_ ( .A(_23354_), .B(_22216_), .S(_05757_), .Y(_23355_) );
  \$mux  #( .WIDTH(32) ) _43576_ ( .A(_23355_), .B(0), .S(_05758_), .Y(_23356_) );
  \$mux  #( .WIDTH(32) ) _43578_ ( .A(_source_stream_conv2d_8_source_33_pat_cur_offset_2), .B(0), .S(_05754_), .Y(_23357_) );
  \$mux  #( .WIDTH(32) ) _43579_ ( .A(_23357_), .B(_22215_), .S(_05756_), .Y(_23358_) );
  \$mux  #( .WIDTH(32) ) _43580_ ( .A(_23358_), .B(0), .S(_05757_), .Y(_23359_) );
  \$mux  #( .WIDTH(32) ) _43582_ ( .A(_source_stream_conv2d_8_source_33_pat_cur_offset_1), .B(0), .S(_05754_), .Y(_23360_) );
  \$mux  #( .WIDTH(32) ) _43583_ ( .A(_23360_), .B(_22214_), .S(_05755_), .Y(_23361_) );
  \$mux  #( .WIDTH(32) ) _43584_ ( .A(_23361_), .B(0), .S(_05756_), .Y(_23362_) );
  \$mux  #( .WIDTH(32) ) _43586_ ( .A(_source_stream_conv2d_8_source_33_pat_cur_offset_0), .B(0), .S(_05754_), .Y(_23363_) );
  \$mux  #( .WIDTH(32) ) _43587_ ( .A(_22213_), .B(_23363_), .S(_05067_), .Y(_23364_) );
  \$mux  #( .WIDTH(32) ) _43588_ ( .A(_23364_), .B(0), .S(_05755_), .Y(_23365_) );
  \$mux  #( .WIDTH(8) ) _43590_ ( .A(__variable_wdata_486), .B(_stream_conv2d_8_source_32_source_ram_rdata), .S(_stream_conv2d_8_source_32_source_ram_rvalid), .Y(_23366_) );
  \$mux  #( .WIDTH(32) ) _43592_ ( .A(_source_stream_conv2d_8_source_32_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_32_pat_stride_3), .S(_05749_), .Y(_23367_) );
  \$mux  #( .WIDTH(32) ) _43594_ ( .A(_source_stream_conv2d_8_source_32_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_32_pat_stride_2), .S(_05749_), .Y(_23368_) );
  \$mux  #( .WIDTH(32) ) _43596_ ( .A(_source_stream_conv2d_8_source_32_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_32_pat_stride_1), .S(_05749_), .Y(_23369_) );
  \$mux  #( .WIDTH(32) ) _43598_ ( .A(_source_stream_conv2d_8_source_32_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_32_pat_stride_0), .S(_05749_), .Y(_23370_) );
  \$mux  #( .WIDTH(33) ) _43600_ ( .A(_source_stream_conv2d_8_source_32_pat_size_buf_3), .B(_source_stream_conv2d_8_source_32_pat_size_3), .S(_05749_), .Y(_23371_) );
  \$mux  #( .WIDTH(33) ) _43602_ ( .A(_source_stream_conv2d_8_source_32_pat_size_buf_2), .B(_source_stream_conv2d_8_source_32_pat_size_2), .S(_05749_), .Y(_23372_) );
  \$mux  #( .WIDTH(33) ) _43604_ ( .A(_source_stream_conv2d_8_source_32_pat_size_buf_1), .B(_source_stream_conv2d_8_source_32_pat_size_1), .S(_05749_), .Y(_23373_) );
  \$mux  #( .WIDTH(33) ) _43606_ ( .A(_source_stream_conv2d_8_source_32_pat_size_buf_0), .B(_source_stream_conv2d_8_source_32_pat_size_0), .S(_05749_), .Y(_23374_) );
  \$mux  #( .WIDTH(33) ) _43608_ ( .A(_source_stream_conv2d_8_source_32_pat_count_3), .B(_26199_), .S(_05749_), .Y(_23375_) );
  \$mux  #( .WIDTH(33) ) _43609_ ( .A(_23375_), .B(_26206_), .S(_05752_), .Y(_23376_) );
  \$mux  #( .WIDTH(33) ) _43610_ ( .A(_23376_), .B(_26207_), .S(_05753_), .Y(_23377_) );
  \$mux  #( .WIDTH(33) ) _43612_ ( .A(_source_stream_conv2d_8_source_32_pat_count_2), .B(_26198_), .S(_05749_), .Y(_23378_) );
  \$mux  #( .WIDTH(33) ) _43613_ ( .A(_23378_), .B(_26204_), .S(_05751_), .Y(_23379_) );
  \$mux  #( .WIDTH(33) ) _43614_ ( .A(_23379_), .B(_26205_), .S(_05752_), .Y(_23380_) );
  \$mux  #( .WIDTH(33) ) _43616_ ( .A(_source_stream_conv2d_8_source_32_pat_count_1), .B(_26197_), .S(_05749_), .Y(_23381_) );
  \$mux  #( .WIDTH(33) ) _43617_ ( .A(_23381_), .B(_26202_), .S(_05750_), .Y(_23382_) );
  \$mux  #( .WIDTH(33) ) _43618_ ( .A(_23382_), .B(_26203_), .S(_05751_), .Y(_23383_) );
  \$mux  #( .WIDTH(33) ) _43620_ ( .A(_source_stream_conv2d_8_source_32_pat_count_0), .B(_26196_), .S(_05749_), .Y(_23384_) );
  \$mux  #( .WIDTH(33) ) _43621_ ( .A(_26200_), .B(_23384_), .S(_05069_), .Y(_23385_) );
  \$mux  #( .WIDTH(33) ) _43622_ ( .A(_23385_), .B(_26201_), .S(_05750_), .Y(_23386_) );
  \$mux  #( .WIDTH(32) ) _43624_ ( .A(_source_stream_conv2d_8_source_32_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23387_) );
  \$mux  #( .WIDTH(32) ) _43626_ ( .A(_source_stream_conv2d_8_source_32_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23388_) );
  \$mux  #( .WIDTH(32) ) _43628_ ( .A(_source_stream_conv2d_8_source_32_pat_stride_1), .B({ 27'h0000000, cparam_conv2d_8_inc_act_laddr_large }), .S(_set_flag_538), .Y(_23389_) );
  \$mux  #( .WIDTH(32) ) _43630_ ( .A(_source_stream_conv2d_8_source_32_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23390_) );
  \$mux  #( .WIDTH(33) ) _43632_ ( .A(_source_stream_conv2d_8_source_32_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23391_) );
  \$mux  #( .WIDTH(33) ) _43634_ ( .A(_source_stream_conv2d_8_source_32_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23392_) );
  \$mux  #( .WIDTH(33) ) _43636_ ( .A(_source_stream_conv2d_8_source_32_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23393_) );
  \$mux  #( .WIDTH(33) ) _43638_ ( .A(_source_stream_conv2d_8_source_32_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23394_) );
  \$mux  #( .WIDTH(32) ) _43640_ ( .A(_source_stream_conv2d_8_source_32_pat_cur_offset_3), .B(0), .S(_05749_), .Y(_23395_) );
  \$mux  #( .WIDTH(32) ) _43641_ ( .A(_23395_), .B(_22212_), .S(_05752_), .Y(_23396_) );
  \$mux  #( .WIDTH(32) ) _43642_ ( .A(_23396_), .B(0), .S(_05753_), .Y(_23397_) );
  \$mux  #( .WIDTH(32) ) _43644_ ( .A(_source_stream_conv2d_8_source_32_pat_cur_offset_2), .B(0), .S(_05749_), .Y(_23398_) );
  \$mux  #( .WIDTH(32) ) _43645_ ( .A(_23398_), .B(_22211_), .S(_05751_), .Y(_23399_) );
  \$mux  #( .WIDTH(32) ) _43646_ ( .A(_23399_), .B(0), .S(_05752_), .Y(_23400_) );
  \$mux  #( .WIDTH(32) ) _43648_ ( .A(_source_stream_conv2d_8_source_32_pat_cur_offset_1), .B(0), .S(_05749_), .Y(_23401_) );
  \$mux  #( .WIDTH(32) ) _43649_ ( .A(_23401_), .B(_22210_), .S(_05750_), .Y(_23402_) );
  \$mux  #( .WIDTH(32) ) _43650_ ( .A(_23402_), .B(0), .S(_05751_), .Y(_23403_) );
  \$mux  #( .WIDTH(32) ) _43652_ ( .A(_source_stream_conv2d_8_source_32_pat_cur_offset_0), .B(0), .S(_05749_), .Y(_23404_) );
  \$mux  #( .WIDTH(32) ) _43653_ ( .A(_22209_), .B(_23404_), .S(_05069_), .Y(_23405_) );
  \$mux  #( .WIDTH(32) ) _43654_ ( .A(_23405_), .B(0), .S(_05750_), .Y(_23406_) );
  \$mux  #( .WIDTH(8) ) _43656_ ( .A(__variable_wdata_485), .B(_stream_conv2d_8_source_31_source_ram_rdata), .S(_stream_conv2d_8_source_31_source_ram_rvalid), .Y(_23407_) );
  \$mux  #( .WIDTH(32) ) _43658_ ( .A(_source_stream_conv2d_8_source_31_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_31_pat_stride_3), .S(_05744_), .Y(_23408_) );
  \$mux  #( .WIDTH(32) ) _43660_ ( .A(_source_stream_conv2d_8_source_31_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_31_pat_stride_2), .S(_05744_), .Y(_23409_) );
  \$mux  #( .WIDTH(32) ) _43662_ ( .A(_source_stream_conv2d_8_source_31_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_31_pat_stride_1), .S(_05744_), .Y(_23410_) );
  \$mux  #( .WIDTH(32) ) _43664_ ( .A(_source_stream_conv2d_8_source_31_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_31_pat_stride_0), .S(_05744_), .Y(_23411_) );
  \$mux  #( .WIDTH(33) ) _43666_ ( .A(_source_stream_conv2d_8_source_31_pat_size_buf_3), .B(_source_stream_conv2d_8_source_31_pat_size_3), .S(_05744_), .Y(_23412_) );
  \$mux  #( .WIDTH(33) ) _43668_ ( .A(_source_stream_conv2d_8_source_31_pat_size_buf_2), .B(_source_stream_conv2d_8_source_31_pat_size_2), .S(_05744_), .Y(_23413_) );
  \$mux  #( .WIDTH(33) ) _43670_ ( .A(_source_stream_conv2d_8_source_31_pat_size_buf_1), .B(_source_stream_conv2d_8_source_31_pat_size_1), .S(_05744_), .Y(_23414_) );
  \$mux  #( .WIDTH(33) ) _43672_ ( .A(_source_stream_conv2d_8_source_31_pat_size_buf_0), .B(_source_stream_conv2d_8_source_31_pat_size_0), .S(_05744_), .Y(_23415_) );
  \$mux  #( .WIDTH(33) ) _43674_ ( .A(_source_stream_conv2d_8_source_31_pat_count_3), .B(_26187_), .S(_05744_), .Y(_23416_) );
  \$mux  #( .WIDTH(33) ) _43675_ ( .A(_23416_), .B(_26194_), .S(_05747_), .Y(_23417_) );
  \$mux  #( .WIDTH(33) ) _43676_ ( .A(_23417_), .B(_26195_), .S(_05748_), .Y(_23418_) );
  \$mux  #( .WIDTH(33) ) _43678_ ( .A(_source_stream_conv2d_8_source_31_pat_count_2), .B(_26186_), .S(_05744_), .Y(_23419_) );
  \$mux  #( .WIDTH(33) ) _43679_ ( .A(_23419_), .B(_26192_), .S(_05746_), .Y(_23420_) );
  \$mux  #( .WIDTH(33) ) _43680_ ( .A(_23420_), .B(_26193_), .S(_05747_), .Y(_23421_) );
  \$mux  #( .WIDTH(33) ) _43682_ ( .A(_source_stream_conv2d_8_source_31_pat_count_1), .B(_26185_), .S(_05744_), .Y(_23422_) );
  \$mux  #( .WIDTH(33) ) _43683_ ( .A(_23422_), .B(_26190_), .S(_05745_), .Y(_23423_) );
  \$mux  #( .WIDTH(33) ) _43684_ ( .A(_23423_), .B(_26191_), .S(_05746_), .Y(_23424_) );
  \$mux  #( .WIDTH(33) ) _43686_ ( .A(_source_stream_conv2d_8_source_31_pat_count_0), .B(_26184_), .S(_05744_), .Y(_23425_) );
  \$mux  #( .WIDTH(33) ) _43687_ ( .A(_26188_), .B(_23425_), .S(_05071_), .Y(_23426_) );
  \$mux  #( .WIDTH(33) ) _43688_ ( .A(_23426_), .B(_26189_), .S(_05745_), .Y(_23427_) );
  \$mux  #( .WIDTH(32) ) _43690_ ( .A(_source_stream_conv2d_8_source_31_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23428_) );
  \$mux  #( .WIDTH(32) ) _43692_ ( .A(_source_stream_conv2d_8_source_31_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23429_) );
  \$mux  #( .WIDTH(32) ) _43694_ ( .A(_source_stream_conv2d_8_source_31_pat_stride_1), .B({ 27'h0000000, cparam_conv2d_8_inc_act_laddr_large }), .S(_set_flag_538), .Y(_23430_) );
  \$mux  #( .WIDTH(32) ) _43696_ ( .A(_source_stream_conv2d_8_source_31_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23431_) );
  \$mux  #( .WIDTH(33) ) _43698_ ( .A(_source_stream_conv2d_8_source_31_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23432_) );
  \$mux  #( .WIDTH(33) ) _43700_ ( .A(_source_stream_conv2d_8_source_31_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23433_) );
  \$mux  #( .WIDTH(33) ) _43702_ ( .A(_source_stream_conv2d_8_source_31_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23434_) );
  \$mux  #( .WIDTH(33) ) _43704_ ( .A(_source_stream_conv2d_8_source_31_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23435_) );
  \$mux  #( .WIDTH(32) ) _43706_ ( .A(_source_stream_conv2d_8_source_31_pat_cur_offset_3), .B(0), .S(_05744_), .Y(_23436_) );
  \$mux  #( .WIDTH(32) ) _43707_ ( .A(_23436_), .B(_22208_), .S(_05747_), .Y(_23437_) );
  \$mux  #( .WIDTH(32) ) _43708_ ( .A(_23437_), .B(0), .S(_05748_), .Y(_23438_) );
  \$mux  #( .WIDTH(32) ) _43710_ ( .A(_source_stream_conv2d_8_source_31_pat_cur_offset_2), .B(0), .S(_05744_), .Y(_23439_) );
  \$mux  #( .WIDTH(32) ) _43711_ ( .A(_23439_), .B(_22207_), .S(_05746_), .Y(_23440_) );
  \$mux  #( .WIDTH(32) ) _43712_ ( .A(_23440_), .B(0), .S(_05747_), .Y(_23441_) );
  \$mux  #( .WIDTH(32) ) _43714_ ( .A(_source_stream_conv2d_8_source_31_pat_cur_offset_1), .B(0), .S(_05744_), .Y(_23442_) );
  \$mux  #( .WIDTH(32) ) _43715_ ( .A(_23442_), .B(_22206_), .S(_05745_), .Y(_23443_) );
  \$mux  #( .WIDTH(32) ) _43716_ ( .A(_23443_), .B(0), .S(_05746_), .Y(_23444_) );
  \$mux  #( .WIDTH(32) ) _43718_ ( .A(_source_stream_conv2d_8_source_31_pat_cur_offset_0), .B(0), .S(_05744_), .Y(_23445_) );
  \$mux  #( .WIDTH(32) ) _43719_ ( .A(_22205_), .B(_23445_), .S(_05071_), .Y(_23446_) );
  \$mux  #( .WIDTH(32) ) _43720_ ( .A(_23446_), .B(0), .S(_05745_), .Y(_23447_) );
  \$mux  #( .WIDTH(8) ) _43722_ ( .A(__variable_wdata_484), .B(_stream_conv2d_8_source_30_source_ram_rdata), .S(_stream_conv2d_8_source_30_source_ram_rvalid), .Y(_23448_) );
  \$mux  #( .WIDTH(32) ) _43724_ ( .A(_source_stream_conv2d_8_source_30_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_30_pat_stride_3), .S(_05739_), .Y(_23449_) );
  \$mux  #( .WIDTH(32) ) _43726_ ( .A(_source_stream_conv2d_8_source_30_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_30_pat_stride_2), .S(_05739_), .Y(_23450_) );
  \$mux  #( .WIDTH(32) ) _43728_ ( .A(_source_stream_conv2d_8_source_30_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_30_pat_stride_1), .S(_05739_), .Y(_23451_) );
  \$mux  #( .WIDTH(32) ) _43730_ ( .A(_source_stream_conv2d_8_source_30_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_30_pat_stride_0), .S(_05739_), .Y(_23452_) );
  \$mux  #( .WIDTH(33) ) _43732_ ( .A(_source_stream_conv2d_8_source_30_pat_size_buf_3), .B(_source_stream_conv2d_8_source_30_pat_size_3), .S(_05739_), .Y(_23453_) );
  \$mux  #( .WIDTH(33) ) _43734_ ( .A(_source_stream_conv2d_8_source_30_pat_size_buf_2), .B(_source_stream_conv2d_8_source_30_pat_size_2), .S(_05739_), .Y(_23454_) );
  \$mux  #( .WIDTH(33) ) _43736_ ( .A(_source_stream_conv2d_8_source_30_pat_size_buf_1), .B(_source_stream_conv2d_8_source_30_pat_size_1), .S(_05739_), .Y(_23455_) );
  \$mux  #( .WIDTH(33) ) _43738_ ( .A(_source_stream_conv2d_8_source_30_pat_size_buf_0), .B(_source_stream_conv2d_8_source_30_pat_size_0), .S(_05739_), .Y(_23456_) );
  \$mux  #( .WIDTH(33) ) _43740_ ( .A(_source_stream_conv2d_8_source_30_pat_count_3), .B(_26175_), .S(_05739_), .Y(_23457_) );
  \$mux  #( .WIDTH(33) ) _43741_ ( .A(_23457_), .B(_26182_), .S(_05742_), .Y(_23458_) );
  \$mux  #( .WIDTH(33) ) _43742_ ( .A(_23458_), .B(_26183_), .S(_05743_), .Y(_23459_) );
  \$mux  #( .WIDTH(33) ) _43744_ ( .A(_source_stream_conv2d_8_source_30_pat_count_2), .B(_26174_), .S(_05739_), .Y(_23460_) );
  \$mux  #( .WIDTH(33) ) _43745_ ( .A(_23460_), .B(_26180_), .S(_05741_), .Y(_23461_) );
  \$mux  #( .WIDTH(33) ) _43746_ ( .A(_23461_), .B(_26181_), .S(_05742_), .Y(_23462_) );
  \$mux  #( .WIDTH(33) ) _43748_ ( .A(_source_stream_conv2d_8_source_30_pat_count_1), .B(_26173_), .S(_05739_), .Y(_23463_) );
  \$mux  #( .WIDTH(33) ) _43749_ ( .A(_23463_), .B(_26178_), .S(_05740_), .Y(_23464_) );
  \$mux  #( .WIDTH(33) ) _43750_ ( .A(_23464_), .B(_26179_), .S(_05741_), .Y(_23465_) );
  \$mux  #( .WIDTH(33) ) _43752_ ( .A(_source_stream_conv2d_8_source_30_pat_count_0), .B(_26172_), .S(_05739_), .Y(_23466_) );
  \$mux  #( .WIDTH(33) ) _43753_ ( .A(_26176_), .B(_23466_), .S(_05073_), .Y(_23467_) );
  \$mux  #( .WIDTH(33) ) _43754_ ( .A(_23467_), .B(_26177_), .S(_05740_), .Y(_23468_) );
  \$mux  #( .WIDTH(32) ) _43756_ ( .A(_source_stream_conv2d_8_source_30_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23469_) );
  \$mux  #( .WIDTH(32) ) _43758_ ( .A(_source_stream_conv2d_8_source_30_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23470_) );
  \$mux  #( .WIDTH(32) ) _43760_ ( .A(_source_stream_conv2d_8_source_30_pat_stride_1), .B({ 27'h0000000, cparam_conv2d_8_inc_act_laddr_large }), .S(_set_flag_538), .Y(_23471_) );
  \$mux  #( .WIDTH(32) ) _43762_ ( .A(_source_stream_conv2d_8_source_30_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23472_) );
  \$mux  #( .WIDTH(33) ) _43764_ ( .A(_source_stream_conv2d_8_source_30_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23473_) );
  \$mux  #( .WIDTH(33) ) _43766_ ( .A(_source_stream_conv2d_8_source_30_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23474_) );
  \$mux  #( .WIDTH(33) ) _43768_ ( .A(_source_stream_conv2d_8_source_30_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23475_) );
  \$mux  #( .WIDTH(33) ) _43770_ ( .A(_source_stream_conv2d_8_source_30_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23476_) );
  \$mux  #( .WIDTH(32) ) _43772_ ( .A(_source_stream_conv2d_8_source_30_pat_cur_offset_3), .B(0), .S(_05739_), .Y(_23477_) );
  \$mux  #( .WIDTH(32) ) _43773_ ( .A(_23477_), .B(_22204_), .S(_05742_), .Y(_23478_) );
  \$mux  #( .WIDTH(32) ) _43774_ ( .A(_23478_), .B(0), .S(_05743_), .Y(_23479_) );
  \$mux  #( .WIDTH(32) ) _43776_ ( .A(_source_stream_conv2d_8_source_30_pat_cur_offset_2), .B(0), .S(_05739_), .Y(_23480_) );
  \$mux  #( .WIDTH(32) ) _43777_ ( .A(_23480_), .B(_22203_), .S(_05741_), .Y(_23481_) );
  \$mux  #( .WIDTH(32) ) _43778_ ( .A(_23481_), .B(0), .S(_05742_), .Y(_23482_) );
  \$mux  #( .WIDTH(32) ) _43780_ ( .A(_source_stream_conv2d_8_source_30_pat_cur_offset_1), .B(0), .S(_05739_), .Y(_23483_) );
  \$mux  #( .WIDTH(32) ) _43781_ ( .A(_23483_), .B(_22202_), .S(_05740_), .Y(_23484_) );
  \$mux  #( .WIDTH(32) ) _43782_ ( .A(_23484_), .B(0), .S(_05741_), .Y(_23485_) );
  \$mux  #( .WIDTH(32) ) _43784_ ( .A(_source_stream_conv2d_8_source_30_pat_cur_offset_0), .B(0), .S(_05739_), .Y(_23486_) );
  \$mux  #( .WIDTH(32) ) _43785_ ( .A(_22201_), .B(_23486_), .S(_05073_), .Y(_23487_) );
  \$mux  #( .WIDTH(32) ) _43786_ ( .A(_23487_), .B(0), .S(_05740_), .Y(_23488_) );
  \$mux  #( .WIDTH(8) ) _43788_ ( .A(__variable_wdata_483), .B(_stream_conv2d_8_source_29_source_ram_rdata), .S(_stream_conv2d_8_source_29_source_ram_rvalid), .Y(_23489_) );
  \$mux  #( .WIDTH(32) ) _43790_ ( .A(_source_stream_conv2d_8_source_29_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_29_pat_stride_3), .S(_05734_), .Y(_23490_) );
  \$mux  #( .WIDTH(32) ) _43792_ ( .A(_source_stream_conv2d_8_source_29_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_29_pat_stride_2), .S(_05734_), .Y(_23491_) );
  \$mux  #( .WIDTH(32) ) _43794_ ( .A(_source_stream_conv2d_8_source_29_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_29_pat_stride_1), .S(_05734_), .Y(_23492_) );
  \$mux  #( .WIDTH(32) ) _43796_ ( .A(_source_stream_conv2d_8_source_29_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_29_pat_stride_0), .S(_05734_), .Y(_23493_) );
  \$mux  #( .WIDTH(33) ) _43798_ ( .A(_source_stream_conv2d_8_source_29_pat_size_buf_3), .B(_source_stream_conv2d_8_source_29_pat_size_3), .S(_05734_), .Y(_23494_) );
  \$mux  #( .WIDTH(33) ) _43800_ ( .A(_source_stream_conv2d_8_source_29_pat_size_buf_2), .B(_source_stream_conv2d_8_source_29_pat_size_2), .S(_05734_), .Y(_23495_) );
  \$mux  #( .WIDTH(33) ) _43802_ ( .A(_source_stream_conv2d_8_source_29_pat_size_buf_1), .B(_source_stream_conv2d_8_source_29_pat_size_1), .S(_05734_), .Y(_23496_) );
  \$mux  #( .WIDTH(33) ) _43804_ ( .A(_source_stream_conv2d_8_source_29_pat_size_buf_0), .B(_source_stream_conv2d_8_source_29_pat_size_0), .S(_05734_), .Y(_23497_) );
  \$mux  #( .WIDTH(33) ) _43806_ ( .A(_source_stream_conv2d_8_source_29_pat_count_3), .B(_26163_), .S(_05734_), .Y(_23498_) );
  \$mux  #( .WIDTH(33) ) _43807_ ( .A(_23498_), .B(_26170_), .S(_05737_), .Y(_23499_) );
  \$mux  #( .WIDTH(33) ) _43808_ ( .A(_23499_), .B(_26171_), .S(_05738_), .Y(_23500_) );
  \$mux  #( .WIDTH(33) ) _43810_ ( .A(_source_stream_conv2d_8_source_29_pat_count_2), .B(_26162_), .S(_05734_), .Y(_23501_) );
  \$mux  #( .WIDTH(33) ) _43811_ ( .A(_23501_), .B(_26168_), .S(_05736_), .Y(_23502_) );
  \$mux  #( .WIDTH(33) ) _43812_ ( .A(_23502_), .B(_26169_), .S(_05737_), .Y(_23503_) );
  \$mux  #( .WIDTH(33) ) _43814_ ( .A(_source_stream_conv2d_8_source_29_pat_count_1), .B(_26161_), .S(_05734_), .Y(_23504_) );
  \$mux  #( .WIDTH(33) ) _43815_ ( .A(_23504_), .B(_26166_), .S(_05735_), .Y(_23505_) );
  \$mux  #( .WIDTH(33) ) _43816_ ( .A(_23505_), .B(_26167_), .S(_05736_), .Y(_23506_) );
  \$mux  #( .WIDTH(33) ) _43818_ ( .A(_source_stream_conv2d_8_source_29_pat_count_0), .B(_26160_), .S(_05734_), .Y(_23507_) );
  \$mux  #( .WIDTH(33) ) _43819_ ( .A(_26164_), .B(_23507_), .S(_05075_), .Y(_23508_) );
  \$mux  #( .WIDTH(33) ) _43820_ ( .A(_23508_), .B(_26165_), .S(_05735_), .Y(_23509_) );
  \$mux  #( .WIDTH(32) ) _43822_ ( .A(_source_stream_conv2d_8_source_29_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23510_) );
  \$mux  #( .WIDTH(32) ) _43824_ ( .A(_source_stream_conv2d_8_source_29_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23511_) );
  \$mux  #( .WIDTH(32) ) _43826_ ( .A(_source_stream_conv2d_8_source_29_pat_stride_1), .B({ 27'h0000000, cparam_conv2d_8_inc_act_laddr_large }), .S(_set_flag_538), .Y(_23512_) );
  \$mux  #( .WIDTH(32) ) _43828_ ( .A(_source_stream_conv2d_8_source_29_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23513_) );
  \$mux  #( .WIDTH(33) ) _43830_ ( .A(_source_stream_conv2d_8_source_29_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23514_) );
  \$mux  #( .WIDTH(33) ) _43832_ ( .A(_source_stream_conv2d_8_source_29_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23515_) );
  \$mux  #( .WIDTH(33) ) _43834_ ( .A(_source_stream_conv2d_8_source_29_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23516_) );
  \$mux  #( .WIDTH(33) ) _43836_ ( .A(_source_stream_conv2d_8_source_29_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23517_) );
  \$mux  #( .WIDTH(32) ) _43838_ ( .A(_source_stream_conv2d_8_source_29_pat_cur_offset_3), .B(0), .S(_05734_), .Y(_23518_) );
  \$mux  #( .WIDTH(32) ) _43839_ ( .A(_23518_), .B(_22200_), .S(_05737_), .Y(_23519_) );
  \$mux  #( .WIDTH(32) ) _43840_ ( .A(_23519_), .B(0), .S(_05738_), .Y(_23520_) );
  \$mux  #( .WIDTH(32) ) _43842_ ( .A(_source_stream_conv2d_8_source_29_pat_cur_offset_2), .B(0), .S(_05734_), .Y(_23521_) );
  \$mux  #( .WIDTH(32) ) _43843_ ( .A(_23521_), .B(_22199_), .S(_05736_), .Y(_23522_) );
  \$mux  #( .WIDTH(32) ) _43844_ ( .A(_23522_), .B(0), .S(_05737_), .Y(_23523_) );
  \$mux  #( .WIDTH(32) ) _43846_ ( .A(_source_stream_conv2d_8_source_29_pat_cur_offset_1), .B(0), .S(_05734_), .Y(_23524_) );
  \$mux  #( .WIDTH(32) ) _43847_ ( .A(_23524_), .B(_22198_), .S(_05735_), .Y(_23525_) );
  \$mux  #( .WIDTH(32) ) _43848_ ( .A(_23525_), .B(0), .S(_05736_), .Y(_23526_) );
  \$mux  #( .WIDTH(32) ) _43850_ ( .A(_source_stream_conv2d_8_source_29_pat_cur_offset_0), .B(0), .S(_05734_), .Y(_23527_) );
  \$mux  #( .WIDTH(32) ) _43851_ ( .A(_22197_), .B(_23527_), .S(_05075_), .Y(_23528_) );
  \$mux  #( .WIDTH(32) ) _43852_ ( .A(_23528_), .B(0), .S(_05735_), .Y(_23529_) );
  \$mux  #( .WIDTH(8) ) _43854_ ( .A(__variable_wdata_482), .B(_stream_conv2d_8_source_28_source_ram_rdata), .S(_stream_conv2d_8_source_28_source_ram_rvalid), .Y(_23530_) );
  \$mux  #( .WIDTH(32) ) _43856_ ( .A(_source_stream_conv2d_8_source_28_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_28_pat_stride_3), .S(_05729_), .Y(_23531_) );
  \$mux  #( .WIDTH(32) ) _43858_ ( .A(_source_stream_conv2d_8_source_28_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_28_pat_stride_2), .S(_05729_), .Y(_23532_) );
  \$mux  #( .WIDTH(32) ) _43860_ ( .A(_source_stream_conv2d_8_source_28_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_28_pat_stride_1), .S(_05729_), .Y(_23533_) );
  \$mux  #( .WIDTH(32) ) _43862_ ( .A(_source_stream_conv2d_8_source_28_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_28_pat_stride_0), .S(_05729_), .Y(_23534_) );
  \$mux  #( .WIDTH(33) ) _43864_ ( .A(_source_stream_conv2d_8_source_28_pat_size_buf_3), .B(_source_stream_conv2d_8_source_28_pat_size_3), .S(_05729_), .Y(_23535_) );
  \$mux  #( .WIDTH(33) ) _43866_ ( .A(_source_stream_conv2d_8_source_28_pat_size_buf_2), .B(_source_stream_conv2d_8_source_28_pat_size_2), .S(_05729_), .Y(_23536_) );
  \$mux  #( .WIDTH(33) ) _43868_ ( .A(_source_stream_conv2d_8_source_28_pat_size_buf_1), .B(_source_stream_conv2d_8_source_28_pat_size_1), .S(_05729_), .Y(_23537_) );
  \$mux  #( .WIDTH(33) ) _43870_ ( .A(_source_stream_conv2d_8_source_28_pat_size_buf_0), .B(_source_stream_conv2d_8_source_28_pat_size_0), .S(_05729_), .Y(_23538_) );
  \$mux  #( .WIDTH(33) ) _43872_ ( .A(_source_stream_conv2d_8_source_28_pat_count_3), .B(_26151_), .S(_05729_), .Y(_23539_) );
  \$mux  #( .WIDTH(33) ) _43873_ ( .A(_23539_), .B(_26158_), .S(_05732_), .Y(_23540_) );
  \$mux  #( .WIDTH(33) ) _43874_ ( .A(_23540_), .B(_26159_), .S(_05733_), .Y(_23541_) );
  \$mux  #( .WIDTH(33) ) _43876_ ( .A(_source_stream_conv2d_8_source_28_pat_count_2), .B(_26150_), .S(_05729_), .Y(_23542_) );
  \$mux  #( .WIDTH(33) ) _43877_ ( .A(_23542_), .B(_26156_), .S(_05731_), .Y(_23543_) );
  \$mux  #( .WIDTH(33) ) _43878_ ( .A(_23543_), .B(_26157_), .S(_05732_), .Y(_23544_) );
  \$mux  #( .WIDTH(33) ) _43880_ ( .A(_source_stream_conv2d_8_source_28_pat_count_1), .B(_26149_), .S(_05729_), .Y(_23545_) );
  \$mux  #( .WIDTH(33) ) _43881_ ( .A(_23545_), .B(_26154_), .S(_05730_), .Y(_23546_) );
  \$mux  #( .WIDTH(33) ) _43882_ ( .A(_23546_), .B(_26155_), .S(_05731_), .Y(_23547_) );
  \$mux  #( .WIDTH(33) ) _43884_ ( .A(_source_stream_conv2d_8_source_28_pat_count_0), .B(_26148_), .S(_05729_), .Y(_23548_) );
  \$mux  #( .WIDTH(33) ) _43885_ ( .A(_26152_), .B(_23548_), .S(_05077_), .Y(_23549_) );
  \$mux  #( .WIDTH(33) ) _43886_ ( .A(_23549_), .B(_26153_), .S(_05730_), .Y(_23550_) );
  \$mux  #( .WIDTH(32) ) _43888_ ( .A(_source_stream_conv2d_8_source_28_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23551_) );
  \$mux  #( .WIDTH(32) ) _43890_ ( .A(_source_stream_conv2d_8_source_28_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23552_) );
  \$mux  #( .WIDTH(32) ) _43892_ ( .A(_source_stream_conv2d_8_source_28_pat_stride_1), .B({ 27'h0000000, cparam_conv2d_8_inc_act_laddr_large }), .S(_set_flag_538), .Y(_23553_) );
  \$mux  #( .WIDTH(32) ) _43894_ ( .A(_source_stream_conv2d_8_source_28_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23554_) );
  \$mux  #( .WIDTH(33) ) _43896_ ( .A(_source_stream_conv2d_8_source_28_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23555_) );
  \$mux  #( .WIDTH(33) ) _43898_ ( .A(_source_stream_conv2d_8_source_28_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23556_) );
  \$mux  #( .WIDTH(33) ) _43900_ ( .A(_source_stream_conv2d_8_source_28_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23557_) );
  \$mux  #( .WIDTH(33) ) _43902_ ( .A(_source_stream_conv2d_8_source_28_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23558_) );
  \$mux  #( .WIDTH(32) ) _43904_ ( .A(_source_stream_conv2d_8_source_28_pat_cur_offset_3), .B(0), .S(_05729_), .Y(_23559_) );
  \$mux  #( .WIDTH(32) ) _43905_ ( .A(_23559_), .B(_22196_), .S(_05732_), .Y(_23560_) );
  \$mux  #( .WIDTH(32) ) _43906_ ( .A(_23560_), .B(0), .S(_05733_), .Y(_23561_) );
  \$mux  #( .WIDTH(32) ) _43908_ ( .A(_source_stream_conv2d_8_source_28_pat_cur_offset_2), .B(0), .S(_05729_), .Y(_23562_) );
  \$mux  #( .WIDTH(32) ) _43909_ ( .A(_23562_), .B(_22195_), .S(_05731_), .Y(_23563_) );
  \$mux  #( .WIDTH(32) ) _43910_ ( .A(_23563_), .B(0), .S(_05732_), .Y(_23564_) );
  \$mux  #( .WIDTH(32) ) _43912_ ( .A(_source_stream_conv2d_8_source_28_pat_cur_offset_1), .B(0), .S(_05729_), .Y(_23565_) );
  \$mux  #( .WIDTH(32) ) _43913_ ( .A(_23565_), .B(_22194_), .S(_05730_), .Y(_23566_) );
  \$mux  #( .WIDTH(32) ) _43914_ ( .A(_23566_), .B(0), .S(_05731_), .Y(_23567_) );
  \$mux  #( .WIDTH(32) ) _43916_ ( .A(_source_stream_conv2d_8_source_28_pat_cur_offset_0), .B(0), .S(_05729_), .Y(_23568_) );
  \$mux  #( .WIDTH(32) ) _43917_ ( .A(_22193_), .B(_23568_), .S(_05077_), .Y(_23569_) );
  \$mux  #( .WIDTH(32) ) _43918_ ( .A(_23569_), .B(0), .S(_05730_), .Y(_23570_) );
  \$mux  #( .WIDTH(8) ) _43920_ ( .A(__variable_wdata_256), .B(_stream_conv2d_8_source_27_source_ram_rdata), .S(_stream_conv2d_8_source_27_source_ram_rvalid), .Y(_23571_) );
  \$mux  #( .WIDTH(32) ) _43922_ ( .A(_source_stream_conv2d_8_source_27_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_27_pat_stride_3), .S(_05724_), .Y(_23572_) );
  \$mux  #( .WIDTH(32) ) _43924_ ( .A(_source_stream_conv2d_8_source_27_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_27_pat_stride_2), .S(_05724_), .Y(_23573_) );
  \$mux  #( .WIDTH(32) ) _43926_ ( .A(_source_stream_conv2d_8_source_27_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_27_pat_stride_1), .S(_05724_), .Y(_23574_) );
  \$mux  #( .WIDTH(32) ) _43928_ ( .A(_source_stream_conv2d_8_source_27_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_27_pat_stride_0), .S(_05724_), .Y(_23575_) );
  \$mux  #( .WIDTH(33) ) _43930_ ( .A(_source_stream_conv2d_8_source_27_pat_size_buf_3), .B(_source_stream_conv2d_8_source_27_pat_size_3), .S(_05724_), .Y(_23576_) );
  \$mux  #( .WIDTH(33) ) _43932_ ( .A(_source_stream_conv2d_8_source_27_pat_size_buf_2), .B(_source_stream_conv2d_8_source_27_pat_size_2), .S(_05724_), .Y(_23577_) );
  \$mux  #( .WIDTH(33) ) _43934_ ( .A(_source_stream_conv2d_8_source_27_pat_size_buf_1), .B(_source_stream_conv2d_8_source_27_pat_size_1), .S(_05724_), .Y(_23578_) );
  \$mux  #( .WIDTH(33) ) _43936_ ( .A(_source_stream_conv2d_8_source_27_pat_size_buf_0), .B(_source_stream_conv2d_8_source_27_pat_size_0), .S(_05724_), .Y(_23579_) );
  \$mux  #( .WIDTH(33) ) _43938_ ( .A(_source_stream_conv2d_8_source_27_pat_count_3), .B(_26139_), .S(_05724_), .Y(_23580_) );
  \$mux  #( .WIDTH(33) ) _43939_ ( .A(_23580_), .B(_26146_), .S(_05727_), .Y(_23581_) );
  \$mux  #( .WIDTH(33) ) _43940_ ( .A(_23581_), .B(_26147_), .S(_05728_), .Y(_23582_) );
  \$mux  #( .WIDTH(33) ) _43942_ ( .A(_source_stream_conv2d_8_source_27_pat_count_2), .B(_26138_), .S(_05724_), .Y(_23583_) );
  \$mux  #( .WIDTH(33) ) _43943_ ( .A(_23583_), .B(_26144_), .S(_05726_), .Y(_23584_) );
  \$mux  #( .WIDTH(33) ) _43944_ ( .A(_23584_), .B(_26145_), .S(_05727_), .Y(_23585_) );
  \$mux  #( .WIDTH(33) ) _43946_ ( .A(_source_stream_conv2d_8_source_27_pat_count_1), .B(_26137_), .S(_05724_), .Y(_23586_) );
  \$mux  #( .WIDTH(33) ) _43947_ ( .A(_23586_), .B(_26142_), .S(_05725_), .Y(_23587_) );
  \$mux  #( .WIDTH(33) ) _43948_ ( .A(_23587_), .B(_26143_), .S(_05726_), .Y(_23588_) );
  \$mux  #( .WIDTH(33) ) _43950_ ( .A(_source_stream_conv2d_8_source_27_pat_count_0), .B(_26136_), .S(_05724_), .Y(_23589_) );
  \$mux  #( .WIDTH(33) ) _43951_ ( .A(_26140_), .B(_23589_), .S(_05079_), .Y(_23590_) );
  \$mux  #( .WIDTH(33) ) _43952_ ( .A(_23590_), .B(_26141_), .S(_05725_), .Y(_23591_) );
  \$mux  #( .WIDTH(32) ) _43954_ ( .A(_source_stream_conv2d_8_source_27_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23592_) );
  \$mux  #( .WIDTH(32) ) _43956_ ( .A(_source_stream_conv2d_8_source_27_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23593_) );
  \$mux  #( .WIDTH(32) ) _43958_ ( .A(_source_stream_conv2d_8_source_27_pat_stride_1), .B(0), .S(_set_flag_538), .Y(_23594_) );
  \$mux  #( .WIDTH(32) ) _43960_ ( .A(_source_stream_conv2d_8_source_27_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23595_) );
  \$mux  #( .WIDTH(33) ) _43962_ ( .A(_source_stream_conv2d_8_source_27_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23596_) );
  \$mux  #( .WIDTH(33) ) _43964_ ( .A(_source_stream_conv2d_8_source_27_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23597_) );
  \$mux  #( .WIDTH(33) ) _43966_ ( .A(_source_stream_conv2d_8_source_27_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23598_) );
  \$mux  #( .WIDTH(33) ) _43968_ ( .A(_source_stream_conv2d_8_source_27_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23599_) );
  \$mux  #( .WIDTH(32) ) _43970_ ( .A(_source_stream_conv2d_8_source_27_pat_cur_offset_3), .B(0), .S(_05724_), .Y(_23600_) );
  \$mux  #( .WIDTH(32) ) _43971_ ( .A(_23600_), .B(_22192_), .S(_05727_), .Y(_23601_) );
  \$mux  #( .WIDTH(32) ) _43972_ ( .A(_23601_), .B(0), .S(_05728_), .Y(_23602_) );
  \$mux  #( .WIDTH(32) ) _43974_ ( .A(_source_stream_conv2d_8_source_27_pat_cur_offset_2), .B(0), .S(_05724_), .Y(_23603_) );
  \$mux  #( .WIDTH(32) ) _43975_ ( .A(_23603_), .B(_22191_), .S(_05726_), .Y(_23604_) );
  \$mux  #( .WIDTH(32) ) _43976_ ( .A(_23604_), .B(0), .S(_05727_), .Y(_23605_) );
  \$mux  #( .WIDTH(32) ) _43978_ ( .A(_source_stream_conv2d_8_source_27_pat_cur_offset_1), .B(0), .S(_05724_), .Y(_23606_) );
  \$mux  #( .WIDTH(32) ) _43979_ ( .A(_23606_), .B(_22190_), .S(_05725_), .Y(_23607_) );
  \$mux  #( .WIDTH(32) ) _43980_ ( .A(_23607_), .B(0), .S(_05726_), .Y(_23608_) );
  \$mux  #( .WIDTH(32) ) _43982_ ( .A(_source_stream_conv2d_8_source_27_pat_cur_offset_0), .B(0), .S(_05724_), .Y(_23609_) );
  \$mux  #( .WIDTH(32) ) _43983_ ( .A(_22189_), .B(_23609_), .S(_05079_), .Y(_23610_) );
  \$mux  #( .WIDTH(32) ) _43984_ ( .A(_23610_), .B(0), .S(_05725_), .Y(_23611_) );
  \$mux  #( .WIDTH(8) ) _43986_ ( .A(__variable_wdata_255), .B(_stream_conv2d_8_source_26_source_ram_rdata), .S(_stream_conv2d_8_source_26_source_ram_rvalid), .Y(_23612_) );
  \$mux  #( .WIDTH(32) ) _43988_ ( .A(_source_stream_conv2d_8_source_26_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_26_pat_stride_3), .S(_05719_), .Y(_23613_) );
  \$mux  #( .WIDTH(32) ) _43990_ ( .A(_source_stream_conv2d_8_source_26_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_26_pat_stride_2), .S(_05719_), .Y(_23614_) );
  \$mux  #( .WIDTH(32) ) _43992_ ( .A(_source_stream_conv2d_8_source_26_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_26_pat_stride_1), .S(_05719_), .Y(_23615_) );
  \$mux  #( .WIDTH(32) ) _43994_ ( .A(_source_stream_conv2d_8_source_26_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_26_pat_stride_0), .S(_05719_), .Y(_23616_) );
  \$mux  #( .WIDTH(33) ) _43996_ ( .A(_source_stream_conv2d_8_source_26_pat_size_buf_3), .B(_source_stream_conv2d_8_source_26_pat_size_3), .S(_05719_), .Y(_23617_) );
  \$mux  #( .WIDTH(33) ) _43998_ ( .A(_source_stream_conv2d_8_source_26_pat_size_buf_2), .B(_source_stream_conv2d_8_source_26_pat_size_2), .S(_05719_), .Y(_23618_) );
  \$mux  #( .WIDTH(33) ) _44000_ ( .A(_source_stream_conv2d_8_source_26_pat_size_buf_1), .B(_source_stream_conv2d_8_source_26_pat_size_1), .S(_05719_), .Y(_23619_) );
  \$mux  #( .WIDTH(33) ) _44002_ ( .A(_source_stream_conv2d_8_source_26_pat_size_buf_0), .B(_source_stream_conv2d_8_source_26_pat_size_0), .S(_05719_), .Y(_23620_) );
  \$mux  #( .WIDTH(33) ) _44004_ ( .A(_source_stream_conv2d_8_source_26_pat_count_3), .B(_26127_), .S(_05719_), .Y(_23621_) );
  \$mux  #( .WIDTH(33) ) _44005_ ( .A(_23621_), .B(_26134_), .S(_05722_), .Y(_23622_) );
  \$mux  #( .WIDTH(33) ) _44006_ ( .A(_23622_), .B(_26135_), .S(_05723_), .Y(_23623_) );
  \$mux  #( .WIDTH(33) ) _44008_ ( .A(_source_stream_conv2d_8_source_26_pat_count_2), .B(_26126_), .S(_05719_), .Y(_23624_) );
  \$mux  #( .WIDTH(33) ) _44009_ ( .A(_23624_), .B(_26132_), .S(_05721_), .Y(_23625_) );
  \$mux  #( .WIDTH(33) ) _44010_ ( .A(_23625_), .B(_26133_), .S(_05722_), .Y(_23626_) );
  \$mux  #( .WIDTH(33) ) _44012_ ( .A(_source_stream_conv2d_8_source_26_pat_count_1), .B(_26125_), .S(_05719_), .Y(_23627_) );
  \$mux  #( .WIDTH(33) ) _44013_ ( .A(_23627_), .B(_26130_), .S(_05720_), .Y(_23628_) );
  \$mux  #( .WIDTH(33) ) _44014_ ( .A(_23628_), .B(_26131_), .S(_05721_), .Y(_23629_) );
  \$mux  #( .WIDTH(33) ) _44016_ ( .A(_source_stream_conv2d_8_source_26_pat_count_0), .B(_26124_), .S(_05719_), .Y(_23630_) );
  \$mux  #( .WIDTH(33) ) _44017_ ( .A(_26128_), .B(_23630_), .S(_05081_), .Y(_23631_) );
  \$mux  #( .WIDTH(33) ) _44018_ ( .A(_23631_), .B(_26129_), .S(_05720_), .Y(_23632_) );
  \$mux  #( .WIDTH(32) ) _44020_ ( .A(_source_stream_conv2d_8_source_26_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23633_) );
  \$mux  #( .WIDTH(32) ) _44022_ ( .A(_source_stream_conv2d_8_source_26_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23634_) );
  \$mux  #( .WIDTH(32) ) _44024_ ( .A(_source_stream_conv2d_8_source_26_pat_stride_1), .B(0), .S(_set_flag_538), .Y(_23635_) );
  \$mux  #( .WIDTH(32) ) _44026_ ( .A(_source_stream_conv2d_8_source_26_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23636_) );
  \$mux  #( .WIDTH(33) ) _44028_ ( .A(_source_stream_conv2d_8_source_26_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23637_) );
  \$mux  #( .WIDTH(33) ) _44030_ ( .A(_source_stream_conv2d_8_source_26_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23638_) );
  \$mux  #( .WIDTH(33) ) _44032_ ( .A(_source_stream_conv2d_8_source_26_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23639_) );
  \$mux  #( .WIDTH(33) ) _44034_ ( .A(_source_stream_conv2d_8_source_26_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23640_) );
  \$mux  #( .WIDTH(32) ) _44036_ ( .A(_source_stream_conv2d_8_source_26_pat_cur_offset_3), .B(0), .S(_05719_), .Y(_23641_) );
  \$mux  #( .WIDTH(32) ) _44037_ ( .A(_23641_), .B(_22187_), .S(_05722_), .Y(_23642_) );
  \$mux  #( .WIDTH(32) ) _44038_ ( .A(_23642_), .B(0), .S(_05723_), .Y(_23643_) );
  \$mux  #( .WIDTH(32) ) _44040_ ( .A(_source_stream_conv2d_8_source_26_pat_cur_offset_2), .B(0), .S(_05719_), .Y(_23644_) );
  \$mux  #( .WIDTH(32) ) _44041_ ( .A(_23644_), .B(_22186_), .S(_05721_), .Y(_23645_) );
  \$mux  #( .WIDTH(32) ) _44042_ ( .A(_23645_), .B(0), .S(_05722_), .Y(_23646_) );
  \$mux  #( .WIDTH(32) ) _44044_ ( .A(_source_stream_conv2d_8_source_26_pat_cur_offset_1), .B(0), .S(_05719_), .Y(_23647_) );
  \$mux  #( .WIDTH(32) ) _44045_ ( .A(_23647_), .B(_22185_), .S(_05720_), .Y(_23648_) );
  \$mux  #( .WIDTH(32) ) _44046_ ( .A(_23648_), .B(0), .S(_05721_), .Y(_23649_) );
  \$mux  #( .WIDTH(32) ) _44048_ ( .A(_source_stream_conv2d_8_source_26_pat_cur_offset_0), .B(0), .S(_05719_), .Y(_23650_) );
  \$mux  #( .WIDTH(32) ) _44049_ ( .A(_22184_), .B(_23650_), .S(_05081_), .Y(_23651_) );
  \$mux  #( .WIDTH(32) ) _44050_ ( .A(_23651_), .B(0), .S(_05720_), .Y(_23652_) );
  \$mux  #( .WIDTH(8) ) _44052_ ( .A(__variable_wdata_254), .B(_stream_conv2d_8_source_25_source_ram_rdata), .S(_stream_conv2d_8_source_25_source_ram_rvalid), .Y(_23653_) );
  \$mux  #( .WIDTH(32) ) _44054_ ( .A(_source_stream_conv2d_8_source_25_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_25_pat_stride_3), .S(_05714_), .Y(_23654_) );
  \$mux  #( .WIDTH(32) ) _44056_ ( .A(_source_stream_conv2d_8_source_25_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_25_pat_stride_2), .S(_05714_), .Y(_23655_) );
  \$mux  #( .WIDTH(32) ) _44058_ ( .A(_source_stream_conv2d_8_source_25_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_25_pat_stride_1), .S(_05714_), .Y(_23656_) );
  \$mux  #( .WIDTH(32) ) _44060_ ( .A(_source_stream_conv2d_8_source_25_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_25_pat_stride_0), .S(_05714_), .Y(_23657_) );
  \$mux  #( .WIDTH(33) ) _44062_ ( .A(_source_stream_conv2d_8_source_25_pat_size_buf_3), .B(_source_stream_conv2d_8_source_25_pat_size_3), .S(_05714_), .Y(_23658_) );
  \$mux  #( .WIDTH(33) ) _44064_ ( .A(_source_stream_conv2d_8_source_25_pat_size_buf_2), .B(_source_stream_conv2d_8_source_25_pat_size_2), .S(_05714_), .Y(_23659_) );
  \$mux  #( .WIDTH(33) ) _44066_ ( .A(_source_stream_conv2d_8_source_25_pat_size_buf_1), .B(_source_stream_conv2d_8_source_25_pat_size_1), .S(_05714_), .Y(_23660_) );
  \$mux  #( .WIDTH(33) ) _44068_ ( .A(_source_stream_conv2d_8_source_25_pat_size_buf_0), .B(_source_stream_conv2d_8_source_25_pat_size_0), .S(_05714_), .Y(_23661_) );
  \$mux  #( .WIDTH(33) ) _44070_ ( .A(_source_stream_conv2d_8_source_25_pat_count_3), .B(_26115_), .S(_05714_), .Y(_23662_) );
  \$mux  #( .WIDTH(33) ) _44071_ ( .A(_23662_), .B(_26122_), .S(_05717_), .Y(_23663_) );
  \$mux  #( .WIDTH(33) ) _44072_ ( .A(_23663_), .B(_26123_), .S(_05718_), .Y(_23664_) );
  \$mux  #( .WIDTH(33) ) _44074_ ( .A(_source_stream_conv2d_8_source_25_pat_count_2), .B(_26114_), .S(_05714_), .Y(_23665_) );
  \$mux  #( .WIDTH(33) ) _44075_ ( .A(_23665_), .B(_26120_), .S(_05716_), .Y(_23666_) );
  \$mux  #( .WIDTH(33) ) _44076_ ( .A(_23666_), .B(_26121_), .S(_05717_), .Y(_23667_) );
  \$mux  #( .WIDTH(33) ) _44078_ ( .A(_source_stream_conv2d_8_source_25_pat_count_1), .B(_26113_), .S(_05714_), .Y(_23668_) );
  \$mux  #( .WIDTH(33) ) _44079_ ( .A(_23668_), .B(_26118_), .S(_05715_), .Y(_23669_) );
  \$mux  #( .WIDTH(33) ) _44080_ ( .A(_23669_), .B(_26119_), .S(_05716_), .Y(_23670_) );
  \$mux  #( .WIDTH(33) ) _44082_ ( .A(_source_stream_conv2d_8_source_25_pat_count_0), .B(_26112_), .S(_05714_), .Y(_23671_) );
  \$mux  #( .WIDTH(33) ) _44083_ ( .A(_26116_), .B(_23671_), .S(_05083_), .Y(_23672_) );
  \$mux  #( .WIDTH(33) ) _44084_ ( .A(_23672_), .B(_26117_), .S(_05715_), .Y(_23673_) );
  \$mux  #( .WIDTH(32) ) _44086_ ( .A(_source_stream_conv2d_8_source_25_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23674_) );
  \$mux  #( .WIDTH(32) ) _44088_ ( .A(_source_stream_conv2d_8_source_25_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23675_) );
  \$mux  #( .WIDTH(32) ) _44090_ ( .A(_source_stream_conv2d_8_source_25_pat_stride_1), .B(0), .S(_set_flag_538), .Y(_23676_) );
  \$mux  #( .WIDTH(32) ) _44092_ ( .A(_source_stream_conv2d_8_source_25_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23677_) );
  \$mux  #( .WIDTH(33) ) _44094_ ( .A(_source_stream_conv2d_8_source_25_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23678_) );
  \$mux  #( .WIDTH(33) ) _44096_ ( .A(_source_stream_conv2d_8_source_25_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23679_) );
  \$mux  #( .WIDTH(33) ) _44098_ ( .A(_source_stream_conv2d_8_source_25_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23680_) );
  \$mux  #( .WIDTH(33) ) _44100_ ( .A(_source_stream_conv2d_8_source_25_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23681_) );
  \$mux  #( .WIDTH(32) ) _44102_ ( .A(_source_stream_conv2d_8_source_25_pat_cur_offset_3), .B(0), .S(_05714_), .Y(_23682_) );
  \$mux  #( .WIDTH(32) ) _44103_ ( .A(_23682_), .B(_22182_), .S(_05717_), .Y(_23683_) );
  \$mux  #( .WIDTH(32) ) _44104_ ( .A(_23683_), .B(0), .S(_05718_), .Y(_23684_) );
  \$mux  #( .WIDTH(32) ) _44106_ ( .A(_source_stream_conv2d_8_source_25_pat_cur_offset_2), .B(0), .S(_05714_), .Y(_23685_) );
  \$mux  #( .WIDTH(32) ) _44107_ ( .A(_23685_), .B(_22181_), .S(_05716_), .Y(_23686_) );
  \$mux  #( .WIDTH(32) ) _44108_ ( .A(_23686_), .B(0), .S(_05717_), .Y(_23687_) );
  \$mux  #( .WIDTH(32) ) _44110_ ( .A(_source_stream_conv2d_8_source_25_pat_cur_offset_1), .B(0), .S(_05714_), .Y(_23688_) );
  \$mux  #( .WIDTH(32) ) _44111_ ( .A(_23688_), .B(_22180_), .S(_05715_), .Y(_23689_) );
  \$mux  #( .WIDTH(32) ) _44112_ ( .A(_23689_), .B(0), .S(_05716_), .Y(_23690_) );
  \$mux  #( .WIDTH(32) ) _44114_ ( .A(_source_stream_conv2d_8_source_25_pat_cur_offset_0), .B(0), .S(_05714_), .Y(_23691_) );
  \$mux  #( .WIDTH(32) ) _44115_ ( .A(_22179_), .B(_23691_), .S(_05083_), .Y(_23692_) );
  \$mux  #( .WIDTH(32) ) _44116_ ( .A(_23692_), .B(0), .S(_05715_), .Y(_23693_) );
  \$mux  #( .WIDTH(8) ) _44118_ ( .A(__variable_wdata_253), .B(_stream_conv2d_8_source_24_source_ram_rdata), .S(_stream_conv2d_8_source_24_source_ram_rvalid), .Y(_23694_) );
  \$mux  #( .WIDTH(32) ) _44120_ ( .A(_source_stream_conv2d_8_source_24_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_24_pat_stride_3), .S(_05709_), .Y(_23695_) );
  \$mux  #( .WIDTH(32) ) _44122_ ( .A(_source_stream_conv2d_8_source_24_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_24_pat_stride_2), .S(_05709_), .Y(_23696_) );
  \$mux  #( .WIDTH(32) ) _44124_ ( .A(_source_stream_conv2d_8_source_24_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_24_pat_stride_1), .S(_05709_), .Y(_23697_) );
  \$mux  #( .WIDTH(32) ) _44126_ ( .A(_source_stream_conv2d_8_source_24_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_24_pat_stride_0), .S(_05709_), .Y(_23698_) );
  \$mux  #( .WIDTH(33) ) _44128_ ( .A(_source_stream_conv2d_8_source_24_pat_size_buf_3), .B(_source_stream_conv2d_8_source_24_pat_size_3), .S(_05709_), .Y(_23699_) );
  \$mux  #( .WIDTH(33) ) _44130_ ( .A(_source_stream_conv2d_8_source_24_pat_size_buf_2), .B(_source_stream_conv2d_8_source_24_pat_size_2), .S(_05709_), .Y(_23700_) );
  \$mux  #( .WIDTH(33) ) _44132_ ( .A(_source_stream_conv2d_8_source_24_pat_size_buf_1), .B(_source_stream_conv2d_8_source_24_pat_size_1), .S(_05709_), .Y(_23701_) );
  \$mux  #( .WIDTH(33) ) _44134_ ( .A(_source_stream_conv2d_8_source_24_pat_size_buf_0), .B(_source_stream_conv2d_8_source_24_pat_size_0), .S(_05709_), .Y(_23702_) );
  \$mux  #( .WIDTH(33) ) _44136_ ( .A(_source_stream_conv2d_8_source_24_pat_count_3), .B(_26103_), .S(_05709_), .Y(_23703_) );
  \$mux  #( .WIDTH(33) ) _44137_ ( .A(_23703_), .B(_26110_), .S(_05712_), .Y(_23704_) );
  \$mux  #( .WIDTH(33) ) _44138_ ( .A(_23704_), .B(_26111_), .S(_05713_), .Y(_23705_) );
  \$mux  #( .WIDTH(33) ) _44140_ ( .A(_source_stream_conv2d_8_source_24_pat_count_2), .B(_26102_), .S(_05709_), .Y(_23706_) );
  \$mux  #( .WIDTH(33) ) _44141_ ( .A(_23706_), .B(_26108_), .S(_05711_), .Y(_23707_) );
  \$mux  #( .WIDTH(33) ) _44142_ ( .A(_23707_), .B(_26109_), .S(_05712_), .Y(_23708_) );
  \$mux  #( .WIDTH(33) ) _44144_ ( .A(_source_stream_conv2d_8_source_24_pat_count_1), .B(_26101_), .S(_05709_), .Y(_23709_) );
  \$mux  #( .WIDTH(33) ) _44145_ ( .A(_23709_), .B(_26106_), .S(_05710_), .Y(_23710_) );
  \$mux  #( .WIDTH(33) ) _44146_ ( .A(_23710_), .B(_26107_), .S(_05711_), .Y(_23711_) );
  \$mux  #( .WIDTH(33) ) _44148_ ( .A(_source_stream_conv2d_8_source_24_pat_count_0), .B(_26100_), .S(_05709_), .Y(_23712_) );
  \$mux  #( .WIDTH(33) ) _44149_ ( .A(_26104_), .B(_23712_), .S(_05085_), .Y(_23713_) );
  \$mux  #( .WIDTH(33) ) _44150_ ( .A(_23713_), .B(_26105_), .S(_05710_), .Y(_23714_) );
  \$mux  #( .WIDTH(32) ) _44152_ ( .A(_source_stream_conv2d_8_source_24_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23715_) );
  \$mux  #( .WIDTH(32) ) _44154_ ( .A(_source_stream_conv2d_8_source_24_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23716_) );
  \$mux  #( .WIDTH(32) ) _44156_ ( .A(_source_stream_conv2d_8_source_24_pat_stride_1), .B(0), .S(_set_flag_538), .Y(_23717_) );
  \$mux  #( .WIDTH(32) ) _44158_ ( .A(_source_stream_conv2d_8_source_24_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23718_) );
  \$mux  #( .WIDTH(33) ) _44160_ ( .A(_source_stream_conv2d_8_source_24_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23719_) );
  \$mux  #( .WIDTH(33) ) _44162_ ( .A(_source_stream_conv2d_8_source_24_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23720_) );
  \$mux  #( .WIDTH(33) ) _44164_ ( .A(_source_stream_conv2d_8_source_24_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23721_) );
  \$mux  #( .WIDTH(33) ) _44166_ ( .A(_source_stream_conv2d_8_source_24_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23722_) );
  \$mux  #( .WIDTH(32) ) _44168_ ( .A(_source_stream_conv2d_8_source_24_pat_cur_offset_3), .B(0), .S(_05709_), .Y(_23723_) );
  \$mux  #( .WIDTH(32) ) _44169_ ( .A(_23723_), .B(_22177_), .S(_05712_), .Y(_23724_) );
  \$mux  #( .WIDTH(32) ) _44170_ ( .A(_23724_), .B(0), .S(_05713_), .Y(_23725_) );
  \$mux  #( .WIDTH(32) ) _44172_ ( .A(_source_stream_conv2d_8_source_24_pat_cur_offset_2), .B(0), .S(_05709_), .Y(_23726_) );
  \$mux  #( .WIDTH(32) ) _44173_ ( .A(_23726_), .B(_22176_), .S(_05711_), .Y(_23727_) );
  \$mux  #( .WIDTH(32) ) _44174_ ( .A(_23727_), .B(0), .S(_05712_), .Y(_23728_) );
  \$mux  #( .WIDTH(32) ) _44176_ ( .A(_source_stream_conv2d_8_source_24_pat_cur_offset_1), .B(0), .S(_05709_), .Y(_23729_) );
  \$mux  #( .WIDTH(32) ) _44177_ ( .A(_23729_), .B(_22175_), .S(_05710_), .Y(_23730_) );
  \$mux  #( .WIDTH(32) ) _44178_ ( .A(_23730_), .B(0), .S(_05711_), .Y(_23731_) );
  \$mux  #( .WIDTH(32) ) _44180_ ( .A(_source_stream_conv2d_8_source_24_pat_cur_offset_0), .B(0), .S(_05709_), .Y(_23732_) );
  \$mux  #( .WIDTH(32) ) _44181_ ( .A(_22174_), .B(_23732_), .S(_05085_), .Y(_23733_) );
  \$mux  #( .WIDTH(32) ) _44182_ ( .A(_23733_), .B(0), .S(_05710_), .Y(_23734_) );
  \$mux  #( .WIDTH(8) ) _44184_ ( .A(__variable_wdata_252), .B(_stream_conv2d_8_source_23_source_ram_rdata), .S(_stream_conv2d_8_source_23_source_ram_rvalid), .Y(_23735_) );
  \$mux  #( .WIDTH(32) ) _44186_ ( .A(_source_stream_conv2d_8_source_23_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_23_pat_stride_3), .S(_05704_), .Y(_23736_) );
  \$mux  #( .WIDTH(32) ) _44188_ ( .A(_source_stream_conv2d_8_source_23_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_23_pat_stride_2), .S(_05704_), .Y(_23737_) );
  \$mux  #( .WIDTH(32) ) _44190_ ( .A(_source_stream_conv2d_8_source_23_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_23_pat_stride_1), .S(_05704_), .Y(_23738_) );
  \$mux  #( .WIDTH(32) ) _44192_ ( .A(_source_stream_conv2d_8_source_23_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_23_pat_stride_0), .S(_05704_), .Y(_23739_) );
  \$mux  #( .WIDTH(33) ) _44194_ ( .A(_source_stream_conv2d_8_source_23_pat_size_buf_3), .B(_source_stream_conv2d_8_source_23_pat_size_3), .S(_05704_), .Y(_23740_) );
  \$mux  #( .WIDTH(33) ) _44196_ ( .A(_source_stream_conv2d_8_source_23_pat_size_buf_2), .B(_source_stream_conv2d_8_source_23_pat_size_2), .S(_05704_), .Y(_23741_) );
  \$mux  #( .WIDTH(33) ) _44198_ ( .A(_source_stream_conv2d_8_source_23_pat_size_buf_1), .B(_source_stream_conv2d_8_source_23_pat_size_1), .S(_05704_), .Y(_23742_) );
  \$mux  #( .WIDTH(33) ) _44200_ ( .A(_source_stream_conv2d_8_source_23_pat_size_buf_0), .B(_source_stream_conv2d_8_source_23_pat_size_0), .S(_05704_), .Y(_23743_) );
  \$mux  #( .WIDTH(33) ) _44202_ ( .A(_source_stream_conv2d_8_source_23_pat_count_3), .B(_26091_), .S(_05704_), .Y(_23744_) );
  \$mux  #( .WIDTH(33) ) _44203_ ( .A(_23744_), .B(_26098_), .S(_05707_), .Y(_23745_) );
  \$mux  #( .WIDTH(33) ) _44204_ ( .A(_23745_), .B(_26099_), .S(_05708_), .Y(_23746_) );
  \$mux  #( .WIDTH(33) ) _44206_ ( .A(_source_stream_conv2d_8_source_23_pat_count_2), .B(_26090_), .S(_05704_), .Y(_23747_) );
  \$mux  #( .WIDTH(33) ) _44207_ ( .A(_23747_), .B(_26096_), .S(_05706_), .Y(_23748_) );
  \$mux  #( .WIDTH(33) ) _44208_ ( .A(_23748_), .B(_26097_), .S(_05707_), .Y(_23749_) );
  \$mux  #( .WIDTH(33) ) _44210_ ( .A(_source_stream_conv2d_8_source_23_pat_count_1), .B(_26089_), .S(_05704_), .Y(_23750_) );
  \$mux  #( .WIDTH(33) ) _44211_ ( .A(_23750_), .B(_26094_), .S(_05705_), .Y(_23751_) );
  \$mux  #( .WIDTH(33) ) _44212_ ( .A(_23751_), .B(_26095_), .S(_05706_), .Y(_23752_) );
  \$mux  #( .WIDTH(33) ) _44214_ ( .A(_source_stream_conv2d_8_source_23_pat_count_0), .B(_26088_), .S(_05704_), .Y(_23753_) );
  \$mux  #( .WIDTH(33) ) _44215_ ( .A(_26092_), .B(_23753_), .S(_05087_), .Y(_23754_) );
  \$mux  #( .WIDTH(33) ) _44216_ ( .A(_23754_), .B(_26093_), .S(_05705_), .Y(_23755_) );
  \$mux  #( .WIDTH(32) ) _44218_ ( .A(_source_stream_conv2d_8_source_23_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23756_) );
  \$mux  #( .WIDTH(32) ) _44220_ ( .A(_source_stream_conv2d_8_source_23_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23757_) );
  \$mux  #( .WIDTH(32) ) _44222_ ( .A(_source_stream_conv2d_8_source_23_pat_stride_1), .B(0), .S(_set_flag_538), .Y(_23758_) );
  \$mux  #( .WIDTH(32) ) _44224_ ( .A(_source_stream_conv2d_8_source_23_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23759_) );
  \$mux  #( .WIDTH(33) ) _44226_ ( .A(_source_stream_conv2d_8_source_23_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23760_) );
  \$mux  #( .WIDTH(33) ) _44228_ ( .A(_source_stream_conv2d_8_source_23_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23761_) );
  \$mux  #( .WIDTH(33) ) _44230_ ( .A(_source_stream_conv2d_8_source_23_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23762_) );
  \$mux  #( .WIDTH(33) ) _44232_ ( .A(_source_stream_conv2d_8_source_23_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23763_) );
  \$mux  #( .WIDTH(32) ) _44234_ ( .A(_source_stream_conv2d_8_source_23_pat_cur_offset_3), .B(0), .S(_05704_), .Y(_23764_) );
  \$mux  #( .WIDTH(32) ) _44235_ ( .A(_23764_), .B(_22172_), .S(_05707_), .Y(_23765_) );
  \$mux  #( .WIDTH(32) ) _44236_ ( .A(_23765_), .B(0), .S(_05708_), .Y(_23766_) );
  \$mux  #( .WIDTH(32) ) _44238_ ( .A(_source_stream_conv2d_8_source_23_pat_cur_offset_2), .B(0), .S(_05704_), .Y(_23767_) );
  \$mux  #( .WIDTH(32) ) _44239_ ( .A(_23767_), .B(_22171_), .S(_05706_), .Y(_23768_) );
  \$mux  #( .WIDTH(32) ) _44240_ ( .A(_23768_), .B(0), .S(_05707_), .Y(_23769_) );
  \$mux  #( .WIDTH(32) ) _44242_ ( .A(_source_stream_conv2d_8_source_23_pat_cur_offset_1), .B(0), .S(_05704_), .Y(_23770_) );
  \$mux  #( .WIDTH(32) ) _44243_ ( .A(_23770_), .B(_22170_), .S(_05705_), .Y(_23771_) );
  \$mux  #( .WIDTH(32) ) _44244_ ( .A(_23771_), .B(0), .S(_05706_), .Y(_23772_) );
  \$mux  #( .WIDTH(32) ) _44246_ ( .A(_source_stream_conv2d_8_source_23_pat_cur_offset_0), .B(0), .S(_05704_), .Y(_23773_) );
  \$mux  #( .WIDTH(32) ) _44247_ ( .A(_22169_), .B(_23773_), .S(_05087_), .Y(_23774_) );
  \$mux  #( .WIDTH(32) ) _44248_ ( .A(_23774_), .B(0), .S(_05705_), .Y(_23775_) );
  \$mux  #( .WIDTH(8) ) _44250_ ( .A(__variable_wdata_251), .B(_stream_conv2d_8_source_22_source_ram_rdata), .S(_stream_conv2d_8_source_22_source_ram_rvalid), .Y(_23776_) );
  \$mux  #( .WIDTH(32) ) _44252_ ( .A(_source_stream_conv2d_8_source_22_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_22_pat_stride_3), .S(_05699_), .Y(_23777_) );
  \$mux  #( .WIDTH(32) ) _44254_ ( .A(_source_stream_conv2d_8_source_22_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_22_pat_stride_2), .S(_05699_), .Y(_23778_) );
  \$mux  #( .WIDTH(32) ) _44256_ ( .A(_source_stream_conv2d_8_source_22_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_22_pat_stride_1), .S(_05699_), .Y(_23779_) );
  \$mux  #( .WIDTH(32) ) _44258_ ( .A(_source_stream_conv2d_8_source_22_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_22_pat_stride_0), .S(_05699_), .Y(_23780_) );
  \$mux  #( .WIDTH(33) ) _44260_ ( .A(_source_stream_conv2d_8_source_22_pat_size_buf_3), .B(_source_stream_conv2d_8_source_22_pat_size_3), .S(_05699_), .Y(_23781_) );
  \$mux  #( .WIDTH(33) ) _44262_ ( .A(_source_stream_conv2d_8_source_22_pat_size_buf_2), .B(_source_stream_conv2d_8_source_22_pat_size_2), .S(_05699_), .Y(_23782_) );
  \$mux  #( .WIDTH(33) ) _44264_ ( .A(_source_stream_conv2d_8_source_22_pat_size_buf_1), .B(_source_stream_conv2d_8_source_22_pat_size_1), .S(_05699_), .Y(_23783_) );
  \$mux  #( .WIDTH(33) ) _44266_ ( .A(_source_stream_conv2d_8_source_22_pat_size_buf_0), .B(_source_stream_conv2d_8_source_22_pat_size_0), .S(_05699_), .Y(_23784_) );
  \$mux  #( .WIDTH(33) ) _44268_ ( .A(_source_stream_conv2d_8_source_22_pat_count_3), .B(_26079_), .S(_05699_), .Y(_23785_) );
  \$mux  #( .WIDTH(33) ) _44269_ ( .A(_23785_), .B(_26086_), .S(_05702_), .Y(_23786_) );
  \$mux  #( .WIDTH(33) ) _44270_ ( .A(_23786_), .B(_26087_), .S(_05703_), .Y(_23787_) );
  \$mux  #( .WIDTH(33) ) _44272_ ( .A(_source_stream_conv2d_8_source_22_pat_count_2), .B(_26078_), .S(_05699_), .Y(_23788_) );
  \$mux  #( .WIDTH(33) ) _44273_ ( .A(_23788_), .B(_26084_), .S(_05701_), .Y(_23789_) );
  \$mux  #( .WIDTH(33) ) _44274_ ( .A(_23789_), .B(_26085_), .S(_05702_), .Y(_23790_) );
  \$mux  #( .WIDTH(33) ) _44276_ ( .A(_source_stream_conv2d_8_source_22_pat_count_1), .B(_26077_), .S(_05699_), .Y(_23791_) );
  \$mux  #( .WIDTH(33) ) _44277_ ( .A(_23791_), .B(_26082_), .S(_05700_), .Y(_23792_) );
  \$mux  #( .WIDTH(33) ) _44278_ ( .A(_23792_), .B(_26083_), .S(_05701_), .Y(_23793_) );
  \$mux  #( .WIDTH(33) ) _44280_ ( .A(_source_stream_conv2d_8_source_22_pat_count_0), .B(_26076_), .S(_05699_), .Y(_23794_) );
  \$mux  #( .WIDTH(33) ) _44281_ ( .A(_26080_), .B(_23794_), .S(_05089_), .Y(_23795_) );
  \$mux  #( .WIDTH(33) ) _44282_ ( .A(_23795_), .B(_26081_), .S(_05700_), .Y(_23796_) );
  \$mux  #( .WIDTH(32) ) _44284_ ( .A(_source_stream_conv2d_8_source_22_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23797_) );
  \$mux  #( .WIDTH(32) ) _44286_ ( .A(_source_stream_conv2d_8_source_22_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23798_) );
  \$mux  #( .WIDTH(32) ) _44288_ ( .A(_source_stream_conv2d_8_source_22_pat_stride_1), .B(0), .S(_set_flag_538), .Y(_23799_) );
  \$mux  #( .WIDTH(32) ) _44290_ ( .A(_source_stream_conv2d_8_source_22_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23800_) );
  \$mux  #( .WIDTH(33) ) _44292_ ( .A(_source_stream_conv2d_8_source_22_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23801_) );
  \$mux  #( .WIDTH(33) ) _44294_ ( .A(_source_stream_conv2d_8_source_22_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23802_) );
  \$mux  #( .WIDTH(33) ) _44296_ ( .A(_source_stream_conv2d_8_source_22_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23803_) );
  \$mux  #( .WIDTH(33) ) _44298_ ( .A(_source_stream_conv2d_8_source_22_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23804_) );
  \$mux  #( .WIDTH(32) ) _44300_ ( .A(_source_stream_conv2d_8_source_22_pat_cur_offset_3), .B(0), .S(_05699_), .Y(_23805_) );
  \$mux  #( .WIDTH(32) ) _44301_ ( .A(_23805_), .B(_22167_), .S(_05702_), .Y(_23806_) );
  \$mux  #( .WIDTH(32) ) _44302_ ( .A(_23806_), .B(0), .S(_05703_), .Y(_23807_) );
  \$mux  #( .WIDTH(32) ) _44304_ ( .A(_source_stream_conv2d_8_source_22_pat_cur_offset_2), .B(0), .S(_05699_), .Y(_23808_) );
  \$mux  #( .WIDTH(32) ) _44305_ ( .A(_23808_), .B(_22166_), .S(_05701_), .Y(_23809_) );
  \$mux  #( .WIDTH(32) ) _44306_ ( .A(_23809_), .B(0), .S(_05702_), .Y(_23810_) );
  \$mux  #( .WIDTH(32) ) _44308_ ( .A(_source_stream_conv2d_8_source_22_pat_cur_offset_1), .B(0), .S(_05699_), .Y(_23811_) );
  \$mux  #( .WIDTH(32) ) _44309_ ( .A(_23811_), .B(_22165_), .S(_05700_), .Y(_23812_) );
  \$mux  #( .WIDTH(32) ) _44310_ ( .A(_23812_), .B(0), .S(_05701_), .Y(_23813_) );
  \$mux  #( .WIDTH(32) ) _44312_ ( .A(_source_stream_conv2d_8_source_22_pat_cur_offset_0), .B(0), .S(_05699_), .Y(_23814_) );
  \$mux  #( .WIDTH(32) ) _44313_ ( .A(_22164_), .B(_23814_), .S(_05089_), .Y(_23815_) );
  \$mux  #( .WIDTH(32) ) _44314_ ( .A(_23815_), .B(0), .S(_05700_), .Y(_23816_) );
  \$mux  #( .WIDTH(8) ) _44316_ ( .A(__variable_wdata_250), .B(_stream_conv2d_8_source_21_source_ram_rdata), .S(_stream_conv2d_8_source_21_source_ram_rvalid), .Y(_23817_) );
  \$mux  #( .WIDTH(32) ) _44318_ ( .A(_source_stream_conv2d_8_source_21_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_21_pat_stride_3), .S(_05694_), .Y(_23818_) );
  \$mux  #( .WIDTH(32) ) _44320_ ( .A(_source_stream_conv2d_8_source_21_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_21_pat_stride_2), .S(_05694_), .Y(_23819_) );
  \$mux  #( .WIDTH(32) ) _44322_ ( .A(_source_stream_conv2d_8_source_21_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_21_pat_stride_1), .S(_05694_), .Y(_23820_) );
  \$mux  #( .WIDTH(32) ) _44324_ ( .A(_source_stream_conv2d_8_source_21_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_21_pat_stride_0), .S(_05694_), .Y(_23821_) );
  \$mux  #( .WIDTH(33) ) _44326_ ( .A(_source_stream_conv2d_8_source_21_pat_size_buf_3), .B(_source_stream_conv2d_8_source_21_pat_size_3), .S(_05694_), .Y(_23822_) );
  \$mux  #( .WIDTH(33) ) _44328_ ( .A(_source_stream_conv2d_8_source_21_pat_size_buf_2), .B(_source_stream_conv2d_8_source_21_pat_size_2), .S(_05694_), .Y(_23823_) );
  \$mux  #( .WIDTH(33) ) _44330_ ( .A(_source_stream_conv2d_8_source_21_pat_size_buf_1), .B(_source_stream_conv2d_8_source_21_pat_size_1), .S(_05694_), .Y(_23824_) );
  \$mux  #( .WIDTH(33) ) _44332_ ( .A(_source_stream_conv2d_8_source_21_pat_size_buf_0), .B(_source_stream_conv2d_8_source_21_pat_size_0), .S(_05694_), .Y(_23825_) );
  \$mux  #( .WIDTH(33) ) _44334_ ( .A(_source_stream_conv2d_8_source_21_pat_count_3), .B(_26067_), .S(_05694_), .Y(_23826_) );
  \$mux  #( .WIDTH(33) ) _44335_ ( .A(_23826_), .B(_26074_), .S(_05697_), .Y(_23827_) );
  \$mux  #( .WIDTH(33) ) _44336_ ( .A(_23827_), .B(_26075_), .S(_05698_), .Y(_23828_) );
  \$mux  #( .WIDTH(33) ) _44338_ ( .A(_source_stream_conv2d_8_source_21_pat_count_2), .B(_26066_), .S(_05694_), .Y(_23829_) );
  \$mux  #( .WIDTH(33) ) _44339_ ( .A(_23829_), .B(_26072_), .S(_05696_), .Y(_23830_) );
  \$mux  #( .WIDTH(33) ) _44340_ ( .A(_23830_), .B(_26073_), .S(_05697_), .Y(_23831_) );
  \$mux  #( .WIDTH(33) ) _44342_ ( .A(_source_stream_conv2d_8_source_21_pat_count_1), .B(_26065_), .S(_05694_), .Y(_23832_) );
  \$mux  #( .WIDTH(33) ) _44343_ ( .A(_23832_), .B(_26070_), .S(_05695_), .Y(_23833_) );
  \$mux  #( .WIDTH(33) ) _44344_ ( .A(_23833_), .B(_26071_), .S(_05696_), .Y(_23834_) );
  \$mux  #( .WIDTH(33) ) _44346_ ( .A(_source_stream_conv2d_8_source_21_pat_count_0), .B(_26064_), .S(_05694_), .Y(_23835_) );
  \$mux  #( .WIDTH(33) ) _44347_ ( .A(_26068_), .B(_23835_), .S(_05091_), .Y(_23836_) );
  \$mux  #( .WIDTH(33) ) _44348_ ( .A(_23836_), .B(_26069_), .S(_05695_), .Y(_23837_) );
  \$mux  #( .WIDTH(32) ) _44350_ ( .A(_source_stream_conv2d_8_source_21_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23838_) );
  \$mux  #( .WIDTH(32) ) _44352_ ( .A(_source_stream_conv2d_8_source_21_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23839_) );
  \$mux  #( .WIDTH(32) ) _44354_ ( .A(_source_stream_conv2d_8_source_21_pat_stride_1), .B(0), .S(_set_flag_538), .Y(_23840_) );
  \$mux  #( .WIDTH(32) ) _44356_ ( .A(_source_stream_conv2d_8_source_21_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23841_) );
  \$mux  #( .WIDTH(33) ) _44358_ ( .A(_source_stream_conv2d_8_source_21_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23842_) );
  \$mux  #( .WIDTH(33) ) _44360_ ( .A(_source_stream_conv2d_8_source_21_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23843_) );
  \$mux  #( .WIDTH(33) ) _44362_ ( .A(_source_stream_conv2d_8_source_21_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23844_) );
  \$mux  #( .WIDTH(33) ) _44364_ ( .A(_source_stream_conv2d_8_source_21_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23845_) );
  \$mux  #( .WIDTH(32) ) _44366_ ( .A(_source_stream_conv2d_8_source_21_pat_cur_offset_3), .B(0), .S(_05694_), .Y(_23846_) );
  \$mux  #( .WIDTH(32) ) _44367_ ( .A(_23846_), .B(_22162_), .S(_05697_), .Y(_23847_) );
  \$mux  #( .WIDTH(32) ) _44368_ ( .A(_23847_), .B(0), .S(_05698_), .Y(_23848_) );
  \$mux  #( .WIDTH(32) ) _44370_ ( .A(_source_stream_conv2d_8_source_21_pat_cur_offset_2), .B(0), .S(_05694_), .Y(_23849_) );
  \$mux  #( .WIDTH(32) ) _44371_ ( .A(_23849_), .B(_22161_), .S(_05696_), .Y(_23850_) );
  \$mux  #( .WIDTH(32) ) _44372_ ( .A(_23850_), .B(0), .S(_05697_), .Y(_23851_) );
  \$mux  #( .WIDTH(32) ) _44374_ ( .A(_source_stream_conv2d_8_source_21_pat_cur_offset_1), .B(0), .S(_05694_), .Y(_23852_) );
  \$mux  #( .WIDTH(32) ) _44375_ ( .A(_23852_), .B(_22160_), .S(_05695_), .Y(_23853_) );
  \$mux  #( .WIDTH(32) ) _44376_ ( .A(_23853_), .B(0), .S(_05696_), .Y(_23854_) );
  \$mux  #( .WIDTH(32) ) _44378_ ( .A(_source_stream_conv2d_8_source_21_pat_cur_offset_0), .B(0), .S(_05694_), .Y(_23855_) );
  \$mux  #( .WIDTH(32) ) _44379_ ( .A(_22159_), .B(_23855_), .S(_05091_), .Y(_23856_) );
  \$mux  #( .WIDTH(32) ) _44380_ ( .A(_23856_), .B(0), .S(_05695_), .Y(_23857_) );
  \$mux  #( .WIDTH(8) ) _44382_ ( .A(__variable_wdata_249), .B(_stream_conv2d_8_source_20_source_ram_rdata), .S(_stream_conv2d_8_source_20_source_ram_rvalid), .Y(_23858_) );
  \$mux  #( .WIDTH(32) ) _44384_ ( .A(_source_stream_conv2d_8_source_20_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_20_pat_stride_3), .S(_05689_), .Y(_23859_) );
  \$mux  #( .WIDTH(32) ) _44386_ ( .A(_source_stream_conv2d_8_source_20_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_20_pat_stride_2), .S(_05689_), .Y(_23860_) );
  \$mux  #( .WIDTH(32) ) _44388_ ( .A(_source_stream_conv2d_8_source_20_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_20_pat_stride_1), .S(_05689_), .Y(_23861_) );
  \$mux  #( .WIDTH(32) ) _44390_ ( .A(_source_stream_conv2d_8_source_20_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_20_pat_stride_0), .S(_05689_), .Y(_23862_) );
  \$mux  #( .WIDTH(33) ) _44392_ ( .A(_source_stream_conv2d_8_source_20_pat_size_buf_3), .B(_source_stream_conv2d_8_source_20_pat_size_3), .S(_05689_), .Y(_23863_) );
  \$mux  #( .WIDTH(33) ) _44394_ ( .A(_source_stream_conv2d_8_source_20_pat_size_buf_2), .B(_source_stream_conv2d_8_source_20_pat_size_2), .S(_05689_), .Y(_23864_) );
  \$mux  #( .WIDTH(33) ) _44396_ ( .A(_source_stream_conv2d_8_source_20_pat_size_buf_1), .B(_source_stream_conv2d_8_source_20_pat_size_1), .S(_05689_), .Y(_23865_) );
  \$mux  #( .WIDTH(33) ) _44398_ ( .A(_source_stream_conv2d_8_source_20_pat_size_buf_0), .B(_source_stream_conv2d_8_source_20_pat_size_0), .S(_05689_), .Y(_23866_) );
  \$mux  #( .WIDTH(33) ) _44400_ ( .A(_source_stream_conv2d_8_source_20_pat_count_3), .B(_26055_), .S(_05689_), .Y(_23867_) );
  \$mux  #( .WIDTH(33) ) _44401_ ( .A(_23867_), .B(_26062_), .S(_05692_), .Y(_23868_) );
  \$mux  #( .WIDTH(33) ) _44402_ ( .A(_23868_), .B(_26063_), .S(_05693_), .Y(_23869_) );
  \$mux  #( .WIDTH(33) ) _44404_ ( .A(_source_stream_conv2d_8_source_20_pat_count_2), .B(_26054_), .S(_05689_), .Y(_23870_) );
  \$mux  #( .WIDTH(33) ) _44405_ ( .A(_23870_), .B(_26060_), .S(_05691_), .Y(_23871_) );
  \$mux  #( .WIDTH(33) ) _44406_ ( .A(_23871_), .B(_26061_), .S(_05692_), .Y(_23872_) );
  \$mux  #( .WIDTH(33) ) _44408_ ( .A(_source_stream_conv2d_8_source_20_pat_count_1), .B(_26053_), .S(_05689_), .Y(_23873_) );
  \$mux  #( .WIDTH(33) ) _44409_ ( .A(_23873_), .B(_26058_), .S(_05690_), .Y(_23874_) );
  \$mux  #( .WIDTH(33) ) _44410_ ( .A(_23874_), .B(_26059_), .S(_05691_), .Y(_23875_) );
  \$mux  #( .WIDTH(33) ) _44412_ ( .A(_source_stream_conv2d_8_source_20_pat_count_0), .B(_26052_), .S(_05689_), .Y(_23876_) );
  \$mux  #( .WIDTH(33) ) _44413_ ( .A(_26056_), .B(_23876_), .S(_05093_), .Y(_23877_) );
  \$mux  #( .WIDTH(33) ) _44414_ ( .A(_23877_), .B(_26057_), .S(_05690_), .Y(_23878_) );
  \$mux  #( .WIDTH(32) ) _44416_ ( .A(_source_stream_conv2d_8_source_20_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23879_) );
  \$mux  #( .WIDTH(32) ) _44418_ ( .A(_source_stream_conv2d_8_source_20_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23880_) );
  \$mux  #( .WIDTH(32) ) _44420_ ( .A(_source_stream_conv2d_8_source_20_pat_stride_1), .B(0), .S(_set_flag_538), .Y(_23881_) );
  \$mux  #( .WIDTH(32) ) _44422_ ( .A(_source_stream_conv2d_8_source_20_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23882_) );
  \$mux  #( .WIDTH(33) ) _44424_ ( .A(_source_stream_conv2d_8_source_20_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23883_) );
  \$mux  #( .WIDTH(33) ) _44426_ ( .A(_source_stream_conv2d_8_source_20_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23884_) );
  \$mux  #( .WIDTH(33) ) _44428_ ( .A(_source_stream_conv2d_8_source_20_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23885_) );
  \$mux  #( .WIDTH(33) ) _44430_ ( .A(_source_stream_conv2d_8_source_20_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23886_) );
  \$mux  #( .WIDTH(32) ) _44432_ ( .A(_source_stream_conv2d_8_source_20_pat_cur_offset_3), .B(0), .S(_05689_), .Y(_23887_) );
  \$mux  #( .WIDTH(32) ) _44433_ ( .A(_23887_), .B(_22157_), .S(_05692_), .Y(_23888_) );
  \$mux  #( .WIDTH(32) ) _44434_ ( .A(_23888_), .B(0), .S(_05693_), .Y(_23889_) );
  \$mux  #( .WIDTH(32) ) _44436_ ( .A(_source_stream_conv2d_8_source_20_pat_cur_offset_2), .B(0), .S(_05689_), .Y(_23890_) );
  \$mux  #( .WIDTH(32) ) _44437_ ( .A(_23890_), .B(_22156_), .S(_05691_), .Y(_23891_) );
  \$mux  #( .WIDTH(32) ) _44438_ ( .A(_23891_), .B(0), .S(_05692_), .Y(_23892_) );
  \$mux  #( .WIDTH(32) ) _44440_ ( .A(_source_stream_conv2d_8_source_20_pat_cur_offset_1), .B(0), .S(_05689_), .Y(_23893_) );
  \$mux  #( .WIDTH(32) ) _44441_ ( .A(_23893_), .B(_22155_), .S(_05690_), .Y(_23894_) );
  \$mux  #( .WIDTH(32) ) _44442_ ( .A(_23894_), .B(0), .S(_05691_), .Y(_23895_) );
  \$mux  #( .WIDTH(32) ) _44444_ ( .A(_source_stream_conv2d_8_source_20_pat_cur_offset_0), .B(0), .S(_05689_), .Y(_23896_) );
  \$mux  #( .WIDTH(32) ) _44445_ ( .A(_22154_), .B(_23896_), .S(_05093_), .Y(_23897_) );
  \$mux  #( .WIDTH(32) ) _44446_ ( .A(_23897_), .B(0), .S(_05690_), .Y(_23898_) );
  \$mux  #( .WIDTH(8) ) _44448_ ( .A(__variable_wdata_248), .B(_stream_conv2d_8_source_19_source_ram_rdata), .S(_stream_conv2d_8_source_19_source_ram_rvalid), .Y(_23899_) );
  \$mux  #( .WIDTH(32) ) _44450_ ( .A(_source_stream_conv2d_8_source_19_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_19_pat_stride_3), .S(_05684_), .Y(_23900_) );
  \$mux  #( .WIDTH(32) ) _44452_ ( .A(_source_stream_conv2d_8_source_19_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_19_pat_stride_2), .S(_05684_), .Y(_23901_) );
  \$mux  #( .WIDTH(32) ) _44454_ ( .A(_source_stream_conv2d_8_source_19_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_19_pat_stride_1), .S(_05684_), .Y(_23902_) );
  \$mux  #( .WIDTH(32) ) _44456_ ( .A(_source_stream_conv2d_8_source_19_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_19_pat_stride_0), .S(_05684_), .Y(_23903_) );
  \$mux  #( .WIDTH(33) ) _44458_ ( .A(_source_stream_conv2d_8_source_19_pat_size_buf_3), .B(_source_stream_conv2d_8_source_19_pat_size_3), .S(_05684_), .Y(_23904_) );
  \$mux  #( .WIDTH(33) ) _44460_ ( .A(_source_stream_conv2d_8_source_19_pat_size_buf_2), .B(_source_stream_conv2d_8_source_19_pat_size_2), .S(_05684_), .Y(_23905_) );
  \$mux  #( .WIDTH(33) ) _44462_ ( .A(_source_stream_conv2d_8_source_19_pat_size_buf_1), .B(_source_stream_conv2d_8_source_19_pat_size_1), .S(_05684_), .Y(_23906_) );
  \$mux  #( .WIDTH(33) ) _44464_ ( .A(_source_stream_conv2d_8_source_19_pat_size_buf_0), .B(_source_stream_conv2d_8_source_19_pat_size_0), .S(_05684_), .Y(_23907_) );
  \$mux  #( .WIDTH(33) ) _44466_ ( .A(_source_stream_conv2d_8_source_19_pat_count_3), .B(_26043_), .S(_05684_), .Y(_23908_) );
  \$mux  #( .WIDTH(33) ) _44467_ ( .A(_23908_), .B(_26050_), .S(_05687_), .Y(_23909_) );
  \$mux  #( .WIDTH(33) ) _44468_ ( .A(_23909_), .B(_26051_), .S(_05688_), .Y(_23910_) );
  \$mux  #( .WIDTH(33) ) _44470_ ( .A(_source_stream_conv2d_8_source_19_pat_count_2), .B(_26042_), .S(_05684_), .Y(_23911_) );
  \$mux  #( .WIDTH(33) ) _44471_ ( .A(_23911_), .B(_26048_), .S(_05686_), .Y(_23912_) );
  \$mux  #( .WIDTH(33) ) _44472_ ( .A(_23912_), .B(_26049_), .S(_05687_), .Y(_23913_) );
  \$mux  #( .WIDTH(33) ) _44474_ ( .A(_source_stream_conv2d_8_source_19_pat_count_1), .B(_26041_), .S(_05684_), .Y(_23914_) );
  \$mux  #( .WIDTH(33) ) _44475_ ( .A(_23914_), .B(_26046_), .S(_05685_), .Y(_23915_) );
  \$mux  #( .WIDTH(33) ) _44476_ ( .A(_23915_), .B(_26047_), .S(_05686_), .Y(_23916_) );
  \$mux  #( .WIDTH(33) ) _44478_ ( .A(_source_stream_conv2d_8_source_19_pat_count_0), .B(_26040_), .S(_05684_), .Y(_23917_) );
  \$mux  #( .WIDTH(33) ) _44479_ ( .A(_26044_), .B(_23917_), .S(_05095_), .Y(_23918_) );
  \$mux  #( .WIDTH(33) ) _44480_ ( .A(_23918_), .B(_26045_), .S(_05685_), .Y(_23919_) );
  \$mux  #( .WIDTH(32) ) _44482_ ( .A(_source_stream_conv2d_8_source_19_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23920_) );
  \$mux  #( .WIDTH(32) ) _44484_ ( .A(_source_stream_conv2d_8_source_19_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23921_) );
  \$mux  #( .WIDTH(32) ) _44486_ ( .A(_source_stream_conv2d_8_source_19_pat_stride_1), .B(0), .S(_set_flag_538), .Y(_23922_) );
  \$mux  #( .WIDTH(32) ) _44488_ ( .A(_source_stream_conv2d_8_source_19_pat_stride_0), .B(1), .S(_set_flag_538), .Y(_23923_) );
  \$mux  #( .WIDTH(33) ) _44490_ ( .A(_source_stream_conv2d_8_source_19_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23924_) );
  \$mux  #( .WIDTH(33) ) _44492_ ( .A(_source_stream_conv2d_8_source_19_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23925_) );
  \$mux  #( .WIDTH(33) ) _44494_ ( .A(_source_stream_conv2d_8_source_19_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23926_) );
  \$mux  #( .WIDTH(33) ) _44496_ ( .A(_source_stream_conv2d_8_source_19_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23927_) );
  \$mux  #( .WIDTH(32) ) _44498_ ( .A(_source_stream_conv2d_8_source_19_pat_cur_offset_3), .B(0), .S(_05684_), .Y(_23928_) );
  \$mux  #( .WIDTH(32) ) _44499_ ( .A(_23928_), .B(_22152_), .S(_05687_), .Y(_23929_) );
  \$mux  #( .WIDTH(32) ) _44500_ ( .A(_23929_), .B(0), .S(_05688_), .Y(_23930_) );
  \$mux  #( .WIDTH(32) ) _44502_ ( .A(_source_stream_conv2d_8_source_19_pat_cur_offset_2), .B(0), .S(_05684_), .Y(_23931_) );
  \$mux  #( .WIDTH(32) ) _44503_ ( .A(_23931_), .B(_22151_), .S(_05686_), .Y(_23932_) );
  \$mux  #( .WIDTH(32) ) _44504_ ( .A(_23932_), .B(0), .S(_05687_), .Y(_23933_) );
  \$mux  #( .WIDTH(32) ) _44506_ ( .A(_source_stream_conv2d_8_source_19_pat_cur_offset_1), .B(0), .S(_05684_), .Y(_23934_) );
  \$mux  #( .WIDTH(32) ) _44507_ ( .A(_23934_), .B(_22150_), .S(_05685_), .Y(_23935_) );
  \$mux  #( .WIDTH(32) ) _44508_ ( .A(_23935_), .B(0), .S(_05686_), .Y(_23936_) );
  \$mux  #( .WIDTH(32) ) _44510_ ( .A(_source_stream_conv2d_8_source_19_pat_cur_offset_0), .B(0), .S(_05684_), .Y(_23937_) );
  \$mux  #( .WIDTH(32) ) _44511_ ( .A(_22149_), .B(_23937_), .S(_05095_), .Y(_23938_) );
  \$mux  #( .WIDTH(32) ) _44512_ ( .A(_23938_), .B(0), .S(_05685_), .Y(_23939_) );
  \$mux  #( .WIDTH(4) ) _44514_ ( .A(__variable_wdata_246), .B(_stream_conv2d_8_constant_17_next_constant_data), .S(_stream_conv2d_8_start), .Y(_23940_) );
  \$mux  #( .WIDTH(1) ) _44516_ ( .A(__variable_wdata_245), .B(_stream_conv2d_8_constant_16_next_constant_data), .S(_stream_conv2d_8_start), .Y(_23941_) );
  \$mux  #( .WIDTH(1) ) _44518_ ( .A(__variable_wdata_244), .B(_stream_conv2d_8_constant_15_next_constant_data), .S(_stream_conv2d_8_start), .Y(_23942_) );
  \$mux  #( .WIDTH(8) ) _44520_ ( .A(__variable_wdata_238), .B(_stream_conv2d_8_source_14_source_empty_data), .S(_stream_conv2d_8_start), .Y(_23943_) );
  \$mux  #( .WIDTH(8) ) _44522_ ( .A(__variable_wdata_231), .B(_stream_conv2d_8_source_12_source_empty_data), .S(_stream_conv2d_8_start), .Y(_23944_) );
  \$mux  #( .WIDTH(8) ) _44524_ ( .A(__variable_wdata_224), .B(_stream_conv2d_8_source_10_source_empty_data), .S(_stream_conv2d_8_start), .Y(_23945_) );
  \$mux  #( .WIDTH(8) ) _44526_ ( .A(__variable_wdata_217), .B(_stream_conv2d_8_source_8_source_ram_rdata), .S(_stream_conv2d_8_source_8_source_ram_rvalid), .Y(_23946_) );
  \$mux  #( .WIDTH(32) ) _44528_ ( .A(_source_stream_conv2d_8_source_8_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_8_pat_stride_3), .S(_05679_), .Y(_23947_) );
  \$mux  #( .WIDTH(32) ) _44530_ ( .A(_source_stream_conv2d_8_source_8_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_8_pat_stride_2), .S(_05679_), .Y(_23948_) );
  \$mux  #( .WIDTH(32) ) _44532_ ( .A(_source_stream_conv2d_8_source_8_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_8_pat_stride_1), .S(_05679_), .Y(_23949_) );
  \$mux  #( .WIDTH(32) ) _44534_ ( .A(_source_stream_conv2d_8_source_8_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_8_pat_stride_0), .S(_05679_), .Y(_23950_) );
  \$mux  #( .WIDTH(33) ) _44536_ ( .A(_source_stream_conv2d_8_source_8_pat_size_buf_3), .B(_source_stream_conv2d_8_source_8_pat_size_3), .S(_05679_), .Y(_23951_) );
  \$mux  #( .WIDTH(33) ) _44538_ ( .A(_source_stream_conv2d_8_source_8_pat_size_buf_2), .B(_source_stream_conv2d_8_source_8_pat_size_2), .S(_05679_), .Y(_23952_) );
  \$mux  #( .WIDTH(33) ) _44540_ ( .A(_source_stream_conv2d_8_source_8_pat_size_buf_1), .B(_source_stream_conv2d_8_source_8_pat_size_1), .S(_05679_), .Y(_23953_) );
  \$mux  #( .WIDTH(33) ) _44542_ ( .A(_source_stream_conv2d_8_source_8_pat_size_buf_0), .B(_source_stream_conv2d_8_source_8_pat_size_0), .S(_05679_), .Y(_23954_) );
  \$mux  #( .WIDTH(33) ) _44544_ ( .A(_source_stream_conv2d_8_source_8_pat_count_3), .B(_26031_), .S(_05679_), .Y(_23955_) );
  \$mux  #( .WIDTH(33) ) _44545_ ( .A(_23955_), .B(_26038_), .S(_05682_), .Y(_23956_) );
  \$mux  #( .WIDTH(33) ) _44546_ ( .A(_23956_), .B(_26039_), .S(_05683_), .Y(_23957_) );
  \$mux  #( .WIDTH(33) ) _44548_ ( .A(_source_stream_conv2d_8_source_8_pat_count_2), .B(_26030_), .S(_05679_), .Y(_23958_) );
  \$mux  #( .WIDTH(33) ) _44549_ ( .A(_23958_), .B(_26036_), .S(_05681_), .Y(_23959_) );
  \$mux  #( .WIDTH(33) ) _44550_ ( .A(_23959_), .B(_26037_), .S(_05682_), .Y(_23960_) );
  \$mux  #( .WIDTH(33) ) _44552_ ( .A(_source_stream_conv2d_8_source_8_pat_count_1), .B(_26029_), .S(_05679_), .Y(_23961_) );
  \$mux  #( .WIDTH(33) ) _44553_ ( .A(_23961_), .B(_26034_), .S(_05680_), .Y(_23962_) );
  \$mux  #( .WIDTH(33) ) _44554_ ( .A(_23962_), .B(_26035_), .S(_05681_), .Y(_23963_) );
  \$mux  #( .WIDTH(33) ) _44556_ ( .A(_source_stream_conv2d_8_source_8_pat_count_0), .B(_26028_), .S(_05679_), .Y(_23964_) );
  \$mux  #( .WIDTH(33) ) _44557_ ( .A(_26032_), .B(_23964_), .S(_05097_), .Y(_23965_) );
  \$mux  #( .WIDTH(33) ) _44558_ ( .A(_23965_), .B(_26033_), .S(_05680_), .Y(_23966_) );
  \$mux  #( .WIDTH(32) ) _44560_ ( .A(_source_stream_conv2d_8_source_8_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_23967_) );
  \$mux  #( .WIDTH(32) ) _44562_ ( .A(_source_stream_conv2d_8_source_8_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_23968_) );
  \$mux  #( .WIDTH(32) ) _44564_ ( .A(_source_stream_conv2d_8_source_8_pat_stride_1), .B(0), .S(_set_flag_538), .Y(_23969_) );
  \$mux  #( .WIDTH(32) ) _44566_ ( .A(_source_stream_conv2d_8_source_8_pat_stride_0), .B(0), .S(_set_flag_538), .Y(_23970_) );
  \$mux  #( .WIDTH(33) ) _44568_ ( .A(_source_stream_conv2d_8_source_8_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_23971_) );
  \$mux  #( .WIDTH(33) ) _44570_ ( .A(_source_stream_conv2d_8_source_8_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_23972_) );
  \$mux  #( .WIDTH(33) ) _44572_ ( .A(_source_stream_conv2d_8_source_8_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_23973_) );
  \$mux  #( .WIDTH(33) ) _44574_ ( .A(_source_stream_conv2d_8_source_8_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_23974_) );
  \$mux  #( .WIDTH(32) ) _44576_ ( .A(_source_stream_conv2d_8_source_8_pat_cur_offset_3), .B(0), .S(_05679_), .Y(_23975_) );
  \$mux  #( .WIDTH(32) ) _44577_ ( .A(_23975_), .B(_22147_), .S(_05682_), .Y(_23976_) );
  \$mux  #( .WIDTH(32) ) _44578_ ( .A(_23976_), .B(0), .S(_05683_), .Y(_23977_) );
  \$mux  #( .WIDTH(32) ) _44580_ ( .A(_source_stream_conv2d_8_source_8_pat_cur_offset_2), .B(0), .S(_05679_), .Y(_23978_) );
  \$mux  #( .WIDTH(32) ) _44581_ ( .A(_23978_), .B(_22146_), .S(_05681_), .Y(_23979_) );
  \$mux  #( .WIDTH(32) ) _44582_ ( .A(_23979_), .B(0), .S(_05682_), .Y(_23980_) );
  \$mux  #( .WIDTH(32) ) _44584_ ( .A(_source_stream_conv2d_8_source_8_pat_cur_offset_1), .B(0), .S(_05679_), .Y(_23981_) );
  \$mux  #( .WIDTH(32) ) _44585_ ( .A(_23981_), .B(_22145_), .S(_05680_), .Y(_23982_) );
  \$mux  #( .WIDTH(32) ) _44586_ ( .A(_23982_), .B(0), .S(_05681_), .Y(_23983_) );
  \$mux  #( .WIDTH(32) ) _44588_ ( .A(_source_stream_conv2d_8_source_8_pat_cur_offset_0), .B(0), .S(_05679_), .Y(_23984_) );
  \$mux  #( .WIDTH(32) ) _44589_ ( .A(_22144_), .B(_23984_), .S(_05097_), .Y(_23985_) );
  \$mux  #( .WIDTH(32) ) _44590_ ( .A(_23985_), .B(0), .S(_05680_), .Y(_23986_) );
  \$mux  #( .WIDTH(32) ) _44592_ ( .A(__variable_wdata_210), .B(_stream_conv2d_8_source_6_source_ram_rdata), .S(_stream_conv2d_8_source_6_source_ram_rvalid), .Y(_23987_) );
  \$mux  #( .WIDTH(32) ) _44594_ ( .A(_source_stream_conv2d_8_source_6_pat_stride_buf_3), .B(_source_stream_conv2d_8_source_6_pat_stride_3), .S(_05674_), .Y(_23988_) );
  \$mux  #( .WIDTH(32) ) _44596_ ( .A(_source_stream_conv2d_8_source_6_pat_stride_buf_2), .B(_source_stream_conv2d_8_source_6_pat_stride_2), .S(_05674_), .Y(_23989_) );
  \$mux  #( .WIDTH(32) ) _44598_ ( .A(_source_stream_conv2d_8_source_6_pat_stride_buf_1), .B(_source_stream_conv2d_8_source_6_pat_stride_1), .S(_05674_), .Y(_23990_) );
  \$mux  #( .WIDTH(32) ) _44600_ ( .A(_source_stream_conv2d_8_source_6_pat_stride_buf_0), .B(_source_stream_conv2d_8_source_6_pat_stride_0), .S(_05674_), .Y(_23991_) );
  \$mux  #( .WIDTH(33) ) _44602_ ( .A(_source_stream_conv2d_8_source_6_pat_size_buf_3), .B(_source_stream_conv2d_8_source_6_pat_size_3), .S(_05674_), .Y(_23992_) );
  \$mux  #( .WIDTH(33) ) _44604_ ( .A(_source_stream_conv2d_8_source_6_pat_size_buf_2), .B(_source_stream_conv2d_8_source_6_pat_size_2), .S(_05674_), .Y(_23993_) );
  \$mux  #( .WIDTH(33) ) _44606_ ( .A(_source_stream_conv2d_8_source_6_pat_size_buf_1), .B(_source_stream_conv2d_8_source_6_pat_size_1), .S(_05674_), .Y(_23994_) );
  \$mux  #( .WIDTH(33) ) _44608_ ( .A(_source_stream_conv2d_8_source_6_pat_size_buf_0), .B(_source_stream_conv2d_8_source_6_pat_size_0), .S(_05674_), .Y(_23995_) );
  \$mux  #( .WIDTH(33) ) _44610_ ( .A(_source_stream_conv2d_8_source_6_pat_count_3), .B(_26019_), .S(_05674_), .Y(_23996_) );
  \$mux  #( .WIDTH(33) ) _44611_ ( .A(_23996_), .B(_26026_), .S(_05677_), .Y(_23997_) );
  \$mux  #( .WIDTH(33) ) _44612_ ( .A(_23997_), .B(_26027_), .S(_05678_), .Y(_23998_) );
  \$mux  #( .WIDTH(33) ) _44614_ ( .A(_source_stream_conv2d_8_source_6_pat_count_2), .B(_26018_), .S(_05674_), .Y(_23999_) );
  \$mux  #( .WIDTH(33) ) _44615_ ( .A(_23999_), .B(_26024_), .S(_05676_), .Y(_24000_) );
  \$mux  #( .WIDTH(33) ) _44616_ ( .A(_24000_), .B(_26025_), .S(_05677_), .Y(_24001_) );
  \$mux  #( .WIDTH(33) ) _44618_ ( .A(_source_stream_conv2d_8_source_6_pat_count_1), .B(_26017_), .S(_05674_), .Y(_24002_) );
  \$mux  #( .WIDTH(33) ) _44619_ ( .A(_24002_), .B(_26022_), .S(_05675_), .Y(_24003_) );
  \$mux  #( .WIDTH(33) ) _44620_ ( .A(_24003_), .B(_26023_), .S(_05676_), .Y(_24004_) );
  \$mux  #( .WIDTH(33) ) _44622_ ( .A(_source_stream_conv2d_8_source_6_pat_count_0), .B(_26016_), .S(_05674_), .Y(_24005_) );
  \$mux  #( .WIDTH(33) ) _44623_ ( .A(_26020_), .B(_24005_), .S(_05099_), .Y(_24006_) );
  \$mux  #( .WIDTH(33) ) _44624_ ( .A(_24006_), .B(_26021_), .S(_05675_), .Y(_24007_) );
  \$mux  #( .WIDTH(32) ) _44626_ ( .A(_source_stream_conv2d_8_source_6_pat_stride_3), .B(0), .S(_set_flag_538), .Y(_24008_) );
  \$mux  #( .WIDTH(32) ) _44628_ ( .A(_source_stream_conv2d_8_source_6_pat_stride_2), .B(0), .S(_set_flag_538), .Y(_24009_) );
  \$mux  #( .WIDTH(32) ) _44630_ ( .A(_source_stream_conv2d_8_source_6_pat_stride_1), .B(_26629_), .S(_set_flag_538), .Y(_24010_) );
  \$mux  #( .WIDTH(32) ) _44632_ ( .A(_source_stream_conv2d_8_source_6_pat_stride_0), .B(0), .S(_set_flag_538), .Y(_24011_) );
  \$mux  #( .WIDTH(33) ) _44634_ ( .A(_source_stream_conv2d_8_source_6_pat_size_3), .B(33'h000000001), .S(_set_flag_538), .Y(_24012_) );
  \$mux  #( .WIDTH(33) ) _44636_ ( .A(_source_stream_conv2d_8_source_6_pat_size_2), .B(33'h000000001), .S(_set_flag_538), .Y(_24013_) );
  \$mux  #( .WIDTH(33) ) _44638_ ( .A(_source_stream_conv2d_8_source_6_pat_size_1), .B({ 1'h0, conv2d_8_next_stream_num_ops }), .S(_set_flag_538), .Y(_24014_) );
  \$mux  #( .WIDTH(33) ) _44640_ ( .A(_source_stream_conv2d_8_source_6_pat_size_0), .B({ 28'h0000000, cparam_conv2d_8_stream_reduce_size }), .S(_set_flag_538), .Y(_24015_) );
  \$mux  #( .WIDTH(32) ) _44642_ ( .A(_source_stream_conv2d_8_source_6_pat_cur_offset_3), .B(0), .S(_05674_), .Y(_24016_) );
  \$mux  #( .WIDTH(32) ) _44643_ ( .A(_24016_), .B(_22143_), .S(_05677_), .Y(_24017_) );
  \$mux  #( .WIDTH(32) ) _44644_ ( .A(_24017_), .B(0), .S(_05678_), .Y(_24018_) );
  \$mux  #( .WIDTH(32) ) _44646_ ( .A(_source_stream_conv2d_8_source_6_pat_cur_offset_2), .B(0), .S(_05674_), .Y(_24019_) );
  \$mux  #( .WIDTH(32) ) _44647_ ( .A(_24019_), .B(_22142_), .S(_05676_), .Y(_24020_) );
  \$mux  #( .WIDTH(32) ) _44648_ ( .A(_24020_), .B(0), .S(_05677_), .Y(_24021_) );
  \$mux  #( .WIDTH(32) ) _44650_ ( .A(_source_stream_conv2d_8_source_6_pat_cur_offset_1), .B(0), .S(_05674_), .Y(_24022_) );
  \$mux  #( .WIDTH(32) ) _44651_ ( .A(_24022_), .B(_22141_), .S(_05675_), .Y(_24023_) );
  \$mux  #( .WIDTH(32) ) _44652_ ( .A(_24023_), .B(0), .S(_05676_), .Y(_24024_) );
  \$mux  #( .WIDTH(32) ) _44654_ ( .A(_source_stream_conv2d_8_source_6_pat_cur_offset_0), .B(0), .S(_05674_), .Y(_24025_) );
  \$mux  #( .WIDTH(32) ) _44655_ ( .A(_22140_), .B(_24025_), .S(_05099_), .Y(_24026_) );
  \$mux  #( .WIDTH(32) ) _44656_ ( .A(_24026_), .B(0), .S(_05675_), .Y(_24027_) );
  \$mux  #( .WIDTH(9) ) _44658_ ( .A(__variable_wdata_197), .B(_stream_conv2d_8_constant_3_next_constant_data), .S(_stream_conv2d_8_start), .Y(_24028_) );
  \$mux  #( .WIDTH(2) ) _44660_ ( .A(__variable_wdata_196), .B(_stream_conv2d_8_constant_2_next_constant_data), .S(_stream_conv2d_8_start), .Y(_24029_) );
  \$mux  #( .WIDTH(2) ) _44662_ ( .A(__variable_wdata_195), .B(_stream_conv2d_8_constant_1_next_constant_data), .S(_stream_conv2d_8_start), .Y(_24030_) );
  \$mux  #( .WIDTH(5) ) _44664_ ( .A(__variable_wdata_194), .B(_stream_conv2d_8_constant_0_next_constant_data), .S(_stream_conv2d_8_start), .Y(_24031_) );
  \$mux  #( .WIDTH(1) ) _44666_ ( .A(1'h1), .B(1'h0), .S(_05101_), .Y(_23201_) );
  \$mux  #( .WIDTH(8) ) _45105_ ( .A(_stream_conv2d_8_sink_37_sink_wdata), .B(_cond_data_755), .S(_05775_), .Y(_24032_) );
  \$mux  #( .WIDTH(1) ) _45107_ ( .A(1'h0), .B(1'h1), .S(_05775_), .Y(_24033_) );
  \$mux  #( .WIDTH(32) ) _45109_ ( .A(_stream_conv2d_8_sink_37_sink_waddr), .B(_26256_), .S(_05774_), .Y(_24034_) );
  \$mux  #( .WIDTH(32) ) _45110_ ( .A(_24034_), .B(_22230_), .S(_05775_), .Y(_24035_) );
  \$mux  #( .WIDTH(8) ) _45112_ ( .A(_stream_conv2d_8_sink_37_sink_ram_sel), .B(8'h15), .S(__set_flag_538_45), .Y(_24036_) );
  \$mux  #( .WIDTH(32) ) _45114_ ( .A(_stream_conv2d_8_sink_37_sink_stride_buf), .B(_stream_conv2d_8_sink_37_sink_stride), .S(_05774_), .Y(_24037_) );
  \$mux  #( .WIDTH(33) ) _45116_ ( .A(_stream_conv2d_8_sink_37_sink_count), .B(_stream_conv2d_8_sink_37_sink_size), .S(_05774_), .Y(_24038_) );
  \$mux  #( .WIDTH(33) ) _45117_ ( .A(_24038_), .B(_26257_), .S(_05775_), .Y(_24039_) );
  \$mux  #( .WIDTH(32) ) _45119_ ( .A(_stream_conv2d_8_sink_37_sink_stride), .B(1), .S(__set_flag_538_45), .Y(_24040_) );
  \$mux  #( .WIDTH(33) ) _45121_ ( .A(_stream_conv2d_8_sink_37_sink_size), .B(__stream_conv2d_8_sink_37_sink_size_1_45), .S(__set_flag_538_45), .Y(_24041_) );
  \$mux  #( .WIDTH(32) ) _45123_ ( .A(_stream_conv2d_8_sink_37_sink_offset), .B(__stream_conv2d_8_sink_37_sink_offset_0_45), .S(__set_flag_538_45), .Y(_24042_) );
  \$mux  #( .WIDTH(3) ) _45125_ ( .A(_stream_conv2d_8_sink_37_sink_mode), .B(3'h1), .S(__set_flag_538_45), .Y(_24043_) );
  \$mux  #( .WIDTH(1) ) _45127_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id9_0_cond_1_1), .Y(_24044_) );
  \$mux  #( .WIDTH(1) ) _45129_ ( .A(1'h1), .B(_stream_conv2d_8_source_36_source_ram_renable), .S(_05061_), .Y(_24045_) );
  \$mux  #( .WIDTH(1) ) _45130_ ( .A(1'h0), .B(_24045_), .S(_05060_), .Y(_24046_) );
  \$mux  #( .WIDTH(32) ) _45132_ ( .A(_stream_conv2d_8_source_36_source_pat_all_offset), .B(_stream_conv2d_8_source_36_source_ram_raddr), .S(_05061_), .Y(_24047_) );
  \$mux  #( .WIDTH(8) ) _45134_ ( .A(_stream_conv2d_8_source_36_source_ram_sel), .B(8'h14), .S(_set_flag_538), .Y(_24048_) );
  \$mux  #( .WIDTH(32) ) _45136_ ( .A(_stream_conv2d_8_source_36_source_offset_buf), .B(_stream_conv2d_8_source_36_source_offset), .S(_05769_), .Y(_24049_) );
  \$mux  #( .WIDTH(32) ) _45138_ ( .A(_stream_conv2d_8_source_36_source_offset), .B(conv2d_8_filter_page_comp_offset_buf), .S(_set_flag_538), .Y(_24050_) );
  \$mux  #( .WIDTH(3) ) _45140_ ( .A(_stream_conv2d_8_source_36_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24051_) );
  \$mux  #( .WIDTH(1) ) _45142_ ( .A(_stream_conv2d_8_source_36_idle), .B(1'h0), .S(_05769_), .Y(_24052_) );
  \$mux  #( .WIDTH(1) ) _45143_ ( .A(1'h1), .B(_24052_), .S(_05060_), .Y(_24053_) );
  \$mux  #( .WIDTH(1) ) _45144_ ( .A(_24053_), .B(1'h1), .S(RST), .Y(_02548_) );
  \$mux  #( .WIDTH(1) ) _45145_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id8_3_cond_1_1), .Y(_24054_) );
  \$mux  #( .WIDTH(1) ) _45147_ ( .A(1'h1), .B(_stream_conv2d_8_source_35_source_ram_renable), .S(_05064_), .Y(_24055_) );
  \$mux  #( .WIDTH(1) ) _45148_ ( .A(1'h0), .B(_24055_), .S(_05062_), .Y(_24056_) );
  \$mux  #( .WIDTH(32) ) _45150_ ( .A(_stream_conv2d_8_source_35_source_pat_all_offset), .B(_stream_conv2d_8_source_35_source_ram_raddr), .S(_05064_), .Y(_24057_) );
  \$mux  #( .WIDTH(8) ) _45152_ ( .A(_stream_conv2d_8_source_35_source_ram_sel), .B(8'h13), .S(_set_flag_538), .Y(_24058_) );
  \$mux  #( .WIDTH(32) ) _45154_ ( .A(_stream_conv2d_8_source_35_source_offset_buf), .B(_stream_conv2d_8_source_35_source_offset), .S(_05764_), .Y(_24059_) );
  \$mux  #( .WIDTH(32) ) _45156_ ( .A(_stream_conv2d_8_source_35_source_offset), .B(conv2d_8_filter_page_comp_offset_buf), .S(_set_flag_538), .Y(_24060_) );
  \$mux  #( .WIDTH(3) ) _45158_ ( .A(_stream_conv2d_8_source_35_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24061_) );
  \$mux  #( .WIDTH(1) ) _45160_ ( .A(_stream_conv2d_8_source_35_idle), .B(1'h0), .S(_05764_), .Y(_24062_) );
  \$mux  #( .WIDTH(1) ) _45161_ ( .A(1'h1), .B(_24062_), .S(_05062_), .Y(_24063_) );
  \$mux  #( .WIDTH(1) ) _45162_ ( .A(_24063_), .B(1'h1), .S(RST), .Y(_02539_) );
  \$mux  #( .WIDTH(1) ) _45163_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id7_3_cond_1_1), .Y(_24064_) );
  \$mux  #( .WIDTH(1) ) _45165_ ( .A(1'h1), .B(_stream_conv2d_8_source_34_source_ram_renable), .S(_05066_), .Y(_24065_) );
  \$mux  #( .WIDTH(1) ) _45166_ ( .A(1'h0), .B(_24065_), .S(_05063_), .Y(_24066_) );
  \$mux  #( .WIDTH(32) ) _45168_ ( .A(_stream_conv2d_8_source_34_source_pat_all_offset), .B(_stream_conv2d_8_source_34_source_ram_raddr), .S(_05066_), .Y(_24067_) );
  \$mux  #( .WIDTH(8) ) _45170_ ( .A(_stream_conv2d_8_source_34_source_ram_sel), .B(8'h12), .S(_set_flag_538), .Y(_24068_) );
  \$mux  #( .WIDTH(32) ) _45172_ ( .A(_stream_conv2d_8_source_34_source_offset_buf), .B(_stream_conv2d_8_source_34_source_offset), .S(_05759_), .Y(_24069_) );
  \$mux  #( .WIDTH(32) ) _45174_ ( .A(_stream_conv2d_8_source_34_source_offset), .B(conv2d_8_filter_page_comp_offset_buf), .S(_set_flag_538), .Y(_24070_) );
  \$mux  #( .WIDTH(3) ) _45176_ ( .A(_stream_conv2d_8_source_34_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24071_) );
  \$mux  #( .WIDTH(1) ) _45178_ ( .A(_stream_conv2d_8_source_34_idle), .B(1'h0), .S(_05759_), .Y(_24072_) );
  \$mux  #( .WIDTH(1) ) _45179_ ( .A(1'h1), .B(_24072_), .S(_05063_), .Y(_24073_) );
  \$mux  #( .WIDTH(1) ) _45180_ ( .A(_24073_), .B(1'h1), .S(RST), .Y(_02530_) );
  \$mux  #( .WIDTH(1) ) _45181_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id6_3_cond_1_1), .Y(_24074_) );
  \$mux  #( .WIDTH(1) ) _45183_ ( .A(1'h1), .B(_stream_conv2d_8_source_33_source_ram_renable), .S(_05067_), .Y(_24075_) );
  \$mux  #( .WIDTH(1) ) _45184_ ( .A(1'h0), .B(_24075_), .S(_05065_), .Y(_24076_) );
  \$mux  #( .WIDTH(32) ) _45186_ ( .A(_stream_conv2d_8_source_33_source_pat_all_offset), .B(_stream_conv2d_8_source_33_source_ram_raddr), .S(_05067_), .Y(_24077_) );
  \$mux  #( .WIDTH(8) ) _45188_ ( .A(_stream_conv2d_8_source_33_source_ram_sel), .B(8'h11), .S(_set_flag_538), .Y(_24078_) );
  \$mux  #( .WIDTH(32) ) _45190_ ( .A(_stream_conv2d_8_source_33_source_offset_buf), .B(_stream_conv2d_8_source_33_source_offset), .S(_05754_), .Y(_24079_) );
  \$mux  #( .WIDTH(32) ) _45192_ ( .A(_stream_conv2d_8_source_33_source_offset), .B(conv2d_8_filter_page_comp_offset_buf), .S(_set_flag_538), .Y(_24080_) );
  \$mux  #( .WIDTH(3) ) _45194_ ( .A(_stream_conv2d_8_source_33_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24081_) );
  \$mux  #( .WIDTH(1) ) _45196_ ( .A(_stream_conv2d_8_source_33_idle), .B(1'h0), .S(_05754_), .Y(_24082_) );
  \$mux  #( .WIDTH(1) ) _45197_ ( .A(1'h1), .B(_24082_), .S(_05065_), .Y(_24083_) );
  \$mux  #( .WIDTH(1) ) _45198_ ( .A(_24083_), .B(1'h1), .S(RST), .Y(_02521_) );
  \$mux  #( .WIDTH(1) ) _45199_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id5_3_cond_1_1), .Y(_24084_) );
  \$mux  #( .WIDTH(1) ) _45201_ ( .A(1'h1), .B(_stream_conv2d_8_source_32_source_ram_renable), .S(_05069_), .Y(_24085_) );
  \$mux  #( .WIDTH(1) ) _45202_ ( .A(1'h0), .B(_24085_), .S(_05068_), .Y(_24086_) );
  \$mux  #( .WIDTH(32) ) _45204_ ( .A(_stream_conv2d_8_source_32_source_pat_all_offset), .B(_stream_conv2d_8_source_32_source_ram_raddr), .S(_05069_), .Y(_24087_) );
  \$mux  #( .WIDTH(8) ) _45206_ ( .A(_stream_conv2d_8_source_32_source_ram_sel), .B(8'h10), .S(_set_flag_538), .Y(_24088_) );
  \$mux  #( .WIDTH(32) ) _45208_ ( .A(_stream_conv2d_8_source_32_source_offset_buf), .B(_stream_conv2d_8_source_32_source_offset), .S(_05749_), .Y(_24089_) );
  \$mux  #( .WIDTH(32) ) _45210_ ( .A(_stream_conv2d_8_source_32_source_offset), .B(conv2d_8_filter_page_comp_offset_buf), .S(_set_flag_538), .Y(_24090_) );
  \$mux  #( .WIDTH(3) ) _45212_ ( .A(_stream_conv2d_8_source_32_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24091_) );
  \$mux  #( .WIDTH(1) ) _45214_ ( .A(_stream_conv2d_8_source_32_idle), .B(1'h0), .S(_05749_), .Y(_24092_) );
  \$mux  #( .WIDTH(1) ) _45215_ ( .A(1'h1), .B(_24092_), .S(_05068_), .Y(_24093_) );
  \$mux  #( .WIDTH(1) ) _45216_ ( .A(_24093_), .B(1'h1), .S(RST), .Y(_02512_) );
  \$mux  #( .WIDTH(1) ) _45217_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id4_3_cond_1_1), .Y(_24094_) );
  \$mux  #( .WIDTH(1) ) _45219_ ( .A(1'h1), .B(_stream_conv2d_8_source_31_source_ram_renable), .S(_05071_), .Y(_24095_) );
  \$mux  #( .WIDTH(1) ) _45220_ ( .A(1'h0), .B(_24095_), .S(_05070_), .Y(_24096_) );
  \$mux  #( .WIDTH(32) ) _45222_ ( .A(_stream_conv2d_8_source_31_source_pat_all_offset), .B(_stream_conv2d_8_source_31_source_ram_raddr), .S(_05071_), .Y(_24097_) );
  \$mux  #( .WIDTH(8) ) _45224_ ( .A(_stream_conv2d_8_source_31_source_ram_sel), .B(8'h0f), .S(_set_flag_538), .Y(_24098_) );
  \$mux  #( .WIDTH(32) ) _45226_ ( .A(_stream_conv2d_8_source_31_source_offset_buf), .B(_stream_conv2d_8_source_31_source_offset), .S(_05744_), .Y(_24099_) );
  \$mux  #( .WIDTH(32) ) _45228_ ( .A(_stream_conv2d_8_source_31_source_offset), .B(conv2d_8_filter_page_comp_offset_buf), .S(_set_flag_538), .Y(_24100_) );
  \$mux  #( .WIDTH(3) ) _45230_ ( .A(_stream_conv2d_8_source_31_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24101_) );
  \$mux  #( .WIDTH(1) ) _45232_ ( .A(_stream_conv2d_8_source_31_idle), .B(1'h0), .S(_05744_), .Y(_24102_) );
  \$mux  #( .WIDTH(1) ) _45233_ ( .A(1'h1), .B(_24102_), .S(_05070_), .Y(_24103_) );
  \$mux  #( .WIDTH(1) ) _45234_ ( .A(_24103_), .B(1'h1), .S(RST), .Y(_02503_) );
  \$mux  #( .WIDTH(1) ) _45235_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id3_3_cond_1_1), .Y(_24104_) );
  \$mux  #( .WIDTH(1) ) _45237_ ( .A(1'h1), .B(_stream_conv2d_8_source_30_source_ram_renable), .S(_05073_), .Y(_24105_) );
  \$mux  #( .WIDTH(1) ) _45238_ ( .A(1'h0), .B(_24105_), .S(_05072_), .Y(_24106_) );
  \$mux  #( .WIDTH(32) ) _45240_ ( .A(_stream_conv2d_8_source_30_source_pat_all_offset), .B(_stream_conv2d_8_source_30_source_ram_raddr), .S(_05073_), .Y(_24107_) );
  \$mux  #( .WIDTH(8) ) _45242_ ( .A(_stream_conv2d_8_source_30_source_ram_sel), .B(8'h0e), .S(_set_flag_538), .Y(_24108_) );
  \$mux  #( .WIDTH(32) ) _45244_ ( .A(_stream_conv2d_8_source_30_source_offset_buf), .B(_stream_conv2d_8_source_30_source_offset), .S(_05739_), .Y(_24109_) );
  \$mux  #( .WIDTH(32) ) _45246_ ( .A(_stream_conv2d_8_source_30_source_offset), .B(conv2d_8_filter_page_comp_offset_buf), .S(_set_flag_538), .Y(_24110_) );
  \$mux  #( .WIDTH(3) ) _45248_ ( .A(_stream_conv2d_8_source_30_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24111_) );
  \$mux  #( .WIDTH(1) ) _45250_ ( .A(_stream_conv2d_8_source_30_idle), .B(1'h0), .S(_05739_), .Y(_24112_) );
  \$mux  #( .WIDTH(1) ) _45251_ ( .A(1'h1), .B(_24112_), .S(_05072_), .Y(_24113_) );
  \$mux  #( .WIDTH(1) ) _45252_ ( .A(_24113_), .B(1'h1), .S(RST), .Y(_02494_) );
  \$mux  #( .WIDTH(1) ) _45253_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id2_3_cond_1_1), .Y(_24114_) );
  \$mux  #( .WIDTH(1) ) _45255_ ( .A(1'h1), .B(_stream_conv2d_8_source_29_source_ram_renable), .S(_05075_), .Y(_24115_) );
  \$mux  #( .WIDTH(1) ) _45256_ ( .A(1'h0), .B(_24115_), .S(_05074_), .Y(_24116_) );
  \$mux  #( .WIDTH(32) ) _45258_ ( .A(_stream_conv2d_8_source_29_source_pat_all_offset), .B(_stream_conv2d_8_source_29_source_ram_raddr), .S(_05075_), .Y(_24117_) );
  \$mux  #( .WIDTH(8) ) _45260_ ( .A(_stream_conv2d_8_source_29_source_ram_sel), .B(8'h0d), .S(_set_flag_538), .Y(_24118_) );
  \$mux  #( .WIDTH(32) ) _45262_ ( .A(_stream_conv2d_8_source_29_source_offset_buf), .B(_stream_conv2d_8_source_29_source_offset), .S(_05734_), .Y(_24119_) );
  \$mux  #( .WIDTH(32) ) _45264_ ( .A(_stream_conv2d_8_source_29_source_offset), .B(conv2d_8_filter_page_comp_offset_buf), .S(_set_flag_538), .Y(_24120_) );
  \$mux  #( .WIDTH(3) ) _45266_ ( .A(_stream_conv2d_8_source_29_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24121_) );
  \$mux  #( .WIDTH(1) ) _45268_ ( .A(_stream_conv2d_8_source_29_idle), .B(1'h0), .S(_05734_), .Y(_24122_) );
  \$mux  #( .WIDTH(1) ) _45269_ ( .A(1'h1), .B(_24122_), .S(_05074_), .Y(_24123_) );
  \$mux  #( .WIDTH(1) ) _45270_ ( .A(_24123_), .B(1'h1), .S(RST), .Y(_02485_) );
  \$mux  #( .WIDTH(1) ) _45271_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id1_3_cond_2_1), .Y(_24124_) );
  \$mux  #( .WIDTH(1) ) _45273_ ( .A(1'h1), .B(_stream_conv2d_8_source_28_source_ram_renable), .S(_05077_), .Y(_24125_) );
  \$mux  #( .WIDTH(1) ) _45274_ ( .A(1'h0), .B(_24125_), .S(_05076_), .Y(_24126_) );
  \$mux  #( .WIDTH(32) ) _45276_ ( .A(_stream_conv2d_8_source_28_source_pat_all_offset), .B(_stream_conv2d_8_source_28_source_ram_raddr), .S(_05077_), .Y(_24127_) );
  \$mux  #( .WIDTH(8) ) _45278_ ( .A(_stream_conv2d_8_source_28_source_ram_sel), .B(8'h0c), .S(_set_flag_538), .Y(_24128_) );
  \$mux  #( .WIDTH(32) ) _45280_ ( .A(_stream_conv2d_8_source_28_source_offset_buf), .B(_stream_conv2d_8_source_28_source_offset), .S(_05729_), .Y(_24129_) );
  \$mux  #( .WIDTH(32) ) _45282_ ( .A(_stream_conv2d_8_source_28_source_offset), .B(conv2d_8_filter_page_comp_offset_buf), .S(_set_flag_538), .Y(_24130_) );
  \$mux  #( .WIDTH(3) ) _45284_ ( .A(_stream_conv2d_8_source_28_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24131_) );
  \$mux  #( .WIDTH(1) ) _45286_ ( .A(_stream_conv2d_8_source_28_idle), .B(1'h0), .S(_05729_), .Y(_24132_) );
  \$mux  #( .WIDTH(1) ) _45287_ ( .A(1'h1), .B(_24132_), .S(_05076_), .Y(_24133_) );
  \$mux  #( .WIDTH(1) ) _45288_ ( .A(_24133_), .B(1'h1), .S(RST), .Y(_02476_) );
  \$mux  #( .WIDTH(1) ) _45289_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id18_0_cond_2_1), .Y(_24134_) );
  \$mux  #( .WIDTH(1) ) _45291_ ( .A(1'h1), .B(_stream_conv2d_8_source_27_source_ram_renable), .S(_05079_), .Y(_24135_) );
  \$mux  #( .WIDTH(1) ) _45292_ ( .A(1'h0), .B(_24135_), .S(_05078_), .Y(_24136_) );
  \$mux  #( .WIDTH(32) ) _45294_ ( .A(_stream_conv2d_8_source_27_source_pat_all_offset), .B(_stream_conv2d_8_source_27_source_ram_raddr), .S(_05079_), .Y(_24137_) );
  \$mux  #( .WIDTH(8) ) _45296_ ( .A(_stream_conv2d_8_source_27_source_ram_sel), .B(8'h0b), .S(_set_flag_538), .Y(_24138_) );
  \$mux  #( .WIDTH(32) ) _45298_ ( .A(_stream_conv2d_8_source_27_source_offset_buf), .B(_stream_conv2d_8_source_27_source_offset), .S(_05724_), .Y(_24139_) );
  \$mux  #( .WIDTH(32) ) _45300_ ( .A(_stream_conv2d_8_source_27_source_offset), .B(_22188_), .S(_set_flag_538), .Y(_24140_) );
  \$mux  #( .WIDTH(3) ) _45302_ ( .A(_stream_conv2d_8_source_27_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24141_) );
  \$mux  #( .WIDTH(1) ) _45304_ ( .A(_stream_conv2d_8_source_27_idle), .B(1'h0), .S(_05724_), .Y(_24142_) );
  \$mux  #( .WIDTH(1) ) _45305_ ( .A(1'h1), .B(_24142_), .S(_05078_), .Y(_24143_) );
  \$mux  #( .WIDTH(1) ) _45306_ ( .A(_24143_), .B(1'h1), .S(RST), .Y(_02467_) );
  \$mux  #( .WIDTH(1) ) _45307_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id17_0_cond_2_1), .Y(_24144_) );
  \$mux  #( .WIDTH(1) ) _45309_ ( .A(1'h1), .B(_stream_conv2d_8_source_26_source_ram_renable), .S(_05081_), .Y(_24145_) );
  \$mux  #( .WIDTH(1) ) _45310_ ( .A(1'h0), .B(_24145_), .S(_05080_), .Y(_24146_) );
  \$mux  #( .WIDTH(32) ) _45312_ ( .A(_stream_conv2d_8_source_26_source_pat_all_offset), .B(_stream_conv2d_8_source_26_source_ram_raddr), .S(_05081_), .Y(_24147_) );
  \$mux  #( .WIDTH(8) ) _45314_ ( .A(_stream_conv2d_8_source_26_source_ram_sel), .B(8'h0a), .S(_set_flag_538), .Y(_24148_) );
  \$mux  #( .WIDTH(32) ) _45316_ ( .A(_stream_conv2d_8_source_26_source_offset_buf), .B(_stream_conv2d_8_source_26_source_offset), .S(_05719_), .Y(_24149_) );
  \$mux  #( .WIDTH(32) ) _45318_ ( .A(_stream_conv2d_8_source_26_source_offset), .B(_22183_), .S(_set_flag_538), .Y(_24150_) );
  \$mux  #( .WIDTH(3) ) _45320_ ( .A(_stream_conv2d_8_source_26_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24151_) );
  \$mux  #( .WIDTH(1) ) _45322_ ( .A(_stream_conv2d_8_source_26_idle), .B(1'h0), .S(_05719_), .Y(_24152_) );
  \$mux  #( .WIDTH(1) ) _45323_ ( .A(1'h1), .B(_24152_), .S(_05080_), .Y(_24153_) );
  \$mux  #( .WIDTH(1) ) _45324_ ( .A(_24153_), .B(1'h1), .S(RST), .Y(_02458_) );
  \$mux  #( .WIDTH(1) ) _45325_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id16_0_cond_3_1), .Y(_24154_) );
  \$mux  #( .WIDTH(1) ) _45327_ ( .A(1'h1), .B(_stream_conv2d_8_source_25_source_ram_renable), .S(_05083_), .Y(_24155_) );
  \$mux  #( .WIDTH(1) ) _45328_ ( .A(1'h0), .B(_24155_), .S(_05082_), .Y(_24156_) );
  \$mux  #( .WIDTH(32) ) _45330_ ( .A(_stream_conv2d_8_source_25_source_pat_all_offset), .B(_stream_conv2d_8_source_25_source_ram_raddr), .S(_05083_), .Y(_24157_) );
  \$mux  #( .WIDTH(8) ) _45332_ ( .A(_stream_conv2d_8_source_25_source_ram_sel), .B(8'h09), .S(_set_flag_538), .Y(_24158_) );
  \$mux  #( .WIDTH(32) ) _45334_ ( .A(_stream_conv2d_8_source_25_source_offset_buf), .B(_stream_conv2d_8_source_25_source_offset), .S(_05714_), .Y(_24159_) );
  \$mux  #( .WIDTH(32) ) _45336_ ( .A(_stream_conv2d_8_source_25_source_offset), .B(_22178_), .S(_set_flag_538), .Y(_24160_) );
  \$mux  #( .WIDTH(3) ) _45338_ ( .A(_stream_conv2d_8_source_25_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24161_) );
  \$mux  #( .WIDTH(1) ) _45340_ ( .A(_stream_conv2d_8_source_25_idle), .B(1'h0), .S(_05714_), .Y(_24162_) );
  \$mux  #( .WIDTH(1) ) _45341_ ( .A(1'h1), .B(_24162_), .S(_05082_), .Y(_24163_) );
  \$mux  #( .WIDTH(1) ) _45342_ ( .A(_24163_), .B(1'h1), .S(RST), .Y(_02449_) );
  \$mux  #( .WIDTH(1) ) _45343_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id15_0_cond_2_1), .Y(_24164_) );
  \$mux  #( .WIDTH(1) ) _45345_ ( .A(1'h1), .B(_stream_conv2d_8_source_24_source_ram_renable), .S(_05085_), .Y(_24165_) );
  \$mux  #( .WIDTH(1) ) _45346_ ( .A(1'h0), .B(_24165_), .S(_05084_), .Y(_24166_) );
  \$mux  #( .WIDTH(32) ) _45348_ ( .A(_stream_conv2d_8_source_24_source_pat_all_offset), .B(_stream_conv2d_8_source_24_source_ram_raddr), .S(_05085_), .Y(_24167_) );
  \$mux  #( .WIDTH(8) ) _45350_ ( .A(_stream_conv2d_8_source_24_source_ram_sel), .B(8'h08), .S(_set_flag_538), .Y(_24168_) );
  \$mux  #( .WIDTH(32) ) _45352_ ( .A(_stream_conv2d_8_source_24_source_offset_buf), .B(_stream_conv2d_8_source_24_source_offset), .S(_05709_), .Y(_24169_) );
  \$mux  #( .WIDTH(32) ) _45354_ ( .A(_stream_conv2d_8_source_24_source_offset), .B(_22173_), .S(_set_flag_538), .Y(_24170_) );
  \$mux  #( .WIDTH(3) ) _45356_ ( .A(_stream_conv2d_8_source_24_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24171_) );
  \$mux  #( .WIDTH(1) ) _45358_ ( .A(_stream_conv2d_8_source_24_idle), .B(1'h0), .S(_05709_), .Y(_24172_) );
  \$mux  #( .WIDTH(1) ) _45359_ ( .A(1'h1), .B(_24172_), .S(_05084_), .Y(_24173_) );
  \$mux  #( .WIDTH(1) ) _45360_ ( .A(_24173_), .B(1'h1), .S(RST), .Y(_02440_) );
  \$mux  #( .WIDTH(1) ) _45361_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id14_0_cond_2_1), .Y(_24174_) );
  \$mux  #( .WIDTH(1) ) _45363_ ( .A(1'h1), .B(_stream_conv2d_8_source_23_source_ram_renable), .S(_05087_), .Y(_24175_) );
  \$mux  #( .WIDTH(1) ) _45364_ ( .A(1'h0), .B(_24175_), .S(_05086_), .Y(_24176_) );
  \$mux  #( .WIDTH(32) ) _45366_ ( .A(_stream_conv2d_8_source_23_source_pat_all_offset), .B(_stream_conv2d_8_source_23_source_ram_raddr), .S(_05087_), .Y(_24177_) );
  \$mux  #( .WIDTH(8) ) _45368_ ( .A(_stream_conv2d_8_source_23_source_ram_sel), .B(8'h07), .S(_set_flag_538), .Y(_24178_) );
  \$mux  #( .WIDTH(32) ) _45370_ ( .A(_stream_conv2d_8_source_23_source_offset_buf), .B(_stream_conv2d_8_source_23_source_offset), .S(_05704_), .Y(_24179_) );
  \$mux  #( .WIDTH(32) ) _45372_ ( .A(_stream_conv2d_8_source_23_source_offset), .B(_22168_), .S(_set_flag_538), .Y(_24180_) );
  \$mux  #( .WIDTH(3) ) _45374_ ( .A(_stream_conv2d_8_source_23_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24181_) );
  \$mux  #( .WIDTH(1) ) _45376_ ( .A(_stream_conv2d_8_source_23_idle), .B(1'h0), .S(_05704_), .Y(_24182_) );
  \$mux  #( .WIDTH(1) ) _45377_ ( .A(1'h1), .B(_24182_), .S(_05086_), .Y(_24183_) );
  \$mux  #( .WIDTH(1) ) _45378_ ( .A(_24183_), .B(1'h1), .S(RST), .Y(_02431_) );
  \$mux  #( .WIDTH(1) ) _45379_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id13_0_cond_3_1), .Y(_24184_) );
  \$mux  #( .WIDTH(1) ) _45381_ ( .A(1'h1), .B(_stream_conv2d_8_source_22_source_ram_renable), .S(_05089_), .Y(_24185_) );
  \$mux  #( .WIDTH(1) ) _45382_ ( .A(1'h0), .B(_24185_), .S(_05088_), .Y(_24186_) );
  \$mux  #( .WIDTH(32) ) _45384_ ( .A(_stream_conv2d_8_source_22_source_pat_all_offset), .B(_stream_conv2d_8_source_22_source_ram_raddr), .S(_05089_), .Y(_24187_) );
  \$mux  #( .WIDTH(8) ) _45386_ ( .A(_stream_conv2d_8_source_22_source_ram_sel), .B(8'h06), .S(_set_flag_538), .Y(_24188_) );
  \$mux  #( .WIDTH(32) ) _45388_ ( .A(_stream_conv2d_8_source_22_source_offset_buf), .B(_stream_conv2d_8_source_22_source_offset), .S(_05699_), .Y(_24189_) );
  \$mux  #( .WIDTH(32) ) _45390_ ( .A(_stream_conv2d_8_source_22_source_offset), .B(_22163_), .S(_set_flag_538), .Y(_24190_) );
  \$mux  #( .WIDTH(3) ) _45392_ ( .A(_stream_conv2d_8_source_22_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24191_) );
  \$mux  #( .WIDTH(1) ) _45394_ ( .A(_stream_conv2d_8_source_22_idle), .B(1'h0), .S(_05699_), .Y(_24192_) );
  \$mux  #( .WIDTH(1) ) _45395_ ( .A(1'h1), .B(_24192_), .S(_05088_), .Y(_24193_) );
  \$mux  #( .WIDTH(1) ) _45396_ ( .A(_24193_), .B(1'h1), .S(RST), .Y(_02422_) );
  \$mux  #( .WIDTH(1) ) _45397_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id12_0_cond_2_1), .Y(_24194_) );
  \$mux  #( .WIDTH(1) ) _45399_ ( .A(1'h1), .B(_stream_conv2d_8_source_21_source_ram_renable), .S(_05091_), .Y(_24195_) );
  \$mux  #( .WIDTH(1) ) _45400_ ( .A(1'h0), .B(_24195_), .S(_05090_), .Y(_24196_) );
  \$mux  #( .WIDTH(32) ) _45402_ ( .A(_stream_conv2d_8_source_21_source_pat_all_offset), .B(_stream_conv2d_8_source_21_source_ram_raddr), .S(_05091_), .Y(_24197_) );
  \$mux  #( .WIDTH(8) ) _45404_ ( .A(_stream_conv2d_8_source_21_source_ram_sel), .B(8'h05), .S(_set_flag_538), .Y(_24198_) );
  \$mux  #( .WIDTH(32) ) _45406_ ( .A(_stream_conv2d_8_source_21_source_offset_buf), .B(_stream_conv2d_8_source_21_source_offset), .S(_05694_), .Y(_24199_) );
  \$mux  #( .WIDTH(32) ) _45408_ ( .A(_stream_conv2d_8_source_21_source_offset), .B(_22158_), .S(_set_flag_538), .Y(_24200_) );
  \$mux  #( .WIDTH(3) ) _45410_ ( .A(_stream_conv2d_8_source_21_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24201_) );
  \$mux  #( .WIDTH(1) ) _45412_ ( .A(_stream_conv2d_8_source_21_idle), .B(1'h0), .S(_05694_), .Y(_24202_) );
  \$mux  #( .WIDTH(1) ) _45413_ ( .A(1'h1), .B(_24202_), .S(_05090_), .Y(_24203_) );
  \$mux  #( .WIDTH(1) ) _45414_ ( .A(_24203_), .B(1'h1), .S(RST), .Y(_02413_) );
  \$mux  #( .WIDTH(1) ) _45415_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id11_0_cond_2_1), .Y(_24204_) );
  \$mux  #( .WIDTH(1) ) _45417_ ( .A(1'h1), .B(_stream_conv2d_8_source_20_source_ram_renable), .S(_05093_), .Y(_24205_) );
  \$mux  #( .WIDTH(1) ) _45418_ ( .A(1'h0), .B(_24205_), .S(_05092_), .Y(_24206_) );
  \$mux  #( .WIDTH(32) ) _45420_ ( .A(_stream_conv2d_8_source_20_source_pat_all_offset), .B(_stream_conv2d_8_source_20_source_ram_raddr), .S(_05093_), .Y(_24207_) );
  \$mux  #( .WIDTH(8) ) _45422_ ( .A(_stream_conv2d_8_source_20_source_ram_sel), .B(8'h04), .S(_set_flag_538), .Y(_24208_) );
  \$mux  #( .WIDTH(32) ) _45424_ ( .A(_stream_conv2d_8_source_20_source_offset_buf), .B(_stream_conv2d_8_source_20_source_offset), .S(_05689_), .Y(_24209_) );
  \$mux  #( .WIDTH(32) ) _45426_ ( .A(_stream_conv2d_8_source_20_source_offset), .B(_22153_), .S(_set_flag_538), .Y(_24210_) );
  \$mux  #( .WIDTH(3) ) _45428_ ( .A(_stream_conv2d_8_source_20_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24211_) );
  \$mux  #( .WIDTH(1) ) _45430_ ( .A(_stream_conv2d_8_source_20_idle), .B(1'h0), .S(_05689_), .Y(_24212_) );
  \$mux  #( .WIDTH(1) ) _45431_ ( .A(1'h1), .B(_24212_), .S(_05092_), .Y(_24213_) );
  \$mux  #( .WIDTH(1) ) _45432_ ( .A(_24213_), .B(1'h1), .S(RST), .Y(_02404_) );
  \$mux  #( .WIDTH(1) ) _45433_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id10_0_cond_3_1), .Y(_24214_) );
  \$mux  #( .WIDTH(1) ) _45435_ ( .A(1'h1), .B(_stream_conv2d_8_source_19_source_ram_renable), .S(_05095_), .Y(_24215_) );
  \$mux  #( .WIDTH(1) ) _45436_ ( .A(1'h0), .B(_24215_), .S(_05094_), .Y(_24216_) );
  \$mux  #( .WIDTH(32) ) _45438_ ( .A(_stream_conv2d_8_source_19_source_pat_all_offset), .B(_stream_conv2d_8_source_19_source_ram_raddr), .S(_05095_), .Y(_24217_) );
  \$mux  #( .WIDTH(8) ) _45440_ ( .A(_stream_conv2d_8_source_19_source_ram_sel), .B(8'h03), .S(_set_flag_538), .Y(_24218_) );
  \$mux  #( .WIDTH(32) ) _45442_ ( .A(_stream_conv2d_8_source_19_source_offset_buf), .B(_stream_conv2d_8_source_19_source_offset), .S(_05684_), .Y(_24219_) );
  \$mux  #( .WIDTH(32) ) _45444_ ( .A(_stream_conv2d_8_source_19_source_offset), .B(_22148_), .S(_set_flag_538), .Y(_24220_) );
  \$mux  #( .WIDTH(3) ) _45446_ ( .A(_stream_conv2d_8_source_19_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24221_) );
  \$mux  #( .WIDTH(1) ) _45448_ ( .A(_stream_conv2d_8_source_19_idle), .B(1'h0), .S(_05684_), .Y(_24222_) );
  \$mux  #( .WIDTH(1) ) _45449_ ( .A(1'h1), .B(_24222_), .S(_05094_), .Y(_24223_) );
  \$mux  #( .WIDTH(1) ) _45450_ ( .A(_24223_), .B(1'h1), .S(RST), .Y(_02395_) );
  \$mux  #( .WIDTH(4) ) _45451_ ( .A(_stream_conv2d_8_constant_17_next_constant_data), .B(cparam_conv2d_8_cshamt_out_value), .S(_set_flag_538), .Y(_24224_) );
  \$mux  #( .WIDTH(1) ) _45453_ ( .A(_stream_conv2d_8_constant_16_next_constant_data), .B(1'h0), .S(_set_flag_538), .Y(_24225_) );
  \$mux  #( .WIDTH(1) ) _45455_ ( .A(_stream_conv2d_8_constant_15_next_constant_data), .B(1'h0), .S(_set_flag_538), .Y(_24226_) );
  \$mux  #( .WIDTH(8) ) _45457_ ( .A(_stream_conv2d_8_source_14_source_empty_data), .B(8'h00), .S(_set_flag_538), .Y(_24227_) );
  \$mux  #( .WIDTH(1) ) _45459_ ( .A(_stream_conv2d_8_source_14_idle), .B(1'h1), .S(_stream_conv2d_8_start), .Y(_24228_) );
  \$mux  #( .WIDTH(1) ) _45460_ ( .A(_24228_), .B(1'h1), .S(RST), .Y(_02393_) );
  \$mux  #( .WIDTH(8) ) _45461_ ( .A(_stream_conv2d_8_source_12_source_empty_data), .B(8'h00), .S(_set_flag_538), .Y(_24229_) );
  \$mux  #( .WIDTH(1) ) _45463_ ( .A(_stream_conv2d_8_source_12_idle), .B(1'h1), .S(_stream_conv2d_8_start), .Y(_24230_) );
  \$mux  #( .WIDTH(1) ) _45464_ ( .A(_24230_), .B(1'h1), .S(RST), .Y(_02391_) );
  \$mux  #( .WIDTH(8) ) _45465_ ( .A(_stream_conv2d_8_source_10_source_empty_data), .B(8'h00), .S(_set_flag_538), .Y(_24231_) );
  \$mux  #( .WIDTH(1) ) _45467_ ( .A(_stream_conv2d_8_source_10_idle), .B(1'h1), .S(_stream_conv2d_8_start), .Y(_24232_) );
  \$mux  #( .WIDTH(1) ) _45468_ ( .A(_24232_), .B(1'h1), .S(RST), .Y(_02389_) );
  \$mux  #( .WIDTH(1) ) _45469_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id0_3_cond_1_1), .Y(_24233_) );
  \$mux  #( .WIDTH(1) ) _45471_ ( .A(1'h1), .B(_stream_conv2d_8_source_8_source_ram_renable), .S(_05097_), .Y(_24234_) );
  \$mux  #( .WIDTH(1) ) _45472_ ( .A(1'h0), .B(_24234_), .S(_05096_), .Y(_24235_) );
  \$mux  #( .WIDTH(32) ) _45474_ ( .A(_stream_conv2d_8_source_8_source_pat_all_offset), .B(_stream_conv2d_8_source_8_source_ram_raddr), .S(_05097_), .Y(_24236_) );
  \$mux  #( .WIDTH(8) ) _45476_ ( .A(_stream_conv2d_8_source_8_source_ram_sel), .B(8'h02), .S(_set_flag_538), .Y(_24237_) );
  \$mux  #( .WIDTH(32) ) _45478_ ( .A(_stream_conv2d_8_source_8_source_offset_buf), .B(_stream_conv2d_8_source_8_source_offset), .S(_05679_), .Y(_24238_) );
  \$mux  #( .WIDTH(32) ) _45480_ ( .A(_stream_conv2d_8_source_8_source_offset), .B(0), .S(_set_flag_538), .Y(_24239_) );
  \$mux  #( .WIDTH(3) ) _45482_ ( .A(_stream_conv2d_8_source_8_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24240_) );
  \$mux  #( .WIDTH(1) ) _45484_ ( .A(_stream_conv2d_8_source_8_idle), .B(1'h0), .S(_05679_), .Y(_24241_) );
  \$mux  #( .WIDTH(1) ) _45485_ ( .A(1'h1), .B(_24241_), .S(_05096_), .Y(_24242_) );
  \$mux  #( .WIDTH(1) ) _45486_ ( .A(_24242_), .B(1'h1), .S(RST), .Y(_02566_) );
  \$mux  #( .WIDTH(1) ) _45487_ ( .A(1'h0), .B(1'h1), .S(_ram_w32_l128_id0_cond_2_1), .Y(_24243_) );
  \$mux  #( .WIDTH(1) ) _45489_ ( .A(1'h1), .B(_stream_conv2d_8_source_6_source_ram_renable), .S(_05099_), .Y(_24244_) );
  \$mux  #( .WIDTH(1) ) _45490_ ( .A(1'h0), .B(_24244_), .S(_05098_), .Y(_24245_) );
  \$mux  #( .WIDTH(32) ) _45492_ ( .A(_stream_conv2d_8_source_6_source_pat_all_offset), .B(_stream_conv2d_8_source_6_source_ram_raddr), .S(_05099_), .Y(_24246_) );
  \$mux  #( .WIDTH(8) ) _45494_ ( .A(_stream_conv2d_8_source_6_source_ram_sel), .B(8'h01), .S(_set_flag_538), .Y(_24247_) );
  \$mux  #( .WIDTH(32) ) _45496_ ( .A(_stream_conv2d_8_source_6_source_offset_buf), .B(_stream_conv2d_8_source_6_source_offset), .S(_05674_), .Y(_24248_) );
  \$mux  #( .WIDTH(32) ) _45498_ ( .A(_stream_conv2d_8_source_6_source_offset), .B(_26628_), .S(_set_flag_538), .Y(_24249_) );
  \$mux  #( .WIDTH(3) ) _45500_ ( .A(_stream_conv2d_8_source_6_source_mode), .B(3'h2), .S(_set_flag_538), .Y(_24250_) );
  \$mux  #( .WIDTH(1) ) _45502_ ( .A(_stream_conv2d_8_source_6_idle), .B(1'h0), .S(_05674_), .Y(_24251_) );
  \$mux  #( .WIDTH(1) ) _45503_ ( .A(1'h1), .B(_24251_), .S(_05098_), .Y(_24252_) );
  \$mux  #( .WIDTH(1) ) _45504_ ( .A(_24252_), .B(1'h1), .S(RST), .Y(_02557_) );
  \$mux  #( .WIDTH(9) ) _45505_ ( .A(_stream_conv2d_8_constant_3_next_constant_data), .B(conv2d_8_stream_pad_masks), .S(_set_flag_538), .Y(_24253_) );
  \$mux  #( .WIDTH(2) ) _45507_ ( .A(_stream_conv2d_8_constant_2_next_constant_data), .B(conv2d_8_row_select_buf), .S(_set_flag_538), .Y(_24254_) );
  \$mux  #( .WIDTH(2) ) _45509_ ( .A(_stream_conv2d_8_constant_1_next_constant_data), .B(conv2d_8_col_select), .S(_set_flag_538), .Y(_24255_) );
  \$mux  #( .WIDTH(5) ) _45511_ ( .A(_stream_conv2d_8_constant_0_next_constant_data), .B(cparam_conv2d_8_stream_reduce_size), .S(_set_flag_538), .Y(_24256_) );
  \$mux  #( .WIDTH(1) ) _45513_ ( .A(_substream__reduce_max_13_size_data_cond_772_43), .B(1'h1), .S(__tmp_884_7), .Y(_24257_) );
  \$mux  #( .WIDTH(1) ) _45514_ ( .A(_24257_), .B(1'h0), .S(__tmp_908_4), .Y(_24258_) );
  \$mux  #( .WIDTH(1) ) _45516_ ( .A(_substream__reduce_max_13_x_data_cond_772_42), .B(1'h1), .S(__tmp_884_7), .Y(_24259_) );
  \$mux  #( .WIDTH(1) ) _45517_ ( .A(_24259_), .B(1'h0), .S(__tmp_908_4), .Y(_24260_) );
  \$mux  #( .WIDTH(1) ) _45519_ ( .A(__reduce_max_13_reduce_reset), .B(1'h0), .S(__tmp_880_9), .Y(_24261_) );
  \$mux  #( .WIDTH(1) ) _45520_ ( .A(_24261_), .B(1'h1), .S(__tmp_908_5), .Y(_24262_) );
  \$mux  #( .WIDTH(1) ) _45521_ ( .A(_24262_), .B(1'h1), .S(RST), .Y(_00620_) );
  \$mux  #( .WIDTH(8) ) _45527_ ( .A(__variable_wdata_188), .B({ 5'h00, __delay_data_1377 }), .S(_substream__reduce_max_13_size_data_cond_772_43), .Y(_24263_) );
  \$mux  #( .WIDTH(8) ) _45529_ ( .A(__variable_wdata_187), .B(_cond_data_771[7:0]), .S(_substream__reduce_max_13_x_data_cond_772_42), .Y(_24264_) );
  \$mux  #( .WIDTH(9) ) _45531_ ( .A(_26541_[8:0]), .B(9'h000), .S(__reduce_max_13_reduce_reset), .Y(_24265_) );
  \$mux  #( .WIDTH(9) ) _45534_ ( .A(_26540_[8:0]), .B(9'h000), .S(__reduce_max_13_reduce_reset), .Y(_24266_) );
  \$mux  #( .WIDTH(32) ) _45536_ ( .A(_26539_), .B({ __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187 }), .S(__reduce_max_13_reduce_reset), .Y(_24267_) );
  \$mux  #( .WIDTH(32) ) _45537_ ( .A({ __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187 }), .B(_24267_), .S(_04892_), .Y(_24268_) );
  \$mux  #( .WIDTH(32) ) _45538_ ( .A(_24268_), .B(-128), .S(RST), .Y(_01714_) );
  \$mux  #( .WIDTH(1) ) _45539_ ( .A(_substream_mul_12_rshift_data_cond_708_26), .B(1'h1), .S(__tmp_627_12), .Y(_24269_) );
  \$mux  #( .WIDTH(1) ) _45540_ ( .A(_24269_), .B(1'h0), .S(__tmp_775_9), .Y(_24270_) );
  \$mux  #( .WIDTH(1) ) _45542_ ( .A(_substream_mul_12_y_data_cond_708_25), .B(1'h1), .S(__tmp_627_12), .Y(_24271_) );
  \$mux  #( .WIDTH(1) ) _45543_ ( .A(_24271_), .B(1'h0), .S(__tmp_775_9), .Y(_24272_) );
  \$mux  #( .WIDTH(1) ) _45545_ ( .A(_substream_mul_12_x_data_cond_708_24), .B(1'h1), .S(__tmp_627_12), .Y(_24273_) );
  \$mux  #( .WIDTH(1) ) _45546_ ( .A(_24273_), .B(1'h0), .S(__tmp_775_9), .Y(_24274_) );
  \$mux  #( .WIDTH(4) ) _45548_ ( .A(__variable_wdata_174), .B(__delay_data_1228[3:0]), .S(_substream_mul_12_rshift_data_cond_708_26), .Y(_24275_) );
  \$mux  #( .WIDTH(8) ) _45550_ ( .A(__variable_wdata_173), .B(__delay_data_1222), .S(_substream_mul_12_y_data_cond_708_25), .Y(_24276_) );
  \$mux  #( .WIDTH(8) ) _45552_ ( .A(__variable_wdata_172), .B(_cond_data_571), .S(_substream_mul_12_x_data_cond_708_24), .Y(_24277_) );
  \$mux  #( .WIDTH(1) ) _45574_ ( .A(_substream_mul_11_rshift_data_cond_691_23), .B(1'h1), .S(__tmp_627_12), .Y(_24278_) );
  \$mux  #( .WIDTH(1) ) _45575_ ( .A(_24278_), .B(1'h0), .S(__tmp_775_9), .Y(_24279_) );
  \$mux  #( .WIDTH(1) ) _45577_ ( .A(_substream_mul_11_y_data_cond_691_22), .B(1'h1), .S(__tmp_627_12), .Y(_24280_) );
  \$mux  #( .WIDTH(1) ) _45578_ ( .A(_24280_), .B(1'h0), .S(__tmp_775_9), .Y(_24281_) );
  \$mux  #( .WIDTH(1) ) _45580_ ( .A(_substream_mul_11_x_data_cond_691_21), .B(1'h1), .S(__tmp_627_12), .Y(_24282_) );
  \$mux  #( .WIDTH(1) ) _45581_ ( .A(_24282_), .B(1'h0), .S(__tmp_775_9), .Y(_24283_) );
  \$mux  #( .WIDTH(4) ) _45583_ ( .A(__variable_wdata_159), .B(__delay_data_1228[3:0]), .S(_substream_mul_11_rshift_data_cond_691_23), .Y(_24284_) );
  \$mux  #( .WIDTH(8) ) _45585_ ( .A(__variable_wdata_158), .B(__delay_data_1189), .S(_substream_mul_11_y_data_cond_691_22), .Y(_24285_) );
  \$mux  #( .WIDTH(8) ) _45587_ ( .A(__variable_wdata_157), .B(_cond_data_569), .S(_substream_mul_11_x_data_cond_691_21), .Y(_24286_) );
  \$mux  #( .WIDTH(1) ) _45609_ ( .A(_substream_mul_10_rshift_data_cond_674_20), .B(1'h1), .S(__tmp_627_12), .Y(_24287_) );
  \$mux  #( .WIDTH(1) ) _45610_ ( .A(_24287_), .B(1'h0), .S(__tmp_775_9), .Y(_24288_) );
  \$mux  #( .WIDTH(1) ) _45612_ ( .A(_substream_mul_10_y_data_cond_674_19), .B(1'h1), .S(__tmp_627_12), .Y(_24289_) );
  \$mux  #( .WIDTH(1) ) _45613_ ( .A(_24289_), .B(1'h0), .S(__tmp_775_9), .Y(_24290_) );
  \$mux  #( .WIDTH(1) ) _45615_ ( .A(_substream_mul_10_x_data_cond_674_18), .B(1'h1), .S(__tmp_627_12), .Y(_24291_) );
  \$mux  #( .WIDTH(1) ) _45616_ ( .A(_24291_), .B(1'h0), .S(__tmp_775_9), .Y(_24292_) );
  \$mux  #( .WIDTH(4) ) _45620_ ( .A(__variable_wdata_144), .B(__delay_data_1228[3:0]), .S(_substream_mul_10_rshift_data_cond_674_20), .Y(_24293_) );
  \$mux  #( .WIDTH(8) ) _45622_ ( .A(__variable_wdata_143), .B(__delay_data_1156), .S(_substream_mul_10_y_data_cond_674_19), .Y(_24294_) );
  \$mux  #( .WIDTH(8) ) _45624_ ( .A(__variable_wdata_142), .B(_cond_data_567), .S(_substream_mul_10_x_data_cond_674_18), .Y(_24295_) );
  \$mux  #( .WIDTH(1) ) _45646_ ( .A(_substream_mul_9_rshift_data_cond_657_17), .B(1'h1), .S(__tmp_627_12), .Y(_24296_) );
  \$mux  #( .WIDTH(1) ) _45647_ ( .A(_24296_), .B(1'h0), .S(__tmp_775_9), .Y(_24297_) );
  \$mux  #( .WIDTH(1) ) _45649_ ( .A(_substream_mul_9_y_data_cond_657_16), .B(1'h1), .S(__tmp_627_12), .Y(_24298_) );
  \$mux  #( .WIDTH(1) ) _45650_ ( .A(_24298_), .B(1'h0), .S(__tmp_775_9), .Y(_24299_) );
  \$mux  #( .WIDTH(1) ) _45652_ ( .A(_substream_mul_9_x_data_cond_657_15), .B(1'h1), .S(__tmp_627_12), .Y(_24300_) );
  \$mux  #( .WIDTH(1) ) _45653_ ( .A(_24300_), .B(1'h0), .S(__tmp_775_9), .Y(_24301_) );
  \$mux  #( .WIDTH(4) ) _45655_ ( .A(__variable_wdata_129), .B(__delay_data_1228[3:0]), .S(_substream_mul_9_rshift_data_cond_657_17), .Y(_24302_) );
  \$mux  #( .WIDTH(8) ) _45657_ ( .A(__variable_wdata_128), .B(__delay_data_1123), .S(_substream_mul_9_y_data_cond_657_16), .Y(_24303_) );
  \$mux  #( .WIDTH(8) ) _45659_ ( .A(__variable_wdata_127), .B(_cond_data_565), .S(_substream_mul_9_x_data_cond_657_15), .Y(_24304_) );
  \$mux  #( .WIDTH(1) ) _45681_ ( .A(_substream_mul_8_rshift_data_cond_640_14), .B(1'h1), .S(__tmp_627_12), .Y(_24305_) );
  \$mux  #( .WIDTH(1) ) _45682_ ( .A(_24305_), .B(1'h0), .S(__tmp_775_9), .Y(_24306_) );
  \$mux  #( .WIDTH(1) ) _45684_ ( .A(_substream_mul_8_y_data_cond_640_13), .B(1'h1), .S(__tmp_627_12), .Y(_24307_) );
  \$mux  #( .WIDTH(1) ) _45685_ ( .A(_24307_), .B(1'h0), .S(__tmp_775_9), .Y(_24308_) );
  \$mux  #( .WIDTH(1) ) _45687_ ( .A(_substream_mul_8_x_data_cond_640_12), .B(1'h1), .S(__tmp_627_12), .Y(_24309_) );
  \$mux  #( .WIDTH(1) ) _45688_ ( .A(_24309_), .B(1'h0), .S(__tmp_775_9), .Y(_24310_) );
  \$mux  #( .WIDTH(4) ) _45690_ ( .A(__variable_wdata_114), .B(__delay_data_1228[3:0]), .S(_substream_mul_8_rshift_data_cond_640_14), .Y(_24311_) );
  \$mux  #( .WIDTH(8) ) _45692_ ( .A(__variable_wdata_113), .B(__delay_data_1089), .S(_substream_mul_8_y_data_cond_640_13), .Y(_24312_) );
  \$mux  #( .WIDTH(8) ) _45694_ ( .A(__variable_wdata_112), .B(_cond_data_563), .S(_substream_mul_8_x_data_cond_640_12), .Y(_24313_) );
  \$mux  #( .WIDTH(1) ) _45716_ ( .A(_substream_mul_7_rshift_data_cond_623_11), .B(1'h1), .S(__tmp_627_12), .Y(_24314_) );
  \$mux  #( .WIDTH(1) ) _45717_ ( .A(_24314_), .B(1'h0), .S(__tmp_775_9), .Y(_24315_) );
  \$mux  #( .WIDTH(1) ) _45719_ ( .A(_substream_mul_7_y_data_cond_623_10), .B(1'h1), .S(__tmp_627_12), .Y(_24316_) );
  \$mux  #( .WIDTH(1) ) _45720_ ( .A(_24316_), .B(1'h0), .S(__tmp_775_9), .Y(_24317_) );
  \$mux  #( .WIDTH(1) ) _45722_ ( .A(_substream_mul_7_x_data_cond_623_9), .B(1'h1), .S(__tmp_627_12), .Y(_24318_) );
  \$mux  #( .WIDTH(1) ) _45723_ ( .A(_24318_), .B(1'h0), .S(__tmp_775_9), .Y(_24319_) );
  \$mux  #( .WIDTH(4) ) _45725_ ( .A(__variable_wdata_99), .B(__delay_data_1228[3:0]), .S(_substream_mul_7_rshift_data_cond_623_11), .Y(_24320_) );
  \$mux  #( .WIDTH(8) ) _45727_ ( .A(__variable_wdata_98), .B(__delay_data_1055), .S(_substream_mul_7_y_data_cond_623_10), .Y(_24321_) );
  \$mux  #( .WIDTH(8) ) _45729_ ( .A(__variable_wdata_97), .B(_cond_data_561), .S(_substream_mul_7_x_data_cond_623_9), .Y(_24322_) );
  \$mux  #( .WIDTH(1) ) _45751_ ( .A(_substream_mul_6_rshift_data_cond_606_8), .B(1'h1), .S(__tmp_627_12), .Y(_24323_) );
  \$mux  #( .WIDTH(1) ) _45752_ ( .A(_24323_), .B(1'h0), .S(__tmp_775_9), .Y(_24324_) );
  \$mux  #( .WIDTH(1) ) _45754_ ( .A(_substream_mul_6_y_data_cond_606_7), .B(1'h1), .S(__tmp_627_12), .Y(_24325_) );
  \$mux  #( .WIDTH(1) ) _45755_ ( .A(_24325_), .B(1'h0), .S(__tmp_775_9), .Y(_24326_) );
  \$mux  #( .WIDTH(1) ) _45757_ ( .A(_substream_mul_6_x_data_cond_606_6), .B(1'h1), .S(__tmp_627_12), .Y(_24327_) );
  \$mux  #( .WIDTH(1) ) _45758_ ( .A(_24327_), .B(1'h0), .S(__tmp_775_9), .Y(_24328_) );
  \$mux  #( .WIDTH(4) ) _45761_ ( .A(__variable_wdata_84), .B(__delay_data_1228[3:0]), .S(_substream_mul_6_rshift_data_cond_606_8), .Y(_24329_) );
  \$mux  #( .WIDTH(8) ) _45763_ ( .A(__variable_wdata_83), .B(__delay_data_1021), .S(_substream_mul_6_y_data_cond_606_7), .Y(_24330_) );
  \$mux  #( .WIDTH(8) ) _45765_ ( .A(__variable_wdata_82), .B(_cond_data_559), .S(_substream_mul_6_x_data_cond_606_6), .Y(_24331_) );
  \$mux  #( .WIDTH(1) ) _45787_ ( .A(_substream_mul_5_rshift_data_cond_589_5), .B(1'h1), .S(__tmp_627_12), .Y(_24332_) );
  \$mux  #( .WIDTH(1) ) _45788_ ( .A(_24332_), .B(1'h0), .S(__tmp_775_9), .Y(_24333_) );
  \$mux  #( .WIDTH(1) ) _45790_ ( .A(_substream_mul_5_y_data_cond_589_4), .B(1'h1), .S(__tmp_627_12), .Y(_24334_) );
  \$mux  #( .WIDTH(1) ) _45791_ ( .A(_24334_), .B(1'h0), .S(__tmp_775_9), .Y(_24335_) );
  \$mux  #( .WIDTH(1) ) _45793_ ( .A(_substream_mul_5_x_data_cond_589_3), .B(1'h1), .S(__tmp_627_12), .Y(_24336_) );
  \$mux  #( .WIDTH(1) ) _45794_ ( .A(_24336_), .B(1'h0), .S(__tmp_775_9), .Y(_24337_) );
  \$mux  #( .WIDTH(4) ) _45796_ ( .A(__variable_wdata_69), .B(__delay_data_1228[3:0]), .S(_substream_mul_5_rshift_data_cond_589_5), .Y(_24338_) );
  \$mux  #( .WIDTH(8) ) _45798_ ( .A(__variable_wdata_68), .B(__delay_data_974), .S(_substream_mul_5_y_data_cond_589_4), .Y(_24339_) );
  \$mux  #( .WIDTH(8) ) _45800_ ( .A(__variable_wdata_67), .B(_cond_data_557), .S(_substream_mul_5_x_data_cond_589_3), .Y(_24340_) );
  \$mux  #( .WIDTH(1) ) _45822_ ( .A(_substream_mul_4_rshift_data_cond_854_46), .B(1'h1), .S(__tmp_1059_8), .Y(_24341_) );
  \$mux  #( .WIDTH(1) ) _45823_ ( .A(_24341_), .B(1'h0), .S(__tmp_1095_5), .Y(_24342_) );
  \$mux  #( .WIDTH(1) ) _45825_ ( .A(_substream_mul_4_y_data_cond_854_45), .B(1'h1), .S(__tmp_1059_8), .Y(_24343_) );
  \$mux  #( .WIDTH(1) ) _45826_ ( .A(_24343_), .B(1'h0), .S(__tmp_1095_5), .Y(_24344_) );
  \$mux  #( .WIDTH(1) ) _45828_ ( .A(_substream_mul_4_x_data_cond_854_44), .B(1'h1), .S(__tmp_1059_8), .Y(_24345_) );
  \$mux  #( .WIDTH(1) ) _45829_ ( .A(_24345_), .B(1'h0), .S(__tmp_1095_5), .Y(_24346_) );
  \$mux  #( .WIDTH(1) ) _45831_ ( .A(_substream_mul_4_rshift_data_cond_572_2), .B(1'h1), .S(__tmp_627_12), .Y(_24347_) );
  \$mux  #( .WIDTH(1) ) _45832_ ( .A(_24347_), .B(1'h0), .S(__tmp_775_9), .Y(_24348_) );
  \$mux  #( .WIDTH(1) ) _45834_ ( .A(_substream_mul_4_y_data_cond_572_1), .B(1'h1), .S(__tmp_627_12), .Y(_24349_) );
  \$mux  #( .WIDTH(1) ) _45835_ ( .A(_24349_), .B(1'h0), .S(__tmp_775_9), .Y(_24350_) );
  \$mux  #( .WIDTH(1) ) _45837_ ( .A(_substream_mul_4_x_data_cond_572_0), .B(1'h1), .S(__tmp_627_12), .Y(_24351_) );
  \$mux  #( .WIDTH(1) ) _45838_ ( .A(_24351_), .B(1'h0), .S(__tmp_775_9), .Y(_24352_) );
  \$mux  #( .WIDTH(4) ) _45840_ ( .A(__variable_wdata_54), .B(__delay_data_1228[3:0]), .S(_substream_mul_4_rshift_data_cond_572_2), .Y(_24353_) );
  \$mux  #( .WIDTH(4) ) _45841_ ( .A(_24353_), .B(__delay_data_1388[3:0]), .S(_substream_mul_4_rshift_data_cond_854_46), .Y(_24354_) );
  \$mux  #( .WIDTH(8) ) _45843_ ( .A(__variable_wdata_53), .B(__delay_data_924), .S(_substream_mul_4_y_data_cond_572_1), .Y(_24355_) );
  \$mux  #( .WIDTH(8) ) _45844_ ( .A(_24355_), .B(__delay_data_1386), .S(_substream_mul_4_y_data_cond_854_45), .Y(_24356_) );
  \$mux  #( .WIDTH(8) ) _45846_ ( .A(__variable_wdata_52), .B(_cond_data_555), .S(_substream_mul_4_x_data_cond_572_0), .Y(_24357_) );
  \$mux  #( .WIDTH(8) ) _45847_ ( .A(_24357_), .B(_cond_data_853), .S(_substream_mul_4_x_data_cond_854_44), .Y(_24358_) );
  \$mux  #( .WIDTH(1) ) _45869_ ( .A(_substream_mul_rshift_clip_3_rshift_data_cond_864_53), .B(1'h1), .S(__tmp_1059_28), .Y(_24359_) );
  \$mux  #( .WIDTH(1) ) _45870_ ( .A(_24359_), .B(1'h0), .S(__tmp_1117_25), .Y(_24360_) );
  \$mux  #( .WIDTH(1) ) _45872_ ( .A(_substream_mul_rshift_clip_3_y_data_cond_864_52), .B(1'h1), .S(__tmp_1059_28), .Y(_24361_) );
  \$mux  #( .WIDTH(1) ) _45873_ ( .A(_24361_), .B(1'h0), .S(__tmp_1117_25), .Y(_24362_) );
  \$mux  #( .WIDTH(1) ) _45875_ ( .A(_substream_mul_rshift_clip_3_x_data_cond_864_51), .B(1'h1), .S(__tmp_1059_28), .Y(_24363_) );
  \$mux  #( .WIDTH(1) ) _45876_ ( .A(_24363_), .B(1'h0), .S(__tmp_1117_25), .Y(_24364_) );
  \$mux  #( .WIDTH(1) ) _45878_ ( .A(_substream_mul_rshift_clip_3_rshift_data_cond_743_41), .B(1'h1), .S(__tmp_627_34), .Y(_24365_) );
  \$mux  #( .WIDTH(1) ) _45879_ ( .A(_24365_), .B(1'h0), .S(__tmp_797_31), .Y(_24366_) );
  \$mux  #( .WIDTH(1) ) _45881_ ( .A(_substream_mul_rshift_clip_3_y_data_cond_743_40), .B(1'h1), .S(__tmp_627_34), .Y(_24367_) );
  \$mux  #( .WIDTH(1) ) _45882_ ( .A(_24367_), .B(1'h0), .S(__tmp_797_31), .Y(_24368_) );
  \$mux  #( .WIDTH(1) ) _45884_ ( .A(_substream_mul_rshift_clip_3_x_data_cond_743_39), .B(1'h1), .S(__tmp_627_34), .Y(_24369_) );
  \$mux  #( .WIDTH(1) ) _45885_ ( .A(_24369_), .B(1'h0), .S(__tmp_797_31), .Y(_24370_) );
  \$mux  #( .WIDTH(6) ) _45900_ ( .A(__variable_wdata_38), .B(__delay_data_1357[5:0]), .S(_substream_mul_rshift_clip_3_rshift_data_cond_743_41), .Y(_24371_) );
  \$mux  #( .WIDTH(6) ) _45901_ ( .A(_24371_), .B(__delay_data_1487[5:0]), .S(_substream_mul_rshift_clip_3_rshift_data_cond_864_53), .Y(_24372_) );
  \$mux  #( .WIDTH(8) ) _45903_ ( .A(__variable_wdata_37), .B(__delay_data_1329), .S(_substream_mul_rshift_clip_3_y_data_cond_743_40), .Y(_24373_) );
  \$mux  #( .WIDTH(8) ) _45904_ ( .A(_24373_), .B(__delay_data_1465), .S(_substream_mul_rshift_clip_3_y_data_cond_864_52), .Y(_24374_) );
  \$mux  #( .WIDTH(32) ) _45906_ ( .A(__variable_wdata_36), .B(_plus_data_742), .S(_substream_mul_rshift_clip_3_x_data_cond_743_39), .Y(_24375_) );
  \$mux  #( .WIDTH(32) ) _45907_ ( .A(_24375_), .B(_plus_data_863), .S(_substream_mul_rshift_clip_3_x_data_cond_864_51), .Y(_24376_) );
  \$mux  #( .WIDTH(1) ) _45923_ ( .A(_substream_add_tree_2_var8_data_cond_725_35), .B(1'h1), .S(__tmp_627_22), .Y(_24377_) );
  \$mux  #( .WIDTH(1) ) _45924_ ( .A(_24377_), .B(1'h0), .S(__tmp_797_19), .Y(_24378_) );
  \$mux  #( .WIDTH(1) ) _45926_ ( .A(_substream_add_tree_2_var7_data_cond_725_34), .B(1'h1), .S(__tmp_627_22), .Y(_24379_) );
  \$mux  #( .WIDTH(1) ) _45927_ ( .A(_24379_), .B(1'h0), .S(__tmp_797_19), .Y(_24380_) );
  \$mux  #( .WIDTH(1) ) _45929_ ( .A(_substream_add_tree_2_var6_data_cond_725_33), .B(1'h1), .S(__tmp_627_22), .Y(_24381_) );
  \$mux  #( .WIDTH(1) ) _45930_ ( .A(_24381_), .B(1'h0), .S(__tmp_797_19), .Y(_24382_) );
  \$mux  #( .WIDTH(1) ) _45932_ ( .A(_substream_add_tree_2_var5_data_cond_725_32), .B(1'h1), .S(__tmp_627_22), .Y(_24383_) );
  \$mux  #( .WIDTH(1) ) _45933_ ( .A(_24383_), .B(1'h0), .S(__tmp_797_19), .Y(_24384_) );
  \$mux  #( .WIDTH(1) ) _45935_ ( .A(_substream_add_tree_2_var4_data_cond_725_31), .B(1'h1), .S(__tmp_627_22), .Y(_24385_) );
  \$mux  #( .WIDTH(1) ) _45936_ ( .A(_24385_), .B(1'h0), .S(__tmp_797_19), .Y(_24386_) );
  \$mux  #( .WIDTH(1) ) _45938_ ( .A(_substream_add_tree_2_var3_data_cond_725_30), .B(1'h1), .S(__tmp_627_22), .Y(_24387_) );
  \$mux  #( .WIDTH(1) ) _45939_ ( .A(_24387_), .B(1'h0), .S(__tmp_797_19), .Y(_24388_) );
  \$mux  #( .WIDTH(1) ) _45941_ ( .A(_substream_add_tree_2_var2_data_cond_725_29), .B(1'h1), .S(__tmp_627_22), .Y(_24389_) );
  \$mux  #( .WIDTH(1) ) _45942_ ( .A(_24389_), .B(1'h0), .S(__tmp_797_19), .Y(_24390_) );
  \$mux  #( .WIDTH(1) ) _45944_ ( .A(_substream_add_tree_2_var1_data_cond_725_28), .B(1'h1), .S(__tmp_627_22), .Y(_24391_) );
  \$mux  #( .WIDTH(1) ) _45945_ ( .A(_24391_), .B(1'h0), .S(__tmp_797_19), .Y(_24392_) );
  \$mux  #( .WIDTH(1) ) _45947_ ( .A(_substream_add_tree_2_var0_data_cond_725_27), .B(1'h1), .S(__tmp_627_22), .Y(_24393_) );
  \$mux  #( .WIDTH(1) ) _45948_ ( .A(_24393_), .B(1'h0), .S(__tmp_797_19), .Y(_24394_) );
  \$mux  #( .WIDTH(32) ) _45950_ ( .A(__variable_wdata_30), .B({ __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724[15], __substreamoutput_data_724 }), .S(_substream_add_tree_2_var8_data_cond_725_35), .Y(_24395_) );
  \$mux  #( .WIDTH(32) ) _45952_ ( .A(__variable_wdata_29), .B({ __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707[15], __substreamoutput_data_707 }), .S(_substream_add_tree_2_var7_data_cond_725_34), .Y(_24396_) );
  \$mux  #( .WIDTH(32) ) _45954_ ( .A(__variable_wdata_28), .B({ __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690[15], __substreamoutput_data_690 }), .S(_substream_add_tree_2_var6_data_cond_725_33), .Y(_24397_) );
  \$mux  #( .WIDTH(32) ) _45956_ ( .A(__variable_wdata_27), .B({ __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673[15], __substreamoutput_data_673 }), .S(_substream_add_tree_2_var5_data_cond_725_32), .Y(_24398_) );
  \$mux  #( .WIDTH(32) ) _45958_ ( .A(__variable_wdata_26), .B({ __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656[15], __substreamoutput_data_656 }), .S(_substream_add_tree_2_var4_data_cond_725_31), .Y(_24399_) );
  \$mux  #( .WIDTH(32) ) _45960_ ( .A(__variable_wdata_25), .B({ __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639[15], __substreamoutput_data_639 }), .S(_substream_add_tree_2_var3_data_cond_725_30), .Y(_24400_) );
  \$mux  #( .WIDTH(32) ) _45962_ ( .A(__variable_wdata_24), .B({ __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622[15], __substreamoutput_data_622 }), .S(_substream_add_tree_2_var2_data_cond_725_29), .Y(_24401_) );
  \$mux  #( .WIDTH(32) ) _45964_ ( .A(__variable_wdata_23), .B({ __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605[15], __substreamoutput_data_605 }), .S(_substream_add_tree_2_var1_data_cond_725_28), .Y(_24402_) );
  \$mux  #( .WIDTH(32) ) _45966_ ( .A(__variable_wdata_22), .B({ __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856 }), .S(_substream_add_tree_2_var0_data_cond_725_27), .Y(_24403_) );
  \$mux  #( .WIDTH(1) ) _45972_ ( .A(_substream_add_tree_1_var0_data_cond_857_47), .B(1'h1), .S(__tmp_1059_18), .Y(_24404_) );
  \$mux  #( .WIDTH(1) ) _45973_ ( .A(_24404_), .B(1'h0), .S(__tmp_1117_15), .Y(_24405_) );
  \$mux  #( .WIDTH(32) ) _45975_ ( .A(__variable_wdata_20), .B({ __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856[15], __substreamoutput_data_856 }), .S(_substream_add_tree_1_var0_data_cond_857_47), .Y(_24406_) );
  \$mux  #( .WIDTH(1) ) _45977_ ( .A(_substream_acc_0_size_data_cond_859_50), .B(1'h1), .S(__tmp_1059_20), .Y(_24407_) );
  \$mux  #( .WIDTH(1) ) _45978_ ( .A(_24407_), .B(1'h0), .S(__tmp_1117_17), .Y(_24408_) );
  \$mux  #( .WIDTH(1) ) _45980_ ( .A(_substream_acc_0_rshift_data_cond_859_49), .B(1'h1), .S(__tmp_1059_20), .Y(_24409_) );
  \$mux  #( .WIDTH(1) ) _45981_ ( .A(_24409_), .B(1'h0), .S(__tmp_1117_17), .Y(_24410_) );
  \$mux  #( .WIDTH(1) ) _45983_ ( .A(_substream_acc_0_x_data_cond_859_48), .B(1'h1), .S(__tmp_1059_20), .Y(_24411_) );
  \$mux  #( .WIDTH(1) ) _45984_ ( .A(_24411_), .B(1'h0), .S(__tmp_1117_17), .Y(_24412_) );
  \$mux  #( .WIDTH(1) ) _45986_ ( .A(_substream_acc_0_size_data_cond_727_38), .B(1'h1), .S(__tmp_627_26), .Y(_24413_) );
  \$mux  #( .WIDTH(1) ) _45987_ ( .A(_24413_), .B(1'h0), .S(__tmp_797_23), .Y(_24414_) );
  \$mux  #( .WIDTH(1) ) _45989_ ( .A(_substream_acc_0_rshift_data_cond_727_37), .B(1'h1), .S(__tmp_627_26), .Y(_24415_) );
  \$mux  #( .WIDTH(1) ) _45990_ ( .A(_24415_), .B(1'h0), .S(__tmp_797_23), .Y(_24416_) );
  \$mux  #( .WIDTH(1) ) _45992_ ( .A(_substream_acc_0_x_data_cond_727_36), .B(1'h1), .S(__tmp_627_26), .Y(_24417_) );
  \$mux  #( .WIDTH(1) ) _45993_ ( .A(_24417_), .B(1'h0), .S(__tmp_797_23), .Y(_24418_) );
  \$mux  #( .WIDTH(1) ) _45995_ ( .A(_acc_0_reduce_reset), .B(1'h0), .S(__tmp_627_28), .Y(_24419_) );
  \$mux  #( .WIDTH(1) ) _45996_ ( .A(_24419_), .B(1'h1), .S(__tmp_797_24), .Y(_24420_) );
  \$mux  #( .WIDTH(1) ) _45997_ ( .A(_24420_), .B(1'h0), .S(__tmp_1059_22), .Y(_24421_) );
  \$mux  #( .WIDTH(1) ) _45998_ ( .A(_24421_), .B(1'h1), .S(__tmp_1117_18), .Y(_24422_) );
  \$mux  #( .WIDTH(1) ) _45999_ ( .A(_24422_), .B(1'h1), .S(RST), .Y(_01356_) );
  \$mux  #( .WIDTH(32) ) _46008_ ( .A(__variable_wdata_2), .B({ 27'h0000000, __delay_data_1271 }), .S(_substream_acc_0_size_data_cond_727_38), .Y(_24423_) );
  \$mux  #( .WIDTH(32) ) _46009_ ( .A(_24423_), .B({ 23'h000000, __delay_data_1419 }), .S(_substream_acc_0_size_data_cond_859_50), .Y(_24424_) );
  \$mux  #( .WIDTH(6) ) _46011_ ( .A(__variable_wdata_1), .B(__delay_data_1249[5:0]), .S(_substream_acc_0_rshift_data_cond_727_37), .Y(_24425_) );
  \$mux  #( .WIDTH(6) ) _46012_ ( .A(_24425_), .B(__delay_data_1403[5:0]), .S(_substream_acc_0_rshift_data_cond_859_49), .Y(_24426_) );
  \$mux  #( .WIDTH(32) ) _46014_ ( .A(__variable_wdata_0), .B(__substreamoutput_data_726), .S(_substream_acc_0_x_data_cond_727_36), .Y(_24427_) );
  \$mux  #( .WIDTH(32) ) _46015_ ( .A(_24427_), .B(__substreamoutput_data_858), .S(_substream_acc_0_x_data_cond_859_48), .Y(_24428_) );
  \$mux  #( .WIDTH(33) ) _46032_ ( .A(_26512_), .B(33'h000000000), .S(_acc_0_reduce_reset), .Y(_24429_) );
  \$mux  #( .WIDTH(33) ) _46035_ ( .A(_26511_), .B(33'h000000000), .S(_acc_0_reduce_reset), .Y(_24430_) );
  \$mux  #( .WIDTH(32) ) _46037_ ( .A(_22122_), .B(__variable_wdata_0), .S(_acc_0_reduce_reset), .Y(_24431_) );
  \$mux  #( .WIDTH(32) ) _46038_ ( .A(__variable_wdata_0), .B(_24431_), .S(_04891_), .Y(_24432_) );
  \$mux  #( .WIDTH(1) ) _46044_ ( .A(_tmp_13), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24433_) );
  \$mux  #( .WIDTH(1) ) _46045_ ( .A(_24433_), .B(1'h1), .S(_05673_), .Y(_24434_) );
  \$mux  #( .WIDTH(34) ) _46047_ ( .A(_tmp_12), .B({ 1'h0, _maxi_read_size }), .S(_05672_), .Y(_24435_) );
  \$mux  #( .WIDTH(34) ) _46048_ ( .A(_24435_), .B(_26005_), .S(_05379_), .Y(_24436_) );
  \$mux  #( .WIDTH(1) ) _46050_ ( .A(ram_w32_l128_id0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24437_) );
  \$mux  #( .WIDTH(1) ) _46051_ ( .A(_24437_), .B(1'h1), .S(_05379_), .Y(_24438_) );
  \$mux  #( .WIDTH(32) ) _46053_ ( .A(ram_w32_l128_id0_1_wdata), .B(_dataflow__delay_data_132), .S(_05379_), .Y(_24439_) );
  \$mux  #( .WIDTH(7) ) _46055_ ( .A(ram_w32_l128_id0_1_addr), .B(_25939_[6:0]), .S(_05672_), .Y(_24440_) );
  \$mux  #( .WIDTH(7) ) _46056_ ( .A(_24440_), .B(_22121_[6:0]), .S(_05379_), .Y(_24441_) );
  \$mux  #( .WIDTH(7) ) _46058_ ( .A(ram_w32_l128_id0_0_addr), .B(_stream_conv2d_8_source_6_source_ram_raddr[6:0]), .S(_tmp_336), .Y(_24442_) );
  \$mux  #( .WIDTH(7) ) _46059_ ( .A(_24442_), .B(_stream_matmul_15_source_6_source_ram_raddr[6:0]), .S(_tmp_992), .Y(_24443_) );
  \$mux  #( .WIDTH(34) ) _46061_ ( .A(_tmp_846), .B(_25945_), .S(_05668_), .Y(_24444_) );
  \$mux  #( .WIDTH(34) ) _46062_ ( .A(_24444_), .B(_26004_), .S(_05669_), .Y(_24445_) );
  \$mux  #( .WIDTH(1) ) _46064_ ( .A(_tmp_845), .B(1'h0), .S(_05666_), .Y(_24446_) );
  \$mux  #( .WIDTH(1) ) _46065_ ( .A(_24446_), .B(_tmp_844), .S(_05667_), .Y(_24447_) );
  \$mux  #( .WIDTH(1) ) _46067_ ( .A(_tmp_844), .B(1'h0), .S(_05667_), .Y(_24448_) );
  \$mux  #( .WIDTH(1) ) _46068_ ( .A(_24448_), .B(_05151_), .S(_05668_), .Y(_24449_) );
  \$mux  #( .WIDTH(1) ) _46069_ ( .A(_24449_), .B(1'h0), .S(_05669_), .Y(_24450_) );
  \$mux  #( .WIDTH(1) ) _46070_ ( .A(_24450_), .B(1'h1), .S(_05670_), .Y(_24451_) );
  \$mux  #( .WIDTH(1) ) _46072_ ( .A(_tmp_843), .B(1'h0), .S(_05666_), .Y(_24452_) );
  \$mux  #( .WIDTH(1) ) _46073_ ( .A(_24452_), .B(1'h1), .S(_05667_), .Y(_24453_) );
  \$mux  #( .WIDTH(1) ) _46075_ ( .A(_tmp_842), .B(1'h0), .S(_05667_), .Y(_24454_) );
  \$mux  #( .WIDTH(1) ) _46076_ ( .A(_24454_), .B(1'h1), .S(_05668_), .Y(_24455_) );
  \$mux  #( .WIDTH(1) ) _46077_ ( .A(_24455_), .B(1'h1), .S(_05669_), .Y(_24456_) );
  \$mux  #( .WIDTH(1) ) _46081_ ( .A(_tmp_835), .B(1'h0), .S(_05666_), .Y(_24457_) );
  \$mux  #( .WIDTH(1) ) _46082_ ( .A(_24457_), .B(1'h1), .S(_05667_), .Y(_24458_) );
  \$mux  #( .WIDTH(9) ) _46085_ ( .A(ram_w8_l2048_id19_3_1_addr), .B(_maxi_write_local_addr[8:0]), .S(_05668_), .Y(_24459_) );
  \$mux  #( .WIDTH(9) ) _46086_ ( .A(_24459_), .B(_22120_[8:0]), .S(_05669_), .Y(_24460_) );
  \$mux  #( .WIDTH(1) ) _46088_ ( .A(ram_w8_l2048_id19_3_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id19_3_cond_0_1), .Y(_24461_) );
  \$mux  #( .WIDTH(1) ) _46089_ ( .A(_24461_), .B(1'h1), .S(_05665_), .Y(_24462_) );
  \$mux  #( .WIDTH(8) ) _46091_ ( .A(ram_w8_l2048_id19_3_0_wdata), .B(_stream_conv2d_8_sink_37_sink_wdata), .S(_05665_), .Y(_24463_) );
  \$mux  #( .WIDTH(9) ) _46093_ ( .A(ram_w8_l2048_id19_3_0_addr), .B(_stream_conv2d_8_sink_37_sink_waddr[10:2]), .S(_05665_), .Y(_24464_) );
  \$mux  #( .WIDTH(34) ) _46095_ ( .A(_tmp_834), .B(_25945_), .S(_05662_), .Y(_24465_) );
  \$mux  #( .WIDTH(34) ) _46096_ ( .A(_24465_), .B(_26003_), .S(_05663_), .Y(_24466_) );
  \$mux  #( .WIDTH(1) ) _46098_ ( .A(_tmp_833), .B(1'h0), .S(_05660_), .Y(_24467_) );
  \$mux  #( .WIDTH(1) ) _46099_ ( .A(_24467_), .B(_tmp_832), .S(_05661_), .Y(_24468_) );
  \$mux  #( .WIDTH(1) ) _46101_ ( .A(_tmp_832), .B(1'h0), .S(_05661_), .Y(_24469_) );
  \$mux  #( .WIDTH(1) ) _46102_ ( .A(_24469_), .B(_05151_), .S(_05662_), .Y(_24470_) );
  \$mux  #( .WIDTH(1) ) _46103_ ( .A(_24470_), .B(1'h0), .S(_05663_), .Y(_24471_) );
  \$mux  #( .WIDTH(1) ) _46104_ ( .A(_24471_), .B(1'h1), .S(_05664_), .Y(_24472_) );
  \$mux  #( .WIDTH(1) ) _46106_ ( .A(_tmp_831), .B(1'h0), .S(_05660_), .Y(_24473_) );
  \$mux  #( .WIDTH(1) ) _46107_ ( .A(_24473_), .B(1'h1), .S(_05661_), .Y(_24474_) );
  \$mux  #( .WIDTH(1) ) _46109_ ( .A(_tmp_830), .B(1'h0), .S(_05661_), .Y(_24475_) );
  \$mux  #( .WIDTH(1) ) _46110_ ( .A(_24475_), .B(1'h1), .S(_05662_), .Y(_24476_) );
  \$mux  #( .WIDTH(1) ) _46111_ ( .A(_24476_), .B(1'h1), .S(_05663_), .Y(_24477_) );
  \$mux  #( .WIDTH(1) ) _46115_ ( .A(_tmp_823), .B(1'h0), .S(_05660_), .Y(_24478_) );
  \$mux  #( .WIDTH(1) ) _46116_ ( .A(_24478_), .B(1'h1), .S(_05661_), .Y(_24479_) );
  \$mux  #( .WIDTH(9) ) _46119_ ( .A(ram_w8_l2048_id19_2_1_addr), .B(_maxi_write_local_addr[8:0]), .S(_05662_), .Y(_24480_) );
  \$mux  #( .WIDTH(9) ) _46120_ ( .A(_24480_), .B(_22119_[8:0]), .S(_05663_), .Y(_24481_) );
  \$mux  #( .WIDTH(1) ) _46122_ ( .A(ram_w8_l2048_id19_2_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id19_2_cond_0_1), .Y(_24482_) );
  \$mux  #( .WIDTH(1) ) _46123_ ( .A(_24482_), .B(1'h1), .S(_05659_), .Y(_24483_) );
  \$mux  #( .WIDTH(8) ) _46125_ ( .A(ram_w8_l2048_id19_2_0_wdata), .B(_stream_conv2d_8_sink_37_sink_wdata), .S(_05659_), .Y(_24484_) );
  \$mux  #( .WIDTH(9) ) _46127_ ( .A(ram_w8_l2048_id19_2_0_addr), .B(_stream_conv2d_8_sink_37_sink_waddr[10:2]), .S(_05659_), .Y(_24485_) );
  \$mux  #( .WIDTH(34) ) _46129_ ( .A(_tmp_822), .B(_25945_), .S(_05656_), .Y(_24486_) );
  \$mux  #( .WIDTH(34) ) _46130_ ( .A(_24486_), .B(_26002_), .S(_05657_), .Y(_24487_) );
  \$mux  #( .WIDTH(1) ) _46132_ ( .A(_tmp_821), .B(1'h0), .S(_05654_), .Y(_24488_) );
  \$mux  #( .WIDTH(1) ) _46133_ ( .A(_24488_), .B(_tmp_820), .S(_05655_), .Y(_24489_) );
  \$mux  #( .WIDTH(1) ) _46135_ ( .A(_tmp_820), .B(1'h0), .S(_05655_), .Y(_24490_) );
  \$mux  #( .WIDTH(1) ) _46136_ ( .A(_24490_), .B(_05151_), .S(_05656_), .Y(_24491_) );
  \$mux  #( .WIDTH(1) ) _46137_ ( .A(_24491_), .B(1'h0), .S(_05657_), .Y(_24492_) );
  \$mux  #( .WIDTH(1) ) _46138_ ( .A(_24492_), .B(1'h1), .S(_05658_), .Y(_24493_) );
  \$mux  #( .WIDTH(1) ) _46140_ ( .A(_tmp_819), .B(1'h0), .S(_05654_), .Y(_24494_) );
  \$mux  #( .WIDTH(1) ) _46141_ ( .A(_24494_), .B(1'h1), .S(_05655_), .Y(_24495_) );
  \$mux  #( .WIDTH(1) ) _46143_ ( .A(_tmp_818), .B(1'h0), .S(_05655_), .Y(_24496_) );
  \$mux  #( .WIDTH(1) ) _46144_ ( .A(_24496_), .B(1'h1), .S(_05656_), .Y(_24497_) );
  \$mux  #( .WIDTH(1) ) _46145_ ( .A(_24497_), .B(1'h1), .S(_05657_), .Y(_24498_) );
  \$mux  #( .WIDTH(1) ) _46149_ ( .A(_tmp_811), .B(1'h0), .S(_05654_), .Y(_24499_) );
  \$mux  #( .WIDTH(1) ) _46150_ ( .A(_24499_), .B(1'h1), .S(_05655_), .Y(_24500_) );
  \$mux  #( .WIDTH(9) ) _46153_ ( .A(ram_w8_l2048_id19_1_1_addr), .B(_maxi_write_local_addr[8:0]), .S(_05656_), .Y(_24501_) );
  \$mux  #( .WIDTH(9) ) _46154_ ( .A(_24501_), .B(_22118_[8:0]), .S(_05657_), .Y(_24502_) );
  \$mux  #( .WIDTH(1) ) _46156_ ( .A(ram_w8_l2048_id19_1_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id19_1_cond_0_1), .Y(_24503_) );
  \$mux  #( .WIDTH(1) ) _46157_ ( .A(_24503_), .B(1'h1), .S(_05653_), .Y(_24504_) );
  \$mux  #( .WIDTH(8) ) _46159_ ( .A(ram_w8_l2048_id19_1_0_wdata), .B(_stream_conv2d_8_sink_37_sink_wdata), .S(_05653_), .Y(_24505_) );
  \$mux  #( .WIDTH(9) ) _46161_ ( .A(ram_w8_l2048_id19_1_0_addr), .B(_stream_conv2d_8_sink_37_sink_waddr[10:2]), .S(_05653_), .Y(_24506_) );
  \$mux  #( .WIDTH(1) ) _46163_ ( .A(_dataflow_cat_valid_74), .B(1'h0), .S(_05274_), .Y(_24507_) );
  \$mux  #( .WIDTH(1) ) _46164_ ( .A(_24507_), .B(_05651_), .S(_05652_), .Y(_24508_) );
  \$mux  #( .WIDTH(32) ) _46166_ ( .A(_dataflow_cat_data_74), .B({ _tmp_841, _tmp_829, _tmp_817, _tmp_805 }), .S(_05652_), .Y(_24509_) );
  \$mux  #( .WIDTH(34) ) _46168_ ( .A(_tmp_810), .B(_25945_), .S(_05648_), .Y(_24510_) );
  \$mux  #( .WIDTH(34) ) _46169_ ( .A(_24510_), .B(_26001_), .S(_05649_), .Y(_24511_) );
  \$mux  #( .WIDTH(1) ) _46171_ ( .A(_tmp_809), .B(1'h0), .S(_05645_), .Y(_24512_) );
  \$mux  #( .WIDTH(1) ) _46172_ ( .A(_24512_), .B(_tmp_808), .S(_05646_), .Y(_24513_) );
  \$mux  #( .WIDTH(1) ) _46174_ ( .A(_tmp_808), .B(1'h0), .S(_05646_), .Y(_24514_) );
  \$mux  #( .WIDTH(1) ) _46175_ ( .A(_24514_), .B(_05151_), .S(_05648_), .Y(_24515_) );
  \$mux  #( .WIDTH(1) ) _46176_ ( .A(_24515_), .B(1'h0), .S(_05649_), .Y(_24516_) );
  \$mux  #( .WIDTH(1) ) _46177_ ( .A(_24516_), .B(1'h1), .S(_05650_), .Y(_24517_) );
  \$mux  #( .WIDTH(1) ) _46179_ ( .A(_tmp_807), .B(1'h0), .S(_05645_), .Y(_24518_) );
  \$mux  #( .WIDTH(1) ) _46180_ ( .A(_24518_), .B(1'h1), .S(_05646_), .Y(_24519_) );
  \$mux  #( .WIDTH(1) ) _46182_ ( .A(_tmp_806), .B(1'h0), .S(_05646_), .Y(_24520_) );
  \$mux  #( .WIDTH(1) ) _46183_ ( .A(_24520_), .B(1'h1), .S(_05648_), .Y(_24521_) );
  \$mux  #( .WIDTH(1) ) _46184_ ( .A(_24521_), .B(1'h1), .S(_05649_), .Y(_24522_) );
  \$mux  #( .WIDTH(1) ) _46188_ ( .A(_tmp_799), .B(1'h0), .S(_05645_), .Y(_24523_) );
  \$mux  #( .WIDTH(1) ) _46189_ ( .A(_24523_), .B(1'h1), .S(_05646_), .Y(_24524_) );
  \$mux  #( .WIDTH(9) ) _46192_ ( .A(ram_w8_l2048_id19_0_1_addr), .B(_maxi_write_local_addr[8:0]), .S(_05648_), .Y(_24525_) );
  \$mux  #( .WIDTH(9) ) _46193_ ( .A(_24525_), .B(_22117_[8:0]), .S(_05649_), .Y(_24526_) );
  \$mux  #( .WIDTH(1) ) _46195_ ( .A(ram_w8_l2048_id19_0_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id19_0_cond_0_1), .Y(_24527_) );
  \$mux  #( .WIDTH(1) ) _46196_ ( .A(_24527_), .B(1'h1), .S(_05644_), .Y(_24528_) );
  \$mux  #( .WIDTH(8) ) _46198_ ( .A(ram_w8_l2048_id19_0_0_wdata), .B(_stream_conv2d_8_sink_37_sink_wdata), .S(_05644_), .Y(_24529_) );
  \$mux  #( .WIDTH(9) ) _46200_ ( .A(ram_w8_l2048_id19_0_0_addr), .B(_stream_conv2d_8_sink_37_sink_waddr[10:2]), .S(_05644_), .Y(_24530_) );
  \$mux  #( .WIDTH(1) ) _46202_ ( .A(ram_w8_l2048_id18_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24531_) );
  \$mux  #( .WIDTH(1) ) _46203_ ( .A(_24531_), .B(_05221_), .S(_05340_), .Y(_24532_) );
  \$mux  #( .WIDTH(8) ) _46205_ ( .A(ram_w8_l2048_id18_3_1_wdata), .B(_dataflow_slice_data_65), .S(_05340_), .Y(_24533_) );
  \$mux  #( .WIDTH(9) ) _46207_ ( .A(ram_w8_l2048_id18_3_1_addr), .B(_tmp_322), .S(_05340_), .Y(_24534_) );
  \$mux  #( .WIDTH(9) ) _46209_ ( .A(ram_w8_l2048_id18_3_0_addr), .B(_stream_conv2d_8_source_27_source_ram_raddr[10:2]), .S(_tmp_447), .Y(_24535_) );
  \$mux  #( .WIDTH(1) ) _46211_ ( .A(ram_w8_l2048_id18_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24536_) );
  \$mux  #( .WIDTH(1) ) _46212_ ( .A(_24536_), .B(_05218_), .S(_05337_), .Y(_24537_) );
  \$mux  #( .WIDTH(8) ) _46214_ ( .A(ram_w8_l2048_id18_2_1_wdata), .B(_dataflow_slice_data_62), .S(_05337_), .Y(_24538_) );
  \$mux  #( .WIDTH(9) ) _46216_ ( .A(ram_w8_l2048_id18_2_1_addr), .B(_tmp_309), .S(_05337_), .Y(_24539_) );
  \$mux  #( .WIDTH(9) ) _46218_ ( .A(ram_w8_l2048_id18_2_0_addr), .B(_stream_conv2d_8_source_27_source_ram_raddr[10:2]), .S(_tmp_447), .Y(_24540_) );
  \$mux  #( .WIDTH(1) ) _46220_ ( .A(ram_w8_l2048_id18_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24541_) );
  \$mux  #( .WIDTH(1) ) _46221_ ( .A(_24541_), .B(_05215_), .S(_05334_), .Y(_24542_) );
  \$mux  #( .WIDTH(8) ) _46223_ ( .A(ram_w8_l2048_id18_1_1_wdata), .B(_dataflow_slice_data_59), .S(_05334_), .Y(_24543_) );
  \$mux  #( .WIDTH(9) ) _46225_ ( .A(ram_w8_l2048_id18_1_1_addr), .B(_tmp_296), .S(_05334_), .Y(_24544_) );
  \$mux  #( .WIDTH(9) ) _46227_ ( .A(ram_w8_l2048_id18_1_0_addr), .B(_stream_conv2d_8_source_27_source_ram_raddr[10:2]), .S(_tmp_447), .Y(_24545_) );
  \$mux  #( .WIDTH(1) ) _46230_ ( .A(ram_w8_l2048_id18_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24546_) );
  \$mux  #( .WIDTH(1) ) _46231_ ( .A(_24546_), .B(_05212_), .S(_05331_), .Y(_24547_) );
  \$mux  #( .WIDTH(8) ) _46233_ ( .A(ram_w8_l2048_id18_0_1_wdata), .B(_dataflow_slice_data_56), .S(_05331_), .Y(_24548_) );
  \$mux  #( .WIDTH(9) ) _46235_ ( .A(ram_w8_l2048_id18_0_1_addr), .B(_tmp_283), .S(_05331_), .Y(_24549_) );
  \$mux  #( .WIDTH(9) ) _46237_ ( .A(ram_w8_l2048_id18_0_0_addr), .B(_stream_conv2d_8_source_27_source_ram_raddr[10:2]), .S(_tmp_447), .Y(_24550_) );
  \$mux  #( .WIDTH(1) ) _46239_ ( .A(ram_w8_l2048_id17_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24551_) );
  \$mux  #( .WIDTH(1) ) _46240_ ( .A(_24551_), .B(_05223_), .S(_05340_), .Y(_24552_) );
  \$mux  #( .WIDTH(8) ) _46242_ ( .A(ram_w8_l2048_id17_3_1_wdata), .B(_dataflow_slice_data_65), .S(_05340_), .Y(_24553_) );
  \$mux  #( .WIDTH(9) ) _46244_ ( .A(ram_w8_l2048_id17_3_1_addr), .B(_tmp_321), .S(_05340_), .Y(_24554_) );
  \$mux  #( .WIDTH(9) ) _46246_ ( .A(ram_w8_l2048_id17_3_0_addr), .B(_stream_conv2d_8_source_26_source_ram_raddr[10:2]), .S(_tmp_437), .Y(_24555_) );
  \$mux  #( .WIDTH(1) ) _46248_ ( .A(ram_w8_l2048_id17_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24556_) );
  \$mux  #( .WIDTH(1) ) _46249_ ( .A(_24556_), .B(_05220_), .S(_05337_), .Y(_24557_) );
  \$mux  #( .WIDTH(8) ) _46251_ ( .A(ram_w8_l2048_id17_2_1_wdata), .B(_dataflow_slice_data_62), .S(_05337_), .Y(_24558_) );
  \$mux  #( .WIDTH(9) ) _46253_ ( .A(ram_w8_l2048_id17_2_1_addr), .B(_tmp_308), .S(_05337_), .Y(_24559_) );
  \$mux  #( .WIDTH(9) ) _46255_ ( .A(ram_w8_l2048_id17_2_0_addr), .B(_stream_conv2d_8_source_26_source_ram_raddr[10:2]), .S(_tmp_437), .Y(_24560_) );
  \$mux  #( .WIDTH(1) ) _46257_ ( .A(ram_w8_l2048_id17_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24561_) );
  \$mux  #( .WIDTH(1) ) _46258_ ( .A(_24561_), .B(_05217_), .S(_05334_), .Y(_24562_) );
  \$mux  #( .WIDTH(8) ) _46260_ ( .A(ram_w8_l2048_id17_1_1_wdata), .B(_dataflow_slice_data_59), .S(_05334_), .Y(_24563_) );
  \$mux  #( .WIDTH(9) ) _46262_ ( .A(ram_w8_l2048_id17_1_1_addr), .B(_tmp_295), .S(_05334_), .Y(_24564_) );
  \$mux  #( .WIDTH(9) ) _46264_ ( .A(ram_w8_l2048_id17_1_0_addr), .B(_stream_conv2d_8_source_26_source_ram_raddr[10:2]), .S(_tmp_437), .Y(_24565_) );
  \$mux  #( .WIDTH(1) ) _46267_ ( .A(ram_w8_l2048_id17_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24566_) );
  \$mux  #( .WIDTH(1) ) _46268_ ( .A(_24566_), .B(_05214_), .S(_05331_), .Y(_24567_) );
  \$mux  #( .WIDTH(8) ) _46270_ ( .A(ram_w8_l2048_id17_0_1_wdata), .B(_dataflow_slice_data_56), .S(_05331_), .Y(_24568_) );
  \$mux  #( .WIDTH(9) ) _46272_ ( .A(ram_w8_l2048_id17_0_1_addr), .B(_tmp_282), .S(_05331_), .Y(_24569_) );
  \$mux  #( .WIDTH(9) ) _46274_ ( .A(ram_w8_l2048_id17_0_0_addr), .B(_stream_conv2d_8_source_26_source_ram_raddr[10:2]), .S(_tmp_437), .Y(_24570_) );
  \$mux  #( .WIDTH(2) ) _46276_ ( .A(_tmp_326), .B(2'h0), .S(_05637_), .Y(_24571_) );
  \$mux  #( .WIDTH(2) ) _46277_ ( .A(_24571_), .B(_22116_[1:0]), .S(_05638_), .Y(_24572_) );
  \$mux  #( .WIDTH(2) ) _46278_ ( .A(_24572_), .B(2'h0), .S(_05639_), .Y(_24573_) );
  \$mux  #( .WIDTH(9) ) _46280_ ( .A(_tmp_319), .B(_25939_[8:0]), .S(_05637_), .Y(_24574_) );
  \$mux  #( .WIDTH(9) ) _46281_ ( .A(_24574_), .B(_tmp_322), .S(_05642_), .Y(_24575_) );
  \$mux  #( .WIDTH(9) ) _46283_ ( .A(_tmp_318), .B(_25939_[8:0]), .S(_05637_), .Y(_24576_) );
  \$mux  #( .WIDTH(9) ) _46284_ ( .A(_24576_), .B(_tmp_321), .S(_05641_), .Y(_24577_) );
  \$mux  #( .WIDTH(9) ) _46286_ ( .A(_tmp_317), .B(_25939_[8:0]), .S(_05637_), .Y(_24578_) );
  \$mux  #( .WIDTH(9) ) _46287_ ( .A(_24578_), .B(_tmp_320), .S(_05640_), .Y(_24579_) );
  \$mux  #( .WIDTH(1) ) _46289_ ( .A(_tmp_316), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24580_) );
  \$mux  #( .WIDTH(1) ) _46290_ ( .A(_24580_), .B(1'h1), .S(_05643_), .Y(_24581_) );
  \$mux  #( .WIDTH(34) ) _46292_ ( .A(_tmp_315), .B({ 1'h0, _maxi_read_size }), .S(_05637_), .Y(_24582_) );
  \$mux  #( .WIDTH(34) ) _46293_ ( .A(_24582_), .B(_26000_), .S(_05340_), .Y(_24583_) );
  \$mux  #( .WIDTH(10) ) _46295_ ( .A(_tmp_314), .B(_25992_[9:0]), .S(_05637_), .Y(_24584_) );
  \$mux  #( .WIDTH(10) ) _46296_ ( .A(_24584_), .B(_25999_[9:0]), .S(_05340_), .Y(_24585_) );
  \$mux  #( .WIDTH(10) ) _46297_ ( .A(_24585_), .B(_25992_[9:0]), .S(_05638_), .Y(_24586_) );
  \$mux  #( .WIDTH(1) ) _46299_ ( .A(ram_w8_l2048_id16_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24587_) );
  \$mux  #( .WIDTH(1) ) _46300_ ( .A(_24587_), .B(_05222_), .S(_05340_), .Y(_24588_) );
  \$mux  #( .WIDTH(8) ) _46302_ ( .A(ram_w8_l2048_id16_3_1_wdata), .B(_dataflow_slice_data_65), .S(_05340_), .Y(_24589_) );
  \$mux  #( .WIDTH(9) ) _46304_ ( .A(ram_w8_l2048_id16_3_1_addr), .B(_tmp_320), .S(_05340_), .Y(_24590_) );
  \$mux  #( .WIDTH(9) ) _46306_ ( .A(ram_w8_l2048_id16_3_0_addr), .B(_stream_conv2d_8_source_25_source_ram_raddr[10:2]), .S(_tmp_427), .Y(_24591_) );
  \$mux  #( .WIDTH(2) ) _46308_ ( .A(_tmp_313), .B(2'h0), .S(_05630_), .Y(_24592_) );
  \$mux  #( .WIDTH(2) ) _46309_ ( .A(_24592_), .B(_22115_[1:0]), .S(_05631_), .Y(_24593_) );
  \$mux  #( .WIDTH(2) ) _46310_ ( .A(_24593_), .B(2'h0), .S(_05632_), .Y(_24594_) );
  \$mux  #( .WIDTH(9) ) _46312_ ( .A(_tmp_306), .B(_25939_[8:0]), .S(_05630_), .Y(_24595_) );
  \$mux  #( .WIDTH(9) ) _46313_ ( .A(_24595_), .B(_tmp_309), .S(_05635_), .Y(_24596_) );
  \$mux  #( .WIDTH(9) ) _46315_ ( .A(_tmp_305), .B(_25939_[8:0]), .S(_05630_), .Y(_24597_) );
  \$mux  #( .WIDTH(9) ) _46316_ ( .A(_24597_), .B(_tmp_308), .S(_05634_), .Y(_24598_) );
  \$mux  #( .WIDTH(9) ) _46318_ ( .A(_tmp_304), .B(_25939_[8:0]), .S(_05630_), .Y(_24599_) );
  \$mux  #( .WIDTH(9) ) _46319_ ( .A(_24599_), .B(_tmp_307), .S(_05633_), .Y(_24600_) );
  \$mux  #( .WIDTH(1) ) _46321_ ( .A(_tmp_303), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24601_) );
  \$mux  #( .WIDTH(1) ) _46322_ ( .A(_24601_), .B(1'h1), .S(_05636_), .Y(_24602_) );
  \$mux  #( .WIDTH(34) ) _46324_ ( .A(_tmp_302), .B({ 1'h0, _maxi_read_size }), .S(_05630_), .Y(_24603_) );
  \$mux  #( .WIDTH(34) ) _46325_ ( .A(_24603_), .B(_25998_), .S(_05337_), .Y(_24604_) );
  \$mux  #( .WIDTH(10) ) _46327_ ( .A(_tmp_301), .B(_25992_[9:0]), .S(_05630_), .Y(_24605_) );
  \$mux  #( .WIDTH(10) ) _46328_ ( .A(_24605_), .B(_25997_[9:0]), .S(_05337_), .Y(_24606_) );
  \$mux  #( .WIDTH(10) ) _46329_ ( .A(_24606_), .B(_25992_[9:0]), .S(_05631_), .Y(_24607_) );
  \$mux  #( .WIDTH(1) ) _46331_ ( .A(ram_w8_l2048_id16_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24608_) );
  \$mux  #( .WIDTH(1) ) _46332_ ( .A(_24608_), .B(_05219_), .S(_05337_), .Y(_24609_) );
  \$mux  #( .WIDTH(8) ) _46334_ ( .A(ram_w8_l2048_id16_2_1_wdata), .B(_dataflow_slice_data_62), .S(_05337_), .Y(_24610_) );
  \$mux  #( .WIDTH(9) ) _46336_ ( .A(ram_w8_l2048_id16_2_1_addr), .B(_tmp_307), .S(_05337_), .Y(_24611_) );
  \$mux  #( .WIDTH(9) ) _46338_ ( .A(ram_w8_l2048_id16_2_0_addr), .B(_stream_conv2d_8_source_25_source_ram_raddr[10:2]), .S(_tmp_427), .Y(_24612_) );
  \$mux  #( .WIDTH(2) ) _46340_ ( .A(_tmp_300), .B(2'h0), .S(_05623_), .Y(_24613_) );
  \$mux  #( .WIDTH(2) ) _46341_ ( .A(_24613_), .B(_22114_[1:0]), .S(_05624_), .Y(_24614_) );
  \$mux  #( .WIDTH(2) ) _46342_ ( .A(_24614_), .B(2'h0), .S(_05625_), .Y(_24615_) );
  \$mux  #( .WIDTH(9) ) _46344_ ( .A(_tmp_293), .B(_25939_[8:0]), .S(_05623_), .Y(_24616_) );
  \$mux  #( .WIDTH(9) ) _46345_ ( .A(_24616_), .B(_tmp_296), .S(_05628_), .Y(_24617_) );
  \$mux  #( .WIDTH(9) ) _46347_ ( .A(_tmp_292), .B(_25939_[8:0]), .S(_05623_), .Y(_24618_) );
  \$mux  #( .WIDTH(9) ) _46348_ ( .A(_24618_), .B(_tmp_295), .S(_05627_), .Y(_24619_) );
  \$mux  #( .WIDTH(9) ) _46350_ ( .A(_tmp_291), .B(_25939_[8:0]), .S(_05623_), .Y(_24620_) );
  \$mux  #( .WIDTH(9) ) _46351_ ( .A(_24620_), .B(_tmp_294), .S(_05626_), .Y(_24621_) );
  \$mux  #( .WIDTH(1) ) _46353_ ( .A(_tmp_290), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24622_) );
  \$mux  #( .WIDTH(1) ) _46354_ ( .A(_24622_), .B(1'h1), .S(_05629_), .Y(_24623_) );
  \$mux  #( .WIDTH(34) ) _46356_ ( .A(_tmp_289), .B({ 1'h0, _maxi_read_size }), .S(_05623_), .Y(_24624_) );
  \$mux  #( .WIDTH(34) ) _46357_ ( .A(_24624_), .B(_25996_), .S(_05334_), .Y(_24625_) );
  \$mux  #( .WIDTH(10) ) _46359_ ( .A(_tmp_288), .B(_25992_[9:0]), .S(_05623_), .Y(_24626_) );
  \$mux  #( .WIDTH(10) ) _46360_ ( .A(_24626_), .B(_25995_[9:0]), .S(_05334_), .Y(_24627_) );
  \$mux  #( .WIDTH(10) ) _46361_ ( .A(_24627_), .B(_25992_[9:0]), .S(_05624_), .Y(_24628_) );
  \$mux  #( .WIDTH(1) ) _46363_ ( .A(ram_w8_l2048_id16_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24629_) );
  \$mux  #( .WIDTH(1) ) _46364_ ( .A(_24629_), .B(_05216_), .S(_05334_), .Y(_24630_) );
  \$mux  #( .WIDTH(8) ) _46366_ ( .A(ram_w8_l2048_id16_1_1_wdata), .B(_dataflow_slice_data_59), .S(_05334_), .Y(_24631_) );
  \$mux  #( .WIDTH(9) ) _46368_ ( .A(ram_w8_l2048_id16_1_1_addr), .B(_tmp_294), .S(_05334_), .Y(_24632_) );
  \$mux  #( .WIDTH(9) ) _46370_ ( .A(ram_w8_l2048_id16_1_0_addr), .B(_stream_conv2d_8_source_25_source_ram_raddr[10:2]), .S(_tmp_427), .Y(_24633_) );
  \$mux  #( .WIDTH(2) ) _46373_ ( .A(_tmp_287), .B(2'h0), .S(_05616_), .Y(_24634_) );
  \$mux  #( .WIDTH(2) ) _46374_ ( .A(_24634_), .B(_22113_[1:0]), .S(_05617_), .Y(_24635_) );
  \$mux  #( .WIDTH(2) ) _46375_ ( .A(_24635_), .B(2'h0), .S(_05618_), .Y(_24636_) );
  \$mux  #( .WIDTH(9) ) _46377_ ( .A(_tmp_280), .B(_25939_[8:0]), .S(_05616_), .Y(_24637_) );
  \$mux  #( .WIDTH(9) ) _46378_ ( .A(_24637_), .B(_tmp_283), .S(_05621_), .Y(_24638_) );
  \$mux  #( .WIDTH(9) ) _46380_ ( .A(_tmp_279), .B(_25939_[8:0]), .S(_05616_), .Y(_24639_) );
  \$mux  #( .WIDTH(9) ) _46381_ ( .A(_24639_), .B(_tmp_282), .S(_05620_), .Y(_24640_) );
  \$mux  #( .WIDTH(9) ) _46383_ ( .A(_tmp_278), .B(_25939_[8:0]), .S(_05616_), .Y(_24641_) );
  \$mux  #( .WIDTH(9) ) _46384_ ( .A(_24641_), .B(_tmp_281), .S(_05619_), .Y(_24642_) );
  \$mux  #( .WIDTH(1) ) _46386_ ( .A(_tmp_277), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24643_) );
  \$mux  #( .WIDTH(1) ) _46387_ ( .A(_24643_), .B(1'h1), .S(_05622_), .Y(_24644_) );
  \$mux  #( .WIDTH(34) ) _46389_ ( .A(_tmp_276), .B({ 1'h0, _maxi_read_size }), .S(_05616_), .Y(_24645_) );
  \$mux  #( .WIDTH(34) ) _46390_ ( .A(_24645_), .B(_25994_), .S(_05331_), .Y(_24646_) );
  \$mux  #( .WIDTH(10) ) _46392_ ( .A(_tmp_275), .B(_25992_[9:0]), .S(_05616_), .Y(_24647_) );
  \$mux  #( .WIDTH(10) ) _46393_ ( .A(_24647_), .B(_25993_[9:0]), .S(_05331_), .Y(_24648_) );
  \$mux  #( .WIDTH(10) ) _46394_ ( .A(_24648_), .B(_25992_[9:0]), .S(_05617_), .Y(_24649_) );
  \$mux  #( .WIDTH(1) ) _46396_ ( .A(ram_w8_l2048_id16_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24650_) );
  \$mux  #( .WIDTH(1) ) _46397_ ( .A(_24650_), .B(_05213_), .S(_05331_), .Y(_24651_) );
  \$mux  #( .WIDTH(8) ) _46399_ ( .A(ram_w8_l2048_id16_0_1_wdata), .B(_dataflow_slice_data_56), .S(_05331_), .Y(_24652_) );
  \$mux  #( .WIDTH(9) ) _46401_ ( .A(ram_w8_l2048_id16_0_1_addr), .B(_tmp_281), .S(_05331_), .Y(_24653_) );
  \$mux  #( .WIDTH(9) ) _46403_ ( .A(ram_w8_l2048_id16_0_0_addr), .B(_stream_conv2d_8_source_25_source_ram_raddr[10:2]), .S(_tmp_427), .Y(_24654_) );
  \$mux  #( .WIDTH(1) ) _46405_ ( .A(ram_w8_l2048_id15_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24655_) );
  \$mux  #( .WIDTH(1) ) _46406_ ( .A(_24655_), .B(_05209_), .S(_05328_), .Y(_24656_) );
  \$mux  #( .WIDTH(8) ) _46408_ ( .A(ram_w8_l2048_id15_3_1_wdata), .B(_dataflow_slice_data_52), .S(_05328_), .Y(_24657_) );
  \$mux  #( .WIDTH(9) ) _46410_ ( .A(ram_w8_l2048_id15_3_1_addr), .B(_tmp_265), .S(_05328_), .Y(_24658_) );
  \$mux  #( .WIDTH(9) ) _46412_ ( .A(ram_w8_l2048_id15_3_0_addr), .B(_stream_conv2d_8_source_24_source_ram_raddr[10:2]), .S(_tmp_417), .Y(_24659_) );
  \$mux  #( .WIDTH(1) ) _46414_ ( .A(ram_w8_l2048_id15_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24660_) );
  \$mux  #( .WIDTH(1) ) _46415_ ( .A(_24660_), .B(_05206_), .S(_05325_), .Y(_24661_) );
  \$mux  #( .WIDTH(8) ) _46417_ ( .A(ram_w8_l2048_id15_2_1_wdata), .B(_dataflow_slice_data_49), .S(_05325_), .Y(_24662_) );
  \$mux  #( .WIDTH(9) ) _46419_ ( .A(ram_w8_l2048_id15_2_1_addr), .B(_tmp_252), .S(_05325_), .Y(_24663_) );
  \$mux  #( .WIDTH(9) ) _46421_ ( .A(ram_w8_l2048_id15_2_0_addr), .B(_stream_conv2d_8_source_24_source_ram_raddr[10:2]), .S(_tmp_417), .Y(_24664_) );
  \$mux  #( .WIDTH(1) ) _46423_ ( .A(ram_w8_l2048_id15_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24665_) );
  \$mux  #( .WIDTH(1) ) _46424_ ( .A(_24665_), .B(_05203_), .S(_05322_), .Y(_24666_) );
  \$mux  #( .WIDTH(8) ) _46426_ ( .A(ram_w8_l2048_id15_1_1_wdata), .B(_dataflow_slice_data_46), .S(_05322_), .Y(_24667_) );
  \$mux  #( .WIDTH(9) ) _46428_ ( .A(ram_w8_l2048_id15_1_1_addr), .B(_tmp_239), .S(_05322_), .Y(_24668_) );
  \$mux  #( .WIDTH(9) ) _46430_ ( .A(ram_w8_l2048_id15_1_0_addr), .B(_stream_conv2d_8_source_24_source_ram_raddr[10:2]), .S(_tmp_417), .Y(_24669_) );
  \$mux  #( .WIDTH(1) ) _46433_ ( .A(ram_w8_l2048_id15_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24670_) );
  \$mux  #( .WIDTH(1) ) _46434_ ( .A(_24670_), .B(_05200_), .S(_05319_), .Y(_24671_) );
  \$mux  #( .WIDTH(8) ) _46436_ ( .A(ram_w8_l2048_id15_0_1_wdata), .B(_dataflow_slice_data_43), .S(_05319_), .Y(_24672_) );
  \$mux  #( .WIDTH(9) ) _46438_ ( .A(ram_w8_l2048_id15_0_1_addr), .B(_tmp_226), .S(_05319_), .Y(_24673_) );
  \$mux  #( .WIDTH(9) ) _46440_ ( .A(ram_w8_l2048_id15_0_0_addr), .B(_stream_conv2d_8_source_24_source_ram_raddr[10:2]), .S(_tmp_417), .Y(_24674_) );
  \$mux  #( .WIDTH(1) ) _46442_ ( .A(ram_w8_l2048_id14_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24675_) );
  \$mux  #( .WIDTH(1) ) _46443_ ( .A(_24675_), .B(_05211_), .S(_05328_), .Y(_24676_) );
  \$mux  #( .WIDTH(8) ) _46445_ ( .A(ram_w8_l2048_id14_3_1_wdata), .B(_dataflow_slice_data_52), .S(_05328_), .Y(_24677_) );
  \$mux  #( .WIDTH(9) ) _46447_ ( .A(ram_w8_l2048_id14_3_1_addr), .B(_tmp_264), .S(_05328_), .Y(_24678_) );
  \$mux  #( .WIDTH(9) ) _46449_ ( .A(ram_w8_l2048_id14_3_0_addr), .B(_stream_conv2d_8_source_23_source_ram_raddr[10:2]), .S(_tmp_407), .Y(_24679_) );
  \$mux  #( .WIDTH(1) ) _46451_ ( .A(ram_w8_l2048_id14_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24680_) );
  \$mux  #( .WIDTH(1) ) _46452_ ( .A(_24680_), .B(_05208_), .S(_05325_), .Y(_24681_) );
  \$mux  #( .WIDTH(8) ) _46454_ ( .A(ram_w8_l2048_id14_2_1_wdata), .B(_dataflow_slice_data_49), .S(_05325_), .Y(_24682_) );
  \$mux  #( .WIDTH(9) ) _46456_ ( .A(ram_w8_l2048_id14_2_1_addr), .B(_tmp_251), .S(_05325_), .Y(_24683_) );
  \$mux  #( .WIDTH(9) ) _46458_ ( .A(ram_w8_l2048_id14_2_0_addr), .B(_stream_conv2d_8_source_23_source_ram_raddr[10:2]), .S(_tmp_407), .Y(_24684_) );
  \$mux  #( .WIDTH(1) ) _46460_ ( .A(ram_w8_l2048_id14_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24685_) );
  \$mux  #( .WIDTH(1) ) _46461_ ( .A(_24685_), .B(_05205_), .S(_05322_), .Y(_24686_) );
  \$mux  #( .WIDTH(8) ) _46463_ ( .A(ram_w8_l2048_id14_1_1_wdata), .B(_dataflow_slice_data_46), .S(_05322_), .Y(_24687_) );
  \$mux  #( .WIDTH(9) ) _46465_ ( .A(ram_w8_l2048_id14_1_1_addr), .B(_tmp_238), .S(_05322_), .Y(_24688_) );
  \$mux  #( .WIDTH(9) ) _46467_ ( .A(ram_w8_l2048_id14_1_0_addr), .B(_stream_conv2d_8_source_23_source_ram_raddr[10:2]), .S(_tmp_407), .Y(_24689_) );
  \$mux  #( .WIDTH(1) ) _46470_ ( .A(ram_w8_l2048_id14_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24690_) );
  \$mux  #( .WIDTH(1) ) _46471_ ( .A(_24690_), .B(_05202_), .S(_05319_), .Y(_24691_) );
  \$mux  #( .WIDTH(8) ) _46473_ ( .A(ram_w8_l2048_id14_0_1_wdata), .B(_dataflow_slice_data_43), .S(_05319_), .Y(_24692_) );
  \$mux  #( .WIDTH(9) ) _46475_ ( .A(ram_w8_l2048_id14_0_1_addr), .B(_tmp_225), .S(_05319_), .Y(_24693_) );
  \$mux  #( .WIDTH(9) ) _46477_ ( .A(ram_w8_l2048_id14_0_0_addr), .B(_stream_conv2d_8_source_23_source_ram_raddr[10:2]), .S(_tmp_407), .Y(_24694_) );
  \$mux  #( .WIDTH(2) ) _46479_ ( .A(_tmp_269), .B(2'h0), .S(_05608_), .Y(_24695_) );
  \$mux  #( .WIDTH(2) ) _46480_ ( .A(_24695_), .B(_22112_[1:0]), .S(_05609_), .Y(_24696_) );
  \$mux  #( .WIDTH(2) ) _46481_ ( .A(_24696_), .B(2'h0), .S(_05610_), .Y(_24697_) );
  \$mux  #( .WIDTH(9) ) _46483_ ( .A(_tmp_262), .B(_25939_[8:0]), .S(_05608_), .Y(_24698_) );
  \$mux  #( .WIDTH(9) ) _46484_ ( .A(_24698_), .B(_tmp_265), .S(_05613_), .Y(_24699_) );
  \$mux  #( .WIDTH(9) ) _46486_ ( .A(_tmp_261), .B(_25939_[8:0]), .S(_05608_), .Y(_24700_) );
  \$mux  #( .WIDTH(9) ) _46487_ ( .A(_24700_), .B(_tmp_264), .S(_05612_), .Y(_24701_) );
  \$mux  #( .WIDTH(9) ) _46489_ ( .A(_tmp_260), .B(_25939_[8:0]), .S(_05608_), .Y(_24702_) );
  \$mux  #( .WIDTH(9) ) _46490_ ( .A(_24702_), .B(_tmp_263), .S(_05611_), .Y(_24703_) );
  \$mux  #( .WIDTH(1) ) _46492_ ( .A(_tmp_259), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24704_) );
  \$mux  #( .WIDTH(1) ) _46493_ ( .A(_24704_), .B(1'h1), .S(_05614_), .Y(_24705_) );
  \$mux  #( .WIDTH(34) ) _46495_ ( .A(_tmp_258), .B({ 1'h0, _maxi_read_size }), .S(_05608_), .Y(_24706_) );
  \$mux  #( .WIDTH(34) ) _46496_ ( .A(_24706_), .B(_25991_), .S(_05328_), .Y(_24707_) );
  \$mux  #( .WIDTH(10) ) _46498_ ( .A(_tmp_257), .B(_25983_[9:0]), .S(_05608_), .Y(_24708_) );
  \$mux  #( .WIDTH(10) ) _46499_ ( .A(_24708_), .B(_25990_[9:0]), .S(_05328_), .Y(_24709_) );
  \$mux  #( .WIDTH(10) ) _46500_ ( .A(_24709_), .B(_25983_[9:0]), .S(_05609_), .Y(_24710_) );
  \$mux  #( .WIDTH(1) ) _46502_ ( .A(ram_w8_l2048_id13_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24711_) );
  \$mux  #( .WIDTH(1) ) _46503_ ( .A(_24711_), .B(_05210_), .S(_05328_), .Y(_24712_) );
  \$mux  #( .WIDTH(8) ) _46505_ ( .A(ram_w8_l2048_id13_3_1_wdata), .B(_dataflow_slice_data_52), .S(_05328_), .Y(_24713_) );
  \$mux  #( .WIDTH(9) ) _46507_ ( .A(ram_w8_l2048_id13_3_1_addr), .B(_tmp_263), .S(_05328_), .Y(_24714_) );
  \$mux  #( .WIDTH(9) ) _46509_ ( .A(ram_w8_l2048_id13_3_0_addr), .B(_stream_conv2d_8_source_22_source_ram_raddr[10:2]), .S(_tmp_397), .Y(_24715_) );
  \$mux  #( .WIDTH(2) ) _46511_ ( .A(_tmp_256), .B(2'h0), .S(_05601_), .Y(_24716_) );
  \$mux  #( .WIDTH(2) ) _46512_ ( .A(_24716_), .B(_22111_[1:0]), .S(_05602_), .Y(_24717_) );
  \$mux  #( .WIDTH(2) ) _46513_ ( .A(_24717_), .B(2'h0), .S(_05603_), .Y(_24718_) );
  \$mux  #( .WIDTH(9) ) _46515_ ( .A(_tmp_249), .B(_25939_[8:0]), .S(_05601_), .Y(_24719_) );
  \$mux  #( .WIDTH(9) ) _46516_ ( .A(_24719_), .B(_tmp_252), .S(_05606_), .Y(_24720_) );
  \$mux  #( .WIDTH(9) ) _46518_ ( .A(_tmp_248), .B(_25939_[8:0]), .S(_05601_), .Y(_24721_) );
  \$mux  #( .WIDTH(9) ) _46519_ ( .A(_24721_), .B(_tmp_251), .S(_05605_), .Y(_24722_) );
  \$mux  #( .WIDTH(9) ) _46521_ ( .A(_tmp_247), .B(_25939_[8:0]), .S(_05601_), .Y(_24723_) );
  \$mux  #( .WIDTH(9) ) _46522_ ( .A(_24723_), .B(_tmp_250), .S(_05604_), .Y(_24724_) );
  \$mux  #( .WIDTH(1) ) _46524_ ( .A(_tmp_246), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24725_) );
  \$mux  #( .WIDTH(1) ) _46525_ ( .A(_24725_), .B(1'h1), .S(_05607_), .Y(_24726_) );
  \$mux  #( .WIDTH(34) ) _46527_ ( .A(_tmp_245), .B({ 1'h0, _maxi_read_size }), .S(_05601_), .Y(_24727_) );
  \$mux  #( .WIDTH(34) ) _46528_ ( .A(_24727_), .B(_25989_), .S(_05325_), .Y(_24728_) );
  \$mux  #( .WIDTH(10) ) _46530_ ( .A(_tmp_244), .B(_25983_[9:0]), .S(_05601_), .Y(_24729_) );
  \$mux  #( .WIDTH(10) ) _46531_ ( .A(_24729_), .B(_25988_[9:0]), .S(_05325_), .Y(_24730_) );
  \$mux  #( .WIDTH(10) ) _46532_ ( .A(_24730_), .B(_25983_[9:0]), .S(_05602_), .Y(_24731_) );
  \$mux  #( .WIDTH(1) ) _46534_ ( .A(ram_w8_l2048_id13_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24732_) );
  \$mux  #( .WIDTH(1) ) _46535_ ( .A(_24732_), .B(_05207_), .S(_05325_), .Y(_24733_) );
  \$mux  #( .WIDTH(8) ) _46537_ ( .A(ram_w8_l2048_id13_2_1_wdata), .B(_dataflow_slice_data_49), .S(_05325_), .Y(_24734_) );
  \$mux  #( .WIDTH(9) ) _46539_ ( .A(ram_w8_l2048_id13_2_1_addr), .B(_tmp_250), .S(_05325_), .Y(_24735_) );
  \$mux  #( .WIDTH(9) ) _46541_ ( .A(ram_w8_l2048_id13_2_0_addr), .B(_stream_conv2d_8_source_22_source_ram_raddr[10:2]), .S(_tmp_397), .Y(_24736_) );
  \$mux  #( .WIDTH(2) ) _46543_ ( .A(_tmp_243), .B(2'h0), .S(_05594_), .Y(_24737_) );
  \$mux  #( .WIDTH(2) ) _46544_ ( .A(_24737_), .B(_22110_[1:0]), .S(_05595_), .Y(_24738_) );
  \$mux  #( .WIDTH(2) ) _46545_ ( .A(_24738_), .B(2'h0), .S(_05596_), .Y(_24739_) );
  \$mux  #( .WIDTH(9) ) _46547_ ( .A(_tmp_236), .B(_25939_[8:0]), .S(_05594_), .Y(_24740_) );
  \$mux  #( .WIDTH(9) ) _46548_ ( .A(_24740_), .B(_tmp_239), .S(_05599_), .Y(_24741_) );
  \$mux  #( .WIDTH(9) ) _46550_ ( .A(_tmp_235), .B(_25939_[8:0]), .S(_05594_), .Y(_24742_) );
  \$mux  #( .WIDTH(9) ) _46551_ ( .A(_24742_), .B(_tmp_238), .S(_05598_), .Y(_24743_) );
  \$mux  #( .WIDTH(9) ) _46553_ ( .A(_tmp_234), .B(_25939_[8:0]), .S(_05594_), .Y(_24744_) );
  \$mux  #( .WIDTH(9) ) _46554_ ( .A(_24744_), .B(_tmp_237), .S(_05597_), .Y(_24745_) );
  \$mux  #( .WIDTH(1) ) _46556_ ( .A(_tmp_233), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24746_) );
  \$mux  #( .WIDTH(1) ) _46557_ ( .A(_24746_), .B(1'h1), .S(_05600_), .Y(_24747_) );
  \$mux  #( .WIDTH(34) ) _46559_ ( .A(_tmp_232), .B({ 1'h0, _maxi_read_size }), .S(_05594_), .Y(_24748_) );
  \$mux  #( .WIDTH(34) ) _46560_ ( .A(_24748_), .B(_25987_), .S(_05322_), .Y(_24749_) );
  \$mux  #( .WIDTH(10) ) _46562_ ( .A(_tmp_231), .B(_25983_[9:0]), .S(_05594_), .Y(_24750_) );
  \$mux  #( .WIDTH(10) ) _46563_ ( .A(_24750_), .B(_25986_[9:0]), .S(_05322_), .Y(_24751_) );
  \$mux  #( .WIDTH(10) ) _46564_ ( .A(_24751_), .B(_25983_[9:0]), .S(_05595_), .Y(_24752_) );
  \$mux  #( .WIDTH(1) ) _46566_ ( .A(ram_w8_l2048_id13_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24753_) );
  \$mux  #( .WIDTH(1) ) _46567_ ( .A(_24753_), .B(_05204_), .S(_05322_), .Y(_24754_) );
  \$mux  #( .WIDTH(8) ) _46569_ ( .A(ram_w8_l2048_id13_1_1_wdata), .B(_dataflow_slice_data_46), .S(_05322_), .Y(_24755_) );
  \$mux  #( .WIDTH(9) ) _46571_ ( .A(ram_w8_l2048_id13_1_1_addr), .B(_tmp_237), .S(_05322_), .Y(_24756_) );
  \$mux  #( .WIDTH(9) ) _46573_ ( .A(ram_w8_l2048_id13_1_0_addr), .B(_stream_conv2d_8_source_22_source_ram_raddr[10:2]), .S(_tmp_397), .Y(_24757_) );
  \$mux  #( .WIDTH(2) ) _46576_ ( .A(_tmp_230), .B(2'h0), .S(_05587_), .Y(_24758_) );
  \$mux  #( .WIDTH(2) ) _46577_ ( .A(_24758_), .B(_22109_[1:0]), .S(_05588_), .Y(_24759_) );
  \$mux  #( .WIDTH(2) ) _46578_ ( .A(_24759_), .B(2'h0), .S(_05589_), .Y(_24760_) );
  \$mux  #( .WIDTH(9) ) _46580_ ( .A(_tmp_223), .B(_25939_[8:0]), .S(_05587_), .Y(_24761_) );
  \$mux  #( .WIDTH(9) ) _46581_ ( .A(_24761_), .B(_tmp_226), .S(_05592_), .Y(_24762_) );
  \$mux  #( .WIDTH(9) ) _46583_ ( .A(_tmp_222), .B(_25939_[8:0]), .S(_05587_), .Y(_24763_) );
  \$mux  #( .WIDTH(9) ) _46584_ ( .A(_24763_), .B(_tmp_225), .S(_05591_), .Y(_24764_) );
  \$mux  #( .WIDTH(9) ) _46586_ ( .A(_tmp_221), .B(_25939_[8:0]), .S(_05587_), .Y(_24765_) );
  \$mux  #( .WIDTH(9) ) _46587_ ( .A(_24765_), .B(_tmp_224), .S(_05590_), .Y(_24766_) );
  \$mux  #( .WIDTH(1) ) _46589_ ( .A(_tmp_220), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24767_) );
  \$mux  #( .WIDTH(1) ) _46590_ ( .A(_24767_), .B(1'h1), .S(_05593_), .Y(_24768_) );
  \$mux  #( .WIDTH(34) ) _46592_ ( .A(_tmp_219), .B({ 1'h0, _maxi_read_size }), .S(_05587_), .Y(_24769_) );
  \$mux  #( .WIDTH(34) ) _46593_ ( .A(_24769_), .B(_25985_), .S(_05319_), .Y(_24770_) );
  \$mux  #( .WIDTH(10) ) _46595_ ( .A(_tmp_218), .B(_25983_[9:0]), .S(_05587_), .Y(_24771_) );
  \$mux  #( .WIDTH(10) ) _46596_ ( .A(_24771_), .B(_25984_[9:0]), .S(_05319_), .Y(_24772_) );
  \$mux  #( .WIDTH(10) ) _46597_ ( .A(_24772_), .B(_25983_[9:0]), .S(_05588_), .Y(_24773_) );
  \$mux  #( .WIDTH(1) ) _46599_ ( .A(ram_w8_l2048_id13_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24774_) );
  \$mux  #( .WIDTH(1) ) _46600_ ( .A(_24774_), .B(_05201_), .S(_05319_), .Y(_24775_) );
  \$mux  #( .WIDTH(8) ) _46602_ ( .A(ram_w8_l2048_id13_0_1_wdata), .B(_dataflow_slice_data_43), .S(_05319_), .Y(_24776_) );
  \$mux  #( .WIDTH(9) ) _46604_ ( .A(ram_w8_l2048_id13_0_1_addr), .B(_tmp_224), .S(_05319_), .Y(_24777_) );
  \$mux  #( .WIDTH(9) ) _46606_ ( .A(ram_w8_l2048_id13_0_0_addr), .B(_stream_conv2d_8_source_22_source_ram_raddr[10:2]), .S(_tmp_397), .Y(_24778_) );
  \$mux  #( .WIDTH(1) ) _46608_ ( .A(ram_w8_l2048_id12_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24779_) );
  \$mux  #( .WIDTH(1) ) _46609_ ( .A(_24779_), .B(_05197_), .S(_05316_), .Y(_24780_) );
  \$mux  #( .WIDTH(8) ) _46611_ ( .A(ram_w8_l2048_id12_3_1_wdata), .B(_dataflow_slice_data_39), .S(_05316_), .Y(_24781_) );
  \$mux  #( .WIDTH(9) ) _46613_ ( .A(ram_w8_l2048_id12_3_1_addr), .B(_tmp_208), .S(_05316_), .Y(_24782_) );
  \$mux  #( .WIDTH(9) ) _46615_ ( .A(ram_w8_l2048_id12_3_0_addr), .B(_stream_conv2d_8_source_21_source_ram_raddr[10:2]), .S(_tmp_387), .Y(_24783_) );
  \$mux  #( .WIDTH(1) ) _46617_ ( .A(ram_w8_l2048_id12_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24784_) );
  \$mux  #( .WIDTH(1) ) _46618_ ( .A(_24784_), .B(_05194_), .S(_05313_), .Y(_24785_) );
  \$mux  #( .WIDTH(8) ) _46620_ ( .A(ram_w8_l2048_id12_2_1_wdata), .B(_dataflow_slice_data_36), .S(_05313_), .Y(_24786_) );
  \$mux  #( .WIDTH(9) ) _46622_ ( .A(ram_w8_l2048_id12_2_1_addr), .B(_tmp_195), .S(_05313_), .Y(_24787_) );
  \$mux  #( .WIDTH(9) ) _46624_ ( .A(ram_w8_l2048_id12_2_0_addr), .B(_stream_conv2d_8_source_21_source_ram_raddr[10:2]), .S(_tmp_387), .Y(_24788_) );
  \$mux  #( .WIDTH(1) ) _46626_ ( .A(ram_w8_l2048_id12_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24789_) );
  \$mux  #( .WIDTH(1) ) _46627_ ( .A(_24789_), .B(_05191_), .S(_05310_), .Y(_24790_) );
  \$mux  #( .WIDTH(8) ) _46629_ ( .A(ram_w8_l2048_id12_1_1_wdata), .B(_dataflow_slice_data_33), .S(_05310_), .Y(_24791_) );
  \$mux  #( .WIDTH(9) ) _46631_ ( .A(ram_w8_l2048_id12_1_1_addr), .B(_tmp_182), .S(_05310_), .Y(_24792_) );
  \$mux  #( .WIDTH(9) ) _46633_ ( .A(ram_w8_l2048_id12_1_0_addr), .B(_stream_conv2d_8_source_21_source_ram_raddr[10:2]), .S(_tmp_387), .Y(_24793_) );
  \$mux  #( .WIDTH(1) ) _46636_ ( .A(ram_w8_l2048_id12_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24794_) );
  \$mux  #( .WIDTH(1) ) _46637_ ( .A(_24794_), .B(_05188_), .S(_05307_), .Y(_24795_) );
  \$mux  #( .WIDTH(8) ) _46639_ ( .A(ram_w8_l2048_id12_0_1_wdata), .B(_dataflow_slice_data_30), .S(_05307_), .Y(_24796_) );
  \$mux  #( .WIDTH(9) ) _46641_ ( .A(ram_w8_l2048_id12_0_1_addr), .B(_tmp_169), .S(_05307_), .Y(_24797_) );
  \$mux  #( .WIDTH(9) ) _46643_ ( .A(ram_w8_l2048_id12_0_0_addr), .B(_stream_conv2d_8_source_21_source_ram_raddr[10:2]), .S(_tmp_387), .Y(_24798_) );
  \$mux  #( .WIDTH(1) ) _46645_ ( .A(ram_w8_l2048_id11_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24799_) );
  \$mux  #( .WIDTH(1) ) _46646_ ( .A(_24799_), .B(_05199_), .S(_05316_), .Y(_24800_) );
  \$mux  #( .WIDTH(8) ) _46648_ ( .A(ram_w8_l2048_id11_3_1_wdata), .B(_dataflow_slice_data_39), .S(_05316_), .Y(_24801_) );
  \$mux  #( .WIDTH(9) ) _46650_ ( .A(ram_w8_l2048_id11_3_1_addr), .B(_tmp_207), .S(_05316_), .Y(_24802_) );
  \$mux  #( .WIDTH(9) ) _46652_ ( .A(ram_w8_l2048_id11_3_0_addr), .B(_stream_conv2d_8_source_20_source_ram_raddr[10:2]), .S(_tmp_377), .Y(_24803_) );
  \$mux  #( .WIDTH(1) ) _46654_ ( .A(ram_w8_l2048_id11_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24804_) );
  \$mux  #( .WIDTH(1) ) _46655_ ( .A(_24804_), .B(_05196_), .S(_05313_), .Y(_24805_) );
  \$mux  #( .WIDTH(8) ) _46657_ ( .A(ram_w8_l2048_id11_2_1_wdata), .B(_dataflow_slice_data_36), .S(_05313_), .Y(_24806_) );
  \$mux  #( .WIDTH(9) ) _46659_ ( .A(ram_w8_l2048_id11_2_1_addr), .B(_tmp_194), .S(_05313_), .Y(_24807_) );
  \$mux  #( .WIDTH(9) ) _46661_ ( .A(ram_w8_l2048_id11_2_0_addr), .B(_stream_conv2d_8_source_20_source_ram_raddr[10:2]), .S(_tmp_377), .Y(_24808_) );
  \$mux  #( .WIDTH(1) ) _46663_ ( .A(ram_w8_l2048_id11_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24809_) );
  \$mux  #( .WIDTH(1) ) _46664_ ( .A(_24809_), .B(_05193_), .S(_05310_), .Y(_24810_) );
  \$mux  #( .WIDTH(8) ) _46666_ ( .A(ram_w8_l2048_id11_1_1_wdata), .B(_dataflow_slice_data_33), .S(_05310_), .Y(_24811_) );
  \$mux  #( .WIDTH(9) ) _46668_ ( .A(ram_w8_l2048_id11_1_1_addr), .B(_tmp_181), .S(_05310_), .Y(_24812_) );
  \$mux  #( .WIDTH(9) ) _46670_ ( .A(ram_w8_l2048_id11_1_0_addr), .B(_stream_conv2d_8_source_20_source_ram_raddr[10:2]), .S(_tmp_377), .Y(_24813_) );
  \$mux  #( .WIDTH(1) ) _46673_ ( .A(ram_w8_l2048_id11_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24814_) );
  \$mux  #( .WIDTH(1) ) _46674_ ( .A(_24814_), .B(_05190_), .S(_05307_), .Y(_24815_) );
  \$mux  #( .WIDTH(8) ) _46676_ ( .A(ram_w8_l2048_id11_0_1_wdata), .B(_dataflow_slice_data_30), .S(_05307_), .Y(_24816_) );
  \$mux  #( .WIDTH(9) ) _46678_ ( .A(ram_w8_l2048_id11_0_1_addr), .B(_tmp_168), .S(_05307_), .Y(_24817_) );
  \$mux  #( .WIDTH(9) ) _46680_ ( .A(ram_w8_l2048_id11_0_0_addr), .B(_stream_conv2d_8_source_20_source_ram_raddr[10:2]), .S(_tmp_377), .Y(_24818_) );
  \$mux  #( .WIDTH(2) ) _46682_ ( .A(_tmp_212), .B(2'h0), .S(_05579_), .Y(_24819_) );
  \$mux  #( .WIDTH(2) ) _46683_ ( .A(_24819_), .B(_22108_[1:0]), .S(_05580_), .Y(_24820_) );
  \$mux  #( .WIDTH(2) ) _46684_ ( .A(_24820_), .B(2'h0), .S(_05581_), .Y(_24821_) );
  \$mux  #( .WIDTH(9) ) _46686_ ( .A(_tmp_205), .B(_25939_[8:0]), .S(_05579_), .Y(_24822_) );
  \$mux  #( .WIDTH(9) ) _46687_ ( .A(_24822_), .B(_tmp_208), .S(_05584_), .Y(_24823_) );
  \$mux  #( .WIDTH(9) ) _46689_ ( .A(_tmp_204), .B(_25939_[8:0]), .S(_05579_), .Y(_24824_) );
  \$mux  #( .WIDTH(9) ) _46690_ ( .A(_24824_), .B(_tmp_207), .S(_05583_), .Y(_24825_) );
  \$mux  #( .WIDTH(9) ) _46692_ ( .A(_tmp_203), .B(_25939_[8:0]), .S(_05579_), .Y(_24826_) );
  \$mux  #( .WIDTH(9) ) _46693_ ( .A(_24826_), .B(_tmp_206), .S(_05582_), .Y(_24827_) );
  \$mux  #( .WIDTH(1) ) _46695_ ( .A(_tmp_202), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24828_) );
  \$mux  #( .WIDTH(1) ) _46696_ ( .A(_24828_), .B(1'h1), .S(_05585_), .Y(_24829_) );
  \$mux  #( .WIDTH(34) ) _46698_ ( .A(_tmp_201), .B({ 1'h0, _maxi_read_size }), .S(_05579_), .Y(_24830_) );
  \$mux  #( .WIDTH(34) ) _46699_ ( .A(_24830_), .B(_25982_), .S(_05316_), .Y(_24831_) );
  \$mux  #( .WIDTH(10) ) _46701_ ( .A(_tmp_200), .B(_25974_[9:0]), .S(_05579_), .Y(_24832_) );
  \$mux  #( .WIDTH(10) ) _46702_ ( .A(_24832_), .B(_25981_[9:0]), .S(_05316_), .Y(_24833_) );
  \$mux  #( .WIDTH(10) ) _46703_ ( .A(_24833_), .B(_25974_[9:0]), .S(_05580_), .Y(_24834_) );
  \$mux  #( .WIDTH(1) ) _46705_ ( .A(ram_w8_l2048_id10_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24835_) );
  \$mux  #( .WIDTH(1) ) _46706_ ( .A(_24835_), .B(_05198_), .S(_05316_), .Y(_24836_) );
  \$mux  #( .WIDTH(8) ) _46708_ ( .A(ram_w8_l2048_id10_3_1_wdata), .B(_dataflow_slice_data_39), .S(_05316_), .Y(_24837_) );
  \$mux  #( .WIDTH(9) ) _46710_ ( .A(ram_w8_l2048_id10_3_1_addr), .B(_tmp_206), .S(_05316_), .Y(_24838_) );
  \$mux  #( .WIDTH(9) ) _46712_ ( .A(ram_w8_l2048_id10_3_0_addr), .B(_stream_conv2d_8_source_19_source_ram_raddr[10:2]), .S(_tmp_367), .Y(_24839_) );
  \$mux  #( .WIDTH(2) ) _46714_ ( .A(_tmp_199), .B(2'h0), .S(_05572_), .Y(_24840_) );
  \$mux  #( .WIDTH(2) ) _46715_ ( .A(_24840_), .B(_22107_[1:0]), .S(_05573_), .Y(_24841_) );
  \$mux  #( .WIDTH(2) ) _46716_ ( .A(_24841_), .B(2'h0), .S(_05574_), .Y(_24842_) );
  \$mux  #( .WIDTH(9) ) _46718_ ( .A(_tmp_192), .B(_25939_[8:0]), .S(_05572_), .Y(_24843_) );
  \$mux  #( .WIDTH(9) ) _46719_ ( .A(_24843_), .B(_tmp_195), .S(_05577_), .Y(_24844_) );
  \$mux  #( .WIDTH(9) ) _46721_ ( .A(_tmp_191), .B(_25939_[8:0]), .S(_05572_), .Y(_24845_) );
  \$mux  #( .WIDTH(9) ) _46722_ ( .A(_24845_), .B(_tmp_194), .S(_05576_), .Y(_24846_) );
  \$mux  #( .WIDTH(9) ) _46724_ ( .A(_tmp_190), .B(_25939_[8:0]), .S(_05572_), .Y(_24847_) );
  \$mux  #( .WIDTH(9) ) _46725_ ( .A(_24847_), .B(_tmp_193), .S(_05575_), .Y(_24848_) );
  \$mux  #( .WIDTH(1) ) _46727_ ( .A(_tmp_189), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24849_) );
  \$mux  #( .WIDTH(1) ) _46728_ ( .A(_24849_), .B(1'h1), .S(_05578_), .Y(_24850_) );
  \$mux  #( .WIDTH(34) ) _46730_ ( .A(_tmp_188), .B({ 1'h0, _maxi_read_size }), .S(_05572_), .Y(_24851_) );
  \$mux  #( .WIDTH(34) ) _46731_ ( .A(_24851_), .B(_25980_), .S(_05313_), .Y(_24852_) );
  \$mux  #( .WIDTH(10) ) _46733_ ( .A(_tmp_187), .B(_25974_[9:0]), .S(_05572_), .Y(_24853_) );
  \$mux  #( .WIDTH(10) ) _46734_ ( .A(_24853_), .B(_25979_[9:0]), .S(_05313_), .Y(_24854_) );
  \$mux  #( .WIDTH(10) ) _46735_ ( .A(_24854_), .B(_25974_[9:0]), .S(_05573_), .Y(_24855_) );
  \$mux  #( .WIDTH(1) ) _46737_ ( .A(ram_w8_l2048_id10_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24856_) );
  \$mux  #( .WIDTH(1) ) _46738_ ( .A(_24856_), .B(_05195_), .S(_05313_), .Y(_24857_) );
  \$mux  #( .WIDTH(8) ) _46740_ ( .A(ram_w8_l2048_id10_2_1_wdata), .B(_dataflow_slice_data_36), .S(_05313_), .Y(_24858_) );
  \$mux  #( .WIDTH(9) ) _46742_ ( .A(ram_w8_l2048_id10_2_1_addr), .B(_tmp_193), .S(_05313_), .Y(_24859_) );
  \$mux  #( .WIDTH(9) ) _46744_ ( .A(ram_w8_l2048_id10_2_0_addr), .B(_stream_conv2d_8_source_19_source_ram_raddr[10:2]), .S(_tmp_367), .Y(_24860_) );
  \$mux  #( .WIDTH(2) ) _46746_ ( .A(_tmp_186), .B(2'h0), .S(_05565_), .Y(_24861_) );
  \$mux  #( .WIDTH(2) ) _46747_ ( .A(_24861_), .B(_22106_[1:0]), .S(_05566_), .Y(_24862_) );
  \$mux  #( .WIDTH(2) ) _46748_ ( .A(_24862_), .B(2'h0), .S(_05567_), .Y(_24863_) );
  \$mux  #( .WIDTH(9) ) _46750_ ( .A(_tmp_179), .B(_25939_[8:0]), .S(_05565_), .Y(_24864_) );
  \$mux  #( .WIDTH(9) ) _46751_ ( .A(_24864_), .B(_tmp_182), .S(_05570_), .Y(_24865_) );
  \$mux  #( .WIDTH(9) ) _46753_ ( .A(_tmp_178), .B(_25939_[8:0]), .S(_05565_), .Y(_24866_) );
  \$mux  #( .WIDTH(9) ) _46754_ ( .A(_24866_), .B(_tmp_181), .S(_05569_), .Y(_24867_) );
  \$mux  #( .WIDTH(9) ) _46756_ ( .A(_tmp_177), .B(_25939_[8:0]), .S(_05565_), .Y(_24868_) );
  \$mux  #( .WIDTH(9) ) _46757_ ( .A(_24868_), .B(_tmp_180), .S(_05568_), .Y(_24869_) );
  \$mux  #( .WIDTH(1) ) _46759_ ( .A(_tmp_176), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24870_) );
  \$mux  #( .WIDTH(1) ) _46760_ ( .A(_24870_), .B(1'h1), .S(_05571_), .Y(_24871_) );
  \$mux  #( .WIDTH(34) ) _46762_ ( .A(_tmp_175), .B({ 1'h0, _maxi_read_size }), .S(_05565_), .Y(_24872_) );
  \$mux  #( .WIDTH(34) ) _46763_ ( .A(_24872_), .B(_25978_), .S(_05310_), .Y(_24873_) );
  \$mux  #( .WIDTH(10) ) _46765_ ( .A(_tmp_174), .B(_25974_[9:0]), .S(_05565_), .Y(_24874_) );
  \$mux  #( .WIDTH(10) ) _46766_ ( .A(_24874_), .B(_25977_[9:0]), .S(_05310_), .Y(_24875_) );
  \$mux  #( .WIDTH(10) ) _46767_ ( .A(_24875_), .B(_25974_[9:0]), .S(_05566_), .Y(_24876_) );
  \$mux  #( .WIDTH(1) ) _46769_ ( .A(ram_w8_l2048_id10_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24877_) );
  \$mux  #( .WIDTH(1) ) _46770_ ( .A(_24877_), .B(_05192_), .S(_05310_), .Y(_24878_) );
  \$mux  #( .WIDTH(8) ) _46772_ ( .A(ram_w8_l2048_id10_1_1_wdata), .B(_dataflow_slice_data_33), .S(_05310_), .Y(_24879_) );
  \$mux  #( .WIDTH(9) ) _46774_ ( .A(ram_w8_l2048_id10_1_1_addr), .B(_tmp_180), .S(_05310_), .Y(_24880_) );
  \$mux  #( .WIDTH(9) ) _46776_ ( .A(ram_w8_l2048_id10_1_0_addr), .B(_stream_conv2d_8_source_19_source_ram_raddr[10:2]), .S(_tmp_367), .Y(_24881_) );
  \$mux  #( .WIDTH(2) ) _46779_ ( .A(_tmp_173), .B(2'h0), .S(_05558_), .Y(_24882_) );
  \$mux  #( .WIDTH(2) ) _46780_ ( .A(_24882_), .B(_22105_[1:0]), .S(_05559_), .Y(_24883_) );
  \$mux  #( .WIDTH(2) ) _46781_ ( .A(_24883_), .B(2'h0), .S(_05560_), .Y(_24884_) );
  \$mux  #( .WIDTH(9) ) _46783_ ( .A(_tmp_166), .B(_25939_[8:0]), .S(_05558_), .Y(_24885_) );
  \$mux  #( .WIDTH(9) ) _46784_ ( .A(_24885_), .B(_tmp_169), .S(_05563_), .Y(_24886_) );
  \$mux  #( .WIDTH(9) ) _46786_ ( .A(_tmp_165), .B(_25939_[8:0]), .S(_05558_), .Y(_24887_) );
  \$mux  #( .WIDTH(9) ) _46787_ ( .A(_24887_), .B(_tmp_168), .S(_05562_), .Y(_24888_) );
  \$mux  #( .WIDTH(9) ) _46789_ ( .A(_tmp_164), .B(_25939_[8:0]), .S(_05558_), .Y(_24889_) );
  \$mux  #( .WIDTH(9) ) _46790_ ( .A(_24889_), .B(_tmp_167), .S(_05561_), .Y(_24890_) );
  \$mux  #( .WIDTH(1) ) _46792_ ( .A(_tmp_163), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24891_) );
  \$mux  #( .WIDTH(1) ) _46793_ ( .A(_24891_), .B(1'h1), .S(_05564_), .Y(_24892_) );
  \$mux  #( .WIDTH(34) ) _46795_ ( .A(_tmp_162), .B({ 1'h0, _maxi_read_size }), .S(_05558_), .Y(_24893_) );
  \$mux  #( .WIDTH(34) ) _46796_ ( .A(_24893_), .B(_25976_), .S(_05307_), .Y(_24894_) );
  \$mux  #( .WIDTH(10) ) _46798_ ( .A(_tmp_161), .B(_25974_[9:0]), .S(_05558_), .Y(_24895_) );
  \$mux  #( .WIDTH(10) ) _46799_ ( .A(_24895_), .B(_25975_[9:0]), .S(_05307_), .Y(_24896_) );
  \$mux  #( .WIDTH(10) ) _46800_ ( .A(_24896_), .B(_25974_[9:0]), .S(_05559_), .Y(_24897_) );
  \$mux  #( .WIDTH(1) ) _46802_ ( .A(ram_w8_l2048_id10_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24898_) );
  \$mux  #( .WIDTH(1) ) _46803_ ( .A(_24898_), .B(_05189_), .S(_05307_), .Y(_24899_) );
  \$mux  #( .WIDTH(8) ) _46805_ ( .A(ram_w8_l2048_id10_0_1_wdata), .B(_dataflow_slice_data_30), .S(_05307_), .Y(_24900_) );
  \$mux  #( .WIDTH(9) ) _46807_ ( .A(ram_w8_l2048_id10_0_1_addr), .B(_tmp_167), .S(_05307_), .Y(_24901_) );
  \$mux  #( .WIDTH(9) ) _46809_ ( .A(ram_w8_l2048_id10_0_0_addr), .B(_stream_conv2d_8_source_19_source_ram_raddr[10:2]), .S(_tmp_367), .Y(_24902_) );
  \$mux  #( .WIDTH(1) ) _46811_ ( .A(ram_w8_l2048_id9_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24903_) );
  \$mux  #( .WIDTH(1) ) _46812_ ( .A(_24903_), .B(_05179_), .S(_05304_), .Y(_24904_) );
  \$mux  #( .WIDTH(8) ) _46814_ ( .A(ram_w8_l2048_id9_3_1_wdata), .B(_dataflow_slice_data_26), .S(_05304_), .Y(_24905_) );
  \$mux  #( .WIDTH(9) ) _46816_ ( .A(ram_w8_l2048_id9_3_1_addr), .B(_tmp_145), .S(_05304_), .Y(_24906_) );
  \$mux  #( .WIDTH(9) ) _46818_ ( .A(ram_w8_l2048_id9_3_0_addr), .B(_stream_conv2d_8_source_36_source_ram_raddr[10:2]), .S(_tmp_537), .Y(_24907_) );
  \$mux  #( .WIDTH(1) ) _46820_ ( .A(ram_w8_l2048_id9_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24908_) );
  \$mux  #( .WIDTH(1) ) _46821_ ( .A(_24908_), .B(_05170_), .S(_05301_), .Y(_24909_) );
  \$mux  #( .WIDTH(8) ) _46823_ ( .A(ram_w8_l2048_id9_2_1_wdata), .B(_dataflow_slice_data_23), .S(_05301_), .Y(_24910_) );
  \$mux  #( .WIDTH(9) ) _46825_ ( .A(ram_w8_l2048_id9_2_1_addr), .B(_tmp_114), .S(_05301_), .Y(_24911_) );
  \$mux  #( .WIDTH(9) ) _46827_ ( .A(ram_w8_l2048_id9_2_0_addr), .B(_stream_conv2d_8_source_36_source_ram_raddr[10:2]), .S(_tmp_537), .Y(_24912_) );
  \$mux  #( .WIDTH(1) ) _46829_ ( .A(ram_w8_l2048_id9_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24913_) );
  \$mux  #( .WIDTH(1) ) _46830_ ( .A(_24913_), .B(_05161_), .S(_05298_), .Y(_24914_) );
  \$mux  #( .WIDTH(8) ) _46832_ ( .A(ram_w8_l2048_id9_1_1_wdata), .B(_dataflow_slice_data_20), .S(_05298_), .Y(_24915_) );
  \$mux  #( .WIDTH(9) ) _46834_ ( .A(ram_w8_l2048_id9_1_1_addr), .B(_tmp_83), .S(_05298_), .Y(_24916_) );
  \$mux  #( .WIDTH(9) ) _46836_ ( .A(ram_w8_l2048_id9_1_0_addr), .B(_stream_conv2d_8_source_36_source_ram_raddr[10:2]), .S(_tmp_537), .Y(_24917_) );
  \$mux  #( .WIDTH(1) ) _46839_ ( .A(ram_w8_l2048_id9_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24918_) );
  \$mux  #( .WIDTH(1) ) _46840_ ( .A(_24918_), .B(_05152_), .S(_05295_), .Y(_24919_) );
  \$mux  #( .WIDTH(8) ) _46842_ ( .A(ram_w8_l2048_id9_0_1_wdata), .B(_dataflow_slice_data_17), .S(_05295_), .Y(_24920_) );
  \$mux  #( .WIDTH(9) ) _46844_ ( .A(ram_w8_l2048_id9_0_1_addr), .B(_tmp_52), .S(_05295_), .Y(_24921_) );
  \$mux  #( .WIDTH(9) ) _46846_ ( .A(ram_w8_l2048_id9_0_0_addr), .B(_stream_conv2d_8_source_36_source_ram_raddr[10:2]), .S(_tmp_537), .Y(_24922_) );
  \$mux  #( .WIDTH(1) ) _46848_ ( .A(ram_w8_l2048_id8_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24923_) );
  \$mux  #( .WIDTH(1) ) _46849_ ( .A(_24923_), .B(_05187_), .S(_05304_), .Y(_24924_) );
  \$mux  #( .WIDTH(8) ) _46851_ ( .A(ram_w8_l2048_id8_3_1_wdata), .B(_dataflow_slice_data_26), .S(_05304_), .Y(_24925_) );
  \$mux  #( .WIDTH(9) ) _46853_ ( .A(ram_w8_l2048_id8_3_1_addr), .B(_tmp_144), .S(_05304_), .Y(_24926_) );
  \$mux  #( .WIDTH(9) ) _46855_ ( .A(ram_w8_l2048_id8_3_0_addr), .B(_stream_conv2d_8_source_35_source_ram_raddr[10:2]), .S(_tmp_527), .Y(_24927_) );
  \$mux  #( .WIDTH(1) ) _46857_ ( .A(ram_w8_l2048_id8_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24928_) );
  \$mux  #( .WIDTH(1) ) _46858_ ( .A(_24928_), .B(_05178_), .S(_05301_), .Y(_24929_) );
  \$mux  #( .WIDTH(8) ) _46860_ ( .A(ram_w8_l2048_id8_2_1_wdata), .B(_dataflow_slice_data_23), .S(_05301_), .Y(_24930_) );
  \$mux  #( .WIDTH(9) ) _46862_ ( .A(ram_w8_l2048_id8_2_1_addr), .B(_tmp_113), .S(_05301_), .Y(_24931_) );
  \$mux  #( .WIDTH(9) ) _46864_ ( .A(ram_w8_l2048_id8_2_0_addr), .B(_stream_conv2d_8_source_35_source_ram_raddr[10:2]), .S(_tmp_527), .Y(_24932_) );
  \$mux  #( .WIDTH(1) ) _46866_ ( .A(ram_w8_l2048_id8_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24933_) );
  \$mux  #( .WIDTH(1) ) _46867_ ( .A(_24933_), .B(_05169_), .S(_05298_), .Y(_24934_) );
  \$mux  #( .WIDTH(8) ) _46869_ ( .A(ram_w8_l2048_id8_1_1_wdata), .B(_dataflow_slice_data_20), .S(_05298_), .Y(_24935_) );
  \$mux  #( .WIDTH(9) ) _46871_ ( .A(ram_w8_l2048_id8_1_1_addr), .B(_tmp_82), .S(_05298_), .Y(_24936_) );
  \$mux  #( .WIDTH(9) ) _46873_ ( .A(ram_w8_l2048_id8_1_0_addr), .B(_stream_conv2d_8_source_35_source_ram_raddr[10:2]), .S(_tmp_527), .Y(_24937_) );
  \$mux  #( .WIDTH(1) ) _46876_ ( .A(ram_w8_l2048_id8_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24938_) );
  \$mux  #( .WIDTH(1) ) _46877_ ( .A(_24938_), .B(_05160_), .S(_05295_), .Y(_24939_) );
  \$mux  #( .WIDTH(8) ) _46879_ ( .A(ram_w8_l2048_id8_0_1_wdata), .B(_dataflow_slice_data_17), .S(_05295_), .Y(_24940_) );
  \$mux  #( .WIDTH(9) ) _46881_ ( .A(ram_w8_l2048_id8_0_1_addr), .B(_tmp_51), .S(_05295_), .Y(_24941_) );
  \$mux  #( .WIDTH(9) ) _46883_ ( .A(ram_w8_l2048_id8_0_0_addr), .B(_stream_conv2d_8_source_35_source_ram_raddr[10:2]), .S(_tmp_527), .Y(_24942_) );
  \$mux  #( .WIDTH(1) ) _46885_ ( .A(ram_w8_l2048_id7_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24943_) );
  \$mux  #( .WIDTH(1) ) _46886_ ( .A(_24943_), .B(_05186_), .S(_05304_), .Y(_24944_) );
  \$mux  #( .WIDTH(8) ) _46888_ ( .A(ram_w8_l2048_id7_3_1_wdata), .B(_dataflow_slice_data_26), .S(_05304_), .Y(_24945_) );
  \$mux  #( .WIDTH(9) ) _46890_ ( .A(ram_w8_l2048_id7_3_1_addr), .B(_tmp_143), .S(_05304_), .Y(_24946_) );
  \$mux  #( .WIDTH(9) ) _46892_ ( .A(ram_w8_l2048_id7_3_0_addr), .B(_stream_conv2d_8_source_34_source_ram_raddr[10:2]), .S(_tmp_517), .Y(_24947_) );
  \$mux  #( .WIDTH(1) ) _46894_ ( .A(ram_w8_l2048_id7_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24948_) );
  \$mux  #( .WIDTH(1) ) _46895_ ( .A(_24948_), .B(_05177_), .S(_05301_), .Y(_24949_) );
  \$mux  #( .WIDTH(8) ) _46897_ ( .A(ram_w8_l2048_id7_2_1_wdata), .B(_dataflow_slice_data_23), .S(_05301_), .Y(_24950_) );
  \$mux  #( .WIDTH(9) ) _46899_ ( .A(ram_w8_l2048_id7_2_1_addr), .B(_tmp_112), .S(_05301_), .Y(_24951_) );
  \$mux  #( .WIDTH(9) ) _46901_ ( .A(ram_w8_l2048_id7_2_0_addr), .B(_stream_conv2d_8_source_34_source_ram_raddr[10:2]), .S(_tmp_517), .Y(_24952_) );
  \$mux  #( .WIDTH(1) ) _46903_ ( .A(ram_w8_l2048_id7_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24953_) );
  \$mux  #( .WIDTH(1) ) _46904_ ( .A(_24953_), .B(_05168_), .S(_05298_), .Y(_24954_) );
  \$mux  #( .WIDTH(8) ) _46906_ ( .A(ram_w8_l2048_id7_1_1_wdata), .B(_dataflow_slice_data_20), .S(_05298_), .Y(_24955_) );
  \$mux  #( .WIDTH(9) ) _46908_ ( .A(ram_w8_l2048_id7_1_1_addr), .B(_tmp_81), .S(_05298_), .Y(_24956_) );
  \$mux  #( .WIDTH(9) ) _46910_ ( .A(ram_w8_l2048_id7_1_0_addr), .B(_stream_conv2d_8_source_34_source_ram_raddr[10:2]), .S(_tmp_517), .Y(_24957_) );
  \$mux  #( .WIDTH(1) ) _46913_ ( .A(ram_w8_l2048_id7_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24958_) );
  \$mux  #( .WIDTH(1) ) _46914_ ( .A(_24958_), .B(_05159_), .S(_05295_), .Y(_24959_) );
  \$mux  #( .WIDTH(8) ) _46916_ ( .A(ram_w8_l2048_id7_0_1_wdata), .B(_dataflow_slice_data_17), .S(_05295_), .Y(_24960_) );
  \$mux  #( .WIDTH(9) ) _46918_ ( .A(ram_w8_l2048_id7_0_1_addr), .B(_tmp_50), .S(_05295_), .Y(_24961_) );
  \$mux  #( .WIDTH(9) ) _46920_ ( .A(ram_w8_l2048_id7_0_0_addr), .B(_stream_conv2d_8_source_34_source_ram_raddr[10:2]), .S(_tmp_517), .Y(_24962_) );
  \$mux  #( .WIDTH(1) ) _46922_ ( .A(ram_w8_l2048_id6_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24963_) );
  \$mux  #( .WIDTH(1) ) _46923_ ( .A(_24963_), .B(_05185_), .S(_05304_), .Y(_24964_) );
  \$mux  #( .WIDTH(8) ) _46925_ ( .A(ram_w8_l2048_id6_3_1_wdata), .B(_dataflow_slice_data_26), .S(_05304_), .Y(_24965_) );
  \$mux  #( .WIDTH(9) ) _46927_ ( .A(ram_w8_l2048_id6_3_1_addr), .B(_tmp_142), .S(_05304_), .Y(_24966_) );
  \$mux  #( .WIDTH(9) ) _46929_ ( .A(ram_w8_l2048_id6_3_0_addr), .B(_stream_conv2d_8_source_33_source_ram_raddr[10:2]), .S(_tmp_507), .Y(_24967_) );
  \$mux  #( .WIDTH(1) ) _46931_ ( .A(ram_w8_l2048_id6_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24968_) );
  \$mux  #( .WIDTH(1) ) _46932_ ( .A(_24968_), .B(_05176_), .S(_05301_), .Y(_24969_) );
  \$mux  #( .WIDTH(8) ) _46934_ ( .A(ram_w8_l2048_id6_2_1_wdata), .B(_dataflow_slice_data_23), .S(_05301_), .Y(_24970_) );
  \$mux  #( .WIDTH(9) ) _46936_ ( .A(ram_w8_l2048_id6_2_1_addr), .B(_tmp_111), .S(_05301_), .Y(_24971_) );
  \$mux  #( .WIDTH(9) ) _46938_ ( .A(ram_w8_l2048_id6_2_0_addr), .B(_stream_conv2d_8_source_33_source_ram_raddr[10:2]), .S(_tmp_507), .Y(_24972_) );
  \$mux  #( .WIDTH(1) ) _46940_ ( .A(ram_w8_l2048_id6_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24973_) );
  \$mux  #( .WIDTH(1) ) _46941_ ( .A(_24973_), .B(_05167_), .S(_05298_), .Y(_24974_) );
  \$mux  #( .WIDTH(8) ) _46943_ ( .A(ram_w8_l2048_id6_1_1_wdata), .B(_dataflow_slice_data_20), .S(_05298_), .Y(_24975_) );
  \$mux  #( .WIDTH(9) ) _46945_ ( .A(ram_w8_l2048_id6_1_1_addr), .B(_tmp_80), .S(_05298_), .Y(_24976_) );
  \$mux  #( .WIDTH(9) ) _46947_ ( .A(ram_w8_l2048_id6_1_0_addr), .B(_stream_conv2d_8_source_33_source_ram_raddr[10:2]), .S(_tmp_507), .Y(_24977_) );
  \$mux  #( .WIDTH(1) ) _46950_ ( .A(ram_w8_l2048_id6_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24978_) );
  \$mux  #( .WIDTH(1) ) _46951_ ( .A(_24978_), .B(_05158_), .S(_05295_), .Y(_24979_) );
  \$mux  #( .WIDTH(8) ) _46953_ ( .A(ram_w8_l2048_id6_0_1_wdata), .B(_dataflow_slice_data_17), .S(_05295_), .Y(_24980_) );
  \$mux  #( .WIDTH(9) ) _46955_ ( .A(ram_w8_l2048_id6_0_1_addr), .B(_tmp_49), .S(_05295_), .Y(_24981_) );
  \$mux  #( .WIDTH(9) ) _46957_ ( .A(ram_w8_l2048_id6_0_0_addr), .B(_stream_conv2d_8_source_33_source_ram_raddr[10:2]), .S(_tmp_507), .Y(_24982_) );
  \$mux  #( .WIDTH(1) ) _46959_ ( .A(ram_w8_l2048_id5_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24983_) );
  \$mux  #( .WIDTH(1) ) _46960_ ( .A(_24983_), .B(_05184_), .S(_05304_), .Y(_24984_) );
  \$mux  #( .WIDTH(8) ) _46962_ ( .A(ram_w8_l2048_id5_3_1_wdata), .B(_dataflow_slice_data_26), .S(_05304_), .Y(_24985_) );
  \$mux  #( .WIDTH(9) ) _46964_ ( .A(ram_w8_l2048_id5_3_1_addr), .B(_tmp_141), .S(_05304_), .Y(_24986_) );
  \$mux  #( .WIDTH(9) ) _46966_ ( .A(ram_w8_l2048_id5_3_0_addr), .B(_stream_conv2d_8_source_32_source_ram_raddr[10:2]), .S(_tmp_497), .Y(_24987_) );
  \$mux  #( .WIDTH(1) ) _46968_ ( .A(ram_w8_l2048_id5_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24988_) );
  \$mux  #( .WIDTH(1) ) _46969_ ( .A(_24988_), .B(_05175_), .S(_05301_), .Y(_24989_) );
  \$mux  #( .WIDTH(8) ) _46971_ ( .A(ram_w8_l2048_id5_2_1_wdata), .B(_dataflow_slice_data_23), .S(_05301_), .Y(_24990_) );
  \$mux  #( .WIDTH(9) ) _46973_ ( .A(ram_w8_l2048_id5_2_1_addr), .B(_tmp_110), .S(_05301_), .Y(_24991_) );
  \$mux  #( .WIDTH(9) ) _46975_ ( .A(ram_w8_l2048_id5_2_0_addr), .B(_stream_conv2d_8_source_32_source_ram_raddr[10:2]), .S(_tmp_497), .Y(_24992_) );
  \$mux  #( .WIDTH(1) ) _46977_ ( .A(ram_w8_l2048_id5_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24993_) );
  \$mux  #( .WIDTH(1) ) _46978_ ( .A(_24993_), .B(_05166_), .S(_05298_), .Y(_24994_) );
  \$mux  #( .WIDTH(8) ) _46980_ ( .A(ram_w8_l2048_id5_1_1_wdata), .B(_dataflow_slice_data_20), .S(_05298_), .Y(_24995_) );
  \$mux  #( .WIDTH(9) ) _46982_ ( .A(ram_w8_l2048_id5_1_1_addr), .B(_tmp_79), .S(_05298_), .Y(_24996_) );
  \$mux  #( .WIDTH(9) ) _46984_ ( .A(ram_w8_l2048_id5_1_0_addr), .B(_stream_conv2d_8_source_32_source_ram_raddr[10:2]), .S(_tmp_497), .Y(_24997_) );
  \$mux  #( .WIDTH(1) ) _46987_ ( .A(ram_w8_l2048_id5_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_24998_) );
  \$mux  #( .WIDTH(1) ) _46988_ ( .A(_24998_), .B(_05157_), .S(_05295_), .Y(_24999_) );
  \$mux  #( .WIDTH(8) ) _46990_ ( .A(ram_w8_l2048_id5_0_1_wdata), .B(_dataflow_slice_data_17), .S(_05295_), .Y(_25000_) );
  \$mux  #( .WIDTH(9) ) _46992_ ( .A(ram_w8_l2048_id5_0_1_addr), .B(_tmp_48), .S(_05295_), .Y(_25001_) );
  \$mux  #( .WIDTH(9) ) _46994_ ( .A(ram_w8_l2048_id5_0_0_addr), .B(_stream_conv2d_8_source_32_source_ram_raddr[10:2]), .S(_tmp_497), .Y(_25002_) );
  \$mux  #( .WIDTH(1) ) _46996_ ( .A(ram_w8_l2048_id4_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25003_) );
  \$mux  #( .WIDTH(1) ) _46997_ ( .A(_25003_), .B(_05183_), .S(_05304_), .Y(_25004_) );
  \$mux  #( .WIDTH(8) ) _46999_ ( .A(ram_w8_l2048_id4_3_1_wdata), .B(_dataflow_slice_data_26), .S(_05304_), .Y(_25005_) );
  \$mux  #( .WIDTH(9) ) _47001_ ( .A(ram_w8_l2048_id4_3_1_addr), .B(_tmp_140), .S(_05304_), .Y(_25006_) );
  \$mux  #( .WIDTH(9) ) _47003_ ( .A(ram_w8_l2048_id4_3_0_addr), .B(_stream_conv2d_8_source_31_source_ram_raddr[10:2]), .S(_tmp_487), .Y(_25007_) );
  \$mux  #( .WIDTH(1) ) _47005_ ( .A(ram_w8_l2048_id4_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25008_) );
  \$mux  #( .WIDTH(1) ) _47006_ ( .A(_25008_), .B(_05174_), .S(_05301_), .Y(_25009_) );
  \$mux  #( .WIDTH(8) ) _47008_ ( .A(ram_w8_l2048_id4_2_1_wdata), .B(_dataflow_slice_data_23), .S(_05301_), .Y(_25010_) );
  \$mux  #( .WIDTH(9) ) _47010_ ( .A(ram_w8_l2048_id4_2_1_addr), .B(_tmp_109), .S(_05301_), .Y(_25011_) );
  \$mux  #( .WIDTH(9) ) _47012_ ( .A(ram_w8_l2048_id4_2_0_addr), .B(_stream_conv2d_8_source_31_source_ram_raddr[10:2]), .S(_tmp_487), .Y(_25012_) );
  \$mux  #( .WIDTH(1) ) _47014_ ( .A(ram_w8_l2048_id4_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25013_) );
  \$mux  #( .WIDTH(1) ) _47015_ ( .A(_25013_), .B(_05165_), .S(_05298_), .Y(_25014_) );
  \$mux  #( .WIDTH(8) ) _47017_ ( .A(ram_w8_l2048_id4_1_1_wdata), .B(_dataflow_slice_data_20), .S(_05298_), .Y(_25015_) );
  \$mux  #( .WIDTH(9) ) _47019_ ( .A(ram_w8_l2048_id4_1_1_addr), .B(_tmp_78), .S(_05298_), .Y(_25016_) );
  \$mux  #( .WIDTH(9) ) _47021_ ( .A(ram_w8_l2048_id4_1_0_addr), .B(_stream_conv2d_8_source_31_source_ram_raddr[10:2]), .S(_tmp_487), .Y(_25017_) );
  \$mux  #( .WIDTH(1) ) _47024_ ( .A(ram_w8_l2048_id4_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25018_) );
  \$mux  #( .WIDTH(1) ) _47025_ ( .A(_25018_), .B(_05156_), .S(_05295_), .Y(_25019_) );
  \$mux  #( .WIDTH(8) ) _47027_ ( .A(ram_w8_l2048_id4_0_1_wdata), .B(_dataflow_slice_data_17), .S(_05295_), .Y(_25020_) );
  \$mux  #( .WIDTH(9) ) _47029_ ( .A(ram_w8_l2048_id4_0_1_addr), .B(_tmp_47), .S(_05295_), .Y(_25021_) );
  \$mux  #( .WIDTH(9) ) _47031_ ( .A(ram_w8_l2048_id4_0_0_addr), .B(_stream_conv2d_8_source_31_source_ram_raddr[10:2]), .S(_tmp_487), .Y(_25022_) );
  \$mux  #( .WIDTH(1) ) _47033_ ( .A(ram_w8_l2048_id3_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25023_) );
  \$mux  #( .WIDTH(1) ) _47034_ ( .A(_25023_), .B(_05182_), .S(_05304_), .Y(_25024_) );
  \$mux  #( .WIDTH(8) ) _47036_ ( .A(ram_w8_l2048_id3_3_1_wdata), .B(_dataflow_slice_data_26), .S(_05304_), .Y(_25025_) );
  \$mux  #( .WIDTH(9) ) _47038_ ( .A(ram_w8_l2048_id3_3_1_addr), .B(_tmp_139), .S(_05304_), .Y(_25026_) );
  \$mux  #( .WIDTH(9) ) _47040_ ( .A(ram_w8_l2048_id3_3_0_addr), .B(_stream_conv2d_8_source_30_source_ram_raddr[10:2]), .S(_tmp_477), .Y(_25027_) );
  \$mux  #( .WIDTH(1) ) _47042_ ( .A(ram_w8_l2048_id3_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25028_) );
  \$mux  #( .WIDTH(1) ) _47043_ ( .A(_25028_), .B(_05173_), .S(_05301_), .Y(_25029_) );
  \$mux  #( .WIDTH(8) ) _47045_ ( .A(ram_w8_l2048_id3_2_1_wdata), .B(_dataflow_slice_data_23), .S(_05301_), .Y(_25030_) );
  \$mux  #( .WIDTH(9) ) _47047_ ( .A(ram_w8_l2048_id3_2_1_addr), .B(_tmp_108), .S(_05301_), .Y(_25031_) );
  \$mux  #( .WIDTH(9) ) _47049_ ( .A(ram_w8_l2048_id3_2_0_addr), .B(_stream_conv2d_8_source_30_source_ram_raddr[10:2]), .S(_tmp_477), .Y(_25032_) );
  \$mux  #( .WIDTH(1) ) _47051_ ( .A(ram_w8_l2048_id3_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25033_) );
  \$mux  #( .WIDTH(1) ) _47052_ ( .A(_25033_), .B(_05164_), .S(_05298_), .Y(_25034_) );
  \$mux  #( .WIDTH(8) ) _47054_ ( .A(ram_w8_l2048_id3_1_1_wdata), .B(_dataflow_slice_data_20), .S(_05298_), .Y(_25035_) );
  \$mux  #( .WIDTH(9) ) _47056_ ( .A(ram_w8_l2048_id3_1_1_addr), .B(_tmp_77), .S(_05298_), .Y(_25036_) );
  \$mux  #( .WIDTH(9) ) _47058_ ( .A(ram_w8_l2048_id3_1_0_addr), .B(_stream_conv2d_8_source_30_source_ram_raddr[10:2]), .S(_tmp_477), .Y(_25037_) );
  \$mux  #( .WIDTH(1) ) _47061_ ( .A(ram_w8_l2048_id3_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25038_) );
  \$mux  #( .WIDTH(1) ) _47062_ ( .A(_25038_), .B(_05155_), .S(_05295_), .Y(_25039_) );
  \$mux  #( .WIDTH(8) ) _47064_ ( .A(ram_w8_l2048_id3_0_1_wdata), .B(_dataflow_slice_data_17), .S(_05295_), .Y(_25040_) );
  \$mux  #( .WIDTH(9) ) _47066_ ( .A(ram_w8_l2048_id3_0_1_addr), .B(_tmp_46), .S(_05295_), .Y(_25041_) );
  \$mux  #( .WIDTH(9) ) _47068_ ( .A(ram_w8_l2048_id3_0_0_addr), .B(_stream_conv2d_8_source_30_source_ram_raddr[10:2]), .S(_tmp_477), .Y(_25042_) );
  \$mux  #( .WIDTH(1) ) _47070_ ( .A(_tmp_982), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25043_) );
  \$mux  #( .WIDTH(1) ) _47071_ ( .A(_25043_), .B(1'h1), .S(_05556_), .Y(_25044_) );
  \$mux  #( .WIDTH(34) ) _47073_ ( .A(_tmp_981), .B({ 1'h0, _maxi_read_size }), .S(_05555_), .Y(_25045_) );
  \$mux  #( .WIDTH(34) ) _47074_ ( .A(_25045_), .B(_25973_), .S(_05376_), .Y(_25046_) );
  \$mux  #( .WIDTH(1) ) _47076_ ( .A(ram_w8_l2048_id2_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25047_) );
  \$mux  #( .WIDTH(1) ) _47077_ ( .A(_25047_), .B(_05181_), .S(_05304_), .Y(_25048_) );
  \$mux  #( .WIDTH(1) ) _47078_ ( .A(_25048_), .B(1'h1), .S(_05376_), .Y(_25049_) );
  \$mux  #( .WIDTH(8) ) _47080_ ( .A(ram_w8_l2048_id2_3_1_wdata), .B(_dataflow_slice_data_26), .S(_05304_), .Y(_25050_) );
  \$mux  #( .WIDTH(8) ) _47081_ ( .A(_25050_), .B(_dataflow_slice_data_122), .S(_05376_), .Y(_25051_) );
  \$mux  #( .WIDTH(9) ) _47083_ ( .A(ram_w8_l2048_id2_3_1_addr), .B(_tmp_138), .S(_05304_), .Y(_25052_) );
  \$mux  #( .WIDTH(9) ) _47084_ ( .A(_25052_), .B(_25939_[8:0]), .S(_05555_), .Y(_25053_) );
  \$mux  #( .WIDTH(9) ) _47085_ ( .A(_25053_), .B(_22104_[8:0]), .S(_05376_), .Y(_25054_) );
  \$mux  #( .WIDTH(9) ) _47087_ ( .A(ram_w8_l2048_id2_3_0_addr), .B(_stream_conv2d_8_source_29_source_ram_raddr[10:2]), .S(_tmp_467), .Y(_25055_) );
  \$mux  #( .WIDTH(9) ) _47088_ ( .A(_25055_), .B(_stream_matmul_15_source_19_source_ram_raddr[10:2]), .S(_tmp_1023), .Y(_25056_) );
  \$mux  #( .WIDTH(1) ) _47090_ ( .A(_tmp_980), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25057_) );
  \$mux  #( .WIDTH(1) ) _47091_ ( .A(_25057_), .B(1'h1), .S(_05554_), .Y(_25058_) );
  \$mux  #( .WIDTH(34) ) _47093_ ( .A(_tmp_979), .B({ 1'h0, _maxi_read_size }), .S(_05553_), .Y(_25059_) );
  \$mux  #( .WIDTH(34) ) _47094_ ( .A(_25059_), .B(_25972_), .S(_05373_), .Y(_25060_) );
  \$mux  #( .WIDTH(1) ) _47096_ ( .A(ram_w8_l2048_id2_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25061_) );
  \$mux  #( .WIDTH(1) ) _47097_ ( .A(_25061_), .B(_05172_), .S(_05301_), .Y(_25062_) );
  \$mux  #( .WIDTH(1) ) _47098_ ( .A(_25062_), .B(1'h1), .S(_05373_), .Y(_25063_) );
  \$mux  #( .WIDTH(8) ) _47100_ ( .A(ram_w8_l2048_id2_2_1_wdata), .B(_dataflow_slice_data_23), .S(_05301_), .Y(_25064_) );
  \$mux  #( .WIDTH(8) ) _47101_ ( .A(_25064_), .B(_dataflow_slice_data_119), .S(_05373_), .Y(_25065_) );
  \$mux  #( .WIDTH(9) ) _47103_ ( .A(ram_w8_l2048_id2_2_1_addr), .B(_tmp_107), .S(_05301_), .Y(_25066_) );
  \$mux  #( .WIDTH(9) ) _47104_ ( .A(_25066_), .B(_25939_[8:0]), .S(_05553_), .Y(_25067_) );
  \$mux  #( .WIDTH(9) ) _47105_ ( .A(_25067_), .B(_22103_[8:0]), .S(_05373_), .Y(_25068_) );
  \$mux  #( .WIDTH(9) ) _47107_ ( .A(ram_w8_l2048_id2_2_0_addr), .B(_stream_conv2d_8_source_29_source_ram_raddr[10:2]), .S(_tmp_467), .Y(_25069_) );
  \$mux  #( .WIDTH(9) ) _47108_ ( .A(_25069_), .B(_stream_matmul_15_source_19_source_ram_raddr[10:2]), .S(_tmp_1023), .Y(_25070_) );
  \$mux  #( .WIDTH(1) ) _47110_ ( .A(_tmp_978), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25071_) );
  \$mux  #( .WIDTH(1) ) _47111_ ( .A(_25071_), .B(1'h1), .S(_05552_), .Y(_25072_) );
  \$mux  #( .WIDTH(34) ) _47113_ ( .A(_tmp_977), .B({ 1'h0, _maxi_read_size }), .S(_05551_), .Y(_25073_) );
  \$mux  #( .WIDTH(34) ) _47114_ ( .A(_25073_), .B(_25971_), .S(_05370_), .Y(_25074_) );
  \$mux  #( .WIDTH(1) ) _47116_ ( .A(ram_w8_l2048_id2_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25075_) );
  \$mux  #( .WIDTH(1) ) _47117_ ( .A(_25075_), .B(_05163_), .S(_05298_), .Y(_25076_) );
  \$mux  #( .WIDTH(1) ) _47118_ ( .A(_25076_), .B(1'h1), .S(_05370_), .Y(_25077_) );
  \$mux  #( .WIDTH(8) ) _47120_ ( .A(ram_w8_l2048_id2_1_1_wdata), .B(_dataflow_slice_data_20), .S(_05298_), .Y(_25078_) );
  \$mux  #( .WIDTH(8) ) _47121_ ( .A(_25078_), .B(_dataflow_slice_data_116), .S(_05370_), .Y(_25079_) );
  \$mux  #( .WIDTH(9) ) _47123_ ( .A(ram_w8_l2048_id2_1_1_addr), .B(_tmp_76), .S(_05298_), .Y(_25080_) );
  \$mux  #( .WIDTH(9) ) _47124_ ( .A(_25080_), .B(_25939_[8:0]), .S(_05551_), .Y(_25081_) );
  \$mux  #( .WIDTH(9) ) _47125_ ( .A(_25081_), .B(_22102_[8:0]), .S(_05370_), .Y(_25082_) );
  \$mux  #( .WIDTH(9) ) _47127_ ( .A(ram_w8_l2048_id2_1_0_addr), .B(_stream_conv2d_8_source_29_source_ram_raddr[10:2]), .S(_tmp_467), .Y(_25083_) );
  \$mux  #( .WIDTH(9) ) _47128_ ( .A(_25083_), .B(_stream_matmul_15_source_19_source_ram_raddr[10:2]), .S(_tmp_1023), .Y(_25084_) );
  \$mux  #( .WIDTH(1) ) _47131_ ( .A(_tmp_976), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25085_) );
  \$mux  #( .WIDTH(1) ) _47132_ ( .A(_25085_), .B(1'h1), .S(_05550_), .Y(_25086_) );
  \$mux  #( .WIDTH(34) ) _47134_ ( .A(_tmp_975), .B({ 1'h0, _maxi_read_size }), .S(_05549_), .Y(_25087_) );
  \$mux  #( .WIDTH(34) ) _47135_ ( .A(_25087_), .B(_25970_), .S(_05367_), .Y(_25088_) );
  \$mux  #( .WIDTH(1) ) _47138_ ( .A(ram_w8_l2048_id2_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25089_) );
  \$mux  #( .WIDTH(1) ) _47139_ ( .A(_25089_), .B(_05154_), .S(_05295_), .Y(_25090_) );
  \$mux  #( .WIDTH(1) ) _47140_ ( .A(_25090_), .B(1'h1), .S(_05367_), .Y(_25091_) );
  \$mux  #( .WIDTH(8) ) _47142_ ( .A(ram_w8_l2048_id2_0_1_wdata), .B(_dataflow_slice_data_17), .S(_05295_), .Y(_25092_) );
  \$mux  #( .WIDTH(8) ) _47143_ ( .A(_25092_), .B(_dataflow_slice_data_113), .S(_05367_), .Y(_25093_) );
  \$mux  #( .WIDTH(9) ) _47145_ ( .A(ram_w8_l2048_id2_0_1_addr), .B(_tmp_45), .S(_05295_), .Y(_25094_) );
  \$mux  #( .WIDTH(9) ) _47146_ ( .A(_25094_), .B(_25939_[8:0]), .S(_05549_), .Y(_25095_) );
  \$mux  #( .WIDTH(9) ) _47147_ ( .A(_25095_), .B(_22101_[8:0]), .S(_05367_), .Y(_25096_) );
  \$mux  #( .WIDTH(9) ) _47149_ ( .A(ram_w8_l2048_id2_0_0_addr), .B(_stream_conv2d_8_source_29_source_ram_raddr[10:2]), .S(_tmp_467), .Y(_25097_) );
  \$mux  #( .WIDTH(9) ) _47150_ ( .A(_25097_), .B(_stream_matmul_15_source_19_source_ram_raddr[10:2]), .S(_tmp_1023), .Y(_25098_) );
  \$mux  #( .WIDTH(34) ) _47152_ ( .A(_tmp_1166), .B(_25945_), .S(_05545_), .Y(_25099_) );
  \$mux  #( .WIDTH(34) ) _47153_ ( .A(_25099_), .B(_25969_), .S(_05546_), .Y(_25100_) );
  \$mux  #( .WIDTH(1) ) _47155_ ( .A(_tmp_1165), .B(1'h0), .S(_05543_), .Y(_25101_) );
  \$mux  #( .WIDTH(1) ) _47156_ ( .A(_25101_), .B(_tmp_1164), .S(_05544_), .Y(_25102_) );
  \$mux  #( .WIDTH(1) ) _47158_ ( .A(_tmp_1164), .B(1'h0), .S(_05544_), .Y(_25103_) );
  \$mux  #( .WIDTH(1) ) _47159_ ( .A(_25103_), .B(_05151_), .S(_05545_), .Y(_25104_) );
  \$mux  #( .WIDTH(1) ) _47160_ ( .A(_25104_), .B(1'h0), .S(_05546_), .Y(_25105_) );
  \$mux  #( .WIDTH(1) ) _47161_ ( .A(_25105_), .B(1'h1), .S(_05547_), .Y(_25106_) );
  \$mux  #( .WIDTH(1) ) _47163_ ( .A(_tmp_1163), .B(1'h0), .S(_05543_), .Y(_25107_) );
  \$mux  #( .WIDTH(1) ) _47164_ ( .A(_25107_), .B(1'h1), .S(_05544_), .Y(_25108_) );
  \$mux  #( .WIDTH(1) ) _47166_ ( .A(_tmp_1162), .B(1'h0), .S(_05544_), .Y(_25109_) );
  \$mux  #( .WIDTH(1) ) _47167_ ( .A(_25109_), .B(1'h1), .S(_05545_), .Y(_25110_) );
  \$mux  #( .WIDTH(1) ) _47168_ ( .A(_25110_), .B(1'h1), .S(_05546_), .Y(_25111_) );
  \$mux  #( .WIDTH(1) ) _47172_ ( .A(_tmp_1155), .B(1'h0), .S(_05543_), .Y(_25112_) );
  \$mux  #( .WIDTH(1) ) _47173_ ( .A(_25112_), .B(1'h1), .S(_05544_), .Y(_25113_) );
  \$mux  #( .WIDTH(1) ) _47176_ ( .A(_tmp_860), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25114_) );
  \$mux  #( .WIDTH(1) ) _47177_ ( .A(_25114_), .B(1'h1), .S(_05541_), .Y(_25115_) );
  \$mux  #( .WIDTH(34) ) _47179_ ( .A(_tmp_859), .B({ 1'h0, _maxi_read_size }), .S(_05540_), .Y(_25116_) );
  \$mux  #( .WIDTH(34) ) _47180_ ( .A(_25116_), .B(_25968_), .S(_05352_), .Y(_25117_) );
  \$mux  #( .WIDTH(4) ) _47182_ ( .A(_tmp_155), .B(4'h0), .S(_05527_), .Y(_25118_) );
  \$mux  #( .WIDTH(4) ) _47183_ ( .A(_25118_), .B(_22098_[3:0]), .S(_05528_), .Y(_25119_) );
  \$mux  #( .WIDTH(4) ) _47184_ ( .A(_25119_), .B(4'h0), .S(_05529_), .Y(_25120_) );
  \$mux  #( .WIDTH(9) ) _47186_ ( .A(_tmp_136), .B(_25939_[8:0]), .S(_05527_), .Y(_25121_) );
  \$mux  #( .WIDTH(9) ) _47187_ ( .A(_25121_), .B(_tmp_145), .S(_05538_), .Y(_25122_) );
  \$mux  #( .WIDTH(9) ) _47189_ ( .A(_tmp_135), .B(_25939_[8:0]), .S(_05527_), .Y(_25123_) );
  \$mux  #( .WIDTH(9) ) _47190_ ( .A(_25123_), .B(_tmp_144), .S(_05537_), .Y(_25124_) );
  \$mux  #( .WIDTH(9) ) _47192_ ( .A(_tmp_134), .B(_25939_[8:0]), .S(_05527_), .Y(_25125_) );
  \$mux  #( .WIDTH(9) ) _47193_ ( .A(_25125_), .B(_tmp_143), .S(_05536_), .Y(_25126_) );
  \$mux  #( .WIDTH(9) ) _47195_ ( .A(_tmp_133), .B(_25939_[8:0]), .S(_05527_), .Y(_25127_) );
  \$mux  #( .WIDTH(9) ) _47196_ ( .A(_25127_), .B(_tmp_142), .S(_05535_), .Y(_25128_) );
  \$mux  #( .WIDTH(9) ) _47198_ ( .A(_tmp_132), .B(_25939_[8:0]), .S(_05527_), .Y(_25129_) );
  \$mux  #( .WIDTH(9) ) _47199_ ( .A(_25129_), .B(_tmp_141), .S(_05534_), .Y(_25130_) );
  \$mux  #( .WIDTH(9) ) _47201_ ( .A(_tmp_131), .B(_25939_[8:0]), .S(_05527_), .Y(_25131_) );
  \$mux  #( .WIDTH(9) ) _47202_ ( .A(_25131_), .B(_tmp_140), .S(_05533_), .Y(_25132_) );
  \$mux  #( .WIDTH(9) ) _47204_ ( .A(_tmp_130), .B(_25939_[8:0]), .S(_05527_), .Y(_25133_) );
  \$mux  #( .WIDTH(9) ) _47205_ ( .A(_25133_), .B(_tmp_139), .S(_05532_), .Y(_25134_) );
  \$mux  #( .WIDTH(9) ) _47207_ ( .A(_tmp_129), .B(_25939_[8:0]), .S(_05527_), .Y(_25135_) );
  \$mux  #( .WIDTH(9) ) _47208_ ( .A(_25135_), .B(_tmp_138), .S(_05531_), .Y(_25136_) );
  \$mux  #( .WIDTH(9) ) _47210_ ( .A(_tmp_128), .B(_25939_[8:0]), .S(_05527_), .Y(_25137_) );
  \$mux  #( .WIDTH(9) ) _47211_ ( .A(_25137_), .B(_tmp_137), .S(_05530_), .Y(_25138_) );
  \$mux  #( .WIDTH(1) ) _47213_ ( .A(_tmp_127), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25139_) );
  \$mux  #( .WIDTH(1) ) _47214_ ( .A(_25139_), .B(1'h1), .S(_05539_), .Y(_25140_) );
  \$mux  #( .WIDTH(34) ) _47216_ ( .A(_tmp_126), .B({ 1'h0, _maxi_read_size }), .S(_05527_), .Y(_25141_) );
  \$mux  #( .WIDTH(34) ) _47217_ ( .A(_25141_), .B(_25967_), .S(_05304_), .Y(_25142_) );
  \$mux  #( .WIDTH(10) ) _47219_ ( .A(_tmp_125), .B(_25953_[9:0]), .S(_05527_), .Y(_25143_) );
  \$mux  #( .WIDTH(10) ) _47220_ ( .A(_25143_), .B(_25966_[9:0]), .S(_05304_), .Y(_25144_) );
  \$mux  #( .WIDTH(10) ) _47221_ ( .A(_25144_), .B(_25953_[9:0]), .S(_05528_), .Y(_25145_) );
  \$mux  #( .WIDTH(1) ) _47223_ ( .A(ram_w8_l2048_id1_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25146_) );
  \$mux  #( .WIDTH(1) ) _47224_ ( .A(_25146_), .B(_05180_), .S(_05304_), .Y(_25147_) );
  \$mux  #( .WIDTH(1) ) _47225_ ( .A(_25147_), .B(1'h1), .S(_05352_), .Y(_25148_) );
  \$mux  #( .WIDTH(8) ) _47227_ ( .A(ram_w8_l2048_id1_3_1_wdata), .B(_dataflow_slice_data_26), .S(_05304_), .Y(_25149_) );
  \$mux  #( .WIDTH(8) ) _47228_ ( .A(_25149_), .B(_dataflow_slice_data_87), .S(_05352_), .Y(_25150_) );
  \$mux  #( .WIDTH(9) ) _47230_ ( .A(ram_w8_l2048_id1_3_1_addr), .B(_tmp_137), .S(_05304_), .Y(_25151_) );
  \$mux  #( .WIDTH(9) ) _47231_ ( .A(_25151_), .B(_25939_[8:0]), .S(_05540_), .Y(_25152_) );
  \$mux  #( .WIDTH(9) ) _47232_ ( .A(_25152_), .B(_22099_[8:0]), .S(_05352_), .Y(_25153_) );
  \$mux  #( .WIDTH(9) ) _47233_ ( .A(_25153_), .B(_maxi_write_local_addr[8:0]), .S(_05545_), .Y(_25154_) );
  \$mux  #( .WIDTH(9) ) _47234_ ( .A(_25154_), .B(_22100_[8:0]), .S(_05546_), .Y(_25155_) );
  \$mux  #( .WIDTH(1) ) _47236_ ( .A(ram_w8_l2048_id1_3_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id1_3_cond_7_1), .Y(_25156_) );
  \$mux  #( .WIDTH(1) ) _47237_ ( .A(_25156_), .B(1'h1), .S(_05542_), .Y(_25157_) );
  \$mux  #( .WIDTH(8) ) _47239_ ( .A(ram_w8_l2048_id1_3_0_wdata), .B(_stream_matmul_15_sink_21_sink_wdata), .S(_05542_), .Y(_25158_) );
  \$mux  #( .WIDTH(9) ) _47241_ ( .A(ram_w8_l2048_id1_3_0_addr), .B(_stream_conv2d_8_source_28_source_ram_raddr[10:2]), .S(_tmp_457), .Y(_25159_) );
  \$mux  #( .WIDTH(9) ) _47242_ ( .A(_25159_), .B(_stream_max_pool_serial_9_source_1_source_ram_raddr[10:2]), .S(_tmp_873), .Y(_25160_) );
  \$mux  #( .WIDTH(9) ) _47243_ ( .A(_25160_), .B(_stream_matmul_15_sink_21_sink_waddr[10:2]), .S(_05542_), .Y(_25161_) );
  \$mux  #( .WIDTH(34) ) _47245_ ( .A(_tmp_1154), .B(_25945_), .S(_05524_), .Y(_25162_) );
  \$mux  #( .WIDTH(34) ) _47246_ ( .A(_25162_), .B(_25965_), .S(_05525_), .Y(_25163_) );
  \$mux  #( .WIDTH(1) ) _47248_ ( .A(_tmp_1153), .B(1'h0), .S(_05522_), .Y(_25164_) );
  \$mux  #( .WIDTH(1) ) _47249_ ( .A(_25164_), .B(_tmp_1152), .S(_05523_), .Y(_25165_) );
  \$mux  #( .WIDTH(1) ) _47251_ ( .A(_tmp_1152), .B(1'h0), .S(_05523_), .Y(_25166_) );
  \$mux  #( .WIDTH(1) ) _47252_ ( .A(_25166_), .B(_05151_), .S(_05524_), .Y(_25167_) );
  \$mux  #( .WIDTH(1) ) _47253_ ( .A(_25167_), .B(1'h0), .S(_05525_), .Y(_25168_) );
  \$mux  #( .WIDTH(1) ) _47254_ ( .A(_25168_), .B(1'h1), .S(_05526_), .Y(_25169_) );
  \$mux  #( .WIDTH(1) ) _47256_ ( .A(_tmp_1151), .B(1'h0), .S(_05522_), .Y(_25170_) );
  \$mux  #( .WIDTH(1) ) _47257_ ( .A(_25170_), .B(1'h1), .S(_05523_), .Y(_25171_) );
  \$mux  #( .WIDTH(1) ) _47259_ ( .A(_tmp_1150), .B(1'h0), .S(_05523_), .Y(_25172_) );
  \$mux  #( .WIDTH(1) ) _47260_ ( .A(_25172_), .B(1'h1), .S(_05524_), .Y(_25173_) );
  \$mux  #( .WIDTH(1) ) _47261_ ( .A(_25173_), .B(1'h1), .S(_05525_), .Y(_25174_) );
  \$mux  #( .WIDTH(1) ) _47265_ ( .A(_tmp_1143), .B(1'h0), .S(_05522_), .Y(_25175_) );
  \$mux  #( .WIDTH(1) ) _47266_ ( .A(_25175_), .B(1'h1), .S(_05523_), .Y(_25176_) );
  \$mux  #( .WIDTH(1) ) _47269_ ( .A(_tmp_858), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25177_) );
  \$mux  #( .WIDTH(1) ) _47270_ ( .A(_25177_), .B(1'h1), .S(_05520_), .Y(_25178_) );
  \$mux  #( .WIDTH(34) ) _47272_ ( .A(_tmp_857), .B({ 1'h0, _maxi_read_size }), .S(_05519_), .Y(_25179_) );
  \$mux  #( .WIDTH(34) ) _47273_ ( .A(_25179_), .B(_25964_), .S(_05349_), .Y(_25180_) );
  \$mux  #( .WIDTH(4) ) _47275_ ( .A(_tmp_124), .B(4'h0), .S(_05506_), .Y(_25181_) );
  \$mux  #( .WIDTH(4) ) _47276_ ( .A(_25181_), .B(_22095_[3:0]), .S(_05507_), .Y(_25182_) );
  \$mux  #( .WIDTH(4) ) _47277_ ( .A(_25182_), .B(4'h0), .S(_05508_), .Y(_25183_) );
  \$mux  #( .WIDTH(9) ) _47279_ ( .A(_tmp_105), .B(_25939_[8:0]), .S(_05506_), .Y(_25184_) );
  \$mux  #( .WIDTH(9) ) _47280_ ( .A(_25184_), .B(_tmp_114), .S(_05517_), .Y(_25185_) );
  \$mux  #( .WIDTH(9) ) _47282_ ( .A(_tmp_104), .B(_25939_[8:0]), .S(_05506_), .Y(_25186_) );
  \$mux  #( .WIDTH(9) ) _47283_ ( .A(_25186_), .B(_tmp_113), .S(_05516_), .Y(_25187_) );
  \$mux  #( .WIDTH(9) ) _47285_ ( .A(_tmp_103), .B(_25939_[8:0]), .S(_05506_), .Y(_25188_) );
  \$mux  #( .WIDTH(9) ) _47286_ ( .A(_25188_), .B(_tmp_112), .S(_05515_), .Y(_25189_) );
  \$mux  #( .WIDTH(9) ) _47288_ ( .A(_tmp_102), .B(_25939_[8:0]), .S(_05506_), .Y(_25190_) );
  \$mux  #( .WIDTH(9) ) _47289_ ( .A(_25190_), .B(_tmp_111), .S(_05514_), .Y(_25191_) );
  \$mux  #( .WIDTH(9) ) _47291_ ( .A(_tmp_101), .B(_25939_[8:0]), .S(_05506_), .Y(_25192_) );
  \$mux  #( .WIDTH(9) ) _47292_ ( .A(_25192_), .B(_tmp_110), .S(_05513_), .Y(_25193_) );
  \$mux  #( .WIDTH(9) ) _47294_ ( .A(_tmp_100), .B(_25939_[8:0]), .S(_05506_), .Y(_25194_) );
  \$mux  #( .WIDTH(9) ) _47295_ ( .A(_25194_), .B(_tmp_109), .S(_05512_), .Y(_25195_) );
  \$mux  #( .WIDTH(9) ) _47297_ ( .A(_tmp_99), .B(_25939_[8:0]), .S(_05506_), .Y(_25196_) );
  \$mux  #( .WIDTH(9) ) _47298_ ( .A(_25196_), .B(_tmp_108), .S(_05511_), .Y(_25197_) );
  \$mux  #( .WIDTH(9) ) _47300_ ( .A(_tmp_98), .B(_25939_[8:0]), .S(_05506_), .Y(_25198_) );
  \$mux  #( .WIDTH(9) ) _47301_ ( .A(_25198_), .B(_tmp_107), .S(_05510_), .Y(_25199_) );
  \$mux  #( .WIDTH(9) ) _47303_ ( .A(_tmp_97), .B(_25939_[8:0]), .S(_05506_), .Y(_25200_) );
  \$mux  #( .WIDTH(9) ) _47304_ ( .A(_25200_), .B(_tmp_106), .S(_05509_), .Y(_25201_) );
  \$mux  #( .WIDTH(1) ) _47306_ ( .A(_tmp_96), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25202_) );
  \$mux  #( .WIDTH(1) ) _47307_ ( .A(_25202_), .B(1'h1), .S(_05518_), .Y(_25203_) );
  \$mux  #( .WIDTH(34) ) _47309_ ( .A(_tmp_95), .B({ 1'h0, _maxi_read_size }), .S(_05506_), .Y(_25204_) );
  \$mux  #( .WIDTH(34) ) _47310_ ( .A(_25204_), .B(_25963_), .S(_05301_), .Y(_25205_) );
  \$mux  #( .WIDTH(10) ) _47312_ ( .A(_tmp_94), .B(_25953_[9:0]), .S(_05506_), .Y(_25206_) );
  \$mux  #( .WIDTH(10) ) _47313_ ( .A(_25206_), .B(_25962_[9:0]), .S(_05301_), .Y(_25207_) );
  \$mux  #( .WIDTH(10) ) _47314_ ( .A(_25207_), .B(_25953_[9:0]), .S(_05507_), .Y(_25208_) );
  \$mux  #( .WIDTH(1) ) _47316_ ( .A(ram_w8_l2048_id1_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25209_) );
  \$mux  #( .WIDTH(1) ) _47317_ ( .A(_25209_), .B(_05171_), .S(_05301_), .Y(_25210_) );
  \$mux  #( .WIDTH(1) ) _47318_ ( .A(_25210_), .B(1'h1), .S(_05349_), .Y(_25211_) );
  \$mux  #( .WIDTH(8) ) _47320_ ( .A(ram_w8_l2048_id1_2_1_wdata), .B(_dataflow_slice_data_23), .S(_05301_), .Y(_25212_) );
  \$mux  #( .WIDTH(8) ) _47321_ ( .A(_25212_), .B(_dataflow_slice_data_84), .S(_05349_), .Y(_25213_) );
  \$mux  #( .WIDTH(9) ) _47323_ ( .A(ram_w8_l2048_id1_2_1_addr), .B(_tmp_106), .S(_05301_), .Y(_25214_) );
  \$mux  #( .WIDTH(9) ) _47324_ ( .A(_25214_), .B(_25939_[8:0]), .S(_05519_), .Y(_25215_) );
  \$mux  #( .WIDTH(9) ) _47325_ ( .A(_25215_), .B(_22096_[8:0]), .S(_05349_), .Y(_25216_) );
  \$mux  #( .WIDTH(9) ) _47326_ ( .A(_25216_), .B(_maxi_write_local_addr[8:0]), .S(_05524_), .Y(_25217_) );
  \$mux  #( .WIDTH(9) ) _47327_ ( .A(_25217_), .B(_22097_[8:0]), .S(_05525_), .Y(_25218_) );
  \$mux  #( .WIDTH(1) ) _47329_ ( .A(ram_w8_l2048_id1_2_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id1_2_cond_7_1), .Y(_25219_) );
  \$mux  #( .WIDTH(1) ) _47330_ ( .A(_25219_), .B(1'h1), .S(_05521_), .Y(_25220_) );
  \$mux  #( .WIDTH(8) ) _47332_ ( .A(ram_w8_l2048_id1_2_0_wdata), .B(_stream_matmul_15_sink_21_sink_wdata), .S(_05521_), .Y(_25221_) );
  \$mux  #( .WIDTH(9) ) _47334_ ( .A(ram_w8_l2048_id1_2_0_addr), .B(_stream_conv2d_8_source_28_source_ram_raddr[10:2]), .S(_tmp_457), .Y(_25222_) );
  \$mux  #( .WIDTH(9) ) _47335_ ( .A(_25222_), .B(_stream_max_pool_serial_9_source_1_source_ram_raddr[10:2]), .S(_tmp_873), .Y(_25223_) );
  \$mux  #( .WIDTH(9) ) _47336_ ( .A(_25223_), .B(_stream_matmul_15_sink_21_sink_waddr[10:2]), .S(_05521_), .Y(_25224_) );
  \$mux  #( .WIDTH(34) ) _47338_ ( .A(_tmp_1142), .B(_25945_), .S(_05503_), .Y(_25225_) );
  \$mux  #( .WIDTH(34) ) _47339_ ( .A(_25225_), .B(_25961_), .S(_05504_), .Y(_25226_) );
  \$mux  #( .WIDTH(1) ) _47341_ ( .A(_tmp_1141), .B(1'h0), .S(_05501_), .Y(_25227_) );
  \$mux  #( .WIDTH(1) ) _47342_ ( .A(_25227_), .B(_tmp_1140), .S(_05502_), .Y(_25228_) );
  \$mux  #( .WIDTH(1) ) _47344_ ( .A(_tmp_1140), .B(1'h0), .S(_05502_), .Y(_25229_) );
  \$mux  #( .WIDTH(1) ) _47345_ ( .A(_25229_), .B(_05151_), .S(_05503_), .Y(_25230_) );
  \$mux  #( .WIDTH(1) ) _47346_ ( .A(_25230_), .B(1'h0), .S(_05504_), .Y(_25231_) );
  \$mux  #( .WIDTH(1) ) _47347_ ( .A(_25231_), .B(1'h1), .S(_05505_), .Y(_25232_) );
  \$mux  #( .WIDTH(1) ) _47349_ ( .A(_tmp_1139), .B(1'h0), .S(_05501_), .Y(_25233_) );
  \$mux  #( .WIDTH(1) ) _47350_ ( .A(_25233_), .B(1'h1), .S(_05502_), .Y(_25234_) );
  \$mux  #( .WIDTH(1) ) _47352_ ( .A(_tmp_1138), .B(1'h0), .S(_05502_), .Y(_25235_) );
  \$mux  #( .WIDTH(1) ) _47353_ ( .A(_25235_), .B(1'h1), .S(_05503_), .Y(_25236_) );
  \$mux  #( .WIDTH(1) ) _47354_ ( .A(_25236_), .B(1'h1), .S(_05504_), .Y(_25237_) );
  \$mux  #( .WIDTH(1) ) _47358_ ( .A(_tmp_1131), .B(1'h0), .S(_05501_), .Y(_25238_) );
  \$mux  #( .WIDTH(1) ) _47359_ ( .A(_25238_), .B(1'h1), .S(_05502_), .Y(_25239_) );
  \$mux  #( .WIDTH(1) ) _47362_ ( .A(_tmp_856), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25240_) );
  \$mux  #( .WIDTH(1) ) _47363_ ( .A(_25240_), .B(1'h1), .S(_05499_), .Y(_25241_) );
  \$mux  #( .WIDTH(34) ) _47365_ ( .A(_tmp_855), .B({ 1'h0, _maxi_read_size }), .S(_05498_), .Y(_25242_) );
  \$mux  #( .WIDTH(34) ) _47366_ ( .A(_25242_), .B(_25960_), .S(_05346_), .Y(_25243_) );
  \$mux  #( .WIDTH(4) ) _47368_ ( .A(_tmp_93), .B(4'h0), .S(_05485_), .Y(_25244_) );
  \$mux  #( .WIDTH(4) ) _47369_ ( .A(_25244_), .B(_22092_[3:0]), .S(_05486_), .Y(_25245_) );
  \$mux  #( .WIDTH(4) ) _47370_ ( .A(_25245_), .B(4'h0), .S(_05487_), .Y(_25246_) );
  \$mux  #( .WIDTH(9) ) _47372_ ( .A(_tmp_74), .B(_25939_[8:0]), .S(_05485_), .Y(_25247_) );
  \$mux  #( .WIDTH(9) ) _47373_ ( .A(_25247_), .B(_tmp_83), .S(_05496_), .Y(_25248_) );
  \$mux  #( .WIDTH(9) ) _47375_ ( .A(_tmp_73), .B(_25939_[8:0]), .S(_05485_), .Y(_25249_) );
  \$mux  #( .WIDTH(9) ) _47376_ ( .A(_25249_), .B(_tmp_82), .S(_05495_), .Y(_25250_) );
  \$mux  #( .WIDTH(9) ) _47378_ ( .A(_tmp_72), .B(_25939_[8:0]), .S(_05485_), .Y(_25251_) );
  \$mux  #( .WIDTH(9) ) _47379_ ( .A(_25251_), .B(_tmp_81), .S(_05494_), .Y(_25252_) );
  \$mux  #( .WIDTH(9) ) _47381_ ( .A(_tmp_71), .B(_25939_[8:0]), .S(_05485_), .Y(_25253_) );
  \$mux  #( .WIDTH(9) ) _47382_ ( .A(_25253_), .B(_tmp_80), .S(_05493_), .Y(_25254_) );
  \$mux  #( .WIDTH(9) ) _47384_ ( .A(_tmp_70), .B(_25939_[8:0]), .S(_05485_), .Y(_25255_) );
  \$mux  #( .WIDTH(9) ) _47385_ ( .A(_25255_), .B(_tmp_79), .S(_05492_), .Y(_25256_) );
  \$mux  #( .WIDTH(9) ) _47387_ ( .A(_tmp_69), .B(_25939_[8:0]), .S(_05485_), .Y(_25257_) );
  \$mux  #( .WIDTH(9) ) _47388_ ( .A(_25257_), .B(_tmp_78), .S(_05491_), .Y(_25258_) );
  \$mux  #( .WIDTH(9) ) _47390_ ( .A(_tmp_68), .B(_25939_[8:0]), .S(_05485_), .Y(_25259_) );
  \$mux  #( .WIDTH(9) ) _47391_ ( .A(_25259_), .B(_tmp_77), .S(_05490_), .Y(_25260_) );
  \$mux  #( .WIDTH(9) ) _47393_ ( .A(_tmp_67), .B(_25939_[8:0]), .S(_05485_), .Y(_25261_) );
  \$mux  #( .WIDTH(9) ) _47394_ ( .A(_25261_), .B(_tmp_76), .S(_05489_), .Y(_25262_) );
  \$mux  #( .WIDTH(9) ) _47396_ ( .A(_tmp_66), .B(_25939_[8:0]), .S(_05485_), .Y(_25263_) );
  \$mux  #( .WIDTH(9) ) _47397_ ( .A(_25263_), .B(_tmp_75), .S(_05488_), .Y(_25264_) );
  \$mux  #( .WIDTH(1) ) _47399_ ( .A(_tmp_65), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25265_) );
  \$mux  #( .WIDTH(1) ) _47400_ ( .A(_25265_), .B(1'h1), .S(_05497_), .Y(_25266_) );
  \$mux  #( .WIDTH(34) ) _47402_ ( .A(_tmp_64), .B({ 1'h0, _maxi_read_size }), .S(_05485_), .Y(_25267_) );
  \$mux  #( .WIDTH(34) ) _47403_ ( .A(_25267_), .B(_25959_), .S(_05298_), .Y(_25268_) );
  \$mux  #( .WIDTH(10) ) _47405_ ( .A(_tmp_63), .B(_25953_[9:0]), .S(_05485_), .Y(_25269_) );
  \$mux  #( .WIDTH(10) ) _47406_ ( .A(_25269_), .B(_25958_[9:0]), .S(_05298_), .Y(_25270_) );
  \$mux  #( .WIDTH(10) ) _47407_ ( .A(_25270_), .B(_25953_[9:0]), .S(_05486_), .Y(_25271_) );
  \$mux  #( .WIDTH(1) ) _47409_ ( .A(ram_w8_l2048_id1_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25272_) );
  \$mux  #( .WIDTH(1) ) _47410_ ( .A(_25272_), .B(_05162_), .S(_05298_), .Y(_25273_) );
  \$mux  #( .WIDTH(1) ) _47411_ ( .A(_25273_), .B(1'h1), .S(_05346_), .Y(_25274_) );
  \$mux  #( .WIDTH(8) ) _47413_ ( .A(ram_w8_l2048_id1_1_1_wdata), .B(_dataflow_slice_data_20), .S(_05298_), .Y(_25275_) );
  \$mux  #( .WIDTH(8) ) _47414_ ( .A(_25275_), .B(_dataflow_slice_data_81), .S(_05346_), .Y(_25276_) );
  \$mux  #( .WIDTH(9) ) _47416_ ( .A(ram_w8_l2048_id1_1_1_addr), .B(_tmp_75), .S(_05298_), .Y(_25277_) );
  \$mux  #( .WIDTH(9) ) _47417_ ( .A(_25277_), .B(_25939_[8:0]), .S(_05498_), .Y(_25278_) );
  \$mux  #( .WIDTH(9) ) _47418_ ( .A(_25278_), .B(_22093_[8:0]), .S(_05346_), .Y(_25279_) );
  \$mux  #( .WIDTH(9) ) _47419_ ( .A(_25279_), .B(_maxi_write_local_addr[8:0]), .S(_05503_), .Y(_25280_) );
  \$mux  #( .WIDTH(9) ) _47420_ ( .A(_25280_), .B(_22094_[8:0]), .S(_05504_), .Y(_25281_) );
  \$mux  #( .WIDTH(1) ) _47422_ ( .A(ram_w8_l2048_id1_1_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id1_1_cond_7_1), .Y(_25282_) );
  \$mux  #( .WIDTH(1) ) _47423_ ( .A(_25282_), .B(1'h1), .S(_05500_), .Y(_25283_) );
  \$mux  #( .WIDTH(8) ) _47425_ ( .A(ram_w8_l2048_id1_1_0_wdata), .B(_stream_matmul_15_sink_21_sink_wdata), .S(_05500_), .Y(_25284_) );
  \$mux  #( .WIDTH(9) ) _47427_ ( .A(ram_w8_l2048_id1_1_0_addr), .B(_stream_conv2d_8_source_28_source_ram_raddr[10:2]), .S(_tmp_457), .Y(_25285_) );
  \$mux  #( .WIDTH(9) ) _47428_ ( .A(_25285_), .B(_stream_max_pool_serial_9_source_1_source_ram_raddr[10:2]), .S(_tmp_873), .Y(_25286_) );
  \$mux  #( .WIDTH(9) ) _47429_ ( .A(_25286_), .B(_stream_matmul_15_sink_21_sink_waddr[10:2]), .S(_05500_), .Y(_25287_) );
  \$mux  #( .WIDTH(1) ) _47431_ ( .A(_dataflow_cat_valid_131), .B(1'h0), .S(_05279_), .Y(_25288_) );
  \$mux  #( .WIDTH(1) ) _47432_ ( .A(_25288_), .B(_05483_), .S(_05484_), .Y(_25289_) );
  \$mux  #( .WIDTH(32) ) _47434_ ( .A(_dataflow_cat_data_131), .B({ _tmp_1161, _tmp_1149, _tmp_1137, _tmp_1125 }), .S(_05484_), .Y(_25290_) );
  \$mux  #( .WIDTH(34) ) _47436_ ( .A(_tmp_1130), .B(_25945_), .S(_05480_), .Y(_25291_) );
  \$mux  #( .WIDTH(34) ) _47437_ ( .A(_25291_), .B(_25957_), .S(_05481_), .Y(_25292_) );
  \$mux  #( .WIDTH(1) ) _47439_ ( .A(_tmp_1129), .B(1'h0), .S(_05477_), .Y(_25293_) );
  \$mux  #( .WIDTH(1) ) _47440_ ( .A(_25293_), .B(_tmp_1128), .S(_05478_), .Y(_25294_) );
  \$mux  #( .WIDTH(1) ) _47442_ ( .A(_tmp_1128), .B(1'h0), .S(_05478_), .Y(_25295_) );
  \$mux  #( .WIDTH(1) ) _47443_ ( .A(_25295_), .B(_05151_), .S(_05480_), .Y(_25296_) );
  \$mux  #( .WIDTH(1) ) _47444_ ( .A(_25296_), .B(1'h0), .S(_05481_), .Y(_25297_) );
  \$mux  #( .WIDTH(1) ) _47445_ ( .A(_25297_), .B(1'h1), .S(_05482_), .Y(_25298_) );
  \$mux  #( .WIDTH(1) ) _47447_ ( .A(_tmp_1127), .B(1'h0), .S(_05477_), .Y(_25299_) );
  \$mux  #( .WIDTH(1) ) _47448_ ( .A(_25299_), .B(1'h1), .S(_05478_), .Y(_25300_) );
  \$mux  #( .WIDTH(1) ) _47450_ ( .A(_tmp_1126), .B(1'h0), .S(_05478_), .Y(_25301_) );
  \$mux  #( .WIDTH(1) ) _47451_ ( .A(_25301_), .B(1'h1), .S(_05480_), .Y(_25302_) );
  \$mux  #( .WIDTH(1) ) _47452_ ( .A(_25302_), .B(1'h1), .S(_05481_), .Y(_25303_) );
  \$mux  #( .WIDTH(1) ) _47456_ ( .A(_tmp_1119), .B(1'h0), .S(_05477_), .Y(_25304_) );
  \$mux  #( .WIDTH(1) ) _47457_ ( .A(_25304_), .B(1'h1), .S(_05478_), .Y(_25305_) );
  \$mux  #( .WIDTH(1) ) _47461_ ( .A(_tmp_854), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25306_) );
  \$mux  #( .WIDTH(1) ) _47462_ ( .A(_25306_), .B(1'h1), .S(_05475_), .Y(_25307_) );
  \$mux  #( .WIDTH(34) ) _47464_ ( .A(_tmp_853), .B({ 1'h0, _maxi_read_size }), .S(_05474_), .Y(_25308_) );
  \$mux  #( .WIDTH(34) ) _47465_ ( .A(_25308_), .B(_25956_), .S(_05343_), .Y(_25309_) );
  \$mux  #( .WIDTH(4) ) _47468_ ( .A(_tmp_62), .B(4'h0), .S(_05460_), .Y(_25310_) );
  \$mux  #( .WIDTH(4) ) _47469_ ( .A(_25310_), .B(_22089_[3:0]), .S(_05461_), .Y(_25311_) );
  \$mux  #( .WIDTH(4) ) _47470_ ( .A(_25311_), .B(4'h0), .S(_05462_), .Y(_25312_) );
  \$mux  #( .WIDTH(9) ) _47472_ ( .A(_tmp_43), .B(_25939_[8:0]), .S(_05460_), .Y(_25313_) );
  \$mux  #( .WIDTH(9) ) _47473_ ( .A(_25313_), .B(_tmp_52), .S(_05471_), .Y(_25314_) );
  \$mux  #( .WIDTH(9) ) _47475_ ( .A(_tmp_42), .B(_25939_[8:0]), .S(_05460_), .Y(_25315_) );
  \$mux  #( .WIDTH(9) ) _47476_ ( .A(_25315_), .B(_tmp_51), .S(_05470_), .Y(_25316_) );
  \$mux  #( .WIDTH(9) ) _47478_ ( .A(_tmp_41), .B(_25939_[8:0]), .S(_05460_), .Y(_25317_) );
  \$mux  #( .WIDTH(9) ) _47479_ ( .A(_25317_), .B(_tmp_50), .S(_05469_), .Y(_25318_) );
  \$mux  #( .WIDTH(9) ) _47481_ ( .A(_tmp_40), .B(_25939_[8:0]), .S(_05460_), .Y(_25319_) );
  \$mux  #( .WIDTH(9) ) _47482_ ( .A(_25319_), .B(_tmp_49), .S(_05468_), .Y(_25320_) );
  \$mux  #( .WIDTH(9) ) _47484_ ( .A(_tmp_39), .B(_25939_[8:0]), .S(_05460_), .Y(_25321_) );
  \$mux  #( .WIDTH(9) ) _47485_ ( .A(_25321_), .B(_tmp_48), .S(_05467_), .Y(_25322_) );
  \$mux  #( .WIDTH(9) ) _47487_ ( .A(_tmp_38), .B(_25939_[8:0]), .S(_05460_), .Y(_25323_) );
  \$mux  #( .WIDTH(9) ) _47488_ ( .A(_25323_), .B(_tmp_47), .S(_05466_), .Y(_25324_) );
  \$mux  #( .WIDTH(9) ) _47490_ ( .A(_tmp_37), .B(_25939_[8:0]), .S(_05460_), .Y(_25325_) );
  \$mux  #( .WIDTH(9) ) _47491_ ( .A(_25325_), .B(_tmp_46), .S(_05465_), .Y(_25326_) );
  \$mux  #( .WIDTH(9) ) _47493_ ( .A(_tmp_36), .B(_25939_[8:0]), .S(_05460_), .Y(_25327_) );
  \$mux  #( .WIDTH(9) ) _47494_ ( .A(_25327_), .B(_tmp_45), .S(_05464_), .Y(_25328_) );
  \$mux  #( .WIDTH(9) ) _47496_ ( .A(_tmp_35), .B(_25939_[8:0]), .S(_05460_), .Y(_25329_) );
  \$mux  #( .WIDTH(9) ) _47497_ ( .A(_25329_), .B(_tmp_44), .S(_05463_), .Y(_25330_) );
  \$mux  #( .WIDTH(1) ) _47499_ ( .A(_tmp_34), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25331_) );
  \$mux  #( .WIDTH(1) ) _47500_ ( .A(_25331_), .B(1'h1), .S(_05472_), .Y(_25332_) );
  \$mux  #( .WIDTH(34) ) _47502_ ( .A(_tmp_33), .B({ 1'h0, _maxi_read_size }), .S(_05460_), .Y(_25333_) );
  \$mux  #( .WIDTH(34) ) _47503_ ( .A(_25333_), .B(_25955_), .S(_05295_), .Y(_25334_) );
  \$mux  #( .WIDTH(10) ) _47505_ ( .A(_tmp_32), .B(_25953_[9:0]), .S(_05460_), .Y(_25335_) );
  \$mux  #( .WIDTH(10) ) _47506_ ( .A(_25335_), .B(_25954_[9:0]), .S(_05295_), .Y(_25336_) );
  \$mux  #( .WIDTH(10) ) _47507_ ( .A(_25336_), .B(_25953_[9:0]), .S(_05461_), .Y(_25337_) );
  \$mux  #( .WIDTH(1) ) _47509_ ( .A(ram_w8_l2048_id1_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25338_) );
  \$mux  #( .WIDTH(1) ) _47510_ ( .A(_25338_), .B(_05153_), .S(_05295_), .Y(_25339_) );
  \$mux  #( .WIDTH(1) ) _47511_ ( .A(_25339_), .B(1'h1), .S(_05343_), .Y(_25340_) );
  \$mux  #( .WIDTH(8) ) _47513_ ( .A(ram_w8_l2048_id1_0_1_wdata), .B(_dataflow_slice_data_17), .S(_05295_), .Y(_25341_) );
  \$mux  #( .WIDTH(8) ) _47514_ ( .A(_25341_), .B(_dataflow_slice_data_78), .S(_05343_), .Y(_25342_) );
  \$mux  #( .WIDTH(9) ) _47516_ ( .A(ram_w8_l2048_id1_0_1_addr), .B(_tmp_44), .S(_05295_), .Y(_25343_) );
  \$mux  #( .WIDTH(9) ) _47517_ ( .A(_25343_), .B(_25939_[8:0]), .S(_05474_), .Y(_25344_) );
  \$mux  #( .WIDTH(9) ) _47518_ ( .A(_25344_), .B(_22090_[8:0]), .S(_05343_), .Y(_25345_) );
  \$mux  #( .WIDTH(9) ) _47519_ ( .A(_25345_), .B(_maxi_write_local_addr[8:0]), .S(_05480_), .Y(_25346_) );
  \$mux  #( .WIDTH(9) ) _47520_ ( .A(_25346_), .B(_22091_[8:0]), .S(_05481_), .Y(_25347_) );
  \$mux  #( .WIDTH(1) ) _47522_ ( .A(ram_w8_l2048_id1_0_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id1_0_cond_7_1), .Y(_25348_) );
  \$mux  #( .WIDTH(1) ) _47523_ ( .A(_25348_), .B(1'h1), .S(_05476_), .Y(_25349_) );
  \$mux  #( .WIDTH(8) ) _47525_ ( .A(ram_w8_l2048_id1_0_0_wdata), .B(_stream_matmul_15_sink_21_sink_wdata), .S(_05476_), .Y(_25350_) );
  \$mux  #( .WIDTH(9) ) _47527_ ( .A(ram_w8_l2048_id1_0_0_addr), .B(_stream_conv2d_8_source_28_source_ram_raddr[10:2]), .S(_tmp_457), .Y(_25351_) );
  \$mux  #( .WIDTH(9) ) _47528_ ( .A(_25351_), .B(_stream_max_pool_serial_9_source_1_source_ram_raddr[10:2]), .S(_tmp_873), .Y(_25352_) );
  \$mux  #( .WIDTH(9) ) _47529_ ( .A(_25352_), .B(_stream_matmul_15_sink_21_sink_waddr[10:2]), .S(_05476_), .Y(_25353_) );
  \$mux  #( .WIDTH(34) ) _47531_ ( .A(_tmp_957), .B(_25945_), .S(_05456_), .Y(_25354_) );
  \$mux  #( .WIDTH(34) ) _47532_ ( .A(_25354_), .B(_25952_), .S(_05457_), .Y(_25355_) );
  \$mux  #( .WIDTH(1) ) _47534_ ( .A(_tmp_956), .B(1'h0), .S(_05454_), .Y(_25356_) );
  \$mux  #( .WIDTH(1) ) _47535_ ( .A(_25356_), .B(_tmp_955), .S(_05455_), .Y(_25357_) );
  \$mux  #( .WIDTH(1) ) _47537_ ( .A(_tmp_955), .B(1'h0), .S(_05455_), .Y(_25358_) );
  \$mux  #( .WIDTH(1) ) _47538_ ( .A(_25358_), .B(_05151_), .S(_05456_), .Y(_25359_) );
  \$mux  #( .WIDTH(1) ) _47539_ ( .A(_25359_), .B(1'h0), .S(_05457_), .Y(_25360_) );
  \$mux  #( .WIDTH(1) ) _47540_ ( .A(_25360_), .B(1'h1), .S(_05458_), .Y(_25361_) );
  \$mux  #( .WIDTH(1) ) _47542_ ( .A(_tmp_954), .B(1'h0), .S(_05454_), .Y(_25362_) );
  \$mux  #( .WIDTH(1) ) _47543_ ( .A(_25362_), .B(1'h1), .S(_05455_), .Y(_25363_) );
  \$mux  #( .WIDTH(1) ) _47545_ ( .A(_tmp_953), .B(1'h0), .S(_05455_), .Y(_25364_) );
  \$mux  #( .WIDTH(1) ) _47546_ ( .A(_25364_), .B(1'h1), .S(_05456_), .Y(_25365_) );
  \$mux  #( .WIDTH(1) ) _47547_ ( .A(_25365_), .B(1'h1), .S(_05457_), .Y(_25366_) );
  \$mux  #( .WIDTH(1) ) _47551_ ( .A(_tmp_946), .B(1'h0), .S(_05454_), .Y(_25367_) );
  \$mux  #( .WIDTH(1) ) _47552_ ( .A(_25367_), .B(1'h1), .S(_05455_), .Y(_25368_) );
  \$mux  #( .WIDTH(1) ) _47555_ ( .A(_tmp_26), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25369_) );
  \$mux  #( .WIDTH(1) ) _47556_ ( .A(_25369_), .B(1'h1), .S(_05452_), .Y(_25370_) );
  \$mux  #( .WIDTH(34) ) _47558_ ( .A(_tmp_25), .B({ 1'h0, _maxi_read_size }), .S(_05451_), .Y(_25371_) );
  \$mux  #( .WIDTH(34) ) _47559_ ( .A(_25371_), .B(_25951_), .S(_05292_), .Y(_25372_) );
  \$mux  #( .WIDTH(1) ) _47561_ ( .A(ram_w8_l2048_id0_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25373_) );
  \$mux  #( .WIDTH(1) ) _47562_ ( .A(_25373_), .B(1'h1), .S(_05292_), .Y(_25374_) );
  \$mux  #( .WIDTH(8) ) _47564_ ( .A(ram_w8_l2048_id0_3_1_wdata), .B(_dataflow_slice_data_13), .S(_05292_), .Y(_25375_) );
  \$mux  #( .WIDTH(9) ) _47566_ ( .A(ram_w8_l2048_id0_3_1_addr), .B(_25939_[8:0]), .S(_05451_), .Y(_25376_) );
  \$mux  #( .WIDTH(9) ) _47567_ ( .A(_25376_), .B(_22087_[8:0]), .S(_05292_), .Y(_25377_) );
  \$mux  #( .WIDTH(9) ) _47568_ ( .A(_25377_), .B(_maxi_write_local_addr[8:0]), .S(_05456_), .Y(_25378_) );
  \$mux  #( .WIDTH(9) ) _47569_ ( .A(_25378_), .B(_22088_[8:0]), .S(_05457_), .Y(_25379_) );
  \$mux  #( .WIDTH(1) ) _47571_ ( .A(ram_w8_l2048_id0_3_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_3_1), .Y(_25380_) );
  \$mux  #( .WIDTH(1) ) _47572_ ( .A(_25380_), .B(1'h1), .S(_05453_), .Y(_25381_) );
  \$mux  #( .WIDTH(8) ) _47574_ ( .A(ram_w8_l2048_id0_3_0_wdata), .B(_stream_max_pool_serial_9_sink_3_sink_wdata), .S(_05453_), .Y(_25382_) );
  \$mux  #( .WIDTH(9) ) _47576_ ( .A(ram_w8_l2048_id0_3_0_addr), .B(_stream_conv2d_8_source_8_source_ram_raddr[10:2]), .S(_tmp_347), .Y(_25383_) );
  \$mux  #( .WIDTH(9) ) _47577_ ( .A(_25383_), .B(_stream_max_pool_serial_9_sink_3_sink_waddr[10:2]), .S(_05453_), .Y(_25384_) );
  \$mux  #( .WIDTH(9) ) _47578_ ( .A(_25384_), .B(_stream_matmul_15_source_8_source_ram_raddr[10:2]), .S(_tmp_1003), .Y(_25385_) );
  \$mux  #( .WIDTH(34) ) _47580_ ( .A(_tmp_945), .B(_25945_), .S(_05448_), .Y(_25386_) );
  \$mux  #( .WIDTH(34) ) _47581_ ( .A(_25386_), .B(_25950_), .S(_05449_), .Y(_25387_) );
  \$mux  #( .WIDTH(1) ) _47583_ ( .A(_tmp_944), .B(1'h0), .S(_05446_), .Y(_25388_) );
  \$mux  #( .WIDTH(1) ) _47584_ ( .A(_25388_), .B(_tmp_943), .S(_05447_), .Y(_25389_) );
  \$mux  #( .WIDTH(1) ) _47586_ ( .A(_tmp_943), .B(1'h0), .S(_05447_), .Y(_25390_) );
  \$mux  #( .WIDTH(1) ) _47587_ ( .A(_25390_), .B(_05151_), .S(_05448_), .Y(_25391_) );
  \$mux  #( .WIDTH(1) ) _47588_ ( .A(_25391_), .B(1'h0), .S(_05449_), .Y(_25392_) );
  \$mux  #( .WIDTH(1) ) _47589_ ( .A(_25392_), .B(1'h1), .S(_05450_), .Y(_25393_) );
  \$mux  #( .WIDTH(1) ) _47591_ ( .A(_tmp_942), .B(1'h0), .S(_05446_), .Y(_25394_) );
  \$mux  #( .WIDTH(1) ) _47592_ ( .A(_25394_), .B(1'h1), .S(_05447_), .Y(_25395_) );
  \$mux  #( .WIDTH(1) ) _47594_ ( .A(_tmp_941), .B(1'h0), .S(_05447_), .Y(_25396_) );
  \$mux  #( .WIDTH(1) ) _47595_ ( .A(_25396_), .B(1'h1), .S(_05448_), .Y(_25397_) );
  \$mux  #( .WIDTH(1) ) _47596_ ( .A(_25397_), .B(1'h1), .S(_05449_), .Y(_25398_) );
  \$mux  #( .WIDTH(1) ) _47600_ ( .A(_tmp_934), .B(1'h0), .S(_05446_), .Y(_25399_) );
  \$mux  #( .WIDTH(1) ) _47601_ ( .A(_25399_), .B(1'h1), .S(_05447_), .Y(_25400_) );
  \$mux  #( .WIDTH(1) ) _47604_ ( .A(_tmp_24), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25401_) );
  \$mux  #( .WIDTH(1) ) _47605_ ( .A(_25401_), .B(1'h1), .S(_05444_), .Y(_25402_) );
  \$mux  #( .WIDTH(34) ) _47607_ ( .A(_tmp_23), .B({ 1'h0, _maxi_read_size }), .S(_05443_), .Y(_25403_) );
  \$mux  #( .WIDTH(34) ) _47608_ ( .A(_25403_), .B(_25949_), .S(_05289_), .Y(_25404_) );
  \$mux  #( .WIDTH(1) ) _47610_ ( .A(ram_w8_l2048_id0_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25405_) );
  \$mux  #( .WIDTH(1) ) _47611_ ( .A(_25405_), .B(1'h1), .S(_05289_), .Y(_25406_) );
  \$mux  #( .WIDTH(8) ) _47613_ ( .A(ram_w8_l2048_id0_2_1_wdata), .B(_dataflow_slice_data_10), .S(_05289_), .Y(_25407_) );
  \$mux  #( .WIDTH(9) ) _47615_ ( .A(ram_w8_l2048_id0_2_1_addr), .B(_25939_[8:0]), .S(_05443_), .Y(_25408_) );
  \$mux  #( .WIDTH(9) ) _47616_ ( .A(_25408_), .B(_22085_[8:0]), .S(_05289_), .Y(_25409_) );
  \$mux  #( .WIDTH(9) ) _47617_ ( .A(_25409_), .B(_maxi_write_local_addr[8:0]), .S(_05448_), .Y(_25410_) );
  \$mux  #( .WIDTH(9) ) _47618_ ( .A(_25410_), .B(_22086_[8:0]), .S(_05449_), .Y(_25411_) );
  \$mux  #( .WIDTH(1) ) _47620_ ( .A(ram_w8_l2048_id0_2_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_2_cond_3_1), .Y(_25412_) );
  \$mux  #( .WIDTH(1) ) _47621_ ( .A(_25412_), .B(1'h1), .S(_05445_), .Y(_25413_) );
  \$mux  #( .WIDTH(8) ) _47623_ ( .A(ram_w8_l2048_id0_2_0_wdata), .B(_stream_max_pool_serial_9_sink_3_sink_wdata), .S(_05445_), .Y(_25414_) );
  \$mux  #( .WIDTH(9) ) _47625_ ( .A(ram_w8_l2048_id0_2_0_addr), .B(_stream_conv2d_8_source_8_source_ram_raddr[10:2]), .S(_tmp_347), .Y(_25415_) );
  \$mux  #( .WIDTH(9) ) _47626_ ( .A(_25415_), .B(_stream_max_pool_serial_9_sink_3_sink_waddr[10:2]), .S(_05445_), .Y(_25416_) );
  \$mux  #( .WIDTH(9) ) _47627_ ( .A(_25416_), .B(_stream_matmul_15_source_8_source_ram_raddr[10:2]), .S(_tmp_1003), .Y(_25417_) );
  \$mux  #( .WIDTH(34) ) _47629_ ( .A(_tmp_933), .B(_25945_), .S(_05440_), .Y(_25418_) );
  \$mux  #( .WIDTH(34) ) _47630_ ( .A(_25418_), .B(_25948_), .S(_05441_), .Y(_25419_) );
  \$mux  #( .WIDTH(1) ) _47632_ ( .A(_tmp_932), .B(1'h0), .S(_05438_), .Y(_25420_) );
  \$mux  #( .WIDTH(1) ) _47633_ ( .A(_25420_), .B(_tmp_931), .S(_05439_), .Y(_25421_) );
  \$mux  #( .WIDTH(1) ) _47635_ ( .A(_tmp_931), .B(1'h0), .S(_05439_), .Y(_25422_) );
  \$mux  #( .WIDTH(1) ) _47636_ ( .A(_25422_), .B(_05151_), .S(_05440_), .Y(_25423_) );
  \$mux  #( .WIDTH(1) ) _47637_ ( .A(_25423_), .B(1'h0), .S(_05441_), .Y(_25424_) );
  \$mux  #( .WIDTH(1) ) _47638_ ( .A(_25424_), .B(1'h1), .S(_05442_), .Y(_25425_) );
  \$mux  #( .WIDTH(1) ) _47640_ ( .A(_tmp_930), .B(1'h0), .S(_05438_), .Y(_25426_) );
  \$mux  #( .WIDTH(1) ) _47641_ ( .A(_25426_), .B(1'h1), .S(_05439_), .Y(_25427_) );
  \$mux  #( .WIDTH(1) ) _47643_ ( .A(_tmp_929), .B(1'h0), .S(_05439_), .Y(_25428_) );
  \$mux  #( .WIDTH(1) ) _47644_ ( .A(_25428_), .B(1'h1), .S(_05440_), .Y(_25429_) );
  \$mux  #( .WIDTH(1) ) _47645_ ( .A(_25429_), .B(1'h1), .S(_05441_), .Y(_25430_) );
  \$mux  #( .WIDTH(1) ) _47649_ ( .A(_tmp_922), .B(1'h0), .S(_05438_), .Y(_25431_) );
  \$mux  #( .WIDTH(1) ) _47650_ ( .A(_25431_), .B(1'h1), .S(_05439_), .Y(_25432_) );
  \$mux  #( .WIDTH(1) ) _47653_ ( .A(_tmp_22), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25433_) );
  \$mux  #( .WIDTH(1) ) _47654_ ( .A(_25433_), .B(1'h1), .S(_05436_), .Y(_25434_) );
  \$mux  #( .WIDTH(34) ) _47656_ ( .A(_tmp_21), .B({ 1'h0, _maxi_read_size }), .S(_05435_), .Y(_25435_) );
  \$mux  #( .WIDTH(34) ) _47657_ ( .A(_25435_), .B(_25947_), .S(_05286_), .Y(_25436_) );
  \$mux  #( .WIDTH(1) ) _47659_ ( .A(ram_w8_l2048_id0_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25437_) );
  \$mux  #( .WIDTH(1) ) _47660_ ( .A(_25437_), .B(1'h1), .S(_05286_), .Y(_25438_) );
  \$mux  #( .WIDTH(8) ) _47662_ ( .A(ram_w8_l2048_id0_1_1_wdata), .B(_dataflow_slice_data_7), .S(_05286_), .Y(_25439_) );
  \$mux  #( .WIDTH(9) ) _47664_ ( .A(ram_w8_l2048_id0_1_1_addr), .B(_25939_[8:0]), .S(_05435_), .Y(_25440_) );
  \$mux  #( .WIDTH(9) ) _47665_ ( .A(_25440_), .B(_22083_[8:0]), .S(_05286_), .Y(_25441_) );
  \$mux  #( .WIDTH(9) ) _47666_ ( .A(_25441_), .B(_maxi_write_local_addr[8:0]), .S(_05440_), .Y(_25442_) );
  \$mux  #( .WIDTH(9) ) _47667_ ( .A(_25442_), .B(_22084_[8:0]), .S(_05441_), .Y(_25443_) );
  \$mux  #( .WIDTH(1) ) _47669_ ( .A(ram_w8_l2048_id0_1_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_1_cond_3_1), .Y(_25444_) );
  \$mux  #( .WIDTH(1) ) _47670_ ( .A(_25444_), .B(1'h1), .S(_05437_), .Y(_25445_) );
  \$mux  #( .WIDTH(8) ) _47672_ ( .A(ram_w8_l2048_id0_1_0_wdata), .B(_stream_max_pool_serial_9_sink_3_sink_wdata), .S(_05437_), .Y(_25446_) );
  \$mux  #( .WIDTH(9) ) _47674_ ( .A(ram_w8_l2048_id0_1_0_addr), .B(_stream_conv2d_8_source_8_source_ram_raddr[10:2]), .S(_tmp_347), .Y(_25447_) );
  \$mux  #( .WIDTH(9) ) _47675_ ( .A(_25447_), .B(_stream_max_pool_serial_9_sink_3_sink_waddr[10:2]), .S(_05437_), .Y(_25448_) );
  \$mux  #( .WIDTH(9) ) _47676_ ( .A(_25448_), .B(_stream_matmul_15_source_8_source_ram_raddr[10:2]), .S(_tmp_1003), .Y(_25449_) );
  \$mux  #( .WIDTH(1) ) _47678_ ( .A(_dataflow_cat_valid_96), .B(1'h0), .S(_05277_), .Y(_25450_) );
  \$mux  #( .WIDTH(1) ) _47679_ ( .A(_25450_), .B(_05433_), .S(_05434_), .Y(_25451_) );
  \$mux  #( .WIDTH(32) ) _47681_ ( .A(_dataflow_cat_data_96), .B({ _tmp_952, _tmp_940, _tmp_928, _tmp_916 }), .S(_05434_), .Y(_25452_) );
  \$mux  #( .WIDTH(34) ) _47684_ ( .A(_tmp_921), .B(_25945_), .S(_05430_), .Y(_25453_) );
  \$mux  #( .WIDTH(34) ) _47685_ ( .A(_25453_), .B(_25946_), .S(_05431_), .Y(_25454_) );
  \$mux  #( .WIDTH(1) ) _47687_ ( .A(_tmp_920), .B(1'h0), .S(_05427_), .Y(_25455_) );
  \$mux  #( .WIDTH(1) ) _47688_ ( .A(_25455_), .B(_tmp_919), .S(_05428_), .Y(_25456_) );
  \$mux  #( .WIDTH(1) ) _47690_ ( .A(_tmp_919), .B(1'h0), .S(_05428_), .Y(_25457_) );
  \$mux  #( .WIDTH(1) ) _47691_ ( .A(_25457_), .B(_05151_), .S(_05430_), .Y(_25458_) );
  \$mux  #( .WIDTH(1) ) _47692_ ( .A(_25458_), .B(1'h0), .S(_05431_), .Y(_25459_) );
  \$mux  #( .WIDTH(1) ) _47693_ ( .A(_25459_), .B(1'h1), .S(_05432_), .Y(_25460_) );
  \$mux  #( .WIDTH(1) ) _47695_ ( .A(_tmp_918), .B(1'h0), .S(_05427_), .Y(_25461_) );
  \$mux  #( .WIDTH(1) ) _47696_ ( .A(_25461_), .B(1'h1), .S(_05428_), .Y(_25462_) );
  \$mux  #( .WIDTH(1) ) _47698_ ( .A(_tmp_917), .B(1'h0), .S(_05428_), .Y(_25463_) );
  \$mux  #( .WIDTH(1) ) _47699_ ( .A(_25463_), .B(1'h1), .S(_05430_), .Y(_25464_) );
  \$mux  #( .WIDTH(1) ) _47700_ ( .A(_25464_), .B(1'h1), .S(_05431_), .Y(_25465_) );
  \$mux  #( .WIDTH(1) ) _47704_ ( .A(_tmp_910), .B(1'h0), .S(_05427_), .Y(_25466_) );
  \$mux  #( .WIDTH(1) ) _47705_ ( .A(_25466_), .B(1'h1), .S(_05428_), .Y(_25467_) );
  \$mux  #( .WIDTH(1) ) _47709_ ( .A(_tmp_20), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25468_) );
  \$mux  #( .WIDTH(1) ) _47710_ ( .A(_25468_), .B(1'h1), .S(_05425_), .Y(_25469_) );
  \$mux  #( .WIDTH(34) ) _47712_ ( .A(_tmp_19), .B({ 1'h0, _maxi_read_size }), .S(_05424_), .Y(_25470_) );
  \$mux  #( .WIDTH(34) ) _47713_ ( .A(_25470_), .B(_25944_), .S(_05283_), .Y(_25471_) );
  \$mux  #( .WIDTH(1) ) _47715_ ( .A(ram_w8_l2048_id0_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25472_) );
  \$mux  #( .WIDTH(1) ) _47716_ ( .A(_25472_), .B(1'h1), .S(_05283_), .Y(_25473_) );
  \$mux  #( .WIDTH(8) ) _47718_ ( .A(ram_w8_l2048_id0_0_1_wdata), .B(_dataflow_slice_data_4), .S(_05283_), .Y(_25474_) );
  \$mux  #( .WIDTH(9) ) _47720_ ( .A(ram_w8_l2048_id0_0_1_addr), .B(_25939_[8:0]), .S(_05424_), .Y(_25475_) );
  \$mux  #( .WIDTH(9) ) _47721_ ( .A(_25475_), .B(_22081_[8:0]), .S(_05283_), .Y(_25476_) );
  \$mux  #( .WIDTH(9) ) _47722_ ( .A(_25476_), .B(_maxi_write_local_addr[8:0]), .S(_05430_), .Y(_25477_) );
  \$mux  #( .WIDTH(9) ) _47723_ ( .A(_25477_), .B(_22082_[8:0]), .S(_05431_), .Y(_25478_) );
  \$mux  #( .WIDTH(1) ) _47725_ ( .A(ram_w8_l2048_id0_0_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_0_cond_3_1), .Y(_25479_) );
  \$mux  #( .WIDTH(1) ) _47726_ ( .A(_25479_), .B(1'h1), .S(_05426_), .Y(_25480_) );
  \$mux  #( .WIDTH(8) ) _47728_ ( .A(ram_w8_l2048_id0_0_0_wdata), .B(_stream_max_pool_serial_9_sink_3_sink_wdata), .S(_05426_), .Y(_25481_) );
  \$mux  #( .WIDTH(9) ) _47730_ ( .A(ram_w8_l2048_id0_0_0_addr), .B(_stream_conv2d_8_source_8_source_ram_raddr[10:2]), .S(_tmp_347), .Y(_25482_) );
  \$mux  #( .WIDTH(9) ) _47731_ ( .A(_25482_), .B(_stream_max_pool_serial_9_sink_3_sink_waddr[10:2]), .S(_05426_), .Y(_25483_) );
  \$mux  #( .WIDTH(9) ) _47732_ ( .A(_25483_), .B(_stream_matmul_15_source_8_source_ram_raddr[10:2]), .S(_tmp_1003), .Y(_25484_) );
  \$mux  #( .WIDTH(1) ) _47734_ ( .A(_tmp_971), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25485_) );
  \$mux  #( .WIDTH(1) ) _47735_ ( .A(_25485_), .B(1'h1), .S(_05422_), .Y(_25486_) );
  \$mux  #( .WIDTH(34) ) _47737_ ( .A(_tmp_970), .B({ 1'h0, _maxi_read_size }), .S(_05421_), .Y(_25487_) );
  \$mux  #( .WIDTH(34) ) _47738_ ( .A(_25487_), .B(_25943_), .S(_05364_), .Y(_25488_) );
  \$mux  #( .WIDTH(1) ) _47740_ ( .A(ram_w8_l4096_id0_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25489_) );
  \$mux  #( .WIDTH(1) ) _47741_ ( .A(_25489_), .B(1'h1), .S(_05364_), .Y(_25490_) );
  \$mux  #( .WIDTH(8) ) _47743_ ( .A(ram_w8_l4096_id0_3_1_wdata), .B(_dataflow_slice_data_109), .S(_05364_), .Y(_25491_) );
  \$mux  #( .WIDTH(10) ) _47745_ ( .A(ram_w8_l4096_id0_3_1_addr), .B(_25939_[9:0]), .S(_05421_), .Y(_25492_) );
  \$mux  #( .WIDTH(10) ) _47746_ ( .A(_25492_), .B(_22080_[9:0]), .S(_05364_), .Y(_25493_) );
  \$mux  #( .WIDTH(10) ) _47748_ ( .A(ram_w8_l4096_id0_3_0_addr), .B(_stream_matmul_15_source_20_source_ram_raddr[11:2]), .S(_tmp_1033), .Y(_25494_) );
  \$mux  #( .WIDTH(1) ) _47750_ ( .A(_tmp_969), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25495_) );
  \$mux  #( .WIDTH(1) ) _47751_ ( .A(_25495_), .B(1'h1), .S(_05420_), .Y(_25496_) );
  \$mux  #( .WIDTH(34) ) _47753_ ( .A(_tmp_968), .B({ 1'h0, _maxi_read_size }), .S(_05419_), .Y(_25497_) );
  \$mux  #( .WIDTH(34) ) _47754_ ( .A(_25497_), .B(_25942_), .S(_05361_), .Y(_25498_) );
  \$mux  #( .WIDTH(1) ) _47756_ ( .A(ram_w8_l4096_id0_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25499_) );
  \$mux  #( .WIDTH(1) ) _47757_ ( .A(_25499_), .B(1'h1), .S(_05361_), .Y(_25500_) );
  \$mux  #( .WIDTH(8) ) _47759_ ( .A(ram_w8_l4096_id0_2_1_wdata), .B(_dataflow_slice_data_106), .S(_05361_), .Y(_25501_) );
  \$mux  #( .WIDTH(10) ) _47761_ ( .A(ram_w8_l4096_id0_2_1_addr), .B(_25939_[9:0]), .S(_05419_), .Y(_25502_) );
  \$mux  #( .WIDTH(10) ) _47762_ ( .A(_25502_), .B(_22079_[9:0]), .S(_05361_), .Y(_25503_) );
  \$mux  #( .WIDTH(10) ) _47764_ ( .A(ram_w8_l4096_id0_2_0_addr), .B(_stream_matmul_15_source_20_source_ram_raddr[11:2]), .S(_tmp_1033), .Y(_25504_) );
  \$mux  #( .WIDTH(1) ) _47766_ ( .A(_tmp_967), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25505_) );
  \$mux  #( .WIDTH(1) ) _47767_ ( .A(_25505_), .B(1'h1), .S(_05418_), .Y(_25506_) );
  \$mux  #( .WIDTH(34) ) _47769_ ( .A(_tmp_966), .B({ 1'h0, _maxi_read_size }), .S(_05417_), .Y(_25507_) );
  \$mux  #( .WIDTH(34) ) _47770_ ( .A(_25507_), .B(_25941_), .S(_05358_), .Y(_25508_) );
  \$mux  #( .WIDTH(1) ) _47772_ ( .A(ram_w8_l4096_id0_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25509_) );
  \$mux  #( .WIDTH(1) ) _47773_ ( .A(_25509_), .B(1'h1), .S(_05358_), .Y(_25510_) );
  \$mux  #( .WIDTH(8) ) _47775_ ( .A(ram_w8_l4096_id0_1_1_wdata), .B(_dataflow_slice_data_103), .S(_05358_), .Y(_25511_) );
  \$mux  #( .WIDTH(10) ) _47777_ ( .A(ram_w8_l4096_id0_1_1_addr), .B(_25939_[9:0]), .S(_05417_), .Y(_25512_) );
  \$mux  #( .WIDTH(10) ) _47778_ ( .A(_25512_), .B(_22078_[9:0]), .S(_05358_), .Y(_25513_) );
  \$mux  #( .WIDTH(10) ) _47780_ ( .A(ram_w8_l4096_id0_1_0_addr), .B(_stream_matmul_15_source_20_source_ram_raddr[11:2]), .S(_tmp_1033), .Y(_25514_) );
  \$mux  #( .WIDTH(1) ) _47784_ ( .A(_tmp_965), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25515_) );
  \$mux  #( .WIDTH(1) ) _47785_ ( .A(_25515_), .B(1'h1), .S(_05416_), .Y(_25516_) );
  \$mux  #( .WIDTH(34) ) _47787_ ( .A(_tmp_964), .B({ 1'h0, _maxi_read_size }), .S(_05415_), .Y(_25517_) );
  \$mux  #( .WIDTH(34) ) _47788_ ( .A(_25517_), .B(_25940_), .S(_05355_), .Y(_25518_) );
  \$mux  #( .WIDTH(1) ) _47790_ ( .A(ram_w8_l4096_id0_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id9_2_cond_0_1), .Y(_25519_) );
  \$mux  #( .WIDTH(1) ) _47791_ ( .A(_25519_), .B(1'h1), .S(_05355_), .Y(_25520_) );
  \$mux  #( .WIDTH(8) ) _47793_ ( .A(ram_w8_l4096_id0_0_1_wdata), .B(_dataflow_slice_data_100), .S(_05355_), .Y(_25521_) );
  \$mux  #( .WIDTH(10) ) _47795_ ( .A(ram_w8_l4096_id0_0_1_addr), .B(_25939_[9:0]), .S(_05415_), .Y(_25522_) );
  \$mux  #( .WIDTH(10) ) _47796_ ( .A(_25522_), .B(_22077_[9:0]), .S(_05355_), .Y(_25523_) );
  \$mux  #( .WIDTH(10) ) _47798_ ( .A(ram_w8_l4096_id0_0_0_addr), .B(_stream_matmul_15_source_20_source_ram_raddr[11:2]), .S(_tmp_1033), .Y(_25524_) );
  \$mux  #( .WIDTH(4) ) _47800_ ( .A(_tmp_5), .B(_tmp_0[5:2]), .S(_05867_), .Y(_25525_) );
  \$mux  #( .WIDTH(4) ) _47801_ ( .A(_25525_), .B(_tmp_5), .S(_04904_), .Y(_25526_) );
  \$mux  #( .WIDTH(4) ) _47802_ ( .A(_25526_), .B(_tmp_5), .S(_RESETN_inv_2), .Y(_02883_) );
  \$mux  #( .WIDTH(32) ) _47803_ ( .A(_saxi_register_fsm), .B(0), .S(_05866_), .Y({ _21737_, _21736_, _21734_, _21733_, _21732_, _21731_, _21730_, _21729_, _21728_, _21727_, _21726_, _21725_, _21723_, _21722_, _21721_, _21720_, _21719_, _21718_, _21717_, _21716_, _21715_, _21714_, _21744_, _21743_, _21742_, _21741_, _21740_, _21739_, _21738_, _21735_, _21724_, _21713_ }) );
  \$mux  #( .WIDTH(32) ) _47804_ ( .A(_saxi_register_fsm), .B(1), .S(_tmp_2), .Y(_25528_) );
  \$mux  #( .WIDTH(32) ) _47805_ ( .A(_25528_), .B(2), .S(_tmp_1), .Y({ _21769_, _21768_, _21766_, _21765_, _21764_, _21763_, _21762_, _21761_, _21760_, _21759_, _21758_, _21757_, _21755_, _21754_, _21753_, _21752_, _21751_, _21750_, _21749_, _21748_, _21747_, _21746_, _21776_, _21775_, _21774_, _21773_, _21772_, _21771_, _21770_, _21767_, _21756_, _21745_ }) );
  \$mux  #( .WIDTH(1) ) _47810_ ( .A(1'h0), .B(1'h1), .S(_05383_), .Y(_25529_) );
  \$mux  #( .WIDTH(1) ) _47811_ ( .A(_25529_), .B(1'h0), .S(_05382_), .Y(_25530_) );
  \$mux  #( .WIDTH(1) ) _47813_ ( .A(1'h0), .B(1'h1), .S(_05382_), .Y(_25531_) );
  \$mux  #( .WIDTH(6) ) _47815_ ( .A(_tmp_0), .B(saxi_araddr), .S(_05383_), .Y(_25532_) );
  \$mux  #( .WIDTH(6) ) _47816_ ( .A(_25532_), .B(saxi_awaddr), .S(_05382_), .Y(_25533_) );
  \$mux  #( .WIDTH(1) ) _47818_ ( .A(_saxi_flag_13), .B(1'h0), .S(_05399_), .Y(_25534_) );
  \$mux  #( .WIDTH(1) ) _47820_ ( .A(_saxi_flag_12), .B(1'h0), .S(_05398_), .Y(_25535_) );
  \$mux  #( .WIDTH(1) ) _47822_ ( .A(_saxi_flag_11), .B(1'h0), .S(_05397_), .Y(_25536_) );
  \$mux  #( .WIDTH(1) ) _47824_ ( .A(_saxi_flag_10), .B(1'h0), .S(_05396_), .Y(_25537_) );
  \$mux  #( .WIDTH(1) ) _47826_ ( .A(_saxi_flag_9), .B(1'h0), .S(_05395_), .Y(_25538_) );
  \$mux  #( .WIDTH(1) ) _47828_ ( .A(_saxi_flag_8), .B(1'h0), .S(_05394_), .Y(_25539_) );
  \$mux  #( .WIDTH(1) ) _47830_ ( .A(_saxi_flag_7), .B(1'h0), .S(_05393_), .Y(_25540_) );
  \$mux  #( .WIDTH(1) ) _47832_ ( .A(_saxi_flag_6), .B(1'h0), .S(_05392_), .Y(_25541_) );
  \$mux  #( .WIDTH(1) ) _47834_ ( .A(_saxi_flag_5), .B(1'h0), .S(_05391_), .Y(_25542_) );
  \$mux  #( .WIDTH(1) ) _47835_ ( .A(1'h0), .B(_25542_), .S(_05150_), .Y(_25543_) );
  \$mux  #( .WIDTH(1) ) _47836_ ( .A(1'h0), .B(_25543_), .S(_05133_), .Y(_25544_) );
  \$mux  #( .WIDTH(1) ) _47838_ ( .A(_saxi_flag_4), .B(1'h0), .S(_05390_), .Y(_25545_) );
  \$mux  #( .WIDTH(1) ) _47839_ ( .A(1'h0), .B(_25545_), .S(_05149_), .Y(_25546_) );
  \$mux  #( .WIDTH(1) ) _47841_ ( .A(_saxi_flag_3), .B(1'h0), .S(_05389_), .Y(_25547_) );
  \$mux  #( .WIDTH(1) ) _47843_ ( .A(_saxi_flag_2), .B(1'h0), .S(_05388_), .Y(_25548_) );
  \$mux  #( .WIDTH(1) ) _47845_ ( .A(_saxi_flag_1), .B(1'h0), .S(_05387_), .Y(_25549_) );
  \$mux  #( .WIDTH(1) ) _47847_ ( .A(_saxi_flag_0), .B(1'h0), .S(_05386_), .Y(_25550_) );
  \$mux  #( .WIDTH(32) ) _47849_ ( .A(_saxi_register_13), .B(_tmp_8), .S(_05399_), .Y(_25551_) );
  \$mux  #( .WIDTH(32) ) _47850_ ( .A(_25551_), .B(saxi_wdata), .S(_05413_), .Y(_25552_) );
  \$mux  #( .WIDTH(32) ) _47851_ ( .A(_25552_), .B(3200), .S(_RESETN_inv_2), .Y(_01733_) );
  \$mux  #( .WIDTH(32) ) _47852_ ( .A(_saxi_register_12), .B(_tmp_8), .S(_05398_), .Y(_25553_) );
  \$mux  #( .WIDTH(32) ) _47853_ ( .A(_25553_), .B(saxi_wdata), .S(_05412_), .Y(_25554_) );
  \$mux  #( .WIDTH(32) ) _47854_ ( .A(_25554_), .B(64), .S(_RESETN_inv_2), .Y(_01732_) );
  \$mux  #( .WIDTH(32) ) _47855_ ( .A(_saxi_register_11), .B(_tmp_8), .S(_05397_), .Y(_25555_) );
  \$mux  #( .WIDTH(32) ) _47856_ ( .A(_25555_), .B(saxi_wdata), .S(_05411_), .Y(_25556_) );
  \$mux  #( .WIDTH(32) ) _47858_ ( .A(_saxi_register_10), .B(_tmp_8), .S(_05396_), .Y(_25557_) );
  \$mux  #( .WIDTH(32) ) _47859_ ( .A(_25557_), .B(saxi_wdata), .S(_05410_), .Y(_25558_) );
  \$mux  #( .WIDTH(32) ) _47860_ ( .A(_25558_), .B(8192), .S(_RESETN_inv_2), .Y(_01730_) );
  \$mux  #( .WIDTH(32) ) _47861_ ( .A(_saxi_register_9), .B(_tmp_8), .S(_05395_), .Y(_25559_) );
  \$mux  #( .WIDTH(32) ) _47862_ ( .A(_25559_), .B(saxi_wdata), .S(_05409_), .Y(_25560_) );
  \$mux  #( .WIDTH(32) ) _47864_ ( .A(_saxi_register_8), .B(_tmp_8), .S(_05394_), .Y(_25561_) );
  \$mux  #( .WIDTH(32) ) _47865_ ( .A(_25561_), .B(saxi_wdata), .S(_05408_), .Y(_25562_) );
  \$mux  #( .WIDTH(32) ) _47867_ ( .A(_saxi_register_7), .B(_tmp_8), .S(_05393_), .Y(_25563_) );
  \$mux  #( .WIDTH(32) ) _47868_ ( .A(_25563_), .B(saxi_wdata), .S(_05407_), .Y(_25564_) );
  \$mux  #( .WIDTH(32) ) _47869_ ( .A(0), .B(_25564_), .S(_04900_), .Y(_25565_) );
  \$mux  #( .WIDTH(32) ) _47871_ ( .A(_saxi_register_6), .B(_tmp_8), .S(_05392_), .Y(_25566_) );
  \$mux  #( .WIDTH(32) ) _47872_ ( .A(_25566_), .B(saxi_wdata), .S(_05406_), .Y(_25567_) );
  \$mux  #( .WIDTH(32) ) _47873_ ( .A(0), .B(_25567_), .S(_04900_), .Y(_25568_) );
  \$mux  #( .WIDTH(32) ) _47875_ ( .A(_saxi_register_5), .B(_tmp_8), .S(_05391_), .Y(_25569_) );
  \$mux  #( .WIDTH(32) ) _47876_ ( .A(_25569_), .B(saxi_wdata), .S(_05405_), .Y(_25570_) );
  \$mux  #( .WIDTH(32) ) _47877_ ( .A(0), .B(_25570_), .S(_04900_), .Y(_25571_) );
  \$mux  #( .WIDTH(32) ) _47878_ ( .A(1), .B(_25571_), .S(_05150_), .Y(_25572_) );
  \$mux  #( .WIDTH(32) ) _47879_ ( .A(0), .B(_25572_), .S(_05133_), .Y(_25573_) );
  \$mux  #( .WIDTH(32) ) _47881_ ( .A(_saxi_register_4), .B(_tmp_8), .S(_05390_), .Y(_25574_) );
  \$mux  #( .WIDTH(32) ) _47882_ ( .A(_25574_), .B(saxi_wdata), .S(_05404_), .Y(_25575_) );
  \$mux  #( .WIDTH(32) ) _47883_ ( .A(0), .B(_25575_), .S(_05149_), .Y(_25576_) );
  \$mux  #( .WIDTH(32) ) _47885_ ( .A(_saxi_register_3), .B(_tmp_8), .S(_05389_), .Y(_25577_) );
  \$mux  #( .WIDTH(32) ) _47886_ ( .A(_25577_), .B(saxi_wdata), .S(_05403_), .Y(_25578_) );
  \$mux  #( .WIDTH(32) ) _47888_ ( .A(_saxi_register_2), .B(_tmp_8), .S(_05388_), .Y(_25579_) );
  \$mux  #( .WIDTH(32) ) _47889_ ( .A(_25579_), .B(saxi_wdata), .S(_05402_), .Y(_25580_) );
  \$mux  #( .WIDTH(32) ) _47891_ ( .A(_saxi_register_1), .B(_tmp_8), .S(_05387_), .Y(_25581_) );
  \$mux  #( .WIDTH(32) ) _47892_ ( .A(_25581_), .B(saxi_wdata), .S(_05401_), .Y(_25582_) );
  \$mux  #( .WIDTH(32) ) _47894_ ( .A(_saxi_register_0), .B(_tmp_8), .S(_05386_), .Y(_25583_) );
  \$mux  #( .WIDTH(32) ) _47895_ ( .A(_25583_), .B(saxi_wdata), .S(_05400_), .Y(_25584_) );
  \$mux  #( .WIDTH(1) ) _47897_ ( .A(saxi_rvalid), .B(1'h0), .S(_saxi_cond_0_1), .Y(_25585_) );
  \$mux  #( .WIDTH(1) ) _47898_ ( .A(_25585_), .B(1'h1), .S(_05384_), .Y(_25586_) );
  \$mux  #( .WIDTH(1) ) _47899_ ( .A(_25586_), .B(saxi_rvalid), .S(_05385_), .Y(_25587_) );
  \$mux  #( .WIDTH(32) ) _47901_ ( .A(saxi_rdata), .B(_tmp_6), .S(_05384_), .Y(_25588_) );
  \$mux  #( .WIDTH(1) ) _47903_ ( .A(saxi_bvalid), .B(1'h0), .S(_05380_), .Y(_25589_) );
  \$mux  #( .WIDTH(1) ) _47904_ ( .A(_25589_), .B(1'h1), .S(_05381_), .Y(_25590_) );
  \$mux  #( .WIDTH(1) ) _47906_ ( .A(_dataflow__delay_valid_132), .B(1'h0), .S(_05379_), .Y(_25591_) );
  \$mux  #( .WIDTH(1) ) _47907_ ( .A(_25591_), .B(_wvalid_11), .S(_05377_), .Y(_25592_) );
  \$mux  #( .WIDTH(32) ) _47909_ ( .A(_dataflow__delay_data_132), .B(_wdata_10), .S(_05378_), .Y(_25593_) );
  \$mux  #( .WIDTH(1) ) _47911_ ( .A(_dataflow_slice_valid_122), .B(1'h0), .S(_05376_), .Y(_25594_) );
  \$mux  #( .WIDTH(1) ) _47912_ ( .A(_25594_), .B(_wvalid_974), .S(_05374_), .Y(_25595_) );
  \$mux  #( .WIDTH(8) ) _47914_ ( .A(_dataflow_slice_data_122), .B(_wdata_973[31:24]), .S(_05375_), .Y(_25596_) );
  \$mux  #( .WIDTH(1) ) _47916_ ( .A(_dataflow_slice_valid_119), .B(1'h0), .S(_05373_), .Y(_25597_) );
  \$mux  #( .WIDTH(1) ) _47917_ ( .A(_25597_), .B(_wvalid_974), .S(_05371_), .Y(_25598_) );
  \$mux  #( .WIDTH(8) ) _47919_ ( .A(_dataflow_slice_data_119), .B(_wdata_973[23:16]), .S(_05372_), .Y(_25599_) );
  \$mux  #( .WIDTH(1) ) _47921_ ( .A(_dataflow_slice_valid_116), .B(1'h0), .S(_05370_), .Y(_25600_) );
  \$mux  #( .WIDTH(1) ) _47922_ ( .A(_25600_), .B(_wvalid_974), .S(_05368_), .Y(_25601_) );
  \$mux  #( .WIDTH(8) ) _47924_ ( .A(_dataflow_slice_data_116), .B(_wdata_973[15:8]), .S(_05369_), .Y(_25602_) );
  \$mux  #( .WIDTH(1) ) _47926_ ( .A(_dataflow_slice_valid_113), .B(1'h0), .S(_05367_), .Y(_25603_) );
  \$mux  #( .WIDTH(1) ) _47927_ ( .A(_25603_), .B(_wvalid_974), .S(_05365_), .Y(_25604_) );
  \$mux  #( .WIDTH(8) ) _47929_ ( .A(_dataflow_slice_data_113), .B(_wdata_973[7:0]), .S(_05366_), .Y(_25605_) );
  \$mux  #( .WIDTH(1) ) _47931_ ( .A(_dataflow_slice_valid_109), .B(1'h0), .S(_05364_), .Y(_25606_) );
  \$mux  #( .WIDTH(1) ) _47932_ ( .A(_25606_), .B(_wvalid_963), .S(_05362_), .Y(_25607_) );
  \$mux  #( .WIDTH(8) ) _47934_ ( .A(_dataflow_slice_data_109), .B(_wdata_962[31:24]), .S(_05363_), .Y(_25608_) );
  \$mux  #( .WIDTH(1) ) _47936_ ( .A(_dataflow_slice_valid_106), .B(1'h0), .S(_05361_), .Y(_25609_) );
  \$mux  #( .WIDTH(1) ) _47937_ ( .A(_25609_), .B(_wvalid_963), .S(_05359_), .Y(_25610_) );
  \$mux  #( .WIDTH(8) ) _47939_ ( .A(_dataflow_slice_data_106), .B(_wdata_962[23:16]), .S(_05360_), .Y(_25611_) );
  \$mux  #( .WIDTH(1) ) _47941_ ( .A(_dataflow_slice_valid_103), .B(1'h0), .S(_05358_), .Y(_25612_) );
  \$mux  #( .WIDTH(1) ) _47942_ ( .A(_25612_), .B(_wvalid_963), .S(_05356_), .Y(_25613_) );
  \$mux  #( .WIDTH(8) ) _47944_ ( .A(_dataflow_slice_data_103), .B(_wdata_962[15:8]), .S(_05357_), .Y(_25614_) );
  \$mux  #( .WIDTH(1) ) _47946_ ( .A(_dataflow_slice_valid_100), .B(1'h0), .S(_05355_), .Y(_25615_) );
  \$mux  #( .WIDTH(1) ) _47947_ ( .A(_25615_), .B(_wvalid_963), .S(_05353_), .Y(_25616_) );
  \$mux  #( .WIDTH(8) ) _47949_ ( .A(_dataflow_slice_data_100), .B(_wdata_962[7:0]), .S(_05354_), .Y(_25617_) );
  \$mux  #( .WIDTH(1) ) _47951_ ( .A(_dataflow_slice_valid_87), .B(1'h0), .S(_05352_), .Y(_25618_) );
  \$mux  #( .WIDTH(1) ) _47952_ ( .A(_25618_), .B(_wvalid_852), .S(_05350_), .Y(_25619_) );
  \$mux  #( .WIDTH(8) ) _47954_ ( .A(_dataflow_slice_data_87), .B(_wdata_851[31:24]), .S(_05351_), .Y(_25620_) );
  \$mux  #( .WIDTH(1) ) _47956_ ( .A(_dataflow_slice_valid_84), .B(1'h0), .S(_05349_), .Y(_25621_) );
  \$mux  #( .WIDTH(1) ) _47957_ ( .A(_25621_), .B(_wvalid_852), .S(_05347_), .Y(_25622_) );
  \$mux  #( .WIDTH(8) ) _47959_ ( .A(_dataflow_slice_data_84), .B(_wdata_851[23:16]), .S(_05348_), .Y(_25623_) );
  \$mux  #( .WIDTH(1) ) _47961_ ( .A(_dataflow_slice_valid_81), .B(1'h0), .S(_05346_), .Y(_25624_) );
  \$mux  #( .WIDTH(1) ) _47962_ ( .A(_25624_), .B(_wvalid_852), .S(_05344_), .Y(_25625_) );
  \$mux  #( .WIDTH(8) ) _47964_ ( .A(_dataflow_slice_data_81), .B(_wdata_851[15:8]), .S(_05345_), .Y(_25626_) );
  \$mux  #( .WIDTH(1) ) _47966_ ( .A(_dataflow_slice_valid_78), .B(1'h0), .S(_05343_), .Y(_25627_) );
  \$mux  #( .WIDTH(1) ) _47967_ ( .A(_25627_), .B(_wvalid_852), .S(_05341_), .Y(_25628_) );
  \$mux  #( .WIDTH(8) ) _47969_ ( .A(_dataflow_slice_data_78), .B(_wdata_851[7:0]), .S(_05342_), .Y(_25629_) );
  \$mux  #( .WIDTH(1) ) _47971_ ( .A(_dataflow_slice_valid_65), .B(1'h0), .S(_05340_), .Y(_25630_) );
  \$mux  #( .WIDTH(1) ) _47972_ ( .A(_25630_), .B(_wvalid_274), .S(_05338_), .Y(_25631_) );
  \$mux  #( .WIDTH(8) ) _47974_ ( .A(_dataflow_slice_data_65), .B(_wdata_273[31:24]), .S(_05339_), .Y(_25632_) );
  \$mux  #( .WIDTH(1) ) _47976_ ( .A(_dataflow_slice_valid_62), .B(1'h0), .S(_05337_), .Y(_25633_) );
  \$mux  #( .WIDTH(1) ) _47977_ ( .A(_25633_), .B(_wvalid_274), .S(_05335_), .Y(_25634_) );
  \$mux  #( .WIDTH(8) ) _47979_ ( .A(_dataflow_slice_data_62), .B(_wdata_273[23:16]), .S(_05336_), .Y(_25635_) );
  \$mux  #( .WIDTH(1) ) _47981_ ( .A(_dataflow_slice_valid_59), .B(1'h0), .S(_05334_), .Y(_25636_) );
  \$mux  #( .WIDTH(1) ) _47982_ ( .A(_25636_), .B(_wvalid_274), .S(_05332_), .Y(_25637_) );
  \$mux  #( .WIDTH(8) ) _47984_ ( .A(_dataflow_slice_data_59), .B(_wdata_273[15:8]), .S(_05333_), .Y(_25638_) );
  \$mux  #( .WIDTH(1) ) _47986_ ( .A(_dataflow_slice_valid_56), .B(1'h0), .S(_05331_), .Y(_25639_) );
  \$mux  #( .WIDTH(1) ) _47987_ ( .A(_25639_), .B(_wvalid_274), .S(_05329_), .Y(_25640_) );
  \$mux  #( .WIDTH(8) ) _47989_ ( .A(_dataflow_slice_data_56), .B(_wdata_273[7:0]), .S(_05330_), .Y(_25641_) );
  \$mux  #( .WIDTH(1) ) _47991_ ( .A(_dataflow_slice_valid_52), .B(1'h0), .S(_05328_), .Y(_25642_) );
  \$mux  #( .WIDTH(1) ) _47992_ ( .A(_25642_), .B(_wvalid_217), .S(_05326_), .Y(_25643_) );
  \$mux  #( .WIDTH(8) ) _47994_ ( .A(_dataflow_slice_data_52), .B(_wdata_216[31:24]), .S(_05327_), .Y(_25644_) );
  \$mux  #( .WIDTH(1) ) _47996_ ( .A(_dataflow_slice_valid_49), .B(1'h0), .S(_05325_), .Y(_25645_) );
  \$mux  #( .WIDTH(1) ) _47997_ ( .A(_25645_), .B(_wvalid_217), .S(_05323_), .Y(_25646_) );
  \$mux  #( .WIDTH(8) ) _47999_ ( .A(_dataflow_slice_data_49), .B(_wdata_216[23:16]), .S(_05324_), .Y(_25647_) );
  \$mux  #( .WIDTH(1) ) _48001_ ( .A(_dataflow_slice_valid_46), .B(1'h0), .S(_05322_), .Y(_25648_) );
  \$mux  #( .WIDTH(1) ) _48002_ ( .A(_25648_), .B(_wvalid_217), .S(_05320_), .Y(_25649_) );
  \$mux  #( .WIDTH(8) ) _48004_ ( .A(_dataflow_slice_data_46), .B(_wdata_216[15:8]), .S(_05321_), .Y(_25650_) );
  \$mux  #( .WIDTH(1) ) _48006_ ( .A(_dataflow_slice_valid_43), .B(1'h0), .S(_05319_), .Y(_25651_) );
  \$mux  #( .WIDTH(1) ) _48007_ ( .A(_25651_), .B(_wvalid_217), .S(_05317_), .Y(_25652_) );
  \$mux  #( .WIDTH(8) ) _48009_ ( .A(_dataflow_slice_data_43), .B(_wdata_216[7:0]), .S(_05318_), .Y(_25653_) );
  \$mux  #( .WIDTH(1) ) _48011_ ( .A(_dataflow_slice_valid_39), .B(1'h0), .S(_05316_), .Y(_25654_) );
  \$mux  #( .WIDTH(1) ) _48012_ ( .A(_25654_), .B(_wvalid_160), .S(_05314_), .Y(_25655_) );
  \$mux  #( .WIDTH(8) ) _48014_ ( .A(_dataflow_slice_data_39), .B(_wdata_159[31:24]), .S(_05315_), .Y(_25656_) );
  \$mux  #( .WIDTH(1) ) _48016_ ( .A(_dataflow_slice_valid_36), .B(1'h0), .S(_05313_), .Y(_25657_) );
  \$mux  #( .WIDTH(1) ) _48017_ ( .A(_25657_), .B(_wvalid_160), .S(_05311_), .Y(_25658_) );
  \$mux  #( .WIDTH(8) ) _48019_ ( .A(_dataflow_slice_data_36), .B(_wdata_159[23:16]), .S(_05312_), .Y(_25659_) );
  \$mux  #( .WIDTH(1) ) _48021_ ( .A(_dataflow_slice_valid_33), .B(1'h0), .S(_05310_), .Y(_25660_) );
  \$mux  #( .WIDTH(1) ) _48022_ ( .A(_25660_), .B(_wvalid_160), .S(_05308_), .Y(_25661_) );
  \$mux  #( .WIDTH(8) ) _48024_ ( .A(_dataflow_slice_data_33), .B(_wdata_159[15:8]), .S(_05309_), .Y(_25662_) );
  \$mux  #( .WIDTH(1) ) _48026_ ( .A(_dataflow_slice_valid_30), .B(1'h0), .S(_05307_), .Y(_25663_) );
  \$mux  #( .WIDTH(1) ) _48027_ ( .A(_25663_), .B(_wvalid_160), .S(_05305_), .Y(_25664_) );
  \$mux  #( .WIDTH(8) ) _48029_ ( .A(_dataflow_slice_data_30), .B(_wdata_159[7:0]), .S(_05306_), .Y(_25665_) );
  \$mux  #( .WIDTH(1) ) _48031_ ( .A(_dataflow_slice_valid_26), .B(1'h0), .S(_05304_), .Y(_25666_) );
  \$mux  #( .WIDTH(1) ) _48032_ ( .A(_25666_), .B(_wvalid_31), .S(_05302_), .Y(_25667_) );
  \$mux  #( .WIDTH(8) ) _48034_ ( .A(_dataflow_slice_data_26), .B(_wdata_30[31:24]), .S(_05303_), .Y(_25668_) );
  \$mux  #( .WIDTH(1) ) _48036_ ( .A(_dataflow_slice_valid_23), .B(1'h0), .S(_05301_), .Y(_25669_) );
  \$mux  #( .WIDTH(1) ) _48037_ ( .A(_25669_), .B(_wvalid_31), .S(_05299_), .Y(_25670_) );
  \$mux  #( .WIDTH(8) ) _48039_ ( .A(_dataflow_slice_data_23), .B(_wdata_30[23:16]), .S(_05300_), .Y(_25671_) );
  \$mux  #( .WIDTH(1) ) _48041_ ( .A(_dataflow_slice_valid_20), .B(1'h0), .S(_05298_), .Y(_25672_) );
  \$mux  #( .WIDTH(1) ) _48042_ ( .A(_25672_), .B(_wvalid_31), .S(_05296_), .Y(_25673_) );
  \$mux  #( .WIDTH(8) ) _48044_ ( .A(_dataflow_slice_data_20), .B(_wdata_30[15:8]), .S(_05297_), .Y(_25674_) );
  \$mux  #( .WIDTH(1) ) _48046_ ( .A(_dataflow_slice_valid_17), .B(1'h0), .S(_05295_), .Y(_25675_) );
  \$mux  #( .WIDTH(1) ) _48047_ ( .A(_25675_), .B(_wvalid_31), .S(_05293_), .Y(_25676_) );
  \$mux  #( .WIDTH(8) ) _48049_ ( .A(_dataflow_slice_data_17), .B(_wdata_30[7:0]), .S(_05294_), .Y(_25677_) );
  \$mux  #( .WIDTH(1) ) _48051_ ( .A(_dataflow_slice_valid_13), .B(1'h0), .S(_05292_), .Y(_25678_) );
  \$mux  #( .WIDTH(1) ) _48052_ ( .A(_25678_), .B(_wvalid_18), .S(_05290_), .Y(_25679_) );
  \$mux  #( .WIDTH(8) ) _48054_ ( .A(_dataflow_slice_data_13), .B(_wdata_17[31:24]), .S(_05291_), .Y(_25680_) );
  \$mux  #( .WIDTH(1) ) _48056_ ( .A(_dataflow_slice_valid_10), .B(1'h0), .S(_05289_), .Y(_25681_) );
  \$mux  #( .WIDTH(1) ) _48057_ ( .A(_25681_), .B(_wvalid_18), .S(_05287_), .Y(_25682_) );
  \$mux  #( .WIDTH(8) ) _48059_ ( .A(_dataflow_slice_data_10), .B(_wdata_17[23:16]), .S(_05288_), .Y(_25683_) );
  \$mux  #( .WIDTH(1) ) _48061_ ( .A(_dataflow_slice_valid_7), .B(1'h0), .S(_05286_), .Y(_25684_) );
  \$mux  #( .WIDTH(1) ) _48062_ ( .A(_25684_), .B(_wvalid_18), .S(_05284_), .Y(_25685_) );
  \$mux  #( .WIDTH(8) ) _48064_ ( .A(_dataflow_slice_data_7), .B(_wdata_17[15:8]), .S(_05285_), .Y(_25686_) );
  \$mux  #( .WIDTH(1) ) _48066_ ( .A(_dataflow_slice_valid_4), .B(1'h0), .S(_05283_), .Y(_25687_) );
  \$mux  #( .WIDTH(1) ) _48067_ ( .A(_25687_), .B(_wvalid_18), .S(_05281_), .Y(_25688_) );
  \$mux  #( .WIDTH(8) ) _48069_ ( .A(_dataflow_slice_data_4), .B(_wdata_17[7:0]), .S(_05282_), .Y(_25689_) );
  \$mux  #( .WIDTH(1) ) _48071_ ( .A(_tmp_1167), .B(1'h0), .S(_saxi_cond_0_1), .Y(_25690_) );
  \$mux  #( .WIDTH(1) ) _48072_ ( .A(_25690_), .B(1'h1), .S(_05280_), .Y(_25691_) );
  \$mux  #( .WIDTH(1) ) _48073_ ( .A(_25691_), .B(_tmp_1167), .S(_05276_), .Y(_25692_) );
  \$mux  #( .WIDTH(32) ) _48075_ ( .A(_maxi_ram_w8_l2048_id1_1_write_local_stride), .B(1), .S(axim_flag_1118), .Y(_25693_) );
  \$mux  #( .WIDTH(33) ) _48077_ ( .A(_maxi_ram_w8_l2048_id1_1_write_size), .B(_22076_), .S(axim_flag_1118), .Y(_25694_) );
  \$mux  #( .WIDTH(32) ) _48079_ ( .A(_maxi_ram_w8_l2048_id1_1_write_global_addr), .B(_22075_), .S(axim_flag_1118), .Y(_25695_) );
  \$mux  #( .WIDTH(32) ) _48081_ ( .A(_maxi_ram_w8_l2048_id1_1_write_local_addr), .B({ 2'h0, _22074_[31:2] }), .S(axim_flag_1118), .Y(_25696_) );
  \$mux  #( .WIDTH(8) ) _48083_ ( .A(_maxi_ram_w8_l2048_id1_1_write_op_sel), .B(8'h03), .S(axim_flag_1118), .Y(_25697_) );
  \$mux  #( .WIDTH(1) ) _48085_ ( .A(1'h0), .B(1'h1), .S(axim_flag_1118), .Y(_25698_) );
  \$mux  #( .WIDTH(32) ) _48087_ ( .A(_maxi_ram_w8_l2048_id2_1_read_local_stride), .B(1), .S(axim_flag_972), .Y(_25699_) );
  \$mux  #( .WIDTH(33) ) _48089_ ( .A(_maxi_ram_w8_l2048_id2_1_read_size), .B(33'h000000048), .S(axim_flag_972), .Y(_25700_) );
  \$mux  #( .WIDTH(32) ) _48091_ ( .A(_maxi_ram_w8_l2048_id2_1_read_global_addr), .B(matmul_15_mux_act_gaddr_0), .S(axim_flag_972), .Y(_25701_) );
  \$mux  #( .WIDTH(32) ) _48093_ ( .A(_maxi_ram_w8_l2048_id2_1_read_local_addr), .B({ 2'h0, matmul_15_act_page_dma_offset_0[31:2] }), .S(axim_flag_972), .Y(_25702_) );
  \$mux  #( .WIDTH(8) ) _48095_ ( .A(_maxi_ram_w8_l2048_id2_1_read_op_sel), .B(8'h09), .S(axim_flag_972), .Y(_25703_) );
  \$mux  #( .WIDTH(1) ) _48097_ ( .A(1'h0), .B(1'h1), .S(axim_flag_972), .Y(_25704_) );
  \$mux  #( .WIDTH(32) ) _48099_ ( .A(_maxi_ram_w8_l4096_id0_1_read_local_stride), .B(1), .S(axim_flag_961), .Y(_25705_) );
  \$mux  #( .WIDTH(33) ) _48101_ ( .A(_maxi_ram_w8_l4096_id0_1_read_size), .B(33'h000000120), .S(axim_flag_961), .Y(_25706_) );
  \$mux  #( .WIDTH(32) ) _48103_ ( .A(_maxi_ram_w8_l4096_id0_1_read_global_addr), .B(_22073_), .S(axim_flag_961), .Y(_25707_) );
  \$mux  #( .WIDTH(32) ) _48105_ ( .A(_maxi_ram_w8_l4096_id0_1_read_local_addr), .B({ 2'h0, matmul_15_filter_page_dma_offset[31:2] }), .S(axim_flag_961), .Y(_25708_) );
  \$mux  #( .WIDTH(8) ) _48107_ ( .A(_maxi_ram_w8_l4096_id0_1_read_op_sel), .B(8'h08), .S(axim_flag_961), .Y(_25709_) );
  \$mux  #( .WIDTH(1) ) _48109_ ( .A(1'h0), .B(1'h1), .S(axim_flag_961), .Y(_25710_) );
  \$mux  #( .WIDTH(1) ) _48111_ ( .A(_tmp_958), .B(1'h0), .S(_saxi_cond_0_1), .Y(_25711_) );
  \$mux  #( .WIDTH(1) ) _48112_ ( .A(_25711_), .B(1'h1), .S(_05278_), .Y(_25712_) );
  \$mux  #( .WIDTH(1) ) _48113_ ( .A(_25712_), .B(_tmp_958), .S(_05276_), .Y(_25713_) );
  \$mux  #( .WIDTH(32) ) _48115_ ( .A(_maxi_ram_w8_l2048_id0_1_write_local_stride), .B(1), .S(axim_flag_909), .Y(_25714_) );
  \$mux  #( .WIDTH(33) ) _48117_ ( .A(_maxi_ram_w8_l2048_id0_1_write_size), .B(_22072_), .S(axim_flag_909), .Y(_25715_) );
  \$mux  #( .WIDTH(32) ) _48119_ ( .A(_maxi_ram_w8_l2048_id0_1_write_global_addr), .B(_22071_), .S(axim_flag_909), .Y(_25716_) );
  \$mux  #( .WIDTH(32) ) _48121_ ( .A(_maxi_ram_w8_l2048_id0_1_write_local_addr), .B({ 2'h0, max_pool_serial_9_out_page_dma_offset[31:2] }), .S(axim_flag_909), .Y(_25717_) );
  \$mux  #( .WIDTH(8) ) _48123_ ( .A(_maxi_ram_w8_l2048_id0_1_write_op_sel), .B(8'h02), .S(axim_flag_909), .Y(_25718_) );
  \$mux  #( .WIDTH(1) ) _48125_ ( .A(1'h0), .B(1'h1), .S(axim_flag_909), .Y(_25719_) );
  \$mux  #( .WIDTH(32) ) _48127_ ( .A(_maxi_ram_w8_l2048_id1_1_read_local_stride), .B(1), .S(axim_flag_850), .Y(_25720_) );
  \$mux  #( .WIDTH(32) ) _48128_ ( .A(_25720_), .B(1), .S(axim_flag_861), .Y(_25721_) );
  \$mux  #( .WIDTH(33) ) _48130_ ( .A(_maxi_ram_w8_l2048_id1_1_read_size), .B(_22067_), .S(axim_flag_850), .Y(_25722_) );
  \$mux  #( .WIDTH(33) ) _48131_ ( .A(_25722_), .B(_22067_), .S(axim_flag_861), .Y(_25723_) );
  \$mux  #( .WIDTH(32) ) _48133_ ( .A(_maxi_ram_w8_l2048_id1_1_read_global_addr), .B(_22066_), .S(axim_flag_850), .Y(_25724_) );
  \$mux  #( .WIDTH(32) ) _48134_ ( .A(_25724_), .B(_22070_), .S(axim_flag_861), .Y(_25725_) );
  \$mux  #( .WIDTH(32) ) _48136_ ( .A(_maxi_ram_w8_l2048_id1_1_read_local_addr), .B({ 2'h0, max_pool_serial_9_act_page_dma_offset[31:2] }), .S(axim_flag_850), .Y(_25726_) );
  \$mux  #( .WIDTH(32) ) _48137_ ( .A(_25726_), .B({ 2'h0, _22068_[31:2] }), .S(axim_flag_861), .Y(_25727_) );
  \$mux  #( .WIDTH(8) ) _48139_ ( .A(_maxi_ram_w8_l2048_id1_1_read_op_sel), .B(8'h07), .S(axim_flag_850), .Y(_25728_) );
  \$mux  #( .WIDTH(8) ) _48140_ ( .A(_25728_), .B(8'h07), .S(axim_flag_861), .Y(_25729_) );
  \$mux  #( .WIDTH(1) ) _48142_ ( .A(1'h0), .B(1'h1), .S(axim_flag_850), .Y(_25730_) );
  \$mux  #( .WIDTH(1) ) _48143_ ( .A(_25730_), .B(1'h1), .S(axim_flag_861), .Y(_25731_) );
  \$mux  #( .WIDTH(1) ) _48145_ ( .A(_tmp_848), .B(1'h0), .S(_saxi_cond_0_1), .Y(_25732_) );
  \$mux  #( .WIDTH(1) ) _48146_ ( .A(_25732_), .B(1'h1), .S(_05275_), .Y(_25733_) );
  \$mux  #( .WIDTH(1) ) _48147_ ( .A(_25733_), .B(_tmp_848), .S(_05276_), .Y(_25734_) );
  \$mux  #( .WIDTH(9) ) _48149_ ( .A(_tmp_847), .B(_maxi_write_cur_size[8:0]), .S(_05271_), .Y(_25735_) );
  \$mux  #( .WIDTH(9) ) _48150_ ( .A(_25735_), .B(_25938_[8:0]), .S(_05274_), .Y(_25736_) );
  \$mux  #( .WIDTH(9) ) _48151_ ( .A(_25736_), .B(_25938_[8:0]), .S(_05277_), .Y(_25737_) );
  \$mux  #( .WIDTH(9) ) _48152_ ( .A(_25737_), .B(_25938_[8:0]), .S(_05279_), .Y(_25738_) );
  \$mux  #( .WIDTH(32) ) _48154_ ( .A(_maxi_ram_w8_l2048_id19_1_write_local_stride), .B(1), .S(axim_flag_798), .Y(_25739_) );
  \$mux  #( .WIDTH(33) ) _48156_ ( .A(_maxi_ram_w8_l2048_id19_1_write_size), .B(_22065_), .S(axim_flag_798), .Y(_25740_) );
  \$mux  #( .WIDTH(32) ) _48158_ ( .A(_maxi_ram_w8_l2048_id19_1_write_global_addr), .B(_22064_), .S(axim_flag_798), .Y(_25741_) );
  \$mux  #( .WIDTH(32) ) _48160_ ( .A(_maxi_ram_w8_l2048_id19_1_write_local_addr), .B({ 2'h0, _22063_[31:2] }), .S(axim_flag_798), .Y(_25742_) );
  \$mux  #( .WIDTH(8) ) _48162_ ( .A(_maxi_ram_w8_l2048_id19_1_write_op_sel), .B(8'h01), .S(axim_flag_798), .Y(_25743_) );
  \$mux  #( .WIDTH(1) ) _48164_ ( .A(1'h0), .B(1'h1), .S(axim_flag_798), .Y(_25744_) );
  \$mux  #( .WIDTH(32) ) _48166_ ( .A(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_local_stride), .B(1), .S(axim_flag_272), .Y(_25745_) );
  \$mux  #( .WIDTH(33) ) _48168_ ( .A(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_size), .B(_22062_), .S(axim_flag_272), .Y(_25746_) );
  \$mux  #( .WIDTH(32) ) _48170_ ( .A(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_global_addr), .B(conv2d_8_mux_act_gaddr_2), .S(axim_flag_272), .Y(_25747_) );
  \$mux  #( .WIDTH(32) ) _48172_ ( .A(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_local_addr), .B({ 2'h0, conv2d_8_act_page_dma_offset_2[31:2] }), .S(axim_flag_272), .Y(_25748_) );
  \$mux  #( .WIDTH(8) ) _48174_ ( .A(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_op_sel), .B(8'h06), .S(axim_flag_272), .Y(_25749_) );
  \$mux  #( .WIDTH(1) ) _48176_ ( .A(1'h0), .B(1'h1), .S(axim_flag_272), .Y(_25750_) );
  \$mux  #( .WIDTH(32) ) _48178_ ( .A(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_local_stride), .B(1), .S(axim_flag_215), .Y(_25751_) );
  \$mux  #( .WIDTH(33) ) _48180_ ( .A(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_size), .B(_22062_), .S(axim_flag_215), .Y(_25752_) );
  \$mux  #( .WIDTH(32) ) _48182_ ( .A(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_global_addr), .B(conv2d_8_mux_act_gaddr_1), .S(axim_flag_215), .Y(_25753_) );
  \$mux  #( .WIDTH(32) ) _48184_ ( .A(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_local_addr), .B({ 2'h0, conv2d_8_act_page_dma_offset_1[31:2] }), .S(axim_flag_215), .Y(_25754_) );
  \$mux  #( .WIDTH(8) ) _48186_ ( .A(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_op_sel), .B(8'h05), .S(axim_flag_215), .Y(_25755_) );
  \$mux  #( .WIDTH(1) ) _48188_ ( .A(1'h0), .B(1'h1), .S(axim_flag_215), .Y(_25756_) );
  \$mux  #( .WIDTH(32) ) _48190_ ( .A(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_local_stride), .B(1), .S(axim_flag_158), .Y(_25757_) );
  \$mux  #( .WIDTH(33) ) _48192_ ( .A(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_size), .B(_22062_), .S(axim_flag_158), .Y(_25758_) );
  \$mux  #( .WIDTH(32) ) _48194_ ( .A(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_global_addr), .B(conv2d_8_mux_act_gaddr_0), .S(axim_flag_158), .Y(_25759_) );
  \$mux  #( .WIDTH(32) ) _48196_ ( .A(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_local_addr), .B({ 2'h0, conv2d_8_act_page_dma_offset_0[31:2] }), .S(axim_flag_158), .Y(_25760_) );
  \$mux  #( .WIDTH(8) ) _48198_ ( .A(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_op_sel), .B(8'h04), .S(axim_flag_158), .Y(_25761_) );
  \$mux  #( .WIDTH(1) ) _48200_ ( .A(1'h0), .B(1'h1), .S(axim_flag_158), .Y(_25762_) );
  \$mux  #( .WIDTH(32) ) _48202_ ( .A(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_local_stride), .B(1), .S(axim_flag_29), .Y(_25763_) );
  \$mux  #( .WIDTH(33) ) _48204_ ( .A(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_size), .B(_22061_), .S(axim_flag_29), .Y(_25764_) );
  \$mux  #( .WIDTH(32) ) _48206_ ( .A(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_global_addr), .B(_22060_), .S(axim_flag_29), .Y(_25765_) );
  \$mux  #( .WIDTH(32) ) _48208_ ( .A(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_local_addr), .B({ 2'h0, conv2d_8_filter_page_dma_offset[31:2] }), .S(axim_flag_29), .Y(_25766_) );
  \$mux  #( .WIDTH(8) ) _48210_ ( .A(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_op_sel), .B(8'h03), .S(axim_flag_29), .Y(_25767_) );
  \$mux  #( .WIDTH(1) ) _48212_ ( .A(1'h0), .B(1'h1), .S(axim_flag_29), .Y(_25768_) );
  \$mux  #( .WIDTH(32) ) _48214_ ( .A(_maxi_ram_w8_l2048_id0_1_read_local_stride), .B(1), .S(axim_flag_16), .Y(_25769_) );
  \$mux  #( .WIDTH(32) ) _48215_ ( .A(_25769_), .B(1), .S(axim_flag_960), .Y(_25770_) );
  \$mux  #( .WIDTH(33) ) _48217_ ( .A(_maxi_ram_w8_l2048_id0_1_read_size), .B(33'h000000001), .S(axim_flag_16), .Y(_25771_) );
  \$mux  #( .WIDTH(33) ) _48218_ ( .A(_25771_), .B(33'h000000001), .S(axim_flag_960), .Y(_25772_) );
  \$mux  #( .WIDTH(32) ) _48220_ ( .A(_maxi_ram_w8_l2048_id0_1_read_global_addr), .B(conv2d_8_arg_objaddr_3), .S(axim_flag_16), .Y(_25773_) );
  \$mux  #( .WIDTH(32) ) _48221_ ( .A(_25773_), .B(matmul_15_arg_objaddr_3), .S(axim_flag_960), .Y(_25774_) );
  \$mux  #( .WIDTH(32) ) _48223_ ( .A(_maxi_ram_w8_l2048_id0_1_read_local_addr), .B(0), .S(axim_flag_16), .Y(_25775_) );
  \$mux  #( .WIDTH(32) ) _48224_ ( .A(_25775_), .B(0), .S(axim_flag_960), .Y(_25776_) );
  \$mux  #( .WIDTH(8) ) _48226_ ( .A(_maxi_ram_w8_l2048_id0_1_read_op_sel), .B(8'h02), .S(axim_flag_16), .Y(_25777_) );
  \$mux  #( .WIDTH(8) ) _48227_ ( .A(_25777_), .B(8'h02), .S(axim_flag_960), .Y(_25778_) );
  \$mux  #( .WIDTH(1) ) _48229_ ( .A(1'h0), .B(1'h1), .S(axim_flag_16), .Y(_25779_) );
  \$mux  #( .WIDTH(1) ) _48230_ ( .A(_25779_), .B(1'h1), .S(axim_flag_960), .Y(_25780_) );
  \$mux  #( .WIDTH(9) ) _48232_ ( .A(_tmp_14), .B(_maxi_read_cur_size[8:0]), .S(_05268_), .Y(_25781_) );
  \$mux  #( .WIDTH(9) ) _48233_ ( .A(_25781_), .B(_25936_[8:0]), .S(_05270_), .Y(_25782_) );
  \$mux  #( .WIDTH(32) ) _48235_ ( .A(_maxi_ram_w32_l128_id0_1_read_local_stride), .B(1), .S(axim_flag_9), .Y(_25783_) );
  \$mux  #( .WIDTH(32) ) _48236_ ( .A(_25783_), .B(1), .S(axim_flag_959), .Y(_25784_) );
  \$mux  #( .WIDTH(33) ) _48238_ ( .A(_maxi_ram_w32_l128_id0_1_read_size), .B({ 28'h0000000, cparam_conv2d_8_bias_num }), .S(axim_flag_9), .Y(_25785_) );
  \$mux  #( .WIDTH(33) ) _48239_ ( .A(_25785_), .B(33'h00000000a), .S(axim_flag_959), .Y(_25786_) );
  \$mux  #( .WIDTH(32) ) _48241_ ( .A(_maxi_ram_w32_l128_id0_1_read_global_addr), .B(conv2d_8_arg_objaddr_2), .S(axim_flag_9), .Y(_25787_) );
  \$mux  #( .WIDTH(32) ) _48242_ ( .A(_25787_), .B(matmul_15_arg_objaddr_2), .S(axim_flag_959), .Y(_25788_) );
  \$mux  #( .WIDTH(32) ) _48244_ ( .A(_maxi_ram_w32_l128_id0_1_read_local_addr), .B(0), .S(axim_flag_9), .Y(_25789_) );
  \$mux  #( .WIDTH(32) ) _48245_ ( .A(_25789_), .B(0), .S(axim_flag_959), .Y(_25790_) );
  \$mux  #( .WIDTH(8) ) _48247_ ( .A(_maxi_ram_w32_l128_id0_1_read_op_sel), .B(8'h01), .S(axim_flag_9), .Y(_25791_) );
  \$mux  #( .WIDTH(8) ) _48248_ ( .A(_25791_), .B(8'h01), .S(axim_flag_959), .Y(_25792_) );
  \$mux  #( .WIDTH(1) ) _48250_ ( .A(1'h0), .B(1'h1), .S(axim_flag_9), .Y(_25793_) );
  \$mux  #( .WIDTH(1) ) _48251_ ( .A(_25793_), .B(1'h1), .S(axim_flag_959), .Y(_25794_) );
  \$mux  #( .WIDTH(1) ) _48254_ ( .A(_maxi_write_idle), .B(1'h0), .S(_maxi_ram_w8_l2048_id19_1_write_start), .Y(_25795_) );
  \$mux  #( .WIDTH(1) ) _48255_ ( .A(_25795_), .B(1'h1), .S(axim_flag_849), .Y(_25796_) );
  \$mux  #( .WIDTH(1) ) _48256_ ( .A(_25796_), .B(1'h0), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_25797_) );
  \$mux  #( .WIDTH(1) ) _48257_ ( .A(_25797_), .B(1'h0), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_25798_) );
  \$mux  #( .WIDTH(1) ) _48258_ ( .A(_25798_), .B(1'h1), .S(_RESETN_inv_2), .Y(_01657_) );
  \$mux  #( .WIDTH(32) ) _48259_ ( .A(_maxi_write_local_stride), .B(_maxi_ram_w8_l2048_id19_1_write_local_stride), .S(_maxi_ram_w8_l2048_id19_1_write_start), .Y(_25799_) );
  \$mux  #( .WIDTH(32) ) _48260_ ( .A(_25799_), .B(_maxi_ram_w8_l2048_id0_1_write_local_stride), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_25800_) );
  \$mux  #( .WIDTH(32) ) _48261_ ( .A(_25800_), .B(_maxi_ram_w8_l2048_id1_1_write_local_stride), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_25801_) );
  \$mux  #( .WIDTH(33) ) _48263_ ( .A(_maxi_write_size), .B(_maxi_ram_w8_l2048_id19_1_write_size), .S(_maxi_ram_w8_l2048_id19_1_write_start), .Y(_25802_) );
  \$mux  #( .WIDTH(33) ) _48264_ ( .A(_25802_), .B(_maxi_ram_w8_l2048_id0_1_write_size), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_25803_) );
  \$mux  #( .WIDTH(33) ) _48265_ ( .A(_25803_), .B(_maxi_ram_w8_l2048_id1_1_write_size), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_25804_) );
  \$mux  #( .WIDTH(32) ) _48267_ ( .A(_maxi_write_global_addr), .B(_maxi_ram_w8_l2048_id19_1_write_global_addr), .S(_maxi_ram_w8_l2048_id19_1_write_start), .Y(_25805_) );
  \$mux  #( .WIDTH(32) ) _48268_ ( .A(_25805_), .B(_maxi_ram_w8_l2048_id0_1_write_global_addr), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_25806_) );
  \$mux  #( .WIDTH(32) ) _48269_ ( .A(_25806_), .B(_maxi_ram_w8_l2048_id1_1_write_global_addr), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_25807_) );
  \$mux  #( .WIDTH(32) ) _48271_ ( .A(_maxi_write_local_addr), .B(_maxi_ram_w8_l2048_id19_1_write_local_addr), .S(_maxi_ram_w8_l2048_id19_1_write_start), .Y(_25808_) );
  \$mux  #( .WIDTH(32) ) _48272_ ( .A(_25808_), .B(_maxi_ram_w8_l2048_id0_1_write_local_addr), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_25809_) );
  \$mux  #( .WIDTH(32) ) _48273_ ( .A(_25809_), .B(_maxi_ram_w8_l2048_id1_1_write_local_addr), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_25810_) );
  \$mux  #( .WIDTH(8) ) _48275_ ( .A(_maxi_write_op_sel), .B(_maxi_ram_w8_l2048_id19_1_write_op_sel), .S(_maxi_ram_w8_l2048_id19_1_write_start), .Y(_25811_) );
  \$mux  #( .WIDTH(8) ) _48276_ ( .A(_25811_), .B(_maxi_ram_w8_l2048_id0_1_write_op_sel), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_25812_) );
  \$mux  #( .WIDTH(8) ) _48277_ ( .A(_25812_), .B(_maxi_ram_w8_l2048_id1_1_write_op_sel), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_25813_) );
  \$mux  #( .WIDTH(1) ) _48279_ ( .A(1'h0), .B(1'h1), .S(_maxi_ram_w8_l2048_id19_1_write_start), .Y(_25814_) );
  \$mux  #( .WIDTH(1) ) _48280_ ( .A(_25814_), .B(1'h1), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_25815_) );
  \$mux  #( .WIDTH(1) ) _48281_ ( .A(_25815_), .B(1'h1), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_25816_) );
  \$mux  #( .WIDTH(1) ) _48283_ ( .A(_maxi_read_idle), .B(1'h0), .S(_maxi_ram_w32_l128_id0_1_read_start), .Y(_25817_) );
  \$mux  #( .WIDTH(1) ) _48284_ ( .A(_25817_), .B(1'h1), .S(axim_flag_15), .Y(_25818_) );
  \$mux  #( .WIDTH(1) ) _48285_ ( .A(_25818_), .B(1'h0), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_25819_) );
  \$mux  #( .WIDTH(1) ) _48286_ ( .A(_25819_), .B(1'h0), .S(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_start), .Y(_25820_) );
  \$mux  #( .WIDTH(1) ) _48287_ ( .A(_25820_), .B(1'h0), .S(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_start), .Y(_25821_) );
  \$mux  #( .WIDTH(1) ) _48288_ ( .A(_25821_), .B(1'h0), .S(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_start), .Y(_25822_) );
  \$mux  #( .WIDTH(1) ) _48289_ ( .A(_25822_), .B(1'h0), .S(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_start), .Y(_25823_) );
  \$mux  #( .WIDTH(1) ) _48290_ ( .A(_25823_), .B(1'h0), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_25824_) );
  \$mux  #( .WIDTH(1) ) _48291_ ( .A(_25824_), .B(1'h0), .S(_maxi_ram_w8_l4096_id0_1_read_start), .Y(_25825_) );
  \$mux  #( .WIDTH(1) ) _48292_ ( .A(_25825_), .B(1'h0), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_25826_) );
  \$mux  #( .WIDTH(1) ) _48293_ ( .A(_25826_), .B(1'h1), .S(_RESETN_inv_2), .Y(_01646_) );
  \$mux  #( .WIDTH(32) ) _48294_ ( .A(_maxi_read_local_stride), .B(_maxi_ram_w32_l128_id0_1_read_local_stride), .S(_maxi_ram_w32_l128_id0_1_read_start), .Y(_25827_) );
  \$mux  #( .WIDTH(32) ) _48295_ ( .A(_25827_), .B(_maxi_ram_w8_l2048_id0_1_read_local_stride), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_25828_) );
  \$mux  #( .WIDTH(32) ) _48296_ ( .A(_25828_), .B(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_local_stride), .S(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_start), .Y(_25829_) );
  \$mux  #( .WIDTH(32) ) _48297_ ( .A(_25829_), .B(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_local_stride), .S(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_start), .Y(_25830_) );
  \$mux  #( .WIDTH(32) ) _48298_ ( .A(_25830_), .B(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_local_stride), .S(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_start), .Y(_25831_) );
  \$mux  #( .WIDTH(32) ) _48299_ ( .A(_25831_), .B(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_local_stride), .S(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_start), .Y(_25832_) );
  \$mux  #( .WIDTH(32) ) _48300_ ( .A(_25832_), .B(_maxi_ram_w8_l2048_id1_1_read_local_stride), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_25833_) );
  \$mux  #( .WIDTH(32) ) _48301_ ( .A(_25833_), .B(_maxi_ram_w8_l4096_id0_1_read_local_stride), .S(_maxi_ram_w8_l4096_id0_1_read_start), .Y(_25834_) );
  \$mux  #( .WIDTH(32) ) _48302_ ( .A(_25834_), .B(_maxi_ram_w8_l2048_id2_1_read_local_stride), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_25835_) );
  \$mux  #( .WIDTH(33) ) _48304_ ( .A(_maxi_read_size), .B(_maxi_ram_w32_l128_id0_1_read_size), .S(_maxi_ram_w32_l128_id0_1_read_start), .Y(_25836_) );
  \$mux  #( .WIDTH(33) ) _48305_ ( .A(_25836_), .B(_maxi_ram_w8_l2048_id0_1_read_size), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_25837_) );
  \$mux  #( .WIDTH(33) ) _48306_ ( .A(_25837_), .B(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_size), .S(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_start), .Y(_25838_) );
  \$mux  #( .WIDTH(33) ) _48307_ ( .A(_25838_), .B(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_size), .S(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_start), .Y(_25839_) );
  \$mux  #( .WIDTH(33) ) _48308_ ( .A(_25839_), .B(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_size), .S(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_start), .Y(_25840_) );
  \$mux  #( .WIDTH(33) ) _48309_ ( .A(_25840_), .B(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_size), .S(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_start), .Y(_25841_) );
  \$mux  #( .WIDTH(33) ) _48310_ ( .A(_25841_), .B(_maxi_ram_w8_l2048_id1_1_read_size), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_25842_) );
  \$mux  #( .WIDTH(33) ) _48311_ ( .A(_25842_), .B(_maxi_ram_w8_l4096_id0_1_read_size), .S(_maxi_ram_w8_l4096_id0_1_read_start), .Y(_25843_) );
  \$mux  #( .WIDTH(33) ) _48312_ ( .A(_25843_), .B(_maxi_ram_w8_l2048_id2_1_read_size), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_25844_) );
  \$mux  #( .WIDTH(32) ) _48314_ ( .A(_maxi_read_global_addr), .B(_maxi_ram_w32_l128_id0_1_read_global_addr), .S(_maxi_ram_w32_l128_id0_1_read_start), .Y(_25845_) );
  \$mux  #( .WIDTH(32) ) _48315_ ( .A(_25845_), .B(_maxi_ram_w8_l2048_id0_1_read_global_addr), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_25846_) );
  \$mux  #( .WIDTH(32) ) _48316_ ( .A(_25846_), .B(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_global_addr), .S(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_start), .Y(_25847_) );
  \$mux  #( .WIDTH(32) ) _48317_ ( .A(_25847_), .B(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_global_addr), .S(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_start), .Y(_25848_) );
  \$mux  #( .WIDTH(32) ) _48318_ ( .A(_25848_), .B(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_global_addr), .S(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_start), .Y(_25849_) );
  \$mux  #( .WIDTH(32) ) _48319_ ( .A(_25849_), .B(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_global_addr), .S(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_start), .Y(_25850_) );
  \$mux  #( .WIDTH(32) ) _48320_ ( .A(_25850_), .B(_maxi_ram_w8_l2048_id1_1_read_global_addr), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_25851_) );
  \$mux  #( .WIDTH(32) ) _48321_ ( .A(_25851_), .B(_maxi_ram_w8_l4096_id0_1_read_global_addr), .S(_maxi_ram_w8_l4096_id0_1_read_start), .Y(_25852_) );
  \$mux  #( .WIDTH(32) ) _48322_ ( .A(_25852_), .B(_maxi_ram_w8_l2048_id2_1_read_global_addr), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_25853_) );
  \$mux  #( .WIDTH(32) ) _48324_ ( .A(_maxi_read_local_addr), .B(_maxi_ram_w32_l128_id0_1_read_local_addr), .S(_maxi_ram_w32_l128_id0_1_read_start), .Y(_25854_) );
  \$mux  #( .WIDTH(32) ) _48325_ ( .A(_25854_), .B(_maxi_ram_w8_l2048_id0_1_read_local_addr), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_25855_) );
  \$mux  #( .WIDTH(32) ) _48326_ ( .A(_25855_), .B(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_local_addr), .S(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_start), .Y(_25856_) );
  \$mux  #( .WIDTH(32) ) _48327_ ( .A(_25856_), .B(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_local_addr), .S(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_start), .Y(_25857_) );
  \$mux  #( .WIDTH(32) ) _48328_ ( .A(_25857_), .B(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_local_addr), .S(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_start), .Y(_25858_) );
  \$mux  #( .WIDTH(32) ) _48329_ ( .A(_25858_), .B(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_local_addr), .S(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_start), .Y(_25859_) );
  \$mux  #( .WIDTH(32) ) _48330_ ( .A(_25859_), .B(_maxi_ram_w8_l2048_id1_1_read_local_addr), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_25860_) );
  \$mux  #( .WIDTH(32) ) _48331_ ( .A(_25860_), .B(_maxi_ram_w8_l4096_id0_1_read_local_addr), .S(_maxi_ram_w8_l4096_id0_1_read_start), .Y(_25861_) );
  \$mux  #( .WIDTH(32) ) _48332_ ( .A(_25861_), .B(_maxi_ram_w8_l2048_id2_1_read_local_addr), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_25862_) );
  \$mux  #( .WIDTH(8) ) _48334_ ( .A(_maxi_read_op_sel), .B(_maxi_ram_w32_l128_id0_1_read_op_sel), .S(_maxi_ram_w32_l128_id0_1_read_start), .Y(_25863_) );
  \$mux  #( .WIDTH(8) ) _48335_ ( .A(_25863_), .B(_maxi_ram_w8_l2048_id0_1_read_op_sel), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_25864_) );
  \$mux  #( .WIDTH(8) ) _48336_ ( .A(_25864_), .B(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_op_sel), .S(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_start), .Y(_25865_) );
  \$mux  #( .WIDTH(8) ) _48337_ ( .A(_25865_), .B(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_op_sel), .S(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_start), .Y(_25866_) );
  \$mux  #( .WIDTH(8) ) _48338_ ( .A(_25866_), .B(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_op_sel), .S(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_start), .Y(_25867_) );
  \$mux  #( .WIDTH(8) ) _48339_ ( .A(_25867_), .B(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_op_sel), .S(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_start), .Y(_25868_) );
  \$mux  #( .WIDTH(8) ) _48340_ ( .A(_25868_), .B(_maxi_ram_w8_l2048_id1_1_read_op_sel), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_25869_) );
  \$mux  #( .WIDTH(8) ) _48341_ ( .A(_25869_), .B(_maxi_ram_w8_l4096_id0_1_read_op_sel), .S(_maxi_ram_w8_l4096_id0_1_read_start), .Y(_25870_) );
  \$mux  #( .WIDTH(8) ) _48342_ ( .A(_25870_), .B(_maxi_ram_w8_l2048_id2_1_read_op_sel), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_25871_) );
  \$mux  #( .WIDTH(1) ) _48344_ ( .A(1'h0), .B(1'h1), .S(_maxi_ram_w32_l128_id0_1_read_start), .Y(_25872_) );
  \$mux  #( .WIDTH(1) ) _48345_ ( .A(_25872_), .B(1'h1), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_25873_) );
  \$mux  #( .WIDTH(1) ) _48346_ ( .A(_25873_), .B(1'h1), .S(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_start), .Y(_25874_) );
  \$mux  #( .WIDTH(1) ) _48347_ ( .A(_25874_), .B(1'h1), .S(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_start), .Y(_25875_) );
  \$mux  #( .WIDTH(1) ) _48348_ ( .A(_25875_), .B(1'h1), .S(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_start), .Y(_25876_) );
  \$mux  #( .WIDTH(1) ) _48349_ ( .A(_25876_), .B(1'h1), .S(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_start), .Y(_25877_) );
  \$mux  #( .WIDTH(1) ) _48350_ ( .A(_25877_), .B(1'h1), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_25878_) );
  \$mux  #( .WIDTH(1) ) _48351_ ( .A(_25878_), .B(1'h1), .S(_maxi_ram_w8_l4096_id0_1_read_start), .Y(_25879_) );
  \$mux  #( .WIDTH(1) ) _48352_ ( .A(_25879_), .B(1'h1), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_25880_) );
  \$mux  #( .WIDTH(1) ) _48354_ ( .A(maxi_arvalid), .B(1'h0), .S(_saxi_cond_0_1), .Y(_25881_) );
  \$mux  #( .WIDTH(1) ) _48355_ ( .A(_25881_), .B(1'h1), .S(_05268_), .Y(_25882_) );
  \$mux  #( .WIDTH(1) ) _48356_ ( .A(_25882_), .B(maxi_arvalid), .S(_05269_), .Y(_25883_) );
  \$mux  #( .WIDTH(8) ) _48358_ ( .A(maxi_arlen), .B(_25935_[7:0]), .S(_05268_), .Y(_25884_) );
  \$mux  #( .WIDTH(32) ) _48360_ ( .A(maxi_araddr), .B(_maxi_read_cur_global_addr), .S(_05268_), .Y(_25885_) );
  \$mux  #( .WIDTH(1) ) _48362_ ( .A(maxi_wvalid), .B(1'h0), .S(_saxi_cond_0_1), .Y(_25886_) );
  \$mux  #( .WIDTH(1) ) _48363_ ( .A(_25886_), .B(1'h1), .S(_05274_), .Y(_25887_) );
  \$mux  #( .WIDTH(1) ) _48364_ ( .A(_25887_), .B(1'h1), .S(_05277_), .Y(_25888_) );
  \$mux  #( .WIDTH(1) ) _48365_ ( .A(_25888_), .B(1'h1), .S(_05279_), .Y(_25889_) );
  \$mux  #( .WIDTH(1) ) _48366_ ( .A(_25889_), .B(maxi_wvalid), .S(_05276_), .Y(_25890_) );
  \$mux  #( .WIDTH(1) ) _48368_ ( .A(maxi_wlast), .B(1'h0), .S(_saxi_cond_0_1), .Y(_25891_) );
  \$mux  #( .WIDTH(1) ) _48369_ ( .A(_25891_), .B(1'h0), .S(_05274_), .Y(_25892_) );
  \$mux  #( .WIDTH(1) ) _48370_ ( .A(_25892_), .B(1'h1), .S(_05275_), .Y(_25893_) );
  \$mux  #( .WIDTH(1) ) _48371_ ( .A(_25893_), .B(1'h0), .S(_05277_), .Y(_25894_) );
  \$mux  #( .WIDTH(1) ) _48372_ ( .A(_25894_), .B(1'h1), .S(_05278_), .Y(_25895_) );
  \$mux  #( .WIDTH(1) ) _48373_ ( .A(_25895_), .B(1'h0), .S(_05279_), .Y(_25896_) );
  \$mux  #( .WIDTH(1) ) _48374_ ( .A(_25896_), .B(1'h1), .S(_05280_), .Y(_25897_) );
  \$mux  #( .WIDTH(1) ) _48375_ ( .A(_25897_), .B(maxi_wlast), .S(_05276_), .Y(_25898_) );
  \$mux  #( .WIDTH(4) ) _48377_ ( .A(maxi_wstrb), .B(4'hf), .S(_05274_), .Y(_25899_) );
  \$mux  #( .WIDTH(4) ) _48378_ ( .A(_25899_), .B(4'hf), .S(_05277_), .Y(_25900_) );
  \$mux  #( .WIDTH(4) ) _48379_ ( .A(_25900_), .B(4'hf), .S(_05279_), .Y(_25901_) );
  \$mux  #( .WIDTH(32) ) _48381_ ( .A(maxi_wdata), .B(_dataflow_cat_data_74), .S(_05274_), .Y(_25902_) );
  \$mux  #( .WIDTH(32) ) _48382_ ( .A(_25902_), .B(_dataflow_cat_data_96), .S(_05277_), .Y(_25903_) );
  \$mux  #( .WIDTH(32) ) _48383_ ( .A(_25903_), .B(_dataflow_cat_data_131), .S(_05279_), .Y(_25904_) );
  \$mux  #( .WIDTH(1) ) _48385_ ( .A(maxi_awvalid), .B(1'h0), .S(_saxi_cond_0_1), .Y(_25905_) );
  \$mux  #( .WIDTH(1) ) _48386_ ( .A(_25905_), .B(1'h1), .S(_05271_), .Y(_25906_) );
  \$mux  #( .WIDTH(1) ) _48387_ ( .A(_25906_), .B(1'h0), .S(_05272_), .Y(_25907_) );
  \$mux  #( .WIDTH(1) ) _48388_ ( .A(_25907_), .B(maxi_awvalid), .S(_05273_), .Y(_25908_) );
  \$mux  #( .WIDTH(8) ) _48390_ ( .A(maxi_awlen), .B(_25937_[7:0]), .S(_05271_), .Y(_25909_) );
  \$mux  #( .WIDTH(32) ) _48392_ ( .A(maxi_awaddr), .B(_maxi_write_cur_global_addr), .S(_05271_), .Y(_25910_) );
  \$mux  #( .WIDTH(32) ) _48792_ ( .A(_stream_matmul_15_sink_21_sink_fsm_4), .B({ _11374_, _11373_, _11371_, _11370_, _11369_, _11368_, _11367_, _11366_, _11365_, _11364_, _11363_, _11362_, _11360_, _11359_, _11358_, _11357_, _11356_, _11355_, _11354_, _11353_, _11352_, _11351_, _11381_, _11380_, _11379_, _11378_, _11377_, _11376_, _11375_, _11372_, _11361_, _11350_ }), .S(_21881_), .Y(_22456_) );
  \$mux  #( .WIDTH(32) ) _48793_ ( .A(_stream_matmul_15_source_20_source_pat_fsm_3), .B({ _11438_, _11437_, _11435_, _11434_, _11433_, _11432_, _11431_, _11430_, _11429_, _11428_, _11427_, _11426_, _11424_, _11423_, _11422_, _11421_, _11420_, _11419_, _11418_, _11417_, _11416_, _11415_, _11445_, _11444_, _11443_, _11442_, _11441_, _11440_, _11439_, _11436_, _11425_, _11414_ }), .S(_21882_), .Y(_22457_) );
  \$mux  #( .WIDTH(32) ) _48794_ ( .A(_stream_matmul_15_source_19_source_pat_fsm_2), .B({ _11534_, _11533_, _11531_, _11530_, _11529_, _11528_, _11527_, _11526_, _11525_, _11524_, _11523_, _11522_, _11520_, _11519_, _11518_, _11517_, _11516_, _11515_, _11514_, _11513_, _11512_, _11511_, _11541_, _11540_, _11539_, _11538_, _11537_, _11536_, _11535_, _11532_, _11521_, _11510_ }), .S(_21883_), .Y(_22458_) );
  \$mux  #( .WIDTH(32) ) _48795_ ( .A(_stream_matmul_15_source_8_source_pat_fsm_1), .B({ _11630_, _11629_, _11627_, _11626_, _11625_, _11624_, _11623_, _11622_, _11621_, _11620_, _11619_, _11618_, _11616_, _11615_, _11614_, _11613_, _11612_, _11611_, _11610_, _11609_, _11608_, _11607_, _11637_, _11636_, _11635_, _11634_, _11633_, _11632_, _11631_, _11628_, _11617_, _11606_ }), .S(_21884_), .Y(_22459_) );
  \$mux  #( .WIDTH(32) ) _48796_ ( .A(_stream_matmul_15_source_6_source_pat_fsm_0), .B({ _11726_, _11725_, _11723_, _11722_, _11721_, _11720_, _11719_, _11718_, _11717_, _11716_, _11715_, _11714_, _11712_, _11711_, _11710_, _11709_, _11708_, _11707_, _11706_, _11705_, _11704_, _11703_, _11733_, _11732_, _11731_, _11730_, _11729_, _11728_, _11727_, _11724_, _11713_, _11702_ }), .S(_21885_), .Y(_22460_) );
  \$mux  #( .WIDTH(32) ) _48797_ ( .A(matmul_15_comp_fsm), .B({ _11822_, _11821_, _11819_, _11818_, _11817_, _11816_, _11815_, _11814_, _11813_, _11812_, _11811_, _11810_, _11808_, _11807_, _11806_, _11805_, _11804_, _11803_, _11802_, _11801_, _11800_, _11799_, _11829_, _11828_, _11827_, _11826_, _11825_, _11824_, _11823_, _11820_, _11809_, _11798_ }), .S(_21886_), .Y(_22468_) );
  \$mux  #( .WIDTH(32) ) _48798_ ( .A(matmul_15_stream_out_local_col), .B(0), .S(_21887_), .Y(_22469_) );
  \$mux  #( .WIDTH(32) ) _48799_ ( .A(matmul_15_stream_act_local_0), .B(0), .S(_21887_), .Y(_22470_) );
  \$mux  #( .WIDTH(1) ) _48800_ ( .A(matmul_15_col_select), .B(1'h0), .S(_21887_), .Y(_22471_) );
  \$mux  #( .WIDTH(32) ) _48801_ ( .A(matmul_15_col_count), .B(0), .S(_21887_), .Y(_22472_) );
  \$mux  #( .WIDTH(1) ) _48802_ ( .A(matmul_15_skip_write_out), .B(_11895_), .S(_04701_), .Y(_22496_) );
  \$mux  #( .WIDTH(1) ) _48803_ ( .A(matmul_15_skip_comp), .B(_11898_), .S(_04701_), .Y(_22497_) );
  \$mux  #( .WIDTH(1) ) _48804_ ( .A(matmul_15_skip_read_act), .B(_11896_), .S(_04701_), .Y(_22498_) );
  \$mux  #( .WIDTH(1) ) _48805_ ( .A(matmul_15_skip_read_filter), .B(_11900_), .S(_04701_), .Y(_22499_) );
  \$mux  #( .WIDTH(32) ) _48806_ ( .A(matmul_15_out_laddr_offset), .B({ _04829_, _04828_, _04825_, _04827_, _04826_, _04824_, _04819_, _04823_, _04822_, _04821_, _04817_, _04820_, _04818_, _04816_, _04811_, _04815_, _04814_, _04813_, _04809_, _04812_, _04810_, _04808_, _04803_, _04807_, _04806_, _04805_, _04801_, _04804_, _04802_, _04800_, _04798_, _04799_ }), .S(_21888_), .Y(_22500_) );
  \$mux  #( .WIDTH(32) ) _48807_ ( .A(matmul_15_out_page_dma_offset), .B({ _12021_, _12020_, _12018_, _12017_, _12016_, _12015_, _12014_, _12013_, _12012_, _12011_, _12010_, _12009_, _12007_, _12006_, _12005_, _12004_, _12003_, _12002_, _12001_, _12000_, _11999_, _11998_, _12028_, _12027_, _12026_, _12025_, _12024_, _12023_, _12022_, _12019_, _12008_, _11997_ }), .S(_04701_), .Y(_22501_) );
  \$mux  #( .WIDTH(32) ) _48808_ ( .A(matmul_15_out_page_comp_offset), .B({ _12085_, _12084_, _12082_, _12081_, _12080_, _12079_, _12078_, _12077_, _12076_, _12075_, _12074_, _12073_, _12071_, _12070_, _12069_, _12068_, _12067_, _12066_, _12065_, _12064_, _12063_, _12062_, _12092_, _12091_, _12090_, _12089_, _12088_, _12087_, _12086_, _12083_, _12072_, _12061_ }), .S(_04701_), .Y(_22502_) );
  \$mux  #( .WIDTH(1) ) _48809_ ( .A(matmul_15_out_page), .B(_12094_), .S(_04701_), .Y(_22503_) );
  \$mux  #( .WIDTH(32) ) _48810_ ( .A(matmul_15_filter_page_dma_offset), .B({ _12151_, _12150_, _12148_, _12147_, _12146_, _12145_, _12144_, _12143_, _12142_, _12141_, _12140_, _12139_, _12137_, _12136_, _12135_, _12134_, _12133_, _12132_, _12131_, _12130_, _12129_, _12128_, _12158_, _12157_, _12156_, _12155_, _12154_, _12153_, _12152_, _12149_, _12138_, _12127_ }), .S(_04701_), .Y(_22504_) );
  \$mux  #( .WIDTH(32) ) _48811_ ( .A(matmul_15_filter_page_comp_offset), .B({ _12215_, _12214_, _12212_, _12211_, _12210_, _12209_, _12208_, _12207_, _12206_, _12205_, _12204_, _12203_, _12201_, _12200_, _12199_, _12198_, _12197_, _12196_, _12195_, _12194_, _12193_, _12192_, _12222_, _12221_, _12220_, _12219_, _12218_, _12217_, _12216_, _12213_, _12202_, _12191_ }), .S(_04701_), .Y(_22505_) );
  \$mux  #( .WIDTH(32) ) _48812_ ( .A(matmul_15_act_page_dma_offset_0), .B(0), .S(_04701_), .Y(_22506_) );
  \$mux  #( .WIDTH(32) ) _48813_ ( .A(matmul_15_act_page_comp_offset_0), .B(0), .S(_04701_), .Y(_22507_) );
  \$mux  #( .WIDTH(32) ) _48814_ ( .A(matmul_15_prev_och_count), .B({ _12247_, _12246_, _12244_, _12243_, _12242_, _12241_, _12240_, _12239_, _12238_, _12237_, _12236_, _12235_, _12233_, _12232_, _12231_, _12230_, _12229_, _12228_, _12227_, _12226_, _12225_, _12224_, _12254_, _12253_, _12252_, _12251_, _12250_, _12249_, _12248_, _12245_, _12234_, _12223_ }), .S(_04701_), .Y(_22509_) );
  \$mux  #( .WIDTH(32) ) _48815_ ( .A(matmul_15_prev_bat_count), .B({ _12279_, _12278_, _12276_, _12275_, _12274_, _12273_, _12272_, _12271_, _12270_, _12269_, _12268_, _12267_, _12265_, _12264_, _12263_, _12262_, _12261_, _12260_, _12259_, _12258_, _12257_, _12256_, _12286_, _12285_, _12284_, _12283_, _12282_, _12281_, _12280_, _12277_, _12266_, _12255_ }), .S(_04701_), .Y(_22510_) );
  \$mux  #( .WIDTH(32) ) _48816_ ( .A(matmul_15_prev_row_count), .B({ _12311_, _12310_, _12308_, _12307_, _12306_, _12305_, _12304_, _12303_, _12302_, _12301_, _12300_, _12299_, _12297_, _12296_, _12295_, _12294_, _12293_, _12292_, _12291_, _12290_, _12289_, _12288_, _12318_, _12317_, _12316_, _12315_, _12314_, _12313_, _12312_, _12309_, _12298_, _12287_ }), .S(_04701_), .Y(_22511_) );
  \$mux  #( .WIDTH(32) ) _48817_ ( .A(matmul_15_out_ram_select), .B({ _04765_, _04764_, _04763_, _04762_, _04761_, _04760_, _04759_, _04758_, _04757_, _04756_, _04755_, _04754_, _04753_, _04752_, _04751_, _04750_, _04749_, _04748_, _04747_, _04746_, _04745_, _04744_, _04743_, _04742_, _04741_, _04740_, _04739_, _04738_, _04737_, _04736_, _04735_, _04734_ }), .S(_21888_), .Y(_22512_) );
  \$mux  #( .WIDTH(32) ) _48818_ ( .A(matmul_15_out_row_count), .B({ _12439_, _12438_, _12436_, _12435_, _12434_, _12433_, _12432_, _12431_, _12430_, _12429_, _12428_, _12427_, _12425_, _12424_, _12423_, _12422_, _12421_, _12420_, _12419_, _12418_, _12417_, _12416_, _12446_, _12445_, _12444_, _12443_, _12442_, _12441_, _12440_, _12437_, _12426_, _12415_ }), .S(_04701_), .Y(_22513_) );
  \$mux  #( .WIDTH(32) ) _48819_ ( .A(matmul_15_och_count), .B({ _12471_, _12470_, _12468_, _12467_, _12466_, _12465_, _12464_, _12463_, _12462_, _12461_, _12460_, _12459_, _12457_, _12456_, _12455_, _12454_, _12453_, _12452_, _12451_, _12450_, _12449_, _12448_, _12478_, _12477_, _12476_, _12475_, _12474_, _12473_, _12472_, _12469_, _12458_, _12447_ }), .S(_04701_), .Y(_22515_) );
  \$mux  #( .WIDTH(32) ) _48820_ ( .A(matmul_15_bat_count), .B(0), .S(_04701_), .Y(_22516_) );
  \$mux  #( .WIDTH(32) ) _48821_ ( .A(matmul_15_row_count), .B(0), .S(_04701_), .Y(_22517_) );
  \$mux  #( .WIDTH(32) ) _48822_ ( .A(matmul_15_sync_out_count), .B({ _12535_, _12534_, _12532_, _12531_, _12530_, _12529_, _12528_, _12527_, _12526_, _12525_, _12524_, _12523_, _12521_, _12520_, _12519_, _12518_, _12517_, _12516_, _12515_, _12514_, _12513_, _12512_, _12542_, _12541_, _12540_, _12539_, _12538_, _12537_, _12536_, _12533_, _12522_, _12511_ }), .S(_21889_), .Y(_22519_) );
  \$mux  #( .WIDTH(32) ) _48823_ ( .A(matmul_15_out_base_offset_och), .B({ _12599_, _12598_, _12596_, _12595_, _12594_, _12593_, _12592_, _12591_, _12590_, _12589_, _12588_, _12587_, _12585_, _12584_, _12583_, _12582_, _12581_, _12580_, _12579_, _12578_, _12577_, _12576_, _12606_, _12605_, _12604_, _12603_, _12602_, _12601_, _12600_, _12597_, _12586_, _12575_ }), .S(_04701_), .Y(_22521_) );
  \$mux  #( .WIDTH(32) ) _48824_ ( .A(matmul_15_out_base_offset_bat), .B({ _12663_, _12662_, _12660_, _12659_, _12658_, _12657_, _12656_, _12655_, _12654_, _12653_, _12652_, _12651_, _12649_, _12648_, _12647_, _12646_, _12645_, _12644_, _12643_, _12642_, _12641_, _12640_, _12670_, _12669_, _12668_, _12667_, _12666_, _12665_, _12664_, _12661_, _12650_, _12639_ }), .S(_04701_), .Y(_22522_) );
  \$mux  #( .WIDTH(32) ) _48825_ ( .A(matmul_15_out_base_offset_row), .B({ _12727_, _12726_, _12724_, _12723_, _12722_, _12721_, _12720_, _12719_, _12718_, _12717_, _12716_, _12715_, _12713_, _12712_, _12711_, _12710_, _12709_, _12708_, _12707_, _12706_, _12705_, _12704_, _12734_, _12733_, _12732_, _12731_, _12730_, _12729_, _12728_, _12725_, _12714_, _12703_ }), .S(_04701_), .Y(_22523_) );
  \$mux  #( .WIDTH(32) ) _48826_ ( .A(matmul_15_out_base_offset_col), .B({ _04733_, _04730_, _04732_, _04728_, _04731_, _04729_, _04726_, _04727_, _04723_, _04725_, _04724_, _04722_, _04716_, _04721_, _04720_, _04712_, _04719_, _04718_, _04717_, _04710_, _04715_, _04714_, _04713_, _04711_, _04709_, _04708_, _04707_, _04706_, _04702_, _04705_, _04704_, _04703_ }), .S(_21888_), .Y(_22524_) );
  \$mux  #( .WIDTH(32) ) _48827_ ( .A(matmul_15_filter_base_offset), .B({ _12791_, _12790_, _12788_, _12787_, _12786_, _12785_, _12784_, _12783_, _12782_, _12781_, _12780_, _12779_, _12777_, _12776_, _12775_, _12774_, _12773_, _12772_, _12771_, _12770_, _12769_, _12768_, _12798_, _12797_, _12796_, _12795_, _12794_, _12793_, _12792_, _12789_, _12778_, _12767_ }), .S(_04701_), .Y(_22526_) );
  \$mux  #( .WIDTH(32) ) _48828_ ( .A(matmul_15_act_base_offset_bat), .B(0), .S(_04701_), .Y(_22527_) );
  \$mux  #( .WIDTH(32) ) _48829_ ( .A(matmul_15_act_base_offset_row), .B(0), .S(_04701_), .Y(_22528_) );
  \$mux  #( .WIDTH(32) ) _48830_ ( .A(control_matmul_15), .B({ _12855_, _12854_, _12852_, _12851_, _12850_, _12849_, _12848_, _12847_, _12846_, _12845_, _12844_, _12843_, _12841_, _12840_, _12839_, _12838_, _12837_, _12836_, _12835_, _12834_, _12833_, _12832_, _12862_, _12861_, _12860_, _12859_, _12858_, _12857_, _12856_, _12853_, _12842_, _12831_ }), .S(_21890_), .Y(_22529_) );
  \$mux  #( .WIDTH(32) ) _48831_ ( .A(_stream_max_pool_serial_9_sink_3_sink_fsm_1), .B({ _13431_, _13430_, _13428_, _13427_, _13426_, _13425_, _13424_, _13423_, _13422_, _13421_, _13420_, _13419_, _13417_, _13416_, _13415_, _13414_, _13413_, _13412_, _13411_, _13410_, _13409_, _13408_, _13438_, _13437_, _13436_, _13435_, _13434_, _13433_, _13432_, _13429_, _13418_, _13407_ }), .S(_21891_), .Y(_22534_) );
  \$mux  #( .WIDTH(32) ) _48832_ ( .A(_stream_max_pool_serial_9_source_1_source_pat_fsm_0), .B({ _13495_, _13494_, _13492_, _13491_, _13490_, _13489_, _13488_, _13487_, _13486_, _13485_, _13484_, _13483_, _13481_, _13480_, _13479_, _13478_, _13477_, _13476_, _13475_, _13474_, _13473_, _13472_, _13502_, _13501_, _13500_, _13499_, _13498_, _13497_, _13496_, _13493_, _13482_, _13471_ }), .S(_21892_), .Y(_22535_) );
  \$mux  #( .WIDTH(32) ) _48833_ ( .A(max_pool_serial_9_comp_fsm), .B({ _13623_, _13622_, _13620_, _13619_, _13618_, _13617_, _13616_, _13615_, _13614_, _13613_, _13612_, _13611_, _13609_, _13608_, _13607_, _13606_, _13605_, _13604_, _13603_, _13602_, _13601_, _13600_, _13630_, _13629_, _13628_, _13627_, _13626_, _13625_, _13624_, _13621_, _13610_, _13599_ }), .S(_21893_), .Y(_22540_) );
  \$mux  #( .WIDTH(32) ) _48834_ ( .A(max_pool_serial_9_stream_out_local), .B({ _13751_, _13750_, _13748_, _13747_, _13746_, _13745_, _13744_, _13743_, _13742_, _13741_, _13740_, _13739_, _13737_, _13736_, _13735_, _13734_, _13733_, _13732_, _13731_, _13730_, _13729_, _13728_, _13758_, _13757_, _13756_, _13755_, _13754_, _13753_, _13752_, _13749_, _13738_, _13727_ }), .S(_21894_), .Y(_22543_) );
  \$mux  #( .WIDTH(32) ) _48835_ ( .A(max_pool_serial_9_stream_act_local), .B({ _13815_, _13814_, _13812_, _13811_, _13810_, _13809_, _13808_, _13807_, _13806_, _13805_, _13804_, _13803_, _13801_, _13800_, _13799_, _13798_, _13797_, _13796_, _13795_, _13794_, _13793_, _13792_, _13822_, _13821_, _13820_, _13819_, _13818_, _13817_, _13816_, _13813_, _13802_, _13791_ }), .S(_21894_), .Y(_22544_) );
  \$mux  #( .WIDTH(32) ) _48836_ ( .A(max_pool_serial_9_col_count), .B({ _13879_, _13878_, _13876_, _13875_, _13874_, _13873_, _13872_, _13871_, _13870_, _13869_, _13868_, _13867_, _13865_, _13864_, _13863_, _13862_, _13861_, _13860_, _13859_, _13858_, _13857_, _13856_, _13886_, _13885_, _13884_, _13883_, _13882_, _13881_, _13880_, _13877_, _13866_, _13855_ }), .S(_21894_), .Y(_22545_) );
  \$mux  #( .WIDTH(32) ) _48837_ ( .A(max_pool_serial_9_out_count), .B({ _13911_, _13910_, _13908_, _13907_, _13906_, _13905_, _13904_, _13903_, _13902_, _13901_, _13900_, _13899_, _13897_, _13896_, _13895_, _13894_, _13893_, _13892_, _13891_, _13890_, _13889_, _13888_, _13918_, _13917_, _13916_, _13915_, _13914_, _13913_, _13912_, _13909_, _13898_, _13887_ }), .S(_21895_), .Y(_22558_) );
  \$mux  #( .WIDTH(1) ) _48838_ ( .A(max_pool_serial_9_skip_write_out), .B(_13920_), .S(_21896_), .Y(_22559_) );
  \$mux  #( .WIDTH(1) ) _48839_ ( .A(max_pool_serial_9_skip_comp), .B(_13922_), .S(_21896_), .Y(_22560_) );
  \$mux  #( .WIDTH(1) ) _48840_ ( .A(max_pool_serial_9_skip_read_act), .B(_13924_), .S(_21896_), .Y(_22561_) );
  \$mux  #( .WIDTH(32) ) _48841_ ( .A(max_pool_serial_9_out_page_dma_offset), .B({ _13981_, _13980_, _13978_, _13977_, _13976_, _13975_, _13974_, _13973_, _13972_, _13971_, _13970_, _13969_, _13967_, _13966_, _13965_, _13964_, _13963_, _13962_, _13961_, _13960_, _13959_, _13958_, _13988_, _13987_, _13986_, _13985_, _13984_, _13983_, _13982_, _13979_, _13968_, _13957_ }), .S(_21896_), .Y(_22562_) );
  \$mux  #( .WIDTH(32) ) _48842_ ( .A(max_pool_serial_9_out_page_comp_offset), .B({ _14045_, _14044_, _14042_, _14041_, _14040_, _14039_, _14038_, _14037_, _14036_, _14035_, _14034_, _14033_, _14031_, _14030_, _14029_, _14028_, _14027_, _14026_, _14025_, _14024_, _14023_, _14022_, _14052_, _14051_, _14050_, _14049_, _14048_, _14047_, _14046_, _14043_, _14032_, _14021_ }), .S(_21896_), .Y(_22563_) );
  \$mux  #( .WIDTH(1) ) _48843_ ( .A(max_pool_serial_9_out_page), .B(_14054_), .S(_21896_), .Y(_22564_) );
  \$mux  #( .WIDTH(32) ) _48844_ ( .A(max_pool_serial_9_act_page_dma_offset), .B({ _14111_, _14110_, _14108_, _14107_, _14106_, _14105_, _14104_, _14103_, _14102_, _14101_, _14100_, _14099_, _14097_, _14096_, _14095_, _14094_, _14093_, _14092_, _14091_, _14090_, _14089_, _14088_, _14118_, _14117_, _14116_, _14115_, _14114_, _14113_, _14112_, _14109_, _14098_, _14087_ }), .S(_21896_), .Y(_22565_) );
  \$mux  #( .WIDTH(32) ) _48845_ ( .A(max_pool_serial_9_act_page_comp_offset), .B({ _14111_, _14110_, _14108_, _14107_, _14106_, _14105_, _14104_, _14103_, _14102_, _14101_, _14100_, _14099_, _14097_, _14096_, _14095_, _14094_, _14093_, _14092_, _14091_, _14090_, _14089_, _14088_, _14118_, _14117_, _14116_, _14115_, _14114_, _14113_, _14112_, _14109_, _14098_, _14087_ }), .S(_21896_), .Y(_22566_) );
  \$mux  #( .WIDTH(1) ) _48846_ ( .A(max_pool_serial_9_act_page), .B(_14120_), .S(_21896_), .Y(_22567_) );
  \$mux  #( .WIDTH(32) ) _48847_ ( .A(max_pool_serial_9_prev_bat_count), .B({ _14145_, _14144_, _14142_, _14141_, _14140_, _14139_, _14138_, _14137_, _14136_, _14135_, _14134_, _14133_, _14131_, _14130_, _14129_, _14128_, _14127_, _14126_, _14125_, _14124_, _14123_, _14122_, _14152_, _14151_, _14150_, _14149_, _14148_, _14147_, _14146_, _14143_, _14132_, _14121_ }), .S(_21896_), .Y(_22568_) );
  \$mux  #( .WIDTH(32) ) _48848_ ( .A(max_pool_serial_9_prev_row_count), .B({ _14177_, _14176_, _14174_, _14173_, _14172_, _14171_, _14170_, _14169_, _14168_, _14167_, _14166_, _14165_, _14163_, _14162_, _14161_, _14160_, _14159_, _14158_, _14157_, _14156_, _14155_, _14154_, _14184_, _14183_, _14182_, _14181_, _14180_, _14179_, _14178_, _14175_, _14164_, _14153_ }), .S(_21896_), .Y(_22569_) );
  \$mux  #( .WIDTH(32) ) _48849_ ( .A(max_pool_serial_9_bat_count), .B({ _14241_, _14240_, _14238_, _14237_, _14236_, _14235_, _14234_, _14233_, _14232_, _14231_, _14230_, _14229_, _14227_, _14226_, _14225_, _14224_, _14223_, _14222_, _14221_, _14220_, _14219_, _14218_, _14248_, _14247_, _14246_, _14245_, _14244_, _14243_, _14242_, _14239_, _14228_, _14217_ }), .S(_21896_), .Y(_22570_) );
  \$mux  #( .WIDTH(32) ) _48850_ ( .A(max_pool_serial_9_row_count), .B({ _14305_, _14304_, _14302_, _14301_, _14300_, _14299_, _14298_, _14297_, _14296_, _14295_, _14294_, _14293_, _14291_, _14290_, _14289_, _14288_, _14287_, _14286_, _14285_, _14284_, _14283_, _14282_, _14312_, _14311_, _14310_, _14309_, _14308_, _14307_, _14306_, _14303_, _14292_, _14281_ }), .S(_21896_), .Y(_22571_) );
  \$mux  #( .WIDTH(32) ) _48851_ ( .A(max_pool_serial_9_out_base_offset_bat), .B({ _14369_, _14368_, _14366_, _14365_, _14364_, _14363_, _14362_, _14361_, _14360_, _14359_, _14358_, _14357_, _14355_, _14354_, _14353_, _14352_, _14351_, _14350_, _14349_, _14348_, _14347_, _14346_, _14376_, _14375_, _14374_, _14373_, _14372_, _14371_, _14370_, _14367_, _14356_, _14345_ }), .S(_21896_), .Y(_22572_) );
  \$mux  #( .WIDTH(32) ) _48852_ ( .A(max_pool_serial_9_out_base_offset_row), .B({ _14433_, _14432_, _14430_, _14429_, _14428_, _14427_, _14426_, _14425_, _14424_, _14423_, _14422_, _14421_, _14419_, _14418_, _14417_, _14416_, _14415_, _14414_, _14413_, _14412_, _14411_, _14410_, _14440_, _14439_, _14438_, _14437_, _14436_, _14435_, _14434_, _14431_, _14420_, _14409_ }), .S(_21896_), .Y(_22574_) );
  \$mux  #( .WIDTH(32) ) _48853_ ( .A(max_pool_serial_9_act_base_offset_bat), .B({ _14497_, _14496_, _14494_, _14493_, _14492_, _14491_, _14490_, _14489_, _14488_, _14487_, _14486_, _14485_, _14483_, _14482_, _14481_, _14480_, _14479_, _14478_, _14477_, _14476_, _14475_, _14474_, _14504_, _14503_, _14502_, _14501_, _14500_, _14499_, _14498_, _14495_, _14484_, _14473_ }), .S(_21896_), .Y(_22575_) );
  \$mux  #( .WIDTH(32) ) _48854_ ( .A(max_pool_serial_9_act_base_offset_row), .B({ _14561_, _14560_, _14558_, _14557_, _14556_, _14555_, _14554_, _14553_, _14552_, _14551_, _14550_, _14549_, _14547_, _14546_, _14545_, _14544_, _14543_, _14542_, _14541_, _14540_, _14539_, _14538_, _14568_, _14567_, _14566_, _14565_, _14564_, _14563_, _14562_, _14559_, _14548_, _14537_ }), .S(_21896_), .Y(_22576_) );
  \$mux  #( .WIDTH(32) ) _48855_ ( .A(control_max_pool_serial_9), .B({ _14625_, _14624_, _14622_, _14621_, _14620_, _14619_, _14618_, _14617_, _14616_, _14615_, _14614_, _14613_, _14611_, _14610_, _14609_, _14608_, _14607_, _14606_, _14605_, _14604_, _14603_, _14602_, _14632_, _14631_, _14630_, _14629_, _14628_, _14627_, _14626_, _14623_, _14612_, _14601_ }), .S(_21897_), .Y(_22578_) );
  \$mux  #( .WIDTH(33) ) _48856_ ( .A(_maxi_write_rest_size), .B({ _15075_, _15074_, _15073_, _15071_, _15070_, _15069_, _15068_, _15067_, _15066_, _15065_, _15064_, _15063_, _15062_, _15060_, _15059_, _15058_, _15057_, _15056_, _15055_, _15054_, _15053_, _15052_, _15051_, _15082_, _15081_, _15080_, _15079_, _15078_, _15077_, _15076_, _15072_, _15061_, _15050_ }), .S(_04832_), .Y(_22588_) );
  \$mux  #( .WIDTH(32) ) _48857_ ( .A(_maxi_write_cur_global_addr), .B({ _15172_, _15171_, _15169_, _15168_, _15167_, _15166_, _15165_, _15164_, _15163_, _15162_, _15161_, _15160_, _15158_, _15157_, _15156_, _15155_, _15154_, _15153_, _15152_, _15151_, _15150_, _15149_, _15179_, _15178_, _15177_, _15176_, _15175_, _15174_, _15173_, _15170_, _15159_, _15148_ }), .S(_21898_), .Y(_22593_) );
  \$mux  #( .WIDTH(32) ) _48858_ ( .A(_maxi_write_fsm), .B({ _15236_, _15235_, _15233_, _15232_, _15231_, _15230_, _15229_, _15228_, _15227_, _15226_, _15225_, _15224_, _15222_, _15221_, _15220_, _15219_, _15218_, _15217_, _15216_, _15215_, _15214_, _15213_, _15243_, _15242_, _15241_, _15240_, _15239_, _15238_, _15237_, _15234_, _15223_, _15212_ }), .S(_21899_), .Y(_22594_) );
  \$mux  #( .WIDTH(32) ) _48859_ ( .A(_stream_conv2d_8_sink_37_sink_fsm_20), .B({ _15396_, _15395_, _15393_, _15392_, _15391_, _15390_, _15389_, _15388_, _15387_, _15386_, _15385_, _15384_, _15382_, _15381_, _15380_, _15379_, _15378_, _15377_, _15376_, _15375_, _15374_, _15373_, _15403_, _15402_, _15401_, _15400_, _15399_, _15398_, _15397_, _15394_, _15383_, _15372_ }), .S(_21900_), .Y(_22599_) );
  \$mux  #( .WIDTH(32) ) _48860_ ( .A(_stream_conv2d_8_source_36_source_pat_fsm_19), .B({ _15460_, _15459_, _15457_, _15456_, _15455_, _15454_, _15453_, _15452_, _15451_, _15450_, _15449_, _15448_, _15446_, _15445_, _15444_, _15443_, _15442_, _15441_, _15440_, _15439_, _15438_, _15437_, _15467_, _15466_, _15465_, _15464_, _15463_, _15462_, _15461_, _15458_, _15447_, _15436_ }), .S(_21901_), .Y(_22600_) );
  \$mux  #( .WIDTH(32) ) _48861_ ( .A(_stream_conv2d_8_source_35_source_pat_fsm_18), .B({ _15556_, _15555_, _15553_, _15552_, _15551_, _15550_, _15549_, _15548_, _15547_, _15546_, _15545_, _15544_, _15542_, _15541_, _15540_, _15539_, _15538_, _15537_, _15536_, _15535_, _15534_, _15533_, _15563_, _15562_, _15561_, _15560_, _15559_, _15558_, _15557_, _15554_, _15543_, _15532_ }), .S(_21902_), .Y(_22601_) );
  \$mux  #( .WIDTH(32) ) _48862_ ( .A(_stream_conv2d_8_source_34_source_pat_fsm_17), .B({ _15652_, _15651_, _15649_, _15648_, _15647_, _15646_, _15645_, _15644_, _15643_, _15642_, _15641_, _15640_, _15638_, _15637_, _15636_, _15635_, _15634_, _15633_, _15632_, _15631_, _15630_, _15629_, _15659_, _15658_, _15657_, _15656_, _15655_, _15654_, _15653_, _15650_, _15639_, _15628_ }), .S(_21903_), .Y(_22602_) );
  \$mux  #( .WIDTH(32) ) _48863_ ( .A(_stream_conv2d_8_source_33_source_pat_fsm_16), .B({ _15748_, _15747_, _15745_, _15744_, _15743_, _15742_, _15741_, _15740_, _15739_, _15738_, _15737_, _15736_, _15734_, _15733_, _15732_, _15731_, _15730_, _15729_, _15728_, _15727_, _15726_, _15725_, _15755_, _15754_, _15753_, _15752_, _15751_, _15750_, _15749_, _15746_, _15735_, _15724_ }), .S(_21904_), .Y(_22603_) );
  \$mux  #( .WIDTH(32) ) _48864_ ( .A(_stream_conv2d_8_source_32_source_pat_fsm_15), .B({ _15844_, _15843_, _15841_, _15840_, _15839_, _15838_, _15837_, _15836_, _15835_, _15834_, _15833_, _15832_, _15830_, _15829_, _15828_, _15827_, _15826_, _15825_, _15824_, _15823_, _15822_, _15821_, _15851_, _15850_, _15849_, _15848_, _15847_, _15846_, _15845_, _15842_, _15831_, _15820_ }), .S(_21905_), .Y(_22604_) );
  \$mux  #( .WIDTH(32) ) _48865_ ( .A(_stream_conv2d_8_source_31_source_pat_fsm_14), .B({ _15940_, _15939_, _15937_, _15936_, _15935_, _15934_, _15933_, _15932_, _15931_, _15930_, _15929_, _15928_, _15926_, _15925_, _15924_, _15923_, _15922_, _15921_, _15920_, _15919_, _15918_, _15917_, _15947_, _15946_, _15945_, _15944_, _15943_, _15942_, _15941_, _15938_, _15927_, _15916_ }), .S(_21906_), .Y(_22605_) );
  \$mux  #( .WIDTH(32) ) _48866_ ( .A(_stream_conv2d_8_source_30_source_pat_fsm_13), .B({ _16036_, _16035_, _16033_, _16032_, _16031_, _16030_, _16029_, _16028_, _16027_, _16026_, _16025_, _16024_, _16022_, _16021_, _16020_, _16019_, _16018_, _16017_, _16016_, _16015_, _16014_, _16013_, _16043_, _16042_, _16041_, _16040_, _16039_, _16038_, _16037_, _16034_, _16023_, _16012_ }), .S(_21907_), .Y(_22606_) );
  \$mux  #( .WIDTH(32) ) _48867_ ( .A(_stream_conv2d_8_source_29_source_pat_fsm_12), .B({ _16132_, _16131_, _16129_, _16128_, _16127_, _16126_, _16125_, _16124_, _16123_, _16122_, _16121_, _16120_, _16118_, _16117_, _16116_, _16115_, _16114_, _16113_, _16112_, _16111_, _16110_, _16109_, _16139_, _16138_, _16137_, _16136_, _16135_, _16134_, _16133_, _16130_, _16119_, _16108_ }), .S(_21908_), .Y(_22607_) );
  \$mux  #( .WIDTH(32) ) _48868_ ( .A(_stream_conv2d_8_source_28_source_pat_fsm_11), .B({ _16228_, _16227_, _16225_, _16224_, _16223_, _16222_, _16221_, _16220_, _16219_, _16218_, _16217_, _16216_, _16214_, _16213_, _16212_, _16211_, _16210_, _16209_, _16208_, _16207_, _16206_, _16205_, _16235_, _16234_, _16233_, _16232_, _16231_, _16230_, _16229_, _16226_, _16215_, _16204_ }), .S(_21909_), .Y(_22608_) );
  \$mux  #( .WIDTH(32) ) _48869_ ( .A(_stream_conv2d_8_source_27_source_pat_fsm_10), .B({ _16324_, _16323_, _16321_, _16320_, _16319_, _16318_, _16317_, _16316_, _16315_, _16314_, _16313_, _16312_, _16310_, _16309_, _16308_, _16307_, _16306_, _16305_, _16304_, _16303_, _16302_, _16301_, _16331_, _16330_, _16329_, _16328_, _16327_, _16326_, _16325_, _16322_, _16311_, _16300_ }), .S(_21910_), .Y(_22609_) );
  \$mux  #( .WIDTH(32) ) _48870_ ( .A(_stream_conv2d_8_source_26_source_pat_fsm_9), .B({ _16420_, _16419_, _16417_, _16416_, _16415_, _16414_, _16413_, _16412_, _16411_, _16410_, _16409_, _16408_, _16406_, _16405_, _16404_, _16403_, _16402_, _16401_, _16400_, _16399_, _16398_, _16397_, _16427_, _16426_, _16425_, _16424_, _16423_, _16422_, _16421_, _16418_, _16407_, _16396_ }), .S(_21911_), .Y(_22610_) );
  \$mux  #( .WIDTH(32) ) _48871_ ( .A(_stream_conv2d_8_source_25_source_pat_fsm_8), .B({ _16516_, _16515_, _16513_, _16512_, _16511_, _16510_, _16509_, _16508_, _16507_, _16506_, _16505_, _16504_, _16502_, _16501_, _16500_, _16499_, _16498_, _16497_, _16496_, _16495_, _16494_, _16493_, _16523_, _16522_, _16521_, _16520_, _16519_, _16518_, _16517_, _16514_, _16503_, _16492_ }), .S(_21912_), .Y(_22611_) );
  \$mux  #( .WIDTH(32) ) _48872_ ( .A(_stream_conv2d_8_source_24_source_pat_fsm_7), .B({ _16612_, _16611_, _16609_, _16608_, _16607_, _16606_, _16605_, _16604_, _16603_, _16602_, _16601_, _16600_, _16598_, _16597_, _16596_, _16595_, _16594_, _16593_, _16592_, _16591_, _16590_, _16589_, _16619_, _16618_, _16617_, _16616_, _16615_, _16614_, _16613_, _16610_, _16599_, _16588_ }), .S(_21913_), .Y(_22612_) );
  \$mux  #( .WIDTH(32) ) _48873_ ( .A(_stream_conv2d_8_source_23_source_pat_fsm_6), .B({ _16708_, _16707_, _16705_, _16704_, _16703_, _16702_, _16701_, _16700_, _16699_, _16698_, _16697_, _16696_, _16694_, _16693_, _16692_, _16691_, _16690_, _16689_, _16688_, _16687_, _16686_, _16685_, _16715_, _16714_, _16713_, _16712_, _16711_, _16710_, _16709_, _16706_, _16695_, _16684_ }), .S(_21914_), .Y(_22613_) );
  \$mux  #( .WIDTH(32) ) _48874_ ( .A(_stream_conv2d_8_source_22_source_pat_fsm_5), .B({ _16804_, _16803_, _16801_, _16800_, _16799_, _16798_, _16797_, _16796_, _16795_, _16794_, _16793_, _16792_, _16790_, _16789_, _16788_, _16787_, _16786_, _16785_, _16784_, _16783_, _16782_, _16781_, _16811_, _16810_, _16809_, _16808_, _16807_, _16806_, _16805_, _16802_, _16791_, _16780_ }), .S(_21915_), .Y(_22614_) );
  \$mux  #( .WIDTH(32) ) _48875_ ( .A(_stream_conv2d_8_source_21_source_pat_fsm_4), .B({ _16900_, _16899_, _16897_, _16896_, _16895_, _16894_, _16893_, _16892_, _16891_, _16890_, _16889_, _16888_, _16886_, _16885_, _16884_, _16883_, _16882_, _16881_, _16880_, _16879_, _16878_, _16877_, _16907_, _16906_, _16905_, _16904_, _16903_, _16902_, _16901_, _16898_, _16887_, _16876_ }), .S(_21916_), .Y(_22615_) );
  \$mux  #( .WIDTH(32) ) _48876_ ( .A(_stream_conv2d_8_source_20_source_pat_fsm_3), .B({ _16996_, _16995_, _16993_, _16992_, _16991_, _16990_, _16989_, _16988_, _16987_, _16986_, _16985_, _16984_, _16982_, _16981_, _16980_, _16979_, _16978_, _16977_, _16976_, _16975_, _16974_, _16973_, _17003_, _17002_, _17001_, _17000_, _16999_, _16998_, _16997_, _16994_, _16983_, _16972_ }), .S(_21917_), .Y(_22616_) );
  \$mux  #( .WIDTH(32) ) _48877_ ( .A(_stream_conv2d_8_source_19_source_pat_fsm_2), .B({ _17092_, _17091_, _17089_, _17088_, _17087_, _17086_, _17085_, _17084_, _17083_, _17082_, _17081_, _17080_, _17078_, _17077_, _17076_, _17075_, _17074_, _17073_, _17072_, _17071_, _17070_, _17069_, _17099_, _17098_, _17097_, _17096_, _17095_, _17094_, _17093_, _17090_, _17079_, _17068_ }), .S(_21918_), .Y(_22617_) );
  \$mux  #( .WIDTH(32) ) _48878_ ( .A(_stream_conv2d_8_source_8_source_pat_fsm_1), .B({ _17188_, _17187_, _17185_, _17184_, _17183_, _17182_, _17181_, _17180_, _17179_, _17178_, _17177_, _17176_, _17174_, _17173_, _17172_, _17171_, _17170_, _17169_, _17168_, _17167_, _17166_, _17165_, _17195_, _17194_, _17193_, _17192_, _17191_, _17190_, _17189_, _17186_, _17175_, _17164_ }), .S(_21919_), .Y(_22618_) );
  \$mux  #( .WIDTH(32) ) _48879_ ( .A(_stream_conv2d_8_source_6_source_pat_fsm_0), .B({ _17284_, _17283_, _17281_, _17280_, _17279_, _17278_, _17277_, _17276_, _17275_, _17274_, _17273_, _17272_, _17270_, _17269_, _17268_, _17267_, _17266_, _17265_, _17264_, _17263_, _17262_, _17261_, _17291_, _17290_, _17289_, _17288_, _17287_, _17286_, _17285_, _17282_, _17271_, _17260_ }), .S(_21920_), .Y(_22619_) );
  \$mux  #( .WIDTH(32) ) _48880_ ( .A(conv2d_8_comp_fsm), .B({ _17412_, _17411_, _17409_, _17408_, _17407_, _17406_, _17405_, _17404_, _17403_, _17402_, _17401_, _17400_, _17398_, _17397_, _17396_, _17395_, _17394_, _17393_, _17392_, _17391_, _17390_, _17389_, _17419_, _17418_, _17417_, _17416_, _17415_, _17414_, _17413_, _17410_, _17399_, _17388_ }), .S(_21921_), .Y(_22629_) );
  \$mux  #( .WIDTH(32) ) _48881_ ( .A(conv2d_8_stream_out_local_col), .B({ _17540_, _17539_, _17537_, _17536_, _17535_, _17534_, _17533_, _17532_, _17531_, _17530_, _17529_, _17528_, _17526_, _17525_, _17524_, _17523_, _17522_, _17521_, _17520_, _17519_, _17518_, _17517_, _17547_, _17546_, _17545_, _17544_, _17543_, _17542_, _17541_, _17538_, _17527_, _17516_ }), .S(_21922_), .Y(_22630_) );
  \$mux  #( .WIDTH(32) ) _48882_ ( .A(conv2d_8_stream_act_local_8), .B({ _17605_, _17604_, _17602_, _17601_, _17600_, _17599_, _17598_, _17597_, _17596_, _17595_, _17594_, _17593_, _17591_, _17590_, _17589_, _17588_, _17587_, _17586_, _17585_, _17584_, _17583_, _17582_, _17612_, _17611_, _17610_, _17609_, _17608_, _17607_, _17606_, _17603_, _17592_, _17581_ }), .S(_21922_), .Y(_22633_) );
  \$mux  #( .WIDTH(32) ) _48883_ ( .A(conv2d_8_stream_act_local_7), .B({ _17702_, _17701_, _17699_, _17698_, _17697_, _17696_, _17695_, _17694_, _17693_, _17692_, _17691_, _17690_, _17688_, _17687_, _17686_, _17685_, _17684_, _17683_, _17682_, _17681_, _17680_, _17679_, _17709_, _17708_, _17707_, _17706_, _17705_, _17704_, _17703_, _17700_, _17689_, _17678_ }), .S(_21922_), .Y(_22635_) );
  \$mux  #( .WIDTH(32) ) _48884_ ( .A(conv2d_8_stream_act_local_6), .B({ _17767_, _17766_, _17764_, _17763_, _17762_, _17761_, _17760_, _17759_, _17758_, _17757_, _17756_, _17755_, _17753_, _17752_, _17751_, _17750_, _17749_, _17748_, _17747_, _17746_, _17745_, _17744_, _17774_, _17773_, _17772_, _17771_, _17770_, _17769_, _17768_, _17765_, _17754_, _17743_ }), .S(_21922_), .Y(_22637_) );
  \$mux  #( .WIDTH(32) ) _48885_ ( .A(conv2d_8_stream_act_local_5), .B({ _17831_, _17830_, _17828_, _17827_, _17826_, _17825_, _17824_, _17823_, _17822_, _17821_, _17820_, _17819_, _17817_, _17816_, _17815_, _17814_, _17813_, _17812_, _17811_, _17810_, _17809_, _17808_, _17838_, _17837_, _17836_, _17835_, _17834_, _17833_, _17832_, _17829_, _17818_, _17807_ }), .S(_21922_), .Y(_22640_) );
  \$mux  #( .WIDTH(32) ) _48886_ ( .A(conv2d_8_stream_act_local_4), .B({ _17895_, _17894_, _17892_, _17891_, _17890_, _17889_, _17888_, _17887_, _17886_, _17885_, _17884_, _17883_, _17881_, _17880_, _17879_, _17878_, _17877_, _17876_, _17875_, _17874_, _17873_, _17872_, _17902_, _17901_, _17900_, _17899_, _17898_, _17897_, _17896_, _17893_, _17882_, _17871_ }), .S(_21922_), .Y(_22642_) );
  \$mux  #( .WIDTH(32) ) _48887_ ( .A(conv2d_8_stream_act_local_3), .B({ _17959_, _17958_, _17956_, _17955_, _17954_, _17953_, _17952_, _17951_, _17950_, _17949_, _17948_, _17947_, _17945_, _17944_, _17943_, _17942_, _17941_, _17940_, _17939_, _17938_, _17937_, _17936_, _17966_, _17965_, _17964_, _17963_, _17962_, _17961_, _17960_, _17957_, _17946_, _17935_ }), .S(_21922_), .Y(_22644_) );
  \$mux  #( .WIDTH(32) ) _48888_ ( .A(conv2d_8_stream_act_local_2), .B({ _18023_, _18022_, _18020_, _18019_, _18018_, _18017_, _18016_, _18015_, _18014_, _18013_, _18012_, _18011_, _18009_, _18008_, _18007_, _18006_, _18005_, _18004_, _18003_, _18002_, _18001_, _18000_, _18030_, _18029_, _18028_, _18027_, _18026_, _18025_, _18024_, _18021_, _18010_, _17999_ }), .S(_21922_), .Y(_22647_) );
  \$mux  #( .WIDTH(32) ) _48889_ ( .A(conv2d_8_stream_act_local_1), .B({ _18087_, _18086_, _18084_, _18083_, _18082_, _18081_, _18080_, _18079_, _18078_, _18077_, _18076_, _18075_, _18073_, _18072_, _18071_, _18070_, _18069_, _18068_, _18067_, _18066_, _18065_, _18064_, _18094_, _18093_, _18092_, _18091_, _18090_, _18089_, _18088_, _18085_, _18074_, _18063_ }), .S(_21922_), .Y(_22649_) );
  \$mux  #( .WIDTH(32) ) _48890_ ( .A(conv2d_8_stream_act_local_0), .B({ _18151_, _18150_, _18148_, _18147_, _18146_, _18145_, _18144_, _18143_, _18142_, _18141_, _18140_, _18139_, _18137_, _18136_, _18135_, _18134_, _18133_, _18132_, _18131_, _18130_, _18129_, _18128_, _18158_, _18157_, _18156_, _18155_, _18154_, _18153_, _18152_, _18149_, _18138_, _18127_ }), .S(_21922_), .Y(_22651_) );
  \$mux  #( .WIDTH(2) ) _48891_ ( .A(conv2d_8_col_select), .B({ _18162_, _18161_ }), .S(_21922_), .Y(_22653_) );
  \$mux  #( .WIDTH(32) ) _48892_ ( .A(conv2d_8_col_count), .B({ _18219_, _18218_, _18216_, _18215_, _18214_, _18213_, _18212_, _18211_, _18210_, _18209_, _18208_, _18207_, _18205_, _18204_, _18203_, _18202_, _18201_, _18200_, _18199_, _18198_, _18197_, _18196_, _18226_, _18225_, _18224_, _18223_, _18222_, _18221_, _18220_, _18217_, _18206_, _18195_ }), .S(_21922_), .Y(_22654_) );
  \$mux  #( .WIDTH(33) ) _48893_ ( .A(_maxi_read_rest_size), .B({ _18285_, _18284_, _18283_, _18281_, _18280_, _18279_, _18278_, _18277_, _18276_, _18275_, _18274_, _18273_, _18272_, _18270_, _18269_, _18268_, _18267_, _18266_, _18265_, _18264_, _18263_, _18262_, _18261_, _18292_, _18291_, _18290_, _18289_, _18288_, _18287_, _18286_, _18282_, _18271_, _18260_ }), .S(_04830_), .Y(_22731_) );
  \$mux  #( .WIDTH(32) ) _48894_ ( .A(_maxi_read_cur_global_addr), .B({ _18382_, _18381_, _18379_, _18378_, _18377_, _18376_, _18375_, _18374_, _18373_, _18372_, _18371_, _18370_, _18368_, _18367_, _18366_, _18365_, _18364_, _18363_, _18362_, _18361_, _18360_, _18359_, _18389_, _18388_, _18387_, _18386_, _18385_, _18384_, _18383_, _18380_, _18369_, _18358_ }), .S(_21923_), .Y(_22736_) );
  \$mux  #( .WIDTH(32) ) _48895_ ( .A(_maxi_read_fsm), .B({ _18446_, _18445_, _18443_, _18442_, _18441_, _18440_, _18439_, _18438_, _18437_, _18436_, _18435_, _18434_, _18432_, _18431_, _18430_, _18429_, _18428_, _18427_, _18426_, _18425_, _18424_, _18423_, _18453_, _18452_, _18451_, _18450_, _18449_, _18448_, _18447_, _18444_, _18433_, _18422_ }), .S(_21924_), .Y(_22737_) );
  \$mux  #( .WIDTH(1) ) _48896_ ( .A(conv2d_8_skip_write_out), .B(_18551_), .S(_04700_), .Y(_22791_) );
  \$mux  #( .WIDTH(1) ) _48897_ ( .A(conv2d_8_skip_comp), .B(_18553_), .S(_04700_), .Y(_22792_) );
  \$mux  #( .WIDTH(1) ) _48898_ ( .A(conv2d_8_skip_read_act), .B(_18555_), .S(_04700_), .Y(_22793_) );
  \$mux  #( .WIDTH(1) ) _48899_ ( .A(conv2d_8_skip_read_filter), .B(_18557_), .S(_04700_), .Y(_22794_) );
  \$mux  #( .WIDTH(32) ) _48900_ ( .A(conv2d_8_out_laddr_offset), .B({ _04833_, _04834_, _04835_, _04836_, _04837_, _04838_, _04839_, _04840_, _04841_, _04842_, _04843_, _04844_, _04845_, _04846_, _04847_, _04848_, _04849_, _04850_, _04851_, _04852_, _04853_, _04854_, _04855_, _04856_, _04857_, _04858_, _04859_, _04860_, _04861_, _04862_, _04863_, _04864_ }), .S(_21925_), .Y(_22795_) );
  \$mux  #( .WIDTH(32) ) _48901_ ( .A(conv2d_8_out_page_dma_offset), .B({ _18678_, _18677_, _18675_, _18674_, _18673_, _18672_, _18671_, _18670_, _18669_, _18668_, _18667_, _18666_, _18664_, _18663_, _18662_, _18661_, _18660_, _18659_, _18658_, _18657_, _18656_, _18655_, _18685_, _18684_, _18683_, _18682_, _18681_, _18680_, _18679_, _18676_, _18665_, _18654_ }), .S(_04700_), .Y(_22796_) );
  \$mux  #( .WIDTH(32) ) _48902_ ( .A(conv2d_8_out_page_comp_offset), .B({ _18742_, _18741_, _18739_, _18738_, _18737_, _18736_, _18735_, _18734_, _18733_, _18732_, _18731_, _18730_, _18728_, _18727_, _18726_, _18725_, _18724_, _18723_, _18722_, _18721_, _18720_, _18719_, _18749_, _18748_, _18747_, _18746_, _18745_, _18744_, _18743_, _18740_, _18729_, _18718_ }), .S(_04700_), .Y(_22797_) );
  \$mux  #( .WIDTH(1) ) _48903_ ( .A(conv2d_8_out_page), .B(_18751_), .S(_04700_), .Y(_22798_) );
  \$mux  #( .WIDTH(32) ) _48904_ ( .A(conv2d_8_filter_page_dma_offset), .B({ _18808_, _18807_, _18805_, _18804_, _18803_, _18802_, _18801_, _18800_, _18799_, _18798_, _18797_, _18796_, _18794_, _18793_, _18792_, _18791_, _18790_, _18789_, _18788_, _18787_, _18786_, _18785_, _18815_, _18814_, _18813_, _18812_, _18811_, _18810_, _18809_, _18806_, _18795_, _18784_ }), .S(_04700_), .Y(_22800_) );
  \$mux  #( .WIDTH(32) ) _48905_ ( .A(conv2d_8_filter_page_comp_offset), .B({ _18872_, _18871_, _18869_, _18868_, _18867_, _18866_, _18865_, _18864_, _18863_, _18862_, _18861_, _18860_, _18858_, _18857_, _18856_, _18855_, _18854_, _18853_, _18852_, _18851_, _18850_, _18849_, _18879_, _18878_, _18877_, _18876_, _18875_, _18874_, _18873_, _18870_, _18859_, _18848_ }), .S(_04700_), .Y(_22802_) );
  \$mux  #( .WIDTH(32) ) _48906_ ( .A(conv2d_8_act_page_dma_offset_2), .B({ _18936_, _18935_, _18933_, _18932_, _18931_, _18930_, _18929_, _18928_, _18927_, _18926_, _18925_, _18924_, _18922_, _18921_, _18920_, _18919_, _18918_, _18917_, _18916_, _18915_, _18914_, _18913_, _18943_, _18942_, _18941_, _18940_, _18939_, _18938_, _18937_, _18934_, _18923_, _18912_ }), .S(_04700_), .Y(_22805_) );
  \$mux  #( .WIDTH(32) ) _48907_ ( .A(conv2d_8_act_page_dma_offset_1), .B({ _19000_, _18999_, _18997_, _18996_, _18995_, _18994_, _18993_, _18992_, _18991_, _18990_, _18989_, _18988_, _18986_, _18985_, _18984_, _18983_, _18982_, _18981_, _18980_, _18979_, _18978_, _18977_, _19007_, _19006_, _19005_, _19004_, _19003_, _19002_, _19001_, _18998_, _18987_, _18976_ }), .S(_04700_), .Y(_22808_) );
  \$mux  #( .WIDTH(32) ) _48908_ ( .A(conv2d_8_act_page_dma_offset_0), .B({ _19064_, _19063_, _19061_, _19060_, _19059_, _19058_, _19057_, _19056_, _19055_, _19054_, _19053_, _19052_, _19050_, _19049_, _19048_, _19047_, _19046_, _19045_, _19044_, _19043_, _19042_, _19041_, _19071_, _19070_, _19069_, _19068_, _19067_, _19066_, _19065_, _19062_, _19051_, _19040_ }), .S(_04700_), .Y(_22811_) );
  \$mux  #( .WIDTH(32) ) _48909_ ( .A(conv2d_8_act_page_comp_offset_2), .B({ _19128_, _19127_, _19125_, _19124_, _19123_, _19122_, _19121_, _19120_, _19119_, _19118_, _19117_, _19116_, _19114_, _19113_, _19112_, _19111_, _19110_, _19109_, _19108_, _19107_, _19106_, _19105_, _19135_, _19134_, _19133_, _19132_, _19131_, _19130_, _19129_, _19126_, _19115_, _19104_ }), .S(_04700_), .Y(_22814_) );
  \$mux  #( .WIDTH(32) ) _48910_ ( .A(conv2d_8_act_page_comp_offset_1), .B({ _19192_, _19191_, _19189_, _19188_, _19187_, _19186_, _19185_, _19184_, _19183_, _19182_, _19181_, _19180_, _19178_, _19177_, _19176_, _19175_, _19174_, _19173_, _19172_, _19171_, _19170_, _19169_, _19199_, _19198_, _19197_, _19196_, _19195_, _19194_, _19193_, _19190_, _19179_, _19168_ }), .S(_04700_), .Y(_22817_) );
  \$mux  #( .WIDTH(32) ) _48911_ ( .A(conv2d_8_act_page_comp_offset_0), .B({ _19256_, _19255_, _19253_, _19252_, _19251_, _19250_, _19249_, _19248_, _19247_, _19246_, _19245_, _19244_, _19242_, _19241_, _19240_, _19239_, _19238_, _19237_, _19236_, _19235_, _19234_, _19233_, _19263_, _19262_, _19261_, _19260_, _19259_, _19258_, _19257_, _19254_, _19243_, _19232_ }), .S(_04700_), .Y(_22820_) );
  \$mux  #( .WIDTH(2) ) _48912_ ( .A(conv2d_8_prev_row_select), .B({ _19267_, _19266_ }), .S(_04700_), .Y(_22821_) );
  \$mux  #( .WIDTH(32) ) _48913_ ( .A(conv2d_8_prev_och_count), .B({ _19292_, _19291_, _19289_, _19288_, _19287_, _19286_, _19285_, _19284_, _19283_, _19282_, _19281_, _19280_, _19278_, _19277_, _19276_, _19275_, _19274_, _19273_, _19272_, _19271_, _19270_, _19269_, _19299_, _19298_, _19297_, _19296_, _19295_, _19294_, _19293_, _19290_, _19279_, _19268_ }), .S(_04700_), .Y(_22822_) );
  \$mux  #( .WIDTH(32) ) _48914_ ( .A(conv2d_8_prev_bat_count), .B({ _19324_, _19323_, _19321_, _19320_, _19319_, _19318_, _19317_, _19316_, _19315_, _19314_, _19313_, _19312_, _19310_, _19309_, _19308_, _19307_, _19306_, _19305_, _19304_, _19303_, _19302_, _19301_, _19331_, _19330_, _19329_, _19328_, _19327_, _19326_, _19325_, _19322_, _19311_, _19300_ }), .S(_04700_), .Y(_22823_) );
  \$mux  #( .WIDTH(32) ) _48915_ ( .A(conv2d_8_prev_row_count), .B({ _19356_, _19355_, _19353_, _19352_, _19351_, _19350_, _19349_, _19348_, _19347_, _19346_, _19345_, _19344_, _19342_, _19341_, _19340_, _19339_, _19338_, _19337_, _19336_, _19335_, _19334_, _19333_, _19363_, _19362_, _19361_, _19360_, _19359_, _19358_, _19357_, _19354_, _19343_, _19332_ }), .S(_04700_), .Y(_22824_) );
  \$mux  #( .WIDTH(32) ) _48916_ ( .A(conv2d_8_out_ram_select), .B({ _04766_, _04767_, _04768_, _04769_, _04770_, _04771_, _04772_, _04773_, _04774_, _04775_, _04776_, _04777_, _04778_, _04779_, _04780_, _04781_, _04782_, _04783_, _04784_, _04785_, _04786_, _04787_, _04788_, _04789_, _04790_, _04792_, _04791_, _04793_, _04794_, _04795_, _04796_, _04797_ }), .S(_21925_), .Y(_22825_) );
  \$mux  #( .WIDTH(32) ) _48917_ ( .A(conv2d_8_out_row_count), .B({ _19484_, _19483_, _19481_, _19480_, _19479_, _19478_, _19477_, _19476_, _19475_, _19474_, _19473_, _19472_, _19470_, _19469_, _19468_, _19467_, _19466_, _19465_, _19464_, _19463_, _19462_, _19461_, _19491_, _19490_, _19489_, _19488_, _19487_, _19486_, _19485_, _19482_, _19471_, _19460_ }), .S(_04700_), .Y(_22827_) );
  \$mux  #( .WIDTH(2) ) _48918_ ( .A(conv2d_8_row_select), .B({ _19495_, _19494_ }), .S(_04700_), .Y(_22829_) );
  \$mux  #( .WIDTH(32) ) _48919_ ( .A(conv2d_8_och_count), .B({ _19552_, _19551_, _19549_, _19548_, _19547_, _19546_, _19545_, _19544_, _19543_, _19542_, _19541_, _19540_, _19538_, _19537_, _19536_, _19535_, _19534_, _19533_, _19532_, _19531_, _19530_, _19529_, _19559_, _19558_, _19557_, _19556_, _19555_, _19554_, _19553_, _19550_, _19539_, _19528_ }), .S(_04700_), .Y(_22830_) );
  \$mux  #( .WIDTH(32) ) _48920_ ( .A(conv2d_8_bat_count), .B({ _19616_, _19615_, _19613_, _19612_, _19611_, _19610_, _19609_, _19608_, _19607_, _19606_, _19605_, _19604_, _19602_, _19601_, _19600_, _19599_, _19598_, _19597_, _19596_, _19595_, _19594_, _19593_, _19623_, _19622_, _19621_, _19620_, _19619_, _19618_, _19617_, _19614_, _19603_, _19592_ }), .S(_04700_), .Y(_22831_) );
  \$mux  #( .WIDTH(32) ) _48921_ ( .A(conv2d_8_row_count), .B({ _19680_, _19679_, _19677_, _19676_, _19675_, _19674_, _19673_, _19672_, _19671_, _19670_, _19669_, _19668_, _19666_, _19665_, _19664_, _19663_, _19662_, _19661_, _19660_, _19659_, _19658_, _19657_, _19687_, _19686_, _19685_, _19684_, _19683_, _19682_, _19681_, _19678_, _19667_, _19656_ }), .S(_04700_), .Y(_22832_) );
  \$mux  #( .WIDTH(32) ) _48922_ ( .A(conv2d_8_sync_out_count), .B({ _19712_, _19711_, _19709_, _19708_, _19707_, _19706_, _19705_, _19704_, _19703_, _19702_, _19701_, _19700_, _19698_, _19697_, _19696_, _19695_, _19694_, _19693_, _19692_, _19691_, _19690_, _19689_, _19719_, _19718_, _19717_, _19716_, _19715_, _19714_, _19713_, _19710_, _19699_, _19688_ }), .S(_21926_), .Y(_22834_) );
  \$mux  #( .WIDTH(1) ) _48923_ ( .A(conv2d_8_dma_flag_2), .B(_19721_), .S(_04700_), .Y(_22835_) );
  \$mux  #( .WIDTH(1) ) _48924_ ( .A(conv2d_8_dma_flag_1), .B(_19721_), .S(_04700_), .Y(_22836_) );
  \$mux  #( .WIDTH(32) ) _48925_ ( .A(conv2d_8_out_base_offset_och), .B({ _19778_, _19777_, _19775_, _19774_, _19773_, _19772_, _19771_, _19770_, _19769_, _19768_, _19767_, _19766_, _19764_, _19763_, _19762_, _19761_, _19760_, _19759_, _19758_, _19757_, _19756_, _19755_, _19785_, _19784_, _19783_, _19782_, _19781_, _19780_, _19779_, _19776_, _19765_, _19754_ }), .S(_04700_), .Y(_22838_) );
  \$mux  #( .WIDTH(32) ) _48926_ ( .A(conv2d_8_out_base_offset_bat), .B({ _19842_, _19841_, _19839_, _19838_, _19837_, _19836_, _19835_, _19834_, _19833_, _19832_, _19831_, _19830_, _19828_, _19827_, _19826_, _19825_, _19824_, _19823_, _19822_, _19821_, _19820_, _19819_, _19849_, _19848_, _19847_, _19846_, _19845_, _19844_, _19843_, _19840_, _19829_, _19818_ }), .S(_04700_), .Y(_22839_) );
  \$mux  #( .WIDTH(32) ) _48927_ ( .A(conv2d_8_out_base_offset_row), .B({ _19906_, _19905_, _19903_, _19902_, _19901_, _19900_, _19899_, _19898_, _19897_, _19896_, _19895_, _19894_, _19892_, _19891_, _19890_, _19889_, _19888_, _19887_, _19886_, _19885_, _19884_, _19883_, _19913_, _19912_, _19911_, _19910_, _19909_, _19908_, _19907_, _19904_, _19893_, _19882_ }), .S(_04700_), .Y(_22841_) );
  \$mux  #( .WIDTH(32) ) _48928_ ( .A(conv2d_8_out_base_offset_col), .B({ _19970_, _19969_, _19967_, _19966_, _19965_, _19964_, _19963_, _19962_, _19961_, _19960_, _19959_, _19958_, _19956_, _19955_, _19954_, _19953_, _19952_, _19951_, _19950_, _19949_, _19948_, _19947_, _19977_, _19976_, _19975_, _19974_, _19973_, _19972_, _19971_, _19968_, _19957_, _19946_ }), .S(_04700_), .Y(_22842_) );
  \$mux  #( .WIDTH(32) ) _48929_ ( .A(conv2d_8_filter_base_offset), .B({ _20034_, _20033_, _20031_, _20030_, _20029_, _20028_, _20027_, _20026_, _20025_, _20024_, _20023_, _20022_, _20020_, _20019_, _20018_, _20017_, _20016_, _20015_, _20014_, _20013_, _20012_, _20011_, _20041_, _20040_, _20039_, _20038_, _20037_, _20036_, _20035_, _20032_, _20021_, _20010_ }), .S(_04700_), .Y(_22844_) );
  \$mux  #( .WIDTH(32) ) _48930_ ( .A(conv2d_8_act_base_offset_bat), .B({ _20098_, _20097_, _20095_, _20094_, _20093_, _20092_, _20091_, _20090_, _20089_, _20088_, _20087_, _20086_, _20084_, _20083_, _20082_, _20081_, _20080_, _20079_, _20078_, _20077_, _20076_, _20075_, _20105_, _20104_, _20103_, _20102_, _20101_, _20100_, _20099_, _20096_, _20085_, _20074_ }), .S(_04700_), .Y(_22845_) );
  \$mux  #( .WIDTH(32) ) _48931_ ( .A(conv2d_8_act_base_offset_row), .B({ _20162_, _20161_, _20159_, _20158_, _20157_, _20156_, _20155_, _20154_, _20153_, _20152_, _20151_, _20150_, _20148_, _20147_, _20146_, _20145_, _20144_, _20143_, _20142_, _20141_, _20140_, _20139_, _20169_, _20168_, _20167_, _20166_, _20165_, _20164_, _20163_, _20160_, _20149_, _20138_ }), .S(_04700_), .Y(_22846_) );
  \$mux  #( .WIDTH(32) ) _48932_ ( .A(control_conv2d_8), .B({ _20226_, _20225_, _20223_, _20222_, _20221_, _20220_, _20219_, _20218_, _20217_, _20216_, _20215_, _20214_, _20212_, _20211_, _20210_, _20209_, _20208_, _20207_, _20206_, _20205_, _20204_, _20203_, _20233_, _20232_, _20231_, _20230_, _20229_, _20228_, _20227_, _20224_, _20213_, _20202_ }), .S(_21927_), .Y(_22848_) );
  \$mux  #( .WIDTH(32) ) _48933_ ( .A(max_pool_serial_9_arg_objaddr_0), .B({ _20962_, _20961_, _20959_, _20958_, _20957_, _20956_, _20955_, _20954_, _20953_, _20952_, _20951_, _20950_, _20948_, _20947_, _20946_, _20945_, _20944_, _20943_, _20942_, _20941_, _20940_, _20939_, _20969_, _20968_, _20967_, _20966_, _20965_, _20964_, _20963_, _20960_, _20949_, _20938_ }), .S(_21928_), .Y(_22859_) );
  \$mux  #( .WIDTH(32) ) _48934_ ( .A(max_pool_serial_9_objaddr), .B({ _20994_, _20993_, _20991_, _20990_, _20989_, _20988_, _20987_, _20986_, _20985_, _20984_, _20983_, _20982_, _20980_, _20979_, _20978_, _20977_, _20976_, _20975_, _20974_, _20973_, _20972_, _20971_, _21001_, _21000_, _20999_, _20998_, _20997_, _20996_, _20995_, _20992_, _20981_, _20970_ }), .S(_21929_), .Y(_22860_) );
  \$mux  #( .WIDTH(32) ) _48935_ ( .A(conv2d_8_arg_objaddr_3), .B({ _21026_, _21025_, _21023_, _21022_, _21021_, _21020_, _21019_, _21018_, _21017_, _21016_, _21015_, _21014_, _21012_, _21011_, _21010_, _21009_, _21008_, _21007_, _21006_, _21005_, _21004_, _21003_, _21033_, _21032_, _21031_, _21030_, _21029_, _21028_, _21027_, _21024_, _21013_, _21002_ }), .S(_21930_), .Y(_22861_) );
  \$mux  #( .WIDTH(32) ) _48936_ ( .A(conv2d_8_arg_objaddr_2), .B({ _21058_, _21057_, _21055_, _21054_, _21053_, _21052_, _21051_, _21050_, _21049_, _21048_, _21047_, _21046_, _21044_, _21043_, _21042_, _21041_, _21040_, _21039_, _21038_, _21037_, _21036_, _21035_, _21065_, _21064_, _21063_, _21062_, _21061_, _21060_, _21059_, _21056_, _21045_, _21034_ }), .S(_21931_), .Y(_22862_) );
  \$mux  #( .WIDTH(32) ) _48937_ ( .A(conv2d_8_arg_objaddr_1), .B({ _21090_, _21089_, _21087_, _21086_, _21085_, _21084_, _21083_, _21082_, _21081_, _21080_, _21079_, _21078_, _21076_, _21075_, _21074_, _21073_, _21072_, _21071_, _21070_, _21069_, _21068_, _21067_, _21097_, _21096_, _21095_, _21094_, _21093_, _21092_, _21091_, _21088_, _21077_, _21066_ }), .S(_21932_), .Y(_22863_) );
  \$mux  #( .WIDTH(32) ) _48938_ ( .A(conv2d_8_arg_objaddr_0), .B({ _21122_, _21121_, _21119_, _21118_, _21117_, _21116_, _21115_, _21114_, _21113_, _21112_, _21111_, _21110_, _21108_, _21107_, _21106_, _21105_, _21104_, _21103_, _21102_, _21101_, _21100_, _21099_, _21129_, _21128_, _21127_, _21126_, _21125_, _21124_, _21123_, _21120_, _21109_, _21098_ }), .S(_21933_), .Y(_22864_) );
  \$mux  #( .WIDTH(32) ) _48939_ ( .A(conv2d_8_objaddr), .B({ _21154_, _21153_, _21151_, _21150_, _21149_, _21148_, _21147_, _21146_, _21145_, _21144_, _21143_, _21142_, _21140_, _21139_, _21138_, _21137_, _21136_, _21135_, _21134_, _21133_, _21132_, _21131_, _21161_, _21160_, _21159_, _21158_, _21157_, _21156_, _21155_, _21152_, _21141_, _21130_ }), .S(_21934_), .Y(_22865_) );
  \$mux  #( .WIDTH(32) ) _48940_ ( .A(main_fsm), .B({ _21187_, _21186_, _21184_, _21183_, _21182_, _21181_, _21180_, _21179_, _21178_, _21177_, _21176_, _21175_, _21173_, _21172_, _21171_, _21170_, _21169_, _21168_, _21167_, _21166_, _21165_, _21164_, _21194_, _21193_, _21192_, _21191_, _21190_, _21189_, _21188_, _21185_, _21174_, _21163_ }), .S(_21935_), .Y(_22866_) );
  \$mux  #( .WIDTH(1) ) _48941_ ( .A(max_pool_serial_9_control_param_index), .B(_04831_), .S(_21936_), .Y(_22867_) );
  \$mux  #( .WIDTH(1) ) _48942_ ( .A(conv2d_8_control_param_index), .B(_21162_), .S(_21937_), .Y(_22868_) );
  \$mux  #( .WIDTH(1) ) _48943_ ( .A(_stream_matmul_15_source_busy), .B(_21387_), .S(_21938_), .Y(_22869_) );
  \$mux  #( .WIDTH(32) ) _48944_ ( .A(_stream_matmul_15_fsm), .B({ _21413_, _21412_, _21410_, _21409_, _21408_, _21407_, _21406_, _21405_, _21404_, _21403_, _21402_, _21401_, _21399_, _21398_, _21397_, _21396_, _21395_, _21394_, _21393_, _21392_, _21391_, _21390_, _21420_, _21419_, _21418_, _21417_, _21416_, _21415_, _21414_, _21411_, _21400_, _21389_ }), .S(_21939_), .Y(_22874_) );
  \$mux  #( .WIDTH(1) ) _48945_ ( .A(_stream_max_pool_serial_9_source_busy), .B(_21485_), .S(_21940_), .Y(_23117_) );
  \$mux  #( .WIDTH(32) ) _48946_ ( .A(_stream_max_pool_serial_9_fsm), .B({ _21511_, _21510_, _21508_, _21507_, _21506_, _21505_, _21504_, _21503_, _21502_, _21501_, _21500_, _21499_, _21497_, _21496_, _21495_, _21494_, _21493_, _21492_, _21491_, _21490_, _21489_, _21488_, _21518_, _21517_, _21516_, _21515_, _21514_, _21513_, _21512_, _21509_, _21498_, _21487_ }), .S(_21941_), .Y(_23122_) );
  \$mux  #( .WIDTH(1) ) _48947_ ( .A(_stream_conv2d_8_source_busy), .B(_21583_), .S(_21942_), .Y(_23195_) );
  \$mux  #( .WIDTH(32) ) _48948_ ( .A(_stream_conv2d_8_fsm), .B({ _21609_, _21608_, _21606_, _21605_, _21604_, _21603_, _21602_, _21601_, _21600_, _21599_, _21598_, _21597_, _21595_, _21594_, _21593_, _21592_, _21591_, _21590_, _21589_, _21588_, _21587_, _21586_, _21616_, _21615_, _21614_, _21613_, _21612_, _21611_, _21610_, _21607_, _21596_, _21585_ }), .S(_21943_), .Y(_23200_) );
  \$mux  #( .WIDTH(32) ) _48949_ ( .A(_saxi_register_fsm), .B({ _21705_, _21704_, _21702_, _21701_, _21700_, _21699_, _21698_, _21697_, _21696_, _21695_, _21694_, _21693_, _21691_, _21690_, _21689_, _21688_, _21687_, _21686_, _21685_, _21684_, _21683_, _21682_, _21712_, _21711_, _21710_, _21709_, _21708_, _21707_, _21706_, _21703_, _21692_, _21681_ }), .S(_21944_), .Y(_25527_) );
  \$mux  #( .WIDTH(2) ) _48950_ ( .A({ 1'hx, _26441_ }), .B({ _26441_, 1'hx }), .S(_counter_data_762[31]), .Y(_25911_) );
  \$mux  #( .WIDTH(66) ) _48951_ ( .A({ _26336_[65:34], _26331_[65:32] }), .B({ _26331_[65:32], 32'h00000000 }), .S(_minus_data_5[5]), .Y(_25912_) );
  \$mux  #( .WIDTH(66) ) _48952_ ( .A({ _26335_[65:50], _26330_[65:16] }), .B({ _26330_[65:16], 16'h0000 }), .S(_minus_data_5[4]), .Y({ _26336_[65:34], _26331_[65:32] }) );
  \$mux  #( .WIDTH(66) ) _48953_ ( .A(_26334_), .B({ _26334_[57:0], 8'h00 }), .S(_minus_data_5[3]), .Y({ _26335_[65:50], _26330_[65:16] }) );
  \$mux  #( .WIDTH(66) ) _48954_ ( .A(_26333_), .B({ _26333_[61:0], 4'h0 }), .S(_minus_data_5[2]), .Y(_26334_) );
  \$mux  #( .WIDTH(66) ) _48955_ ( .A(_26332_), .B({ _26332_[63:0], 2'h0 }), .S(_minus_data_5[1]), .Y(_26333_) );
  \$mux  #( .WIDTH(66) ) _48956_ ( .A(66'h00000000000000001), .B(66'h00000000000000002), .S(_minus_data_5[0]), .Y(_26332_) );
  \$mux  #( .WIDTH(18) ) _48957_ ( .A(_26339_), .B({ _26339_[9:0], 8'h00 }), .S(_minus_data_57[3]), .Y(_25913_) );
  \$mux  #( .WIDTH(18) ) _48958_ ( .A(_26338_), .B({ _26338_[13:0], 4'h0 }), .S(_minus_data_57[2]), .Y(_26339_) );
  \$mux  #( .WIDTH(18) ) _48959_ ( .A(_26337_), .B({ _26337_[15:0], 2'h0 }), .S(_minus_data_57[1]), .Y(_26338_) );
  \$mux  #( .WIDTH(18) ) _48960_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_57[0]), .Y(_26337_) );
  \$mux  #( .WIDTH(18) ) _48961_ ( .A(_26342_), .B({ _26342_[9:0], 8'h00 }), .S(_minus_data_72[3]), .Y(_25914_) );
  \$mux  #( .WIDTH(18) ) _48962_ ( .A(_26341_), .B({ _26341_[13:0], 4'h0 }), .S(_minus_data_72[2]), .Y(_26342_) );
  \$mux  #( .WIDTH(18) ) _48963_ ( .A(_26340_), .B({ _26340_[15:0], 2'h0 }), .S(_minus_data_72[1]), .Y(_26341_) );
  \$mux  #( .WIDTH(18) ) _48964_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_72[0]), .Y(_26340_) );
  \$mux  #( .WIDTH(18) ) _48965_ ( .A(_26345_), .B({ _26345_[9:0], 8'h00 }), .S(_minus_data_87[3]), .Y(_25915_) );
  \$mux  #( .WIDTH(18) ) _48966_ ( .A(_26344_), .B({ _26344_[13:0], 4'h0 }), .S(_minus_data_87[2]), .Y(_26345_) );
  \$mux  #( .WIDTH(18) ) _48967_ ( .A(_26343_), .B({ _26343_[15:0], 2'h0 }), .S(_minus_data_87[1]), .Y(_26344_) );
  \$mux  #( .WIDTH(18) ) _48968_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_87[0]), .Y(_26343_) );
  \$mux  #( .WIDTH(18) ) _48969_ ( .A(_26348_), .B({ _26348_[9:0], 8'h00 }), .S(_minus_data_102[3]), .Y(_25916_) );
  \$mux  #( .WIDTH(18) ) _48970_ ( .A(_26347_), .B({ _26347_[13:0], 4'h0 }), .S(_minus_data_102[2]), .Y(_26348_) );
  \$mux  #( .WIDTH(18) ) _48971_ ( .A(_26346_), .B({ _26346_[15:0], 2'h0 }), .S(_minus_data_102[1]), .Y(_26347_) );
  \$mux  #( .WIDTH(18) ) _48972_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_102[0]), .Y(_26346_) );
  \$mux  #( .WIDTH(18) ) _48973_ ( .A(_26351_), .B({ _26351_[9:0], 8'h00 }), .S(_minus_data_117[3]), .Y(_25917_) );
  \$mux  #( .WIDTH(18) ) _48974_ ( .A(_26350_), .B({ _26350_[13:0], 4'h0 }), .S(_minus_data_117[2]), .Y(_26351_) );
  \$mux  #( .WIDTH(18) ) _48975_ ( .A(_26349_), .B({ _26349_[15:0], 2'h0 }), .S(_minus_data_117[1]), .Y(_26350_) );
  \$mux  #( .WIDTH(18) ) _48976_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_117[0]), .Y(_26349_) );
  \$mux  #( .WIDTH(18) ) _48977_ ( .A(_26354_), .B({ _26354_[9:0], 8'h00 }), .S(_minus_data_132[3]), .Y(_25918_) );
  \$mux  #( .WIDTH(18) ) _48978_ ( .A(_26353_), .B({ _26353_[13:0], 4'h0 }), .S(_minus_data_132[2]), .Y(_26354_) );
  \$mux  #( .WIDTH(18) ) _48979_ ( .A(_26352_), .B({ _26352_[15:0], 2'h0 }), .S(_minus_data_132[1]), .Y(_26353_) );
  \$mux  #( .WIDTH(18) ) _48980_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_132[0]), .Y(_26352_) );
  \$mux  #( .WIDTH(18) ) _48981_ ( .A(_26357_), .B({ _26357_[9:0], 8'h00 }), .S(_minus_data_147[3]), .Y(_25919_) );
  \$mux  #( .WIDTH(18) ) _48982_ ( .A(_26356_), .B({ _26356_[13:0], 4'h0 }), .S(_minus_data_147[2]), .Y(_26357_) );
  \$mux  #( .WIDTH(18) ) _48983_ ( .A(_26355_), .B({ _26355_[15:0], 2'h0 }), .S(_minus_data_147[1]), .Y(_26356_) );
  \$mux  #( .WIDTH(18) ) _48984_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_147[0]), .Y(_26355_) );
  \$mux  #( .WIDTH(18) ) _48985_ ( .A(_26360_), .B({ _26360_[9:0], 8'h00 }), .S(_minus_data_162[3]), .Y(_25920_) );
  \$mux  #( .WIDTH(18) ) _48986_ ( .A(_26359_), .B({ _26359_[13:0], 4'h0 }), .S(_minus_data_162[2]), .Y(_26360_) );
  \$mux  #( .WIDTH(18) ) _48987_ ( .A(_26358_), .B({ _26358_[15:0], 2'h0 }), .S(_minus_data_162[1]), .Y(_26359_) );
  \$mux  #( .WIDTH(18) ) _48988_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_162[0]), .Y(_26358_) );
  \$mux  #( .WIDTH(18) ) _48989_ ( .A(_26363_), .B({ _26363_[9:0], 8'h00 }), .S(_minus_data_177[3]), .Y(_25921_) );
  \$mux  #( .WIDTH(18) ) _48990_ ( .A(_26362_), .B({ _26362_[13:0], 4'h0 }), .S(_minus_data_177[2]), .Y(_26363_) );
  \$mux  #( .WIDTH(18) ) _48991_ ( .A(_26361_), .B({ _26361_[15:0], 2'h0 }), .S(_minus_data_177[1]), .Y(_26362_) );
  \$mux  #( .WIDTH(18) ) _48992_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_177[0]), .Y(_26361_) );
  \$mux  #( .WIDTH(32) ) _48993_ ( .A(_26366_), .B({ _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31], _26366_[31] }), .S(__delay_data_734[5]), .Y(_25924_) );
  \$mux  #( .WIDTH(32) ) _48994_ ( .A(_26364_), .B({ _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31], _26364_[31:16] }), .S(__delay_data_734[4]), .Y(_26366_) );
  \$mux  #( .WIDTH(32) ) _48995_ ( .A({ _26365_[31], _26365_[22:0], _26369_[7:0] }), .B({ _26365_[31], _26365_[31], _26365_[31], _26365_[31], _26365_[31], _26365_[31], _26365_[31], _26365_[31], _26365_[31], _26365_[22:0] }), .S(__delay_data_734[3]), .Y(_26364_) );
  \$mux  #( .WIDTH(32) ) _48996_ ( .A(_26368_), .B({ _26368_[31], _26368_[31], _26368_[31], _26368_[31], _26368_[31:4] }), .S(__delay_data_734[2]), .Y({ _26365_[31], _26365_[22:0], _26369_[7:0] }) );
  \$mux  #( .WIDTH(32) ) _48997_ ( .A(_26367_), .B({ _26367_[31], _26367_[31], _26367_[31:2] }), .S(__delay_data_734[1]), .Y(_26368_) );
  \$mux  #( .WIDTH(32) ) _48998_ ( .A(_plus_data_18), .B({ _plus_data_18[31], _plus_data_18[31:1] }), .S(__delay_data_734[0]), .Y(_26367_) );
  \$mux  #( .WIDTH(40) ) _48999_ ( .A(_26372_), .B({ _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39], _26372_[39:32] }), .S(__delay_data_747[5]), .Y(_25925_) );
  \$mux  #( .WIDTH(40) ) _49000_ ( .A(_26370_), .B({ _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39], _26370_[39:16] }), .S(__delay_data_747[4]), .Y(_26372_) );
  \$mux  #( .WIDTH(40) ) _49001_ ( .A({ _26371_[39], _26371_[30:0], _26375_[7:0] }), .B({ _26371_[39], _26371_[39], _26371_[39], _26371_[39], _26371_[39], _26371_[39], _26371_[39], _26371_[39], _26371_[39], _26371_[30:0] }), .S(__delay_data_747[3]), .Y(_26370_) );
  \$mux  #( .WIDTH(40) ) _49002_ ( .A(_26374_), .B({ _26374_[39], _26374_[39], _26374_[39], _26374_[39], _26374_[39:4] }), .S(__delay_data_747[2]), .Y({ _26371_[39], _26371_[30:0], _26375_[7:0] }) );
  \$mux  #( .WIDTH(40) ) _49003_ ( .A(_26373_), .B({ _26373_[39], _26373_[39], _26373_[39:2] }), .S(__delay_data_747[1]), .Y(_26374_) );
  \$mux  #( .WIDTH(40) ) _49004_ ( .A(_times_mul_odata_reg_39), .B({ _times_mul_odata_reg_39[39], _times_mul_odata_reg_39[39:1] }), .S(__delay_data_747[0]), .Y(_26373_) );
  \$mux  #( .WIDTH(16) ) _49005_ ( .A({ _26376_[15], _26376_[6:0], _26379_[7:0] }), .B({ _26376_[15], _26376_[15], _26376_[15], _26376_[15], _26376_[15], _26376_[15], _26376_[15], _26376_[15], _26376_[15], _26376_[6:0] }), .S(__delay_data_586[3]), .Y(_25926_) );
  \$mux  #( .WIDTH(16) ) _49006_ ( .A(_26378_), .B({ _26378_[15], _26378_[15], _26378_[15], _26378_[15], _26378_[15:4] }), .S(__delay_data_586[2]), .Y({ _26376_[15], _26376_[6:0], _26379_[7:0] }) );
  \$mux  #( .WIDTH(16) ) _49007_ ( .A(_26377_), .B({ _26377_[15], _26377_[15], _26377_[15:2] }), .S(__delay_data_586[1]), .Y(_26378_) );
  \$mux  #( .WIDTH(16) ) _49008_ ( .A(__muladd_madd_odata_reg_65), .B({ __muladd_madd_odata_reg_65[15], __muladd_madd_odata_reg_65[15:1] }), .S(__delay_data_586[0]), .Y(_26377_) );
  \$mux  #( .WIDTH(16) ) _49009_ ( .A({ _26380_[15], _26380_[6:0], _26383_[7:0] }), .B({ _26380_[15], _26380_[15], _26380_[15], _26380_[15], _26380_[15], _26380_[15], _26380_[15], _26380_[15], _26380_[15], _26380_[6:0] }), .S(__delay_data_603[3]), .Y(_25927_) );
  \$mux  #( .WIDTH(16) ) _49010_ ( .A(_26382_), .B({ _26382_[15], _26382_[15], _26382_[15], _26382_[15], _26382_[15:4] }), .S(__delay_data_603[2]), .Y({ _26380_[15], _26380_[6:0], _26383_[7:0] }) );
  \$mux  #( .WIDTH(16) ) _49011_ ( .A(_26381_), .B({ _26381_[15], _26381_[15], _26381_[15:2] }), .S(__delay_data_603[1]), .Y(_26382_) );
  \$mux  #( .WIDTH(16) ) _49012_ ( .A(__muladd_madd_odata_reg_80), .B({ __muladd_madd_odata_reg_80[15], __muladd_madd_odata_reg_80[15:1] }), .S(__delay_data_603[0]), .Y(_26381_) );
  \$mux  #( .WIDTH(16) ) _49013_ ( .A({ _26384_[15], _26384_[6:0], _26387_[7:0] }), .B({ _26384_[15], _26384_[15], _26384_[15], _26384_[15], _26384_[15], _26384_[15], _26384_[15], _26384_[15], _26384_[15], _26384_[6:0] }), .S(__delay_data_620[3]), .Y(_25928_) );
  \$mux  #( .WIDTH(16) ) _49014_ ( .A(_26386_), .B({ _26386_[15], _26386_[15], _26386_[15], _26386_[15], _26386_[15:4] }), .S(__delay_data_620[2]), .Y({ _26384_[15], _26384_[6:0], _26387_[7:0] }) );
  \$mux  #( .WIDTH(16) ) _49015_ ( .A(_26385_), .B({ _26385_[15], _26385_[15], _26385_[15:2] }), .S(__delay_data_620[1]), .Y(_26386_) );
  \$mux  #( .WIDTH(16) ) _49016_ ( .A(__muladd_madd_odata_reg_95), .B({ __muladd_madd_odata_reg_95[15], __muladd_madd_odata_reg_95[15:1] }), .S(__delay_data_620[0]), .Y(_26385_) );
  \$mux  #( .WIDTH(16) ) _49017_ ( .A({ _26388_[15], _26388_[6:0], _26391_[7:0] }), .B({ _26388_[15], _26388_[15], _26388_[15], _26388_[15], _26388_[15], _26388_[15], _26388_[15], _26388_[15], _26388_[15], _26388_[6:0] }), .S(__delay_data_637[3]), .Y(_25929_) );
  \$mux  #( .WIDTH(16) ) _49018_ ( .A(_26390_), .B({ _26390_[15], _26390_[15], _26390_[15], _26390_[15], _26390_[15:4] }), .S(__delay_data_637[2]), .Y({ _26388_[15], _26388_[6:0], _26391_[7:0] }) );
  \$mux  #( .WIDTH(16) ) _49019_ ( .A(_26389_), .B({ _26389_[15], _26389_[15], _26389_[15:2] }), .S(__delay_data_637[1]), .Y(_26390_) );
  \$mux  #( .WIDTH(16) ) _49020_ ( .A(__muladd_madd_odata_reg_110), .B({ __muladd_madd_odata_reg_110[15], __muladd_madd_odata_reg_110[15:1] }), .S(__delay_data_637[0]), .Y(_26389_) );
  \$mux  #( .WIDTH(16) ) _49021_ ( .A({ _26392_[15], _26392_[6:0], _26395_[7:0] }), .B({ _26392_[15], _26392_[15], _26392_[15], _26392_[15], _26392_[15], _26392_[15], _26392_[15], _26392_[15], _26392_[15], _26392_[6:0] }), .S(__delay_data_654[3]), .Y(_25930_) );
  \$mux  #( .WIDTH(16) ) _49022_ ( .A(_26394_), .B({ _26394_[15], _26394_[15], _26394_[15], _26394_[15], _26394_[15:4] }), .S(__delay_data_654[2]), .Y({ _26392_[15], _26392_[6:0], _26395_[7:0] }) );
  \$mux  #( .WIDTH(16) ) _49023_ ( .A(_26393_), .B({ _26393_[15], _26393_[15], _26393_[15:2] }), .S(__delay_data_654[1]), .Y(_26394_) );
  \$mux  #( .WIDTH(16) ) _49024_ ( .A(__muladd_madd_odata_reg_125), .B({ __muladd_madd_odata_reg_125[15], __muladd_madd_odata_reg_125[15:1] }), .S(__delay_data_654[0]), .Y(_26393_) );
  \$mux  #( .WIDTH(16) ) _49025_ ( .A({ _26396_[15], _26396_[6:0], _26399_[7:0] }), .B({ _26396_[15], _26396_[15], _26396_[15], _26396_[15], _26396_[15], _26396_[15], _26396_[15], _26396_[15], _26396_[15], _26396_[6:0] }), .S(__delay_data_671[3]), .Y(_25931_) );
  \$mux  #( .WIDTH(16) ) _49026_ ( .A(_26398_), .B({ _26398_[15], _26398_[15], _26398_[15], _26398_[15], _26398_[15:4] }), .S(__delay_data_671[2]), .Y({ _26396_[15], _26396_[6:0], _26399_[7:0] }) );
  \$mux  #( .WIDTH(16) ) _49027_ ( .A(_26397_), .B({ _26397_[15], _26397_[15], _26397_[15:2] }), .S(__delay_data_671[1]), .Y(_26398_) );
  \$mux  #( .WIDTH(16) ) _49028_ ( .A(__muladd_madd_odata_reg_140), .B({ __muladd_madd_odata_reg_140[15], __muladd_madd_odata_reg_140[15:1] }), .S(__delay_data_671[0]), .Y(_26397_) );
  \$mux  #( .WIDTH(16) ) _49029_ ( .A({ _26400_[15], _26400_[6:0], _26403_[7:0] }), .B({ _26400_[15], _26400_[15], _26400_[15], _26400_[15], _26400_[15], _26400_[15], _26400_[15], _26400_[15], _26400_[15], _26400_[6:0] }), .S(__delay_data_688[3]), .Y(_25932_) );
  \$mux  #( .WIDTH(16) ) _49030_ ( .A(_26402_), .B({ _26402_[15], _26402_[15], _26402_[15], _26402_[15], _26402_[15:4] }), .S(__delay_data_688[2]), .Y({ _26400_[15], _26400_[6:0], _26403_[7:0] }) );
  \$mux  #( .WIDTH(16) ) _49031_ ( .A(_26401_), .B({ _26401_[15], _26401_[15], _26401_[15:2] }), .S(__delay_data_688[1]), .Y(_26402_) );
  \$mux  #( .WIDTH(16) ) _49032_ ( .A(__muladd_madd_odata_reg_155), .B({ __muladd_madd_odata_reg_155[15], __muladd_madd_odata_reg_155[15:1] }), .S(__delay_data_688[0]), .Y(_26401_) );
  \$mux  #( .WIDTH(16) ) _49033_ ( .A({ _26404_[15], _26404_[6:0], _26407_[7:0] }), .B({ _26404_[15], _26404_[15], _26404_[15], _26404_[15], _26404_[15], _26404_[15], _26404_[15], _26404_[15], _26404_[15], _26404_[6:0] }), .S(__delay_data_705[3]), .Y(_25933_) );
  \$mux  #( .WIDTH(16) ) _49034_ ( .A(_26406_), .B({ _26406_[15], _26406_[15], _26406_[15], _26406_[15], _26406_[15:4] }), .S(__delay_data_705[2]), .Y({ _26404_[15], _26404_[6:0], _26407_[7:0] }) );
  \$mux  #( .WIDTH(16) ) _49035_ ( .A(_26405_), .B({ _26405_[15], _26405_[15], _26405_[15:2] }), .S(__delay_data_705[1]), .Y(_26406_) );
  \$mux  #( .WIDTH(16) ) _49036_ ( .A(__muladd_madd_odata_reg_170), .B({ __muladd_madd_odata_reg_170[15], __muladd_madd_odata_reg_170[15:1] }), .S(__delay_data_705[0]), .Y(_26405_) );
  \$mux  #( .WIDTH(16) ) _49037_ ( .A({ _26408_[15], _26408_[6:0], _26411_[7:0] }), .B({ _26408_[15], _26408_[15], _26408_[15], _26408_[15], _26408_[15], _26408_[15], _26408_[15], _26408_[15], _26408_[15], _26408_[6:0] }), .S(__delay_data_722[3]), .Y(_25934_) );
  \$mux  #( .WIDTH(16) ) _49038_ ( .A(_26410_), .B({ _26410_[15], _26410_[15], _26410_[15], _26410_[15], _26410_[15:4] }), .S(__delay_data_722[2]), .Y({ _26408_[15], _26408_[6:0], _26411_[7:0] }) );
  \$mux  #( .WIDTH(16) ) _49039_ ( .A(_26409_), .B({ _26409_[15], _26409_[15], _26409_[15:2] }), .S(__delay_data_722[1]), .Y(_26410_) );
  \$mux  #( .WIDTH(16) ) _49040_ ( .A(__muladd_madd_odata_reg_185), .B({ __muladd_madd_odata_reg_185[15], __muladd_madd_odata_reg_185[15:1] }), .S(__delay_data_722[0]), .Y(_26409_) );
  \$mux  #( .WIDTH(1) ) _49041_ ( .A(_26442_), .B(_26443_), .S(_counter_data_762[1]), .Y(_26412_) );
  \$mux  #( .WIDTH(1) ) _49042_ ( .A(_26412_), .B(1'hx), .S(_counter_data_762[2]), .Y(_26413_) );
  \$mux  #( .WIDTH(1) ) _49043_ ( .A(_26413_), .B(1'hx), .S(_counter_data_762[3]), .Y(_26414_) );
  \$mux  #( .WIDTH(1) ) _49044_ ( .A(_26414_), .B(1'hx), .S(_counter_data_762[4]), .Y(_26415_) );
  \$mux  #( .WIDTH(1) ) _49045_ ( .A(_26415_), .B(1'hx), .S(_counter_data_762[5]), .Y(_26416_) );
  \$mux  #( .WIDTH(1) ) _49046_ ( .A(_26416_), .B(1'hx), .S(_counter_data_762[6]), .Y(_26417_) );
  \$mux  #( .WIDTH(1) ) _49047_ ( .A(_26417_), .B(1'hx), .S(_counter_data_762[7]), .Y(_26418_) );
  \$mux  #( .WIDTH(1) ) _49048_ ( .A(_26418_), .B(1'hx), .S(_counter_data_762[8]), .Y(_26419_) );
  \$mux  #( .WIDTH(1) ) _49049_ ( .A(_26419_), .B(1'hx), .S(_counter_data_762[9]), .Y(_26420_) );
  \$mux  #( .WIDTH(1) ) _49050_ ( .A(_26420_), .B(1'hx), .S(_counter_data_762[10]), .Y(_26421_) );
  \$mux  #( .WIDTH(1) ) _49051_ ( .A(_26421_), .B(1'hx), .S(_counter_data_762[11]), .Y(_26422_) );
  \$mux  #( .WIDTH(1) ) _49052_ ( .A(_26422_), .B(1'hx), .S(_counter_data_762[12]), .Y(_26423_) );
  \$mux  #( .WIDTH(1) ) _49053_ ( .A(_26423_), .B(1'hx), .S(_counter_data_762[13]), .Y(_26424_) );
  \$mux  #( .WIDTH(1) ) _49054_ ( .A(_26424_), .B(1'hx), .S(_counter_data_762[14]), .Y(_26425_) );
  \$mux  #( .WIDTH(1) ) _49055_ ( .A(_26425_), .B(1'hx), .S(_counter_data_762[15]), .Y(_26426_) );
  \$mux  #( .WIDTH(1) ) _49056_ ( .A(_26426_), .B(1'hx), .S(_counter_data_762[16]), .Y(_26427_) );
  \$mux  #( .WIDTH(1) ) _49057_ ( .A(_26427_), .B(1'hx), .S(_counter_data_762[17]), .Y(_26428_) );
  \$mux  #( .WIDTH(1) ) _49058_ ( .A(_26428_), .B(1'hx), .S(_counter_data_762[18]), .Y(_26429_) );
  \$mux  #( .WIDTH(1) ) _49059_ ( .A(_26429_), .B(1'hx), .S(_counter_data_762[19]), .Y(_26430_) );
  \$mux  #( .WIDTH(1) ) _49060_ ( .A(_26430_), .B(1'hx), .S(_counter_data_762[20]), .Y(_26431_) );
  \$mux  #( .WIDTH(1) ) _49061_ ( .A(_26431_), .B(1'hx), .S(_counter_data_762[21]), .Y(_26432_) );
  \$mux  #( .WIDTH(1) ) _49062_ ( .A(_26432_), .B(1'hx), .S(_counter_data_762[22]), .Y(_26433_) );
  \$mux  #( .WIDTH(1) ) _49063_ ( .A(_26433_), .B(1'hx), .S(_counter_data_762[23]), .Y(_26434_) );
  \$mux  #( .WIDTH(1) ) _49064_ ( .A(_26434_), .B(1'hx), .S(_counter_data_762[24]), .Y(_26435_) );
  \$mux  #( .WIDTH(1) ) _49065_ ( .A(_26435_), .B(1'hx), .S(_counter_data_762[25]), .Y(_26436_) );
  \$mux  #( .WIDTH(1) ) _49066_ ( .A(_26436_), .B(1'hx), .S(_counter_data_762[26]), .Y(_26437_) );
  \$mux  #( .WIDTH(1) ) _49067_ ( .A(_26437_), .B(1'hx), .S(_counter_data_762[27]), .Y(_26438_) );
  \$mux  #( .WIDTH(1) ) _49068_ ( .A(_26438_), .B(1'hx), .S(_counter_data_762[28]), .Y(_26439_) );
  \$mux  #( .WIDTH(1) ) _49069_ ( .A(_26439_), .B(1'hx), .S(_counter_data_762[29]), .Y(_26440_) );
  \$mux  #( .WIDTH(1) ) _49070_ ( .A(_26440_), .B(1'hx), .S(_counter_data_762[30]), .Y(_26441_) );
  \$mux  #( .WIDTH(1) ) _49071_ ( .A(__delay_data_1372[0]), .B(__delay_data_1372[1]), .S(_counter_data_762[0]), .Y(_26442_) );
  \$mux  #( .WIDTH(1) ) _49072_ ( .A(__delay_data_1372[2]), .B(__delay_data_1372[3]), .S(_counter_data_762[0]), .Y(_26443_) );
  \$mux  #( .WIDTH(8) ) _49141_ ( .A(__tmp_805_1), .B(ram_w8_l2048_id19_0_1_rdata), .S(__tmp_804_1), .Y(_tmp_805) );
  \$mux  #( .WIDTH(8) ) _49142_ ( .A(__tmp_817_1), .B(ram_w8_l2048_id19_1_1_rdata), .S(__tmp_816_1), .Y(_tmp_817) );
  \$mux  #( .WIDTH(8) ) _49143_ ( .A(__tmp_829_1), .B(ram_w8_l2048_id19_2_1_rdata), .S(__tmp_828_1), .Y(_tmp_829) );
  \$mux  #( .WIDTH(8) ) _49144_ ( .A(__tmp_841_1), .B(ram_w8_l2048_id19_3_1_rdata), .S(__tmp_840_1), .Y(_tmp_841) );
  \$mux  #( .WIDTH(32) ) _49145_ ( .A(_26444_), .B(_26445_), .S(_04964_), .Y(_26446_) );
  \$mux  #( .WIDTH(32) ) _49146_ ( .A(1), .B(_26446_), .S(_04885_), .Y({ _26447_[31:1], conv2d_8_mux_next_dma_flag_0 }) );
  \$mux  #( .WIDTH(32) ) _49147_ ( .A(_26444_), .B(0), .S(_04965_), .Y(_26445_) );
  \$mux  #( .WIDTH(32) ) _49148_ ( .A(1), .B(_26445_), .S(_04964_), .Y(_26448_) );
  \$mux  #( .WIDTH(32) ) _49149_ ( .A(_26444_), .B(_26448_), .S(_04885_), .Y({ _26449_[31:1], conv2d_8_mux_next_dma_flag_1 }) );
  \$mux  #( .WIDTH(32) ) _49150_ ( .A(0), .B(1), .S(conv2d_8_update_filter), .Y(_26444_) );
  \$mux  #( .WIDTH(32) ) _49151_ ( .A(1), .B(0), .S(_04965_), .Y(_26450_) );
  \$mux  #( .WIDTH(32) ) _49152_ ( .A(_26444_), .B(_26450_), .S(_04964_), .Y(_26451_) );
  \$mux  #( .WIDTH(32) ) _49153_ ( .A(_26444_), .B(_26451_), .S(_04885_), .Y({ _26452_[31:1], conv2d_8_mux_next_dma_flag_2 }) );
  \$mux  #( .WIDTH(32) ) _49154_ ( .A({ 24'h000000, ram_w8_l2048_id1_3_0_rdata }), .B(0), .S(_04968_), .Y(_26453_) );
  \$mux  #( .WIDTH(32) ) _49155_ ( .A({ 24'h000000, ram_w8_l2048_id1_2_0_rdata }), .B(_26453_), .S(_04967_), .Y(_26454_) );
  \$mux  #( .WIDTH(32) ) _49156_ ( .A({ 24'h000000, ram_w8_l2048_id1_1_0_rdata }), .B(_26454_), .S(_04966_), .Y(_26455_) );
  \$mux  #( .WIDTH(32) ) _49157_ ( .A({ 24'h000000, ram_w8_l2048_id1_0_0_rdata }), .B(_26455_), .S(_04886_), .Y({ _26456_[31:8], _tmp_870 }) );
  \$mux  #( .WIDTH(32) ) _49158_ ( .A({ _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870[7], _tmp_870 }), .B(0), .S(_04995_), .Y({ _26457_[31:8], _stream_max_pool_serial_9_source_1_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49159_ ( .A(0), .B(1), .S(_set_flag_876), .Y({ _26458_[31:1], _stream_max_pool_serial_9_start_flag }) );
  \$mux  #( .WIDTH(8) ) _49160_ ( .A(__tmp_916_1), .B(ram_w8_l2048_id0_0_1_rdata), .S(__tmp_915_1), .Y(_tmp_916) );
  \$mux  #( .WIDTH(8) ) _49161_ ( .A(__tmp_928_1), .B(ram_w8_l2048_id0_1_1_rdata), .S(__tmp_927_1), .Y(_tmp_928) );
  \$mux  #( .WIDTH(8) ) _49162_ ( .A(__tmp_940_1), .B(ram_w8_l2048_id0_2_1_rdata), .S(__tmp_939_1), .Y(_tmp_940) );
  \$mux  #( .WIDTH(8) ) _49163_ ( .A(__tmp_952_1), .B(ram_w8_l2048_id0_3_1_rdata), .S(__tmp_951_1), .Y(_tmp_952) );
  \$mux  #( .WIDTH(32) ) _49164_ ( .A(_22047_), .B(0), .S(matmul_15_row_select), .Y(matmul_15_mux_act_gaddr_0) );
  \$mux  #( .WIDTH(1) ) _49165_ ( .A(matmul_15_dma_pad_mask_0), .B(1'h0), .S(matmul_15_row_select), .Y(matmul_15_mux_dma_pad_mask_0) );
  \$mux  #( .WIDTH(1) ) _49166_ ( .A(matmul_15_dma_flag_0), .B(1'h0), .S(matmul_15_prev_row_select), .Y(matmul_15_mux_dma_flag_0) );
  \$mux  #( .WIDTH(32) ) _49167_ ( .A(ram_w32_l128_id0_0_rdata), .B(0), .S(_05015_), .Y(_stream_matmul_15_source_6_source_ram_rdata) );
  \$mux  #( .WIDTH(32) ) _49168_ ( .A({ 24'h000000, ram_w8_l2048_id0_3_0_rdata }), .B(0), .S(_04971_), .Y(_26459_) );
  \$mux  #( .WIDTH(32) ) _49169_ ( .A({ 24'h000000, ram_w8_l2048_id0_2_0_rdata }), .B(_26459_), .S(_04970_), .Y(_26460_) );
  \$mux  #( .WIDTH(32) ) _49170_ ( .A({ 24'h000000, ram_w8_l2048_id0_1_0_rdata }), .B(_26460_), .S(_04969_), .Y(_26461_) );
  \$mux  #( .WIDTH(32) ) _49171_ ( .A({ 24'h000000, ram_w8_l2048_id0_0_0_rdata }), .B(_26461_), .S(_04887_), .Y({ _26462_[31:8], _tmp_1000 }) );
  \$mux  #( .WIDTH(32) ) _49172_ ( .A({ _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000[7], _tmp_1000 }), .B(0), .S(_04993_), .Y({ _26463_[31:8], _stream_matmul_15_source_8_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49173_ ( .A({ 24'h000000, ram_w8_l2048_id2_3_0_rdata }), .B(0), .S(_04974_), .Y(_26464_) );
  \$mux  #( .WIDTH(32) ) _49174_ ( .A({ 24'h000000, ram_w8_l2048_id2_2_0_rdata }), .B(_26464_), .S(_04973_), .Y(_26465_) );
  \$mux  #( .WIDTH(32) ) _49175_ ( .A({ 24'h000000, ram_w8_l2048_id2_1_0_rdata }), .B(_26465_), .S(_04972_), .Y(_26466_) );
  \$mux  #( .WIDTH(32) ) _49176_ ( .A({ 24'h000000, ram_w8_l2048_id2_0_0_rdata }), .B(_26466_), .S(_04888_), .Y({ _26467_[31:8], _tmp_1020 }) );
  \$mux  #( .WIDTH(32) ) _49177_ ( .A({ _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020[7], _tmp_1020 }), .B(0), .S(_04997_), .Y({ _26468_[31:8], _stream_matmul_15_source_19_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49178_ ( .A({ 24'h000000, ram_w8_l4096_id0_3_0_rdata }), .B(0), .S(_04977_), .Y(_26469_) );
  \$mux  #( .WIDTH(32) ) _49179_ ( .A({ 24'h000000, ram_w8_l4096_id0_2_0_rdata }), .B(_26469_), .S(_04976_), .Y(_26470_) );
  \$mux  #( .WIDTH(32) ) _49180_ ( .A({ 24'h000000, ram_w8_l4096_id0_1_0_rdata }), .B(_26470_), .S(_04975_), .Y(_26471_) );
  \$mux  #( .WIDTH(32) ) _49181_ ( .A({ 24'h000000, ram_w8_l4096_id0_0_0_rdata }), .B(_26471_), .S(_04889_), .Y({ _26472_[31:8], _tmp_1030 }) );
  \$mux  #( .WIDTH(32) ) _49182_ ( .A({ _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030[7], _tmp_1030 }), .B(0), .S(_04991_), .Y({ _26473_[31:8], _stream_matmul_15_source_20_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49183_ ( .A(0), .B(1), .S(_05264_), .Y({ _26474_[31:1], _stream_matmul_15_start_flag }) );
  \$mux  #( .WIDTH(8) ) _49184_ ( .A(__tmp_1125_1), .B(ram_w8_l2048_id1_0_1_rdata), .S(__tmp_1124_1), .Y(_tmp_1125) );
  \$mux  #( .WIDTH(8) ) _49185_ ( .A(__tmp_1137_1), .B(ram_w8_l2048_id1_1_1_rdata), .S(__tmp_1136_1), .Y(_tmp_1137) );
  \$mux  #( .WIDTH(8) ) _49186_ ( .A(__tmp_1149_1), .B(ram_w8_l2048_id1_2_1_rdata), .S(__tmp_1148_1), .Y(_tmp_1149) );
  \$mux  #( .WIDTH(8) ) _49187_ ( .A(__tmp_1161_1), .B(ram_w8_l2048_id1_3_1_rdata), .S(__tmp_1160_1), .Y(_tmp_1161) );
  \$mux  #( .WIDTH(32) ) _49188_ ( .A(0), .B(1), .S(_05267_), .Y(_26475_) );
  \$mux  #( .WIDTH(32) ) _49189_ ( .A(_26475_), .B(1), .S(_05266_), .Y(_26476_) );
  \$mux  #( .WIDTH(32) ) _49190_ ( .A(_26476_), .B(1), .S(_05265_), .Y({ _26477_[31:1], _maxi_write_data_done }) );
  \$mux  #( .WIDTH(32) ) _49191_ ( .A(1), .B(0), .S(_21874_), .Y(_26478_) );
  \$mux  #( .WIDTH(32) ) _49192_ ( .A(1), .B(0), .S(_21875_), .Y(_26479_) );
  \$mux  #( .WIDTH(32) ) _49193_ ( .A(1), .B(0), .S(_21876_), .Y(_26480_) );
  \$mux  #( .WIDTH(32) ) _49194_ ( .A(1), .B(0), .S(_21877_), .Y(_26481_) );
  \$mux  #( .WIDTH(32) ) _49195_ ( .A(1), .B(0), .S(_21878_), .Y(_26482_) );
  \$mux  #( .WIDTH(32) ) _49196_ ( .A(1), .B(0), .S(_21879_), .Y(_26483_) );
  \$mux  #( .WIDTH(32) ) _49197_ ( .A(_saxi_register_13), .B(32'hxxxxxxxx), .S(_04990_), .Y(_26484_) );
  \$mux  #( .WIDTH(32) ) _49198_ ( .A(_saxi_register_12), .B(_26484_), .S(_04989_), .Y(_26485_) );
  \$mux  #( .WIDTH(32) ) _49199_ ( .A(_saxi_register_11), .B(_26485_), .S(_04988_), .Y(_26486_) );
  \$mux  #( .WIDTH(32) ) _49200_ ( .A(_saxi_register_10), .B(_26486_), .S(_04987_), .Y(_26487_) );
  \$mux  #( .WIDTH(32) ) _49201_ ( .A(_saxi_register_9), .B(_26487_), .S(_04986_), .Y(_26488_) );
  \$mux  #( .WIDTH(32) ) _49202_ ( .A(_saxi_register_8), .B(_26488_), .S(_04985_), .Y(_26489_) );
  \$mux  #( .WIDTH(32) ) _49203_ ( .A(_saxi_register_7), .B(_26489_), .S(_04984_), .Y(_26490_) );
  \$mux  #( .WIDTH(32) ) _49204_ ( .A(_saxi_register_6), .B(_26490_), .S(_04983_), .Y(_26491_) );
  \$mux  #( .WIDTH(32) ) _49205_ ( .A(_saxi_register_5), .B(_26491_), .S(_04982_), .Y(_26492_) );
  \$mux  #( .WIDTH(32) ) _49206_ ( .A(_saxi_register_4), .B(_26492_), .S(_04981_), .Y(_26493_) );
  \$mux  #( .WIDTH(32) ) _49207_ ( .A(_saxi_register_3), .B(_26493_), .S(_04980_), .Y(_26494_) );
  \$mux  #( .WIDTH(32) ) _49208_ ( .A(_saxi_register_2), .B(_26494_), .S(_04979_), .Y(_26495_) );
  \$mux  #( .WIDTH(32) ) _49209_ ( .A(_saxi_register_1), .B(_26495_), .S(_04978_), .Y(_26496_) );
  \$mux  #( .WIDTH(32) ) _49210_ ( .A(_saxi_register_0), .B(_26496_), .S(_04890_), .Y(_tmp_6) );
  \$mux  #( .WIDTH(32) ) _49211_ ( .A({ 31'h00000000, _saxi_flag_13 }), .B(32'hxxxxxxxx), .S(_04990_), .Y(_26497_) );
  \$mux  #( .WIDTH(32) ) _49212_ ( .A({ 31'h00000000, _saxi_flag_12 }), .B(_26497_), .S(_04989_), .Y(_26498_) );
  \$mux  #( .WIDTH(32) ) _49213_ ( .A({ 31'h00000000, _saxi_flag_11 }), .B(_26498_), .S(_04988_), .Y(_26499_) );
  \$mux  #( .WIDTH(32) ) _49214_ ( .A({ 31'h00000000, _saxi_flag_10 }), .B(_26499_), .S(_04987_), .Y(_26500_) );
  \$mux  #( .WIDTH(32) ) _49215_ ( .A({ 31'h00000000, _saxi_flag_9 }), .B(_26500_), .S(_04986_), .Y(_26501_) );
  \$mux  #( .WIDTH(32) ) _49216_ ( .A({ 31'h00000000, _saxi_flag_8 }), .B(_26501_), .S(_04985_), .Y(_26502_) );
  \$mux  #( .WIDTH(32) ) _49217_ ( .A({ 31'h00000000, _saxi_flag_7 }), .B(_26502_), .S(_04984_), .Y(_26503_) );
  \$mux  #( .WIDTH(32) ) _49218_ ( .A({ 31'h00000000, _saxi_flag_6 }), .B(_26503_), .S(_04983_), .Y(_26504_) );
  \$mux  #( .WIDTH(32) ) _49219_ ( .A({ 31'h00000000, _saxi_flag_5 }), .B(_26504_), .S(_04982_), .Y(_26505_) );
  \$mux  #( .WIDTH(32) ) _49220_ ( .A({ 31'h00000000, _saxi_flag_4 }), .B(_26505_), .S(_04981_), .Y(_26506_) );
  \$mux  #( .WIDTH(32) ) _49221_ ( .A({ 31'h00000000, _saxi_flag_3 }), .B(_26506_), .S(_04980_), .Y(_26507_) );
  \$mux  #( .WIDTH(32) ) _49222_ ( .A({ 31'h00000000, _saxi_flag_2 }), .B(_26507_), .S(_04979_), .Y(_26508_) );
  \$mux  #( .WIDTH(32) ) _49223_ ( .A({ 31'h00000000, _saxi_flag_1 }), .B(_26508_), .S(_04978_), .Y(_26509_) );
  \$mux  #( .WIDTH(32) ) _49224_ ( .A({ 31'h00000000, _saxi_flag_0 }), .B(_26509_), .S(_04890_), .Y({ _26510_[31:1], _tmp_7 }) );
  \$mux  #( .WIDTH(33) ) _49225_ ( .A(_22123_), .B(33'h000000000), .S(_05233_), .Y(_26511_) );
  \$mux  #( .WIDTH(33) ) _49226_ ( .A(_22124_), .B(33'h000000000), .S(_05234_), .Y(_26512_) );
  \$mux  #( .WIDTH(66) ) _49227_ ( .A(66'h00000000000000000), .B(_sll_data_7), .S(__delay_data_728), .Y(_26513_) );
  \$mux  #( .WIDTH(40) ) _49228_ ( .A(__delay_data_748), .B(40'h000000007f), .S(_greaterthan_data_41), .Y(_26514_) );
  \$mux  #( .WIDTH(40) ) _49229_ ( .A(__delay_data_748), .B(40'hffffffff81), .S(_lessthan_data_45), .Y(_26515_) );
  \$mux  #( .WIDTH(40) ) _49230_ ( .A(_cond_data_47), .B(_cond_data_43), .S(__delay_data_749), .Y(_26516_) );
  \$mux  #( .WIDTH(32) ) _49231_ ( .A(_saxi_resetval_13), .B(32'hxxxxxxxx), .S(_04990_), .Y(_26517_) );
  \$mux  #( .WIDTH(32) ) _49232_ ( .A(_saxi_resetval_12), .B(_26517_), .S(_04989_), .Y(_26518_) );
  \$mux  #( .WIDTH(32) ) _49233_ ( .A(_saxi_resetval_11), .B(_26518_), .S(_04988_), .Y(_26519_) );
  \$mux  #( .WIDTH(32) ) _49234_ ( .A(_saxi_resetval_10), .B(_26519_), .S(_04987_), .Y(_26520_) );
  \$mux  #( .WIDTH(32) ) _49235_ ( .A(_saxi_resetval_9), .B(_26520_), .S(_04986_), .Y(_26521_) );
  \$mux  #( .WIDTH(32) ) _49236_ ( .A(_saxi_resetval_8), .B(_26521_), .S(_04985_), .Y(_26522_) );
  \$mux  #( .WIDTH(32) ) _49237_ ( .A(_saxi_resetval_7), .B(_26522_), .S(_04984_), .Y(_26523_) );
  \$mux  #( .WIDTH(32) ) _49238_ ( .A(_saxi_resetval_6), .B(_26523_), .S(_04983_), .Y(_26524_) );
  \$mux  #( .WIDTH(32) ) _49239_ ( .A(_saxi_resetval_5), .B(_26524_), .S(_04982_), .Y(_26525_) );
  \$mux  #( .WIDTH(32) ) _49240_ ( .A(_saxi_resetval_4), .B(_26525_), .S(_04981_), .Y(_26526_) );
  \$mux  #( .WIDTH(32) ) _49241_ ( .A(_saxi_resetval_3), .B(_26526_), .S(_04980_), .Y(_26527_) );
  \$mux  #( .WIDTH(32) ) _49242_ ( .A(_saxi_resetval_2), .B(_26527_), .S(_04979_), .Y(_26528_) );
  \$mux  #( .WIDTH(32) ) _49243_ ( .A(_saxi_resetval_1), .B(_26528_), .S(_04978_), .Y(_26529_) );
  \$mux  #( .WIDTH(32) ) _49244_ ( .A(_saxi_resetval_0), .B(_26529_), .S(_04890_), .Y(_tmp_8) );
  \$mux  #( .WIDTH(18) ) _49245_ ( .A(18'h00000), .B(_sll_data_59), .S(__delay_data_573), .Y(_26530_) );
  \$mux  #( .WIDTH(18) ) _49246_ ( .A(18'h00000), .B(_sll_data_74), .S(__delay_data_590), .Y(_26531_) );
  \$mux  #( .WIDTH(18) ) _49247_ ( .A(18'h00000), .B(_sll_data_89), .S(__delay_data_607), .Y(_26532_) );
  \$mux  #( .WIDTH(18) ) _49248_ ( .A(18'h00000), .B(_sll_data_104), .S(__delay_data_624), .Y(_26533_) );
  \$mux  #( .WIDTH(18) ) _49249_ ( .A(18'h00000), .B(_sll_data_119), .S(__delay_data_641), .Y(_26534_) );
  \$mux  #( .WIDTH(18) ) _49250_ ( .A(18'h00000), .B(_sll_data_134), .S(__delay_data_658), .Y(_26535_) );
  \$mux  #( .WIDTH(18) ) _49251_ ( .A(18'h00000), .B(_sll_data_149), .S(__delay_data_675), .Y(_26536_) );
  \$mux  #( .WIDTH(18) ) _49252_ ( .A(18'h00000), .B(_sll_data_164), .S(__delay_data_692), .Y(_26537_) );
  \$mux  #( .WIDTH(18) ) _49253_ ( .A(18'h00000), .B(_sll_data_179), .S(__delay_data_709), .Y(_26538_) );
  \$mux  #( .WIDTH(32) ) _49254_ ( .A({ __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187[7], __variable_wdata_187 }), .B(_reducecustom_data_191), .S(_05260_), .Y(_26539_) );
  \$mux  #( .WIDTH(32) ) _49255_ ( .A(_22134_), .B(0), .S(_05236_), .Y(_26540_) );
  \$mux  #( .WIDTH(32) ) _49256_ ( .A(_22135_), .B(0), .S(_05237_), .Y(_26541_) );
  \$mux  #( .WIDTH(32) ) _49257_ ( .A(28), .B(14), .S(conv2d_8_control_param_index), .Y({ _26542_[31:5], cparam_conv2d_8_act_num_row }) );
  \$mux  #( .WIDTH(32) ) _49258_ ( .A(8), .B(6), .S(conv2d_8_control_param_index), .Y({ _26544_[31:4], cparam_conv2d_8_cshamt_out_value }) );
  \$mux  #( .WIDTH(32) ) _49259_ ( .A(27), .B(11), .S(conv2d_8_control_param_index), .Y({ _26547_[31:5], cparam_conv2d_8_max_col_count }) );
  \$mux  #( .WIDTH(32) ) _49260_ ( .A(36), .B(64), .S(conv2d_8_control_param_index), .Y({ _26548_[31:7], cparam_conv2d_8_och_count_step }) );
  \$mux  #( .WIDTH(32) ) _49261_ ( .A(-112), .B(0), .S(conv2d_8_control_param_index), .Y(cparam_conv2d_8_act_offset_values_0) );
  \$mux  #( .WIDTH(32) ) _49262_ ( .A(0), .B(224), .S(conv2d_8_control_param_index), .Y(cparam_conv2d_8_act_offset_values_1) );
  \$mux  #( .WIDTH(32) ) _49263_ ( .A(112), .B(448), .S(conv2d_8_control_param_index), .Y(cparam_conv2d_8_act_offset_values_2) );
  \$mux  #( .WIDTH(32) ) _49264_ ( .A(112), .B(224), .S(conv2d_8_control_param_index), .Y({ _26549_[31:8], cparam_conv2d_8_act_read_size }) );
  \$mux  #( .WIDTH(32) ) _49265_ ( .A(40), .B(80), .S(conv2d_8_control_param_index), .Y({ _26551_[31:7], cparam_conv2d_8_act_read_step }) );
  \$mux  #( .WIDTH(32) ) _49266_ ( .A(576), .B(1152), .S(conv2d_8_control_param_index), .Y({ _26552_[31:11], cparam_conv2d_8_filter_base_step }) );
  \$mux  #( .WIDTH(32) ) _49267_ ( .A(64), .B(128), .S(conv2d_8_control_param_index), .Y({ _26553_[31:8], cparam_conv2d_8_filter_read_step }) );
  \$mux  #( .WIDTH(32) ) _49268_ ( .A(448), .B(96), .S(conv2d_8_control_param_index), .Y({ _26554_[31:9], cparam_conv2d_8_out_row_step }) );
  \$mux  #( .WIDTH(32) ) _49269_ ( .A(1), .B(16), .S(conv2d_8_control_param_index), .Y({ _26555_[31:5], cparam_conv2d_8_stream_reduce_size }) );
  \$mux  #( .WIDTH(32) ) _49270_ ( .A(2), .B(0), .S(conv2d_8_control_param_index), .Y({ _26556_[31:2], cparam_conv2d_8_col_select_initval }) );
  \$mux  #( .WIDTH(32) ) _49271_ ( .A(4), .B(16), .S(conv2d_8_control_param_index), .Y({ _26550_[31:5], cparam_conv2d_8_inc_act_laddr_large }) );
  \$mux  #( .WIDTH(32) ) _49272_ ( .A(16), .B(8), .S(conv2d_8_control_param_index), .Y({ _26543_[31:5], cparam_conv2d_8_bias_num }) );
  \$mux  #( .WIDTH(32) ) _49273_ ( .A(-4), .B(0), .S(conv2d_8_control_param_index), .Y({ _26557_[31:4], cparam_conv2d_8_stream_act_local_large_offset }) );
  \$mux  #( .WIDTH(32) ) _49274_ ( .A(1), .B(0), .S(conv2d_8_control_param_index), .Y({ _26546_[31:1], cparam_conv2d_8_pad_col_left }) );
  \$mux  #( .WIDTH(32) ) _49275_ ( .A(28), .B(12), .S(conv2d_8_control_param_index), .Y({ _26545_[31:5], cparam_conv2d_8_inc_sync_out }) );
  \$mux  #( .WIDTH(32) ) _49276_ ( .A(28), .B(12), .S(max_pool_serial_9_control_param_index), .Y({ _26558_[31:5], cparam_max_pool_serial_9_act_num_col }) );
  \$mux  #( .WIDTH(32) ) _49277_ ( .A(25), .B(9), .S(max_pool_serial_9_control_param_index), .Y({ _26559_[31:5], cparam_max_pool_serial_9_max_col_count }) );
  \$mux  #( .WIDTH(32) ) _49278_ ( .A(896), .B(192), .S(max_pool_serial_9_control_param_index), .Y({ _26560_[31:10], cparam_max_pool_serial_9_act_row_step }) );
  \$mux  #( .WIDTH(32) ) _49279_ ( .A(448), .B(96), .S(max_pool_serial_9_control_param_index), .Y(cparam_max_pool_serial_9_act_offset_values_1) );
  \$mux  #( .WIDTH(32) ) _49280_ ( .A(224), .B(48), .S(max_pool_serial_9_control_param_index), .Y({ _26562_[31:8], cparam_max_pool_serial_9_out_row_step }) );
  \$mux  #( .WIDTH(32) ) _49281_ ( .A(32), .B(16), .S(max_pool_serial_9_control_param_index), .Y({ _26563_[31:6], cparam_max_pool_serial_9_inc_act_laddr }) );
  \$mux  #( .WIDTH(32) ) _49282_ ( .A(16), .B(8), .S(max_pool_serial_9_control_param_index), .Y({ _26561_[31:5], cparam_max_pool_serial_9_inc_out_laddr }) );
  \$mux  #( .WIDTH(8) ) _49283_ ( .A(8'h00), .B(__delay_data_868), .S(_eq_data_337), .Y(_26564_) );
  \$mux  #( .WIDTH(8) ) _49284_ ( .A(8'h00), .B(__delay_data_874), .S(_eq_data_337), .Y(_26565_) );
  \$mux  #( .WIDTH(8) ) _49285_ ( .A(8'h00), .B(__delay_data_870), .S(_eq_data_337), .Y(_26566_) );
  \$mux  #( .WIDTH(8) ) _49286_ ( .A(8'h00), .B(__delay_data_877), .S(_eq_data_337), .Y(_26567_) );
  \$mux  #( .WIDTH(8) ) _49287_ ( .A(8'h00), .B(__delay_data_883), .S(_eq_data_337), .Y(_26568_) );
  \$mux  #( .WIDTH(8) ) _49288_ ( .A(8'h00), .B(__delay_data_879), .S(_eq_data_337), .Y(_26569_) );
  \$mux  #( .WIDTH(8) ) _49289_ ( .A(8'h00), .B(__delay_data_886), .S(_eq_data_337), .Y(_26570_) );
  \$mux  #( .WIDTH(8) ) _49290_ ( .A(8'h00), .B(__delay_data_892), .S(_eq_data_337), .Y(_26571_) );
  \$mux  #( .WIDTH(8) ) _49291_ ( .A(8'h00), .B(__delay_data_888), .S(_eq_data_337), .Y(_26572_) );
  \$mux  #( .WIDTH(8) ) _49292_ ( .A(_cond_data_259), .B(__delay_data_871), .S(__delay_data_869), .Y(_26573_) );
  \$mux  #( .WIDTH(8) ) _49293_ ( .A(_cond_data_269), .B(__delay_data_932), .S(__delay_data_869), .Y(_26574_) );
  \$mux  #( .WIDTH(8) ) _49294_ ( .A(_cond_data_279), .B(__delay_data_875), .S(__delay_data_869), .Y(_26575_) );
  \$mux  #( .WIDTH(8) ) _49295_ ( .A(_cond_data_289), .B(__delay_data_880), .S(__delay_data_869), .Y(_26576_) );
  \$mux  #( .WIDTH(8) ) _49296_ ( .A(_cond_data_299), .B(__delay_data_937), .S(__delay_data_869), .Y(_26577_) );
  \$mux  #( .WIDTH(8) ) _49297_ ( .A(_cond_data_309), .B(__delay_data_884), .S(__delay_data_869), .Y(_26578_) );
  \$mux  #( .WIDTH(8) ) _49298_ ( .A(_cond_data_319), .B(__delay_data_889), .S(__delay_data_869), .Y(_26579_) );
  \$mux  #( .WIDTH(8) ) _49299_ ( .A(_cond_data_329), .B(__delay_data_942), .S(__delay_data_869), .Y(_26580_) );
  \$mux  #( .WIDTH(8) ) _49300_ ( .A(_cond_data_339), .B(__delay_data_893), .S(__delay_data_869), .Y(_26581_) );
  \$mux  #( .WIDTH(8) ) _49301_ ( .A(_cond_data_263), .B(__delay_data_876), .S(__delay_data_991), .Y(_26582_) );
  \$mux  #( .WIDTH(8) ) _49302_ ( .A(_cond_data_273), .B(__delay_data_935), .S(__delay_data_991), .Y(_26583_) );
  \$mux  #( .WIDTH(8) ) _49303_ ( .A(_cond_data_283), .B(__delay_data_984), .S(__delay_data_991), .Y(_26584_) );
  \$mux  #( .WIDTH(8) ) _49304_ ( .A(_cond_data_293), .B(__delay_data_885), .S(__delay_data_991), .Y(_26585_) );
  \$mux  #( .WIDTH(8) ) _49305_ ( .A(_cond_data_303), .B(__delay_data_940), .S(__delay_data_991), .Y(_26586_) );
  \$mux  #( .WIDTH(8) ) _49306_ ( .A(_cond_data_313), .B(__delay_data_988), .S(__delay_data_991), .Y(_26587_) );
  \$mux  #( .WIDTH(8) ) _49307_ ( .A(_cond_data_323), .B(__delay_data_894), .S(__delay_data_991), .Y(_26588_) );
  \$mux  #( .WIDTH(8) ) _49308_ ( .A(_cond_data_333), .B(__delay_data_945), .S(__delay_data_991), .Y(_26589_) );
  \$mux  #( .WIDTH(8) ) _49309_ ( .A(_cond_data_343), .B(__delay_data_992), .S(__delay_data_991), .Y(_26590_) );
  \$mux  #( .WIDTH(8) ) _49310_ ( .A(8'h00), .B(_cond_data_326), .S(__delay_data_1198), .Y(_26591_) );
  \$mux  #( .WIDTH(8) ) _49311_ ( .A(8'h00), .B(_cond_data_266), .S(__delay_data_1198), .Y(_26592_) );
  \$mux  #( .WIDTH(8) ) _49312_ ( .A(8'h00), .B(_cond_data_296), .S(__delay_data_1198), .Y(_26593_) );
  \$mux  #( .WIDTH(8) ) _49313_ ( .A(8'h00), .B(_cond_data_336), .S(__delay_data_1198), .Y(_26594_) );
  \$mux  #( .WIDTH(8) ) _49314_ ( .A(8'h00), .B(_cond_data_276), .S(__delay_data_1198), .Y(_26595_) );
  \$mux  #( .WIDTH(8) ) _49315_ ( .A(8'h00), .B(_cond_data_306), .S(__delay_data_1198), .Y(_26596_) );
  \$mux  #( .WIDTH(8) ) _49316_ ( .A(8'h00), .B(_cond_data_346), .S(__delay_data_1198), .Y(_26597_) );
  \$mux  #( .WIDTH(8) ) _49317_ ( .A(8'h00), .B(_cond_data_286), .S(__delay_data_1198), .Y(_26598_) );
  \$mux  #( .WIDTH(8) ) _49318_ ( .A(8'h00), .B(_cond_data_316), .S(__delay_data_1198), .Y(_26599_) );
  \$mux  #( .WIDTH(8) ) _49319_ ( .A(_cond_data_349), .B(__delay_data_902), .S(__delay_data_1202), .Y(_26600_) );
  \$mux  #( .WIDTH(8) ) _49320_ ( .A(_cond_data_359), .B(__delay_data_1035), .S(__delay_data_1202), .Y(_26601_) );
  \$mux  #( .WIDTH(8) ) _49321_ ( .A(_cond_data_369), .B(__delay_data_908), .S(__delay_data_1202), .Y(_26602_) );
  \$mux  #( .WIDTH(8) ) _49322_ ( .A(_cond_data_379), .B(__delay_data_953), .S(__delay_data_1202), .Y(_26603_) );
  \$mux  #( .WIDTH(8) ) _49323_ ( .A(_cond_data_389), .B(__delay_data_1069), .S(__delay_data_1202), .Y(_26604_) );
  \$mux  #( .WIDTH(8) ) _49324_ ( .A(_cond_data_399), .B(__delay_data_959), .S(__delay_data_1202), .Y(_26605_) );
  \$mux  #( .WIDTH(8) ) _49325_ ( .A(_cond_data_409), .B(__delay_data_1000), .S(__delay_data_1202), .Y(_26606_) );
  \$mux  #( .WIDTH(8) ) _49326_ ( .A(_cond_data_419), .B(__delay_data_1103), .S(__delay_data_1202), .Y(_26607_) );
  \$mux  #( .WIDTH(8) ) _49327_ ( .A(_cond_data_429), .B(__delay_data_1006), .S(__delay_data_1202), .Y(_26608_) );
  \$mux  #( .WIDTH(8) ) _49328_ ( .A(_cond_data_353), .B(__delay_data_909), .S(__delay_data_1207), .Y(_26609_) );
  \$mux  #( .WIDTH(8) ) _49329_ ( .A(_cond_data_363), .B(__delay_data_1041), .S(__delay_data_1207), .Y(_26610_) );
  \$mux  #( .WIDTH(8) ) _49330_ ( .A(_cond_data_373), .B(__delay_data_1142), .S(__delay_data_1207), .Y(_26611_) );
  \$mux  #( .WIDTH(8) ) _49331_ ( .A(_cond_data_383), .B(__delay_data_960), .S(__delay_data_1207), .Y(_26612_) );
  \$mux  #( .WIDTH(8) ) _49332_ ( .A(_cond_data_393), .B(__delay_data_1075), .S(__delay_data_1207), .Y(_26613_) );
  \$mux  #( .WIDTH(8) ) _49333_ ( .A(_cond_data_403), .B(__delay_data_1175), .S(__delay_data_1207), .Y(_26614_) );
  \$mux  #( .WIDTH(8) ) _49334_ ( .A(_cond_data_413), .B(__delay_data_1007), .S(__delay_data_1207), .Y(_26615_) );
  \$mux  #( .WIDTH(8) ) _49335_ ( .A(_cond_data_423), .B(__delay_data_1109), .S(__delay_data_1207), .Y(_26616_) );
  \$mux  #( .WIDTH(8) ) _49336_ ( .A(_cond_data_433), .B(__delay_data_1208), .S(__delay_data_1207), .Y(_26617_) );
  \$mux  #( .WIDTH(8) ) _49337_ ( .A(_cond_data_356), .B(8'h00), .S(__delay_data_915), .Y(_26618_) );
  \$mux  #( .WIDTH(8) ) _49338_ ( .A(_cond_data_386), .B(8'h00), .S(__delay_data_966), .Y(_26619_) );
  \$mux  #( .WIDTH(8) ) _49339_ ( .A(_cond_data_416), .B(8'h00), .S(__delay_data_1013), .Y(_26620_) );
  \$mux  #( .WIDTH(8) ) _49340_ ( .A(_cond_data_366), .B(8'h00), .S(__delay_data_1047), .Y(_26621_) );
  \$mux  #( .WIDTH(8) ) _49341_ ( .A(_cond_data_396), .B(8'h00), .S(__delay_data_1081), .Y(_26622_) );
  \$mux  #( .WIDTH(8) ) _49342_ ( .A(_cond_data_426), .B(8'h00), .S(__delay_data_1115), .Y(_26623_) );
  \$mux  #( .WIDTH(8) ) _49343_ ( .A(_cond_data_376), .B(8'h00), .S(__delay_data_1148), .Y(_26624_) );
  \$mux  #( .WIDTH(8) ) _49344_ ( .A(_cond_data_406), .B(8'h00), .S(__delay_data_1181), .Y(_26625_) );
  \$mux  #( .WIDTH(8) ) _49345_ ( .A(_cond_data_436), .B(8'h00), .S(__delay_data_1214), .Y(_26626_) );
  \$mux  #( .WIDTH(8) ) _49346_ ( .A(8'h00), .B(__delay_data_1358), .S(_greaterthan_data_753), .Y(_26627_) );
  \$mux  #( .WIDTH(32) ) _49347_ ( .A(0), .B(conv2d_8_och_count_buf), .S(_05016_), .Y(_26628_) );
  \$mux  #( .WIDTH(32) ) _49348_ ( .A(0), .B(1), .S(_05016_), .Y(_26629_) );
  \$mux  #( .WIDTH(32) ) _49349_ ( .A(_22232_), .B(0), .S(_05238_), .Y(_26630_) );
  \$mux  #( .WIDTH(9) ) _49350_ ( .A({ __delay_data_1374[7], __delay_data_1374 }), .B(9'h180), .S(_pointer_data_764), .Y(_26631_) );
  \$mux  #( .WIDTH(8) ) _49351_ ( .A(8'h00), .B(__delay_data_1378), .S(_eq_data_831), .Y(_26632_) );
  \$mux  #( .WIDTH(8) ) _49352_ ( .A(8'h00), .B(_cond_data_833), .S(__delay_data_1379), .Y(_26633_) );
  \$mux  #( .WIDTH(8) ) _49353_ ( .A(_cond_data_837), .B(8'h00), .S(__delay_data_1381), .Y(_26634_) );
  \$mux  #( .WIDTH(32) ) _49354_ ( .A(1), .B(0), .S(_04895_), .Y({ _21969_, _21968_, _21966_, _21965_, _21964_, _21963_, _21962_, _21961_, _21960_, _21959_, _21958_, _21957_, _21955_, _21954_, _21953_, _21952_, _21951_, _21950_, _21949_, _21948_, _21947_, _21946_, _21976_, _21975_, _21974_, _21973_, _21972_, _21971_, _21970_, _21967_, _21956_, _21945_ }) );
  \$mux  #( .WIDTH(32) ) _49355_ ( .A(1), .B(0), .S(_05017_), .Y(_26635_) );
  \$mux  #( .WIDTH(32) ) _49356_ ( .A(0), .B(_26635_), .S(_04895_), .Y({ _22001_, _22000_, _21998_, _21997_, _21996_, _21995_, _21994_, _21993_, _21992_, _21991_, _21990_, _21989_, _21987_, _21986_, _21985_, _21984_, _21983_, _21982_, _21981_, _21980_, _21979_, _21978_, _22008_, _22007_, _22006_, _22005_, _22004_, _22003_, _22002_, _21999_, _21988_, _21977_ }) );
  \$mux  #( .WIDTH(32) ) _49357_ ( .A(1), .B(0), .S(_05018_), .Y(_26636_) );
  \$mux  #( .WIDTH(32) ) _49358_ ( .A(0), .B(_26636_), .S(_05017_), .Y(_26637_) );
  \$mux  #( .WIDTH(32) ) _49359_ ( .A(0), .B(_26637_), .S(_04895_), .Y({ _22033_, _22032_, _22030_, _22029_, _22028_, _22027_, _22026_, _22025_, _22024_, _22023_, _22022_, _22021_, _22019_, _22018_, _22017_, _22016_, _22015_, _22014_, _22013_, _22012_, _22011_, _22010_, _22040_, _22039_, _22038_, _22037_, _22036_, _22035_, _22034_, _22031_, _22020_, _22009_ }) );
  \$mux  #( .WIDTH(32) ) _49360_ ( .A(_22358_), .B(0), .S(_04965_), .Y(_26638_) );
  \$mux  #( .WIDTH(32) ) _49361_ ( .A(_22356_), .B(_26638_), .S(_04964_), .Y(_26639_) );
  \$mux  #( .WIDTH(32) ) _49362_ ( .A(_22354_), .B(_26639_), .S(_04885_), .Y(conv2d_8_mux_act_gaddr_0) );
  \$mux  #( .WIDTH(32) ) _49363_ ( .A(_22356_), .B(0), .S(_04965_), .Y(_26640_) );
  \$mux  #( .WIDTH(32) ) _49364_ ( .A(_22354_), .B(_26640_), .S(_04964_), .Y(_26641_) );
  \$mux  #( .WIDTH(32) ) _49365_ ( .A(_22358_), .B(_26641_), .S(_04885_), .Y(conv2d_8_mux_act_gaddr_1) );
  \$mux  #( .WIDTH(32) ) _49366_ ( .A(_22354_), .B(0), .S(_04965_), .Y(_26642_) );
  \$mux  #( .WIDTH(32) ) _49367_ ( .A(_22358_), .B(_26642_), .S(_04964_), .Y(_26643_) );
  \$mux  #( .WIDTH(32) ) _49368_ ( .A(_22356_), .B(_26643_), .S(_04885_), .Y(conv2d_8_mux_act_gaddr_2) );
  \$mux  #( .WIDTH(1) ) _49369_ ( .A(conv2d_8_dma_pad_mask_1), .B(1'h0), .S(_04965_), .Y(_26644_) );
  \$mux  #( .WIDTH(1) ) _49370_ ( .A(conv2d_8_dma_pad_mask_2), .B(_26644_), .S(_04964_), .Y(_26645_) );
  \$mux  #( .WIDTH(1) ) _49371_ ( .A(conv2d_8_dma_pad_mask_0), .B(_26645_), .S(_04885_), .Y(conv2d_8_mux_dma_pad_mask_0) );
  \$mux  #( .WIDTH(1) ) _49372_ ( .A(conv2d_8_dma_pad_mask_2), .B(1'h0), .S(_04965_), .Y(_26646_) );
  \$mux  #( .WIDTH(1) ) _49373_ ( .A(conv2d_8_dma_pad_mask_0), .B(_26646_), .S(_04964_), .Y(_26647_) );
  \$mux  #( .WIDTH(1) ) _49374_ ( .A(conv2d_8_dma_pad_mask_1), .B(_26647_), .S(_04885_), .Y(conv2d_8_mux_dma_pad_mask_1) );
  \$mux  #( .WIDTH(1) ) _49375_ ( .A(conv2d_8_dma_pad_mask_0), .B(1'h0), .S(_04965_), .Y(_26648_) );
  \$mux  #( .WIDTH(1) ) _49376_ ( .A(conv2d_8_dma_pad_mask_1), .B(_26648_), .S(_04964_), .Y(_26649_) );
  \$mux  #( .WIDTH(1) ) _49377_ ( .A(conv2d_8_dma_pad_mask_2), .B(_26649_), .S(_04885_), .Y(conv2d_8_mux_dma_pad_mask_2) );
  \$mux  #( .WIDTH(1) ) _49378_ ( .A(conv2d_8_dma_flag_1), .B(1'h0), .S(_04906_), .Y(_26650_) );
  \$mux  #( .WIDTH(1) ) _49379_ ( .A(conv2d_8_dma_flag_2), .B(_26650_), .S(_04905_), .Y(_26651_) );
  \$mux  #( .WIDTH(1) ) _49380_ ( .A(conv2d_8_dma_flag_0), .B(_26651_), .S(_04865_), .Y(conv2d_8_mux_dma_flag_0) );
  \$mux  #( .WIDTH(1) ) _49381_ ( .A(conv2d_8_dma_flag_2), .B(1'h0), .S(_04906_), .Y(_26652_) );
  \$mux  #( .WIDTH(1) ) _49382_ ( .A(conv2d_8_dma_flag_0), .B(_26652_), .S(_04905_), .Y(_26653_) );
  \$mux  #( .WIDTH(1) ) _49383_ ( .A(conv2d_8_dma_flag_1), .B(_26653_), .S(_04865_), .Y(conv2d_8_mux_dma_flag_1) );
  \$mux  #( .WIDTH(1) ) _49384_ ( .A(conv2d_8_dma_flag_0), .B(1'h0), .S(_04906_), .Y(_26654_) );
  \$mux  #( .WIDTH(1) ) _49385_ ( .A(conv2d_8_dma_flag_1), .B(_26654_), .S(_04905_), .Y(_26655_) );
  \$mux  #( .WIDTH(1) ) _49386_ ( .A(conv2d_8_dma_flag_2), .B(_26655_), .S(_04865_), .Y(conv2d_8_mux_dma_flag_2) );
  \$mux  #( .WIDTH(32) ) _49387_ ( .A(ram_w32_l128_id0_0_rdata), .B(0), .S(_05014_), .Y(_stream_conv2d_8_source_6_source_ram_rdata) );
  \$mux  #( .WIDTH(32) ) _49388_ ( .A({ 24'h000000, ram_w8_l2048_id0_3_0_rdata }), .B(0), .S(_04909_), .Y(_26656_) );
  \$mux  #( .WIDTH(32) ) _49389_ ( .A({ 24'h000000, ram_w8_l2048_id0_2_0_rdata }), .B(_26656_), .S(_04908_), .Y(_26657_) );
  \$mux  #( .WIDTH(32) ) _49390_ ( .A({ 24'h000000, ram_w8_l2048_id0_1_0_rdata }), .B(_26657_), .S(_04907_), .Y(_26658_) );
  \$mux  #( .WIDTH(32) ) _49391_ ( .A({ 24'h000000, ram_w8_l2048_id0_0_0_rdata }), .B(_26658_), .S(_04866_), .Y({ _26659_[31:8], _tmp_344 }) );
  \$mux  #( .WIDTH(32) ) _49392_ ( .A({ _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344[7], _tmp_344 }), .B(0), .S(_04992_), .Y({ _26660_[31:8], _stream_conv2d_8_source_8_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49393_ ( .A({ 24'h000000, ram_w8_l2048_id10_3_0_rdata }), .B(0), .S(_04912_), .Y(_26661_) );
  \$mux  #( .WIDTH(32) ) _49394_ ( .A({ 24'h000000, ram_w8_l2048_id10_2_0_rdata }), .B(_26661_), .S(_04911_), .Y(_26662_) );
  \$mux  #( .WIDTH(32) ) _49395_ ( .A({ 24'h000000, ram_w8_l2048_id10_1_0_rdata }), .B(_26662_), .S(_04910_), .Y(_26663_) );
  \$mux  #( .WIDTH(32) ) _49396_ ( .A({ 24'h000000, ram_w8_l2048_id10_0_0_rdata }), .B(_26663_), .S(_04867_), .Y({ _26664_[31:8], _tmp_364 }) );
  \$mux  #( .WIDTH(32) ) _49397_ ( .A({ _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364[7], _tmp_364 }), .B(0), .S(_05005_), .Y({ _26665_[31:8], _stream_conv2d_8_source_19_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49398_ ( .A({ 24'h000000, ram_w8_l2048_id11_3_0_rdata }), .B(0), .S(_04915_), .Y(_26666_) );
  \$mux  #( .WIDTH(32) ) _49399_ ( .A({ 24'h000000, ram_w8_l2048_id11_2_0_rdata }), .B(_26666_), .S(_04914_), .Y(_26667_) );
  \$mux  #( .WIDTH(32) ) _49400_ ( .A({ 24'h000000, ram_w8_l2048_id11_1_0_rdata }), .B(_26667_), .S(_04913_), .Y(_26668_) );
  \$mux  #( .WIDTH(32) ) _49401_ ( .A({ 24'h000000, ram_w8_l2048_id11_0_0_rdata }), .B(_26668_), .S(_04868_), .Y({ _26669_[31:8], _tmp_374 }) );
  \$mux  #( .WIDTH(32) ) _49402_ ( .A({ _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374[7], _tmp_374 }), .B(0), .S(_05006_), .Y({ _26670_[31:8], _stream_conv2d_8_source_20_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49403_ ( .A({ 24'h000000, ram_w8_l2048_id12_3_0_rdata }), .B(0), .S(_04918_), .Y(_26671_) );
  \$mux  #( .WIDTH(32) ) _49404_ ( .A({ 24'h000000, ram_w8_l2048_id12_2_0_rdata }), .B(_26671_), .S(_04917_), .Y(_26672_) );
  \$mux  #( .WIDTH(32) ) _49405_ ( .A({ 24'h000000, ram_w8_l2048_id12_1_0_rdata }), .B(_26672_), .S(_04916_), .Y(_26673_) );
  \$mux  #( .WIDTH(32) ) _49406_ ( .A({ 24'h000000, ram_w8_l2048_id12_0_0_rdata }), .B(_26673_), .S(_04869_), .Y({ _26674_[31:8], _tmp_384 }) );
  \$mux  #( .WIDTH(32) ) _49407_ ( .A({ _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384[7], _tmp_384 }), .B(0), .S(_05007_), .Y({ _26675_[31:8], _stream_conv2d_8_source_21_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49408_ ( .A({ 24'h000000, ram_w8_l2048_id13_3_0_rdata }), .B(0), .S(_04921_), .Y(_26676_) );
  \$mux  #( .WIDTH(32) ) _49409_ ( .A({ 24'h000000, ram_w8_l2048_id13_2_0_rdata }), .B(_26676_), .S(_04920_), .Y(_26677_) );
  \$mux  #( .WIDTH(32) ) _49410_ ( .A({ 24'h000000, ram_w8_l2048_id13_1_0_rdata }), .B(_26677_), .S(_04919_), .Y(_26678_) );
  \$mux  #( .WIDTH(32) ) _49411_ ( .A({ 24'h000000, ram_w8_l2048_id13_0_0_rdata }), .B(_26678_), .S(_04870_), .Y({ _26679_[31:8], _tmp_394 }) );
  \$mux  #( .WIDTH(32) ) _49412_ ( .A({ _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394[7], _tmp_394 }), .B(0), .S(_05008_), .Y({ _26680_[31:8], _stream_conv2d_8_source_22_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49413_ ( .A({ 24'h000000, ram_w8_l2048_id14_3_0_rdata }), .B(0), .S(_04924_), .Y(_26681_) );
  \$mux  #( .WIDTH(32) ) _49414_ ( .A({ 24'h000000, ram_w8_l2048_id14_2_0_rdata }), .B(_26681_), .S(_04923_), .Y(_26682_) );
  \$mux  #( .WIDTH(32) ) _49415_ ( .A({ 24'h000000, ram_w8_l2048_id14_1_0_rdata }), .B(_26682_), .S(_04922_), .Y(_26683_) );
  \$mux  #( .WIDTH(32) ) _49416_ ( .A({ 24'h000000, ram_w8_l2048_id14_0_0_rdata }), .B(_26683_), .S(_04871_), .Y({ _26684_[31:8], _tmp_404 }) );
  \$mux  #( .WIDTH(32) ) _49417_ ( .A({ _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404[7], _tmp_404 }), .B(0), .S(_05009_), .Y({ _26685_[31:8], _stream_conv2d_8_source_23_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49418_ ( .A({ 24'h000000, ram_w8_l2048_id15_3_0_rdata }), .B(0), .S(_04927_), .Y(_26686_) );
  \$mux  #( .WIDTH(32) ) _49419_ ( .A({ 24'h000000, ram_w8_l2048_id15_2_0_rdata }), .B(_26686_), .S(_04926_), .Y(_26687_) );
  \$mux  #( .WIDTH(32) ) _49420_ ( .A({ 24'h000000, ram_w8_l2048_id15_1_0_rdata }), .B(_26687_), .S(_04925_), .Y(_26688_) );
  \$mux  #( .WIDTH(32) ) _49421_ ( .A({ 24'h000000, ram_w8_l2048_id15_0_0_rdata }), .B(_26688_), .S(_04872_), .Y({ _26689_[31:8], _tmp_414 }) );
  \$mux  #( .WIDTH(32) ) _49422_ ( .A({ _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414[7], _tmp_414 }), .B(0), .S(_05010_), .Y({ _26690_[31:8], _stream_conv2d_8_source_24_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49423_ ( .A({ 24'h000000, ram_w8_l2048_id16_3_0_rdata }), .B(0), .S(_04930_), .Y(_26691_) );
  \$mux  #( .WIDTH(32) ) _49424_ ( .A({ 24'h000000, ram_w8_l2048_id16_2_0_rdata }), .B(_26691_), .S(_04929_), .Y(_26692_) );
  \$mux  #( .WIDTH(32) ) _49425_ ( .A({ 24'h000000, ram_w8_l2048_id16_1_0_rdata }), .B(_26692_), .S(_04928_), .Y(_26693_) );
  \$mux  #( .WIDTH(32) ) _49426_ ( .A({ 24'h000000, ram_w8_l2048_id16_0_0_rdata }), .B(_26693_), .S(_04873_), .Y({ _26694_[31:8], _tmp_424 }) );
  \$mux  #( .WIDTH(32) ) _49427_ ( .A({ _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424[7], _tmp_424 }), .B(0), .S(_05011_), .Y({ _26695_[31:8], _stream_conv2d_8_source_25_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49428_ ( .A({ 24'h000000, ram_w8_l2048_id17_3_0_rdata }), .B(0), .S(_04933_), .Y(_26696_) );
  \$mux  #( .WIDTH(32) ) _49429_ ( .A({ 24'h000000, ram_w8_l2048_id17_2_0_rdata }), .B(_26696_), .S(_04932_), .Y(_26697_) );
  \$mux  #( .WIDTH(32) ) _49430_ ( .A({ 24'h000000, ram_w8_l2048_id17_1_0_rdata }), .B(_26697_), .S(_04931_), .Y(_26698_) );
  \$mux  #( .WIDTH(32) ) _49431_ ( .A({ 24'h000000, ram_w8_l2048_id17_0_0_rdata }), .B(_26698_), .S(_04874_), .Y({ _26699_[31:8], _tmp_434 }) );
  \$mux  #( .WIDTH(32) ) _49432_ ( .A({ _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434[7], _tmp_434 }), .B(0), .S(_05012_), .Y({ _26700_[31:8], _stream_conv2d_8_source_26_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49433_ ( .A({ 24'h000000, ram_w8_l2048_id18_3_0_rdata }), .B(0), .S(_04936_), .Y(_26701_) );
  \$mux  #( .WIDTH(32) ) _49434_ ( .A({ 24'h000000, ram_w8_l2048_id18_2_0_rdata }), .B(_26701_), .S(_04935_), .Y(_26702_) );
  \$mux  #( .WIDTH(32) ) _49435_ ( .A({ 24'h000000, ram_w8_l2048_id18_1_0_rdata }), .B(_26702_), .S(_04934_), .Y(_26703_) );
  \$mux  #( .WIDTH(32) ) _49436_ ( .A({ 24'h000000, ram_w8_l2048_id18_0_0_rdata }), .B(_26703_), .S(_04875_), .Y({ _26704_[31:8], _tmp_444 }) );
  \$mux  #( .WIDTH(32) ) _49437_ ( .A({ _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444[7], _tmp_444 }), .B(0), .S(_05013_), .Y({ _26705_[31:8], _stream_conv2d_8_source_27_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49438_ ( .A({ 24'h000000, ram_w8_l2048_id1_3_0_rdata }), .B(0), .S(_04939_), .Y(_26706_) );
  \$mux  #( .WIDTH(32) ) _49439_ ( .A({ 24'h000000, ram_w8_l2048_id1_2_0_rdata }), .B(_26706_), .S(_04938_), .Y(_26707_) );
  \$mux  #( .WIDTH(32) ) _49440_ ( .A({ 24'h000000, ram_w8_l2048_id1_1_0_rdata }), .B(_26707_), .S(_04937_), .Y(_26708_) );
  \$mux  #( .WIDTH(32) ) _49441_ ( .A({ 24'h000000, ram_w8_l2048_id1_0_0_rdata }), .B(_26708_), .S(_04876_), .Y({ _26709_[31:8], _tmp_454 }) );
  \$mux  #( .WIDTH(32) ) _49442_ ( .A({ _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454[7], _tmp_454 }), .B(0), .S(_04994_), .Y({ _26710_[31:8], _stream_conv2d_8_source_28_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49443_ ( .A({ 24'h000000, ram_w8_l2048_id2_3_0_rdata }), .B(0), .S(_04942_), .Y(_26711_) );
  \$mux  #( .WIDTH(32) ) _49444_ ( .A({ 24'h000000, ram_w8_l2048_id2_2_0_rdata }), .B(_26711_), .S(_04941_), .Y(_26712_) );
  \$mux  #( .WIDTH(32) ) _49445_ ( .A({ 24'h000000, ram_w8_l2048_id2_1_0_rdata }), .B(_26712_), .S(_04940_), .Y(_26713_) );
  \$mux  #( .WIDTH(32) ) _49446_ ( .A({ 24'h000000, ram_w8_l2048_id2_0_0_rdata }), .B(_26713_), .S(_04877_), .Y({ _26714_[31:8], _tmp_464 }) );
  \$mux  #( .WIDTH(32) ) _49447_ ( .A({ _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464[7], _tmp_464 }), .B(0), .S(_04996_), .Y({ _26715_[31:8], _stream_conv2d_8_source_29_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49448_ ( .A({ 24'h000000, ram_w8_l2048_id3_1_0_rdata }), .B(_26719_), .S(_04943_), .Y(_26716_) );
  \$mux  #( .WIDTH(32) ) _49449_ ( .A({ 24'h000000, ram_w8_l2048_id3_0_0_rdata }), .B(_26716_), .S(_04878_), .Y({ _26717_[31:8], _tmp_474 }) );
  \$mux  #( .WIDTH(32) ) _49450_ ( .A({ 24'h000000, ram_w8_l2048_id3_3_0_rdata }), .B(0), .S(_04945_), .Y(_26718_) );
  \$mux  #( .WIDTH(32) ) _49451_ ( .A({ 24'h000000, ram_w8_l2048_id3_2_0_rdata }), .B(_26718_), .S(_04944_), .Y(_26719_) );
  \$mux  #( .WIDTH(32) ) _49452_ ( .A({ _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474[7], _tmp_474 }), .B(0), .S(_04998_), .Y({ _26720_[31:8], _stream_conv2d_8_source_30_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49453_ ( .A({ 24'h000000, ram_w8_l2048_id4_3_0_rdata }), .B(0), .S(_04948_), .Y(_26721_) );
  \$mux  #( .WIDTH(32) ) _49454_ ( .A({ 24'h000000, ram_w8_l2048_id4_2_0_rdata }), .B(_26721_), .S(_04947_), .Y(_26722_) );
  \$mux  #( .WIDTH(32) ) _49455_ ( .A({ 24'h000000, ram_w8_l2048_id4_1_0_rdata }), .B(_26722_), .S(_04946_), .Y(_26723_) );
  \$mux  #( .WIDTH(32) ) _49456_ ( .A({ 24'h000000, ram_w8_l2048_id4_0_0_rdata }), .B(_26723_), .S(_04879_), .Y({ _26724_[31:8], _tmp_484 }) );
  \$mux  #( .WIDTH(32) ) _49457_ ( .A({ _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484[7], _tmp_484 }), .B(0), .S(_04999_), .Y({ _26725_[31:8], _stream_conv2d_8_source_31_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49458_ ( .A({ 24'h000000, ram_w8_l2048_id5_3_0_rdata }), .B(0), .S(_04951_), .Y(_26726_) );
  \$mux  #( .WIDTH(32) ) _49459_ ( .A({ 24'h000000, ram_w8_l2048_id5_2_0_rdata }), .B(_26726_), .S(_04950_), .Y(_26727_) );
  \$mux  #( .WIDTH(32) ) _49460_ ( .A({ 24'h000000, ram_w8_l2048_id5_1_0_rdata }), .B(_26727_), .S(_04949_), .Y(_26728_) );
  \$mux  #( .WIDTH(32) ) _49461_ ( .A({ 24'h000000, ram_w8_l2048_id5_0_0_rdata }), .B(_26728_), .S(_04880_), .Y({ _26729_[31:8], _tmp_494 }) );
  \$mux  #( .WIDTH(32) ) _49462_ ( .A({ _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494[7], _tmp_494 }), .B(0), .S(_05000_), .Y({ _26730_[31:8], _stream_conv2d_8_source_32_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49463_ ( .A({ 24'h000000, ram_w8_l2048_id6_3_0_rdata }), .B(0), .S(_04954_), .Y(_26731_) );
  \$mux  #( .WIDTH(32) ) _49464_ ( .A({ 24'h000000, ram_w8_l2048_id6_2_0_rdata }), .B(_26731_), .S(_04953_), .Y(_26732_) );
  \$mux  #( .WIDTH(32) ) _49465_ ( .A({ 24'h000000, ram_w8_l2048_id6_1_0_rdata }), .B(_26732_), .S(_04952_), .Y(_26733_) );
  \$mux  #( .WIDTH(32) ) _49466_ ( .A({ 24'h000000, ram_w8_l2048_id6_0_0_rdata }), .B(_26733_), .S(_04881_), .Y({ _26734_[31:8], _tmp_504 }) );
  \$mux  #( .WIDTH(32) ) _49467_ ( .A({ _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504[7], _tmp_504 }), .B(0), .S(_05001_), .Y({ _26735_[31:8], _stream_conv2d_8_source_33_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49468_ ( .A({ 24'h000000, ram_w8_l2048_id7_3_0_rdata }), .B(0), .S(_04957_), .Y(_26736_) );
  \$mux  #( .WIDTH(32) ) _49469_ ( .A({ 24'h000000, ram_w8_l2048_id7_2_0_rdata }), .B(_26736_), .S(_04956_), .Y(_26737_) );
  \$mux  #( .WIDTH(32) ) _49470_ ( .A({ 24'h000000, ram_w8_l2048_id7_1_0_rdata }), .B(_26737_), .S(_04955_), .Y(_26738_) );
  \$mux  #( .WIDTH(32) ) _49471_ ( .A({ 24'h000000, ram_w8_l2048_id7_0_0_rdata }), .B(_26738_), .S(_04882_), .Y({ _26739_[31:8], _tmp_514 }) );
  \$mux  #( .WIDTH(32) ) _49472_ ( .A({ _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514[7], _tmp_514 }), .B(0), .S(_05002_), .Y({ _26740_[31:8], _stream_conv2d_8_source_34_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49473_ ( .A({ 24'h000000, ram_w8_l2048_id8_3_0_rdata }), .B(0), .S(_04960_), .Y(_26741_) );
  \$mux  #( .WIDTH(32) ) _49474_ ( .A({ 24'h000000, ram_w8_l2048_id8_2_0_rdata }), .B(_26741_), .S(_04959_), .Y(_26742_) );
  \$mux  #( .WIDTH(32) ) _49475_ ( .A({ 24'h000000, ram_w8_l2048_id8_1_0_rdata }), .B(_26742_), .S(_04958_), .Y(_26743_) );
  \$mux  #( .WIDTH(32) ) _49476_ ( .A({ 24'h000000, ram_w8_l2048_id8_0_0_rdata }), .B(_26743_), .S(_04883_), .Y({ _26744_[31:8], _tmp_524 }) );
  \$mux  #( .WIDTH(32) ) _49477_ ( .A({ _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524[7], _tmp_524 }), .B(0), .S(_05003_), .Y({ _26745_[31:8], _stream_conv2d_8_source_35_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49478_ ( .A({ 24'h000000, ram_w8_l2048_id9_3_0_rdata }), .B(0), .S(_04963_), .Y(_26746_) );
  \$mux  #( .WIDTH(32) ) _49479_ ( .A({ 24'h000000, ram_w8_l2048_id9_2_0_rdata }), .B(_26746_), .S(_04962_), .Y(_26747_) );
  \$mux  #( .WIDTH(32) ) _49480_ ( .A({ 24'h000000, ram_w8_l2048_id9_1_0_rdata }), .B(_26747_), .S(_04961_), .Y(_26748_) );
  \$mux  #( .WIDTH(32) ) _49481_ ( .A({ 24'h000000, ram_w8_l2048_id9_0_0_rdata }), .B(_26748_), .S(_04884_), .Y({ _26749_[31:8], _tmp_534 }) );
  \$mux  #( .WIDTH(32) ) _49482_ ( .A({ _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534[7], _tmp_534 }), .B(0), .S(_05004_), .Y({ _26750_[31:8], _stream_conv2d_8_source_36_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _49483_ ( .A(0), .B(1), .S(_05863_), .Y({ _26751_[31:1], _stream_conv2d_8_start_flag }) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37773_ ( .CLK(CLK), .D(_22456_), .Q(_stream_matmul_15_sink_21_sink_fsm_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37774_ ( .CLK(CLK), .D(_22457_), .Q(_stream_matmul_15_source_20_source_pat_fsm_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37775_ ( .CLK(CLK), .D(_stream_matmul_15_source_20_source_ram_raddr[1:0]), .Q(__tmp_1025_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37776_ ( .CLK(CLK), .D(__tmp_1025_1), .Q(__tmp_1025_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37777_ ( .CLK(CLK), .D(_22458_), .Q(_stream_matmul_15_source_19_source_pat_fsm_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37778_ ( .CLK(CLK), .D(_22459_), .Q(_stream_matmul_15_source_8_source_pat_fsm_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37779_ ( .CLK(CLK), .D(_22460_), .Q(_stream_matmul_15_source_6_source_pat_fsm_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37780_ ( .CLK(CLK), .D(_22475_), .Q(matmul_15_next_stream_num_ops), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37781_ ( .CLK(CLK), .D(_22474_), .Q(matmul_15_sync_comp_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37782_ ( .CLK(CLK), .D(_22472_), .Q(matmul_15_col_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) matmul_15_col_select_reg ( .CLK(CLK), .D(_22471_), .Q(matmul_15_col_select), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37784_ ( .CLK(CLK), .D(_22470_), .Q(matmul_15_stream_act_local_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37785_ ( .CLK(CLK), .D(_22469_), .Q(matmul_15_stream_out_local_col), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37786_ ( .CLK(CLK), .D(_22468_), .Q(matmul_15_comp_fsm), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37787_ ( .CLK(CLK), .D(_22467_), .Q(matmul_15_filter_page_comp_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37788_ ( .CLK(CLK), .D(_22466_), .Q(matmul_15_act_page_comp_offset_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37789_ ( .CLK(CLK), .D(_22465_), .Q(matmul_15_out_page_comp_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37790_ ( .CLK(CLK), .D(_22464_), .Q(matmul_15_row_count_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) matmul_15_row_select_buf_reg ( .CLK(CLK), .D(_22463_), .Q(matmul_15_row_select_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37792_ ( .CLK(CLK), .D(_22462_), .Q(matmul_15_och_count_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) matmul_15_stream_pad_masks_reg ( .CLK(CLK), .D(_22461_), .Q(matmul_15_stream_pad_masks), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37794_ ( .CLK(CLK), .D(_22529_), .Q(control_matmul_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37795_ ( .CLK(CLK), .D(_22528_), .Q(matmul_15_act_base_offset_row), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37796_ ( .CLK(CLK), .D(_22527_), .Q(matmul_15_act_base_offset_bat), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37797_ ( .CLK(CLK), .D(_22526_), .Q(matmul_15_filter_base_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37798_ ( .CLK(CLK), .D(_22525_), .Q(matmul_15_out_base_offset_val), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37799_ ( .CLK(CLK), .D(_22524_), .Q(matmul_15_out_base_offset_col), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37800_ ( .CLK(CLK), .D(_22523_), .Q(matmul_15_out_base_offset_row), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37801_ ( .CLK(CLK), .D(_22522_), .Q(matmul_15_out_base_offset_bat), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37802_ ( .CLK(CLK), .D(_22521_), .Q(matmul_15_out_base_offset_och), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) matmul_15_dma_flag_0_reg ( .CLK(CLK), .D(_22520_), .Q(matmul_15_dma_flag_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37804_ ( .CLK(CLK), .D(_22519_), .Q(matmul_15_sync_out_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37805_ ( .CLK(CLK), .D(_22518_), .Q(matmul_15_next_out_write_size), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37806_ ( .CLK(CLK), .D(_22517_), .Q(matmul_15_row_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37807_ ( .CLK(CLK), .D(_22516_), .Q(matmul_15_bat_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37808_ ( .CLK(CLK), .D(_22515_), .Q(matmul_15_och_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) matmul_15_row_select_reg ( .CLK(CLK), .D(_22514_), .Q(matmul_15_row_select), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37810_ ( .CLK(CLK), .D(_22513_), .Q(matmul_15_out_row_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37811_ ( .CLK(CLK), .D(_22512_), .Q(matmul_15_out_ram_select), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37812_ ( .CLK(CLK), .D(_22511_), .Q(matmul_15_prev_row_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37813_ ( .CLK(CLK), .D(_22510_), .Q(matmul_15_prev_bat_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37814_ ( .CLK(CLK), .D(_22509_), .Q(matmul_15_prev_och_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) matmul_15_prev_row_select_reg ( .CLK(CLK), .D(_22508_), .Q(matmul_15_prev_row_select), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37816_ ( .CLK(CLK), .D(_22507_), .Q(matmul_15_act_page_comp_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37817_ ( .CLK(CLK), .D(_22506_), .Q(matmul_15_act_page_dma_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37818_ ( .CLK(CLK), .D(_22505_), .Q(matmul_15_filter_page_comp_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37819_ ( .CLK(CLK), .D(_22504_), .Q(matmul_15_filter_page_dma_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) matmul_15_out_page_reg ( .CLK(CLK), .D(_22503_), .Q(matmul_15_out_page), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37821_ ( .CLK(CLK), .D(_22502_), .Q(matmul_15_out_page_comp_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37822_ ( .CLK(CLK), .D(_22501_), .Q(matmul_15_out_page_dma_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37823_ ( .CLK(CLK), .D(_22500_), .Q(matmul_15_out_laddr_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) matmul_15_skip_read_filter_reg ( .CLK(CLK), .D(_22499_), .Q(matmul_15_skip_read_filter), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) matmul_15_skip_read_act_reg ( .CLK(CLK), .D(_22498_), .Q(matmul_15_skip_read_act), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) matmul_15_skip_comp_reg ( .CLK(CLK), .D(_22497_), .Q(matmul_15_skip_comp), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) matmul_15_skip_write_out_reg  ( .CLK(CLK), .D(_03133_), .Q(matmul_15_skip_write_out) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_959_reg ( .CLK(CLK), .D(_22495_), .Q(axim_flag_959), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37829_ ( .CLK(CLK), .D(control_matmul_15), .Q(_d1_control_matmul_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_matmul_15_cond_3_0_1_reg ( .CLK(CLK), .D(_22492_), .Q(_control_matmul_15_cond_3_0_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_960_reg ( .CLK(CLK), .D(_22491_), .Q(axim_flag_960), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_matmul_15_cond_8_1_1_reg ( .CLK(CLK), .D(_22488_), .Q(_control_matmul_15_cond_8_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_961_reg ( .CLK(CLK), .D(_22487_), .Q(axim_flag_961), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_matmul_15_cond_14_2_1_reg ( .CLK(CLK), .D(_22484_), .Q(_control_matmul_15_cond_14_2_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_972_reg ( .CLK(CLK), .D(_22483_), .Q(axim_flag_972), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_matmul_15_cond_22_3_1_reg ( .CLK(CLK), .D(_22480_), .Q(_control_matmul_15_cond_22_3_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_1118_reg ( .CLK(CLK), .D(_22479_), .Q(axim_flag_1118), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_matmul_15_cond_32_4_1_reg ( .CLK(CLK), .D(_22476_), .Q(_control_matmul_15_cond_32_4_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37839_ ( .CLK(CLK), .D(_22534_), .Q(_stream_max_pool_serial_9_sink_3_sink_fsm_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37840_ ( .CLK(CLK), .D(_22535_), .Q(_stream_max_pool_serial_9_source_1_source_pat_fsm_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37841_ ( .CLK(CLK), .D(_22545_), .Q(max_pool_serial_9_col_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37842_ ( .CLK(CLK), .D(_22544_), .Q(max_pool_serial_9_stream_act_local), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37843_ ( .CLK(CLK), .D(_22543_), .Q(max_pool_serial_9_stream_out_local), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37844_ ( .CLK(CLK), .D(_22542_), .Q(max_pool_serial_9_comp_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37845_ ( .CLK(CLK), .D(_22540_), .Q(max_pool_serial_9_comp_fsm), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37846_ ( .CLK(CLK), .D(_22539_), .Q(max_pool_serial_9_act_page_comp_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37847_ ( .CLK(CLK), .D(_22538_), .Q(max_pool_serial_9_out_page_comp_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37848_ ( .CLK(CLK), .D(_22537_), .Q(max_pool_serial_9_row_count_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _37849_ ( .CLK(CLK), .D(_22536_), .Q(max_pool_serial_9_stream_pad_masks), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37850_ ( .CLK(CLK), .D(_22578_), .Q(control_max_pool_serial_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37851_ ( .CLK(CLK), .D(_22576_), .Q(max_pool_serial_9_act_base_offset_row), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37852_ ( .CLK(CLK), .D(_22575_), .Q(max_pool_serial_9_act_base_offset_bat), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37853_ ( .CLK(CLK), .D(_22574_), .Q(max_pool_serial_9_out_base_offset_row), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37854_ ( .CLK(CLK), .D(_22572_), .Q(max_pool_serial_9_out_base_offset_bat), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37855_ ( .CLK(CLK), .D(_22571_), .Q(max_pool_serial_9_row_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37856_ ( .CLK(CLK), .D(_22570_), .Q(max_pool_serial_9_bat_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37857_ ( .CLK(CLK), .D(_22569_), .Q(max_pool_serial_9_prev_row_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37858_ ( .CLK(CLK), .D(_22568_), .Q(max_pool_serial_9_prev_bat_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) max_pool_serial_9_act_page_reg ( .CLK(CLK), .D(_22567_), .Q(max_pool_serial_9_act_page), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37860_ ( .CLK(CLK), .D(_22566_), .Q(max_pool_serial_9_act_page_comp_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37861_ ( .CLK(CLK), .D(_22565_), .Q(max_pool_serial_9_act_page_dma_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) max_pool_serial_9_out_page_reg ( .CLK(CLK), .D(_22564_), .Q(max_pool_serial_9_out_page), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37863_ ( .CLK(CLK), .D(_22563_), .Q(max_pool_serial_9_out_page_comp_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37864_ ( .CLK(CLK), .D(_22562_), .Q(max_pool_serial_9_out_page_dma_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) max_pool_serial_9_skip_read_act_reg ( .CLK(CLK), .D(_22561_), .Q(max_pool_serial_9_skip_read_act), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) max_pool_serial_9_skip_comp_reg ( .CLK(CLK), .D(_22560_), .Q(max_pool_serial_9_skip_comp), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) max_pool_serial_9_skip_write_out_reg ( .CLK(CLK), .D(_22559_), .Q(max_pool_serial_9_skip_write_out), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37868_ ( .CLK(CLK), .D(_22558_), .Q(max_pool_serial_9_out_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_850_reg ( .CLK(CLK), .D(_22557_), .Q(axim_flag_850), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37870_ ( .CLK(CLK), .D(control_max_pool_serial_9), .Q(_d1_control_max_pool_serial_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_max_pool_serial_9_cond_5_0_1_reg ( .CLK(CLK), .D(_22554_), .Q(_control_max_pool_serial_9_cond_5_0_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_861_reg ( .CLK(CLK), .D(_22553_), .Q(axim_flag_861), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_max_pool_serial_9_cond_11_1_1_reg ( .CLK(CLK), .D(_22550_), .Q(_control_max_pool_serial_9_cond_11_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_909_reg ( .CLK(CLK), .D(_22549_), .Q(axim_flag_909), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_max_pool_serial_9_cond_19_2_1_reg ( .CLK(CLK), .D(_22546_), .Q(_control_max_pool_serial_9_cond_19_2_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37876_ ( .CLK(CLK), .D(_22594_), .Q(_maxi_write_fsm), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37877_ ( .CLK(CLK), .D(_22593_), .Q(_maxi_write_cur_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _37878_ ( .CLK(CLK), .D(_22592_), .Q(_maxi_write_cur_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _37879_ ( .CLK(CLK), .D(_22588_), .Q(_maxi_write_rest_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_849_reg ( .CLK(CLK), .D(_22585_), .Q(axim_flag_849), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37881_ ( .CLK(CLK), .D(_maxi_write_fsm), .Q(_d1__maxi_write_fsm), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __maxi_write_fsm_cond_4_0_1_reg ( .CLK(CLK), .D(_22582_), .Q(__maxi_write_fsm_cond_4_0_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37883_ ( .CLK(CLK), .D(_22599_), .Q(_stream_conv2d_8_sink_37_sink_fsm_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37884_ ( .CLK(CLK), .D(_22600_), .Q(_stream_conv2d_8_source_36_source_pat_fsm_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37885_ ( .CLK(CLK), .D(_stream_conv2d_8_source_36_source_ram_raddr[1:0]), .Q(__tmp_529_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37886_ ( .CLK(CLK), .D(__tmp_529_1), .Q(__tmp_529_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37887_ ( .CLK(CLK), .D(_22601_), .Q(_stream_conv2d_8_source_35_source_pat_fsm_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37888_ ( .CLK(CLK), .D(_stream_conv2d_8_source_35_source_ram_raddr[1:0]), .Q(__tmp_519_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37889_ ( .CLK(CLK), .D(__tmp_519_1), .Q(__tmp_519_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37890_ ( .CLK(CLK), .D(_22602_), .Q(_stream_conv2d_8_source_34_source_pat_fsm_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37891_ ( .CLK(CLK), .D(_stream_conv2d_8_source_34_source_ram_raddr[1:0]), .Q(__tmp_509_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37892_ ( .CLK(CLK), .D(__tmp_509_1), .Q(__tmp_509_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37893_ ( .CLK(CLK), .D(_22603_), .Q(_stream_conv2d_8_source_33_source_pat_fsm_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37894_ ( .CLK(CLK), .D(_stream_conv2d_8_source_33_source_ram_raddr[1:0]), .Q(__tmp_499_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37895_ ( .CLK(CLK), .D(__tmp_499_1), .Q(__tmp_499_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37896_ ( .CLK(CLK), .D(_22604_), .Q(_stream_conv2d_8_source_32_source_pat_fsm_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37897_ ( .CLK(CLK), .D(_stream_conv2d_8_source_32_source_ram_raddr[1:0]), .Q(__tmp_489_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37898_ ( .CLK(CLK), .D(__tmp_489_1), .Q(__tmp_489_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37899_ ( .CLK(CLK), .D(_22605_), .Q(_stream_conv2d_8_source_31_source_pat_fsm_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37900_ ( .CLK(CLK), .D(_stream_conv2d_8_source_31_source_ram_raddr[1:0]), .Q(__tmp_479_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37901_ ( .CLK(CLK), .D(__tmp_479_1), .Q(__tmp_479_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37902_ ( .CLK(CLK), .D(_22606_), .Q(_stream_conv2d_8_source_30_source_pat_fsm_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37903_ ( .CLK(CLK), .D(_stream_conv2d_8_source_30_source_ram_raddr[1:0]), .Q(__tmp_469_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37904_ ( .CLK(CLK), .D(__tmp_469_1), .Q(__tmp_469_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37905_ ( .CLK(CLK), .D(_22607_), .Q(_stream_conv2d_8_source_29_source_pat_fsm_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37906_ ( .CLK(CLK), .D(_stream_conv2d_8_source_29_source_ram_raddr[1:0]), .Q(__tmp_459_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37907_ ( .CLK(CLK), .D(__tmp_459_1), .Q(__tmp_459_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37908_ ( .CLK(CLK), .D(_stream_matmul_15_source_19_source_ram_raddr[1:0]), .Q(__tmp_1015_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37909_ ( .CLK(CLK), .D(__tmp_1015_1), .Q(__tmp_1015_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37910_ ( .CLK(CLK), .D(_22608_), .Q(_stream_conv2d_8_source_28_source_pat_fsm_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37911_ ( .CLK(CLK), .D(_stream_conv2d_8_source_28_source_ram_raddr[1:0]), .Q(__tmp_449_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37912_ ( .CLK(CLK), .D(__tmp_449_1), .Q(__tmp_449_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37913_ ( .CLK(CLK), .D(_stream_max_pool_serial_9_source_1_source_ram_raddr[1:0]), .Q(__tmp_865_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37914_ ( .CLK(CLK), .D(__tmp_865_1), .Q(__tmp_865_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37915_ ( .CLK(CLK), .D(_22609_), .Q(_stream_conv2d_8_source_27_source_pat_fsm_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37916_ ( .CLK(CLK), .D(_stream_conv2d_8_source_27_source_ram_raddr[1:0]), .Q(__tmp_439_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37917_ ( .CLK(CLK), .D(__tmp_439_1), .Q(__tmp_439_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37918_ ( .CLK(CLK), .D(_22610_), .Q(_stream_conv2d_8_source_26_source_pat_fsm_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37919_ ( .CLK(CLK), .D(_stream_conv2d_8_source_26_source_ram_raddr[1:0]), .Q(__tmp_429_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37920_ ( .CLK(CLK), .D(__tmp_429_1), .Q(__tmp_429_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37921_ ( .CLK(CLK), .D(_22611_), .Q(_stream_conv2d_8_source_25_source_pat_fsm_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37922_ ( .CLK(CLK), .D(_stream_conv2d_8_source_25_source_ram_raddr[1:0]), .Q(__tmp_419_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37923_ ( .CLK(CLK), .D(__tmp_419_1), .Q(__tmp_419_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37924_ ( .CLK(CLK), .D(_22612_), .Q(_stream_conv2d_8_source_24_source_pat_fsm_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37925_ ( .CLK(CLK), .D(_stream_conv2d_8_source_24_source_ram_raddr[1:0]), .Q(__tmp_409_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37926_ ( .CLK(CLK), .D(__tmp_409_1), .Q(__tmp_409_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37927_ ( .CLK(CLK), .D(_22613_), .Q(_stream_conv2d_8_source_23_source_pat_fsm_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37928_ ( .CLK(CLK), .D(_stream_conv2d_8_source_23_source_ram_raddr[1:0]), .Q(__tmp_399_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37929_ ( .CLK(CLK), .D(__tmp_399_1), .Q(__tmp_399_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37930_ ( .CLK(CLK), .D(_22614_), .Q(_stream_conv2d_8_source_22_source_pat_fsm_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37931_ ( .CLK(CLK), .D(_stream_conv2d_8_source_22_source_ram_raddr[1:0]), .Q(__tmp_389_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37932_ ( .CLK(CLK), .D(__tmp_389_1), .Q(__tmp_389_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37933_ ( .CLK(CLK), .D(_22615_), .Q(_stream_conv2d_8_source_21_source_pat_fsm_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37934_ ( .CLK(CLK), .D(_stream_conv2d_8_source_21_source_ram_raddr[1:0]), .Q(__tmp_379_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37935_ ( .CLK(CLK), .D(__tmp_379_1), .Q(__tmp_379_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37936_ ( .CLK(CLK), .D(_22616_), .Q(_stream_conv2d_8_source_20_source_pat_fsm_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37937_ ( .CLK(CLK), .D(_stream_conv2d_8_source_20_source_ram_raddr[1:0]), .Q(__tmp_369_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37938_ ( .CLK(CLK), .D(__tmp_369_1), .Q(__tmp_369_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37939_ ( .CLK(CLK), .D(_22617_), .Q(_stream_conv2d_8_source_19_source_pat_fsm_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37940_ ( .CLK(CLK), .D(_stream_conv2d_8_source_19_source_ram_raddr[1:0]), .Q(__tmp_359_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37941_ ( .CLK(CLK), .D(__tmp_359_1), .Q(__tmp_359_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37942_ ( .CLK(CLK), .D(_22618_), .Q(_stream_conv2d_8_source_8_source_pat_fsm_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37943_ ( .CLK(CLK), .D(_stream_conv2d_8_source_8_source_ram_raddr[1:0]), .Q(__tmp_339_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37944_ ( .CLK(CLK), .D(__tmp_339_1), .Q(__tmp_339_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37945_ ( .CLK(CLK), .D(_stream_matmul_15_source_8_source_ram_raddr[1:0]), .Q(__tmp_995_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37946_ ( .CLK(CLK), .D(__tmp_995_1), .Q(__tmp_995_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37947_ ( .CLK(CLK), .D(_22619_), .Q(_stream_conv2d_8_source_6_source_pat_fsm_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37948_ ( .CLK(CLK), .D(_22657_), .Q(conv2d_8_next_stream_num_ops), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37949_ ( .CLK(CLK), .D(_22656_), .Q(conv2d_8_sync_comp_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37950_ ( .CLK(CLK), .D(_22654_), .Q(conv2d_8_col_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37951_ ( .CLK(CLK), .D(_22653_), .Q(conv2d_8_col_select), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37952_ ( .CLK(CLK), .D(_22651_), .Q(conv2d_8_stream_act_local_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37953_ ( .CLK(CLK), .D(_22649_), .Q(conv2d_8_stream_act_local_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37954_ ( .CLK(CLK), .D(_22647_), .Q(conv2d_8_stream_act_local_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37955_ ( .CLK(CLK), .D(_22644_), .Q(conv2d_8_stream_act_local_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37956_ ( .CLK(CLK), .D(_22642_), .Q(conv2d_8_stream_act_local_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37957_ ( .CLK(CLK), .D(_22640_), .Q(conv2d_8_stream_act_local_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37958_ ( .CLK(CLK), .D(_22637_), .Q(conv2d_8_stream_act_local_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37959_ ( .CLK(CLK), .D(_22635_), .Q(conv2d_8_stream_act_local_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37960_ ( .CLK(CLK), .D(_22633_), .Q(conv2d_8_stream_act_local_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37961_ ( .CLK(CLK), .D(_22630_), .Q(conv2d_8_stream_out_local_col), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37962_ ( .CLK(CLK), .D(_22629_), .Q(conv2d_8_comp_fsm), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37963_ ( .CLK(CLK), .D(_22628_), .Q(conv2d_8_filter_page_comp_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37964_ ( .CLK(CLK), .D(_22627_), .Q(conv2d_8_act_page_comp_offset_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37965_ ( .CLK(CLK), .D(_22626_), .Q(conv2d_8_act_page_comp_offset_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37966_ ( .CLK(CLK), .D(_22625_), .Q(conv2d_8_act_page_comp_offset_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37967_ ( .CLK(CLK), .D(_22624_), .Q(conv2d_8_out_page_comp_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37968_ ( .CLK(CLK), .D(_22623_), .Q(conv2d_8_row_count_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _37969_ ( .CLK(CLK), .D(_22622_), .Q(conv2d_8_row_select_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37970_ ( .CLK(CLK), .D(_22621_), .Q(conv2d_8_och_count_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _37971_ ( .CLK(CLK), .D(_22620_), .Q(conv2d_8_stream_pad_masks), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _37972_ ( .CLK(CLK), .D(_22658_), .Q(req_block_size_270), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _37973_ ( .CLK(CLK), .D(_22659_), .Q(req_block_size_213), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _37974_ ( .CLK(CLK), .D(_22660_), .Q(req_block_size_156), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _37975_ ( .CLK(CLK), .D(_22661_), .Q(req_block_size_27), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37976_ ( .CLK(CLK), .D(_22737_), .Q(_maxi_read_fsm), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37977_ ( .CLK(CLK), .D(_22736_), .Q(_maxi_read_cur_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _37978_ ( .CLK(CLK), .D(_22735_), .Q(_maxi_read_cur_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _37979_ ( .CLK(CLK), .D(_22731_), .Q(_maxi_read_rest_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37980_ ( .CLK(CLK), .D(_22728_), .Q(_wdata_10), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _wvalid_11_reg ( .CLK(CLK), .D(_22726_), .Q(_wvalid_11), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37982_ ( .CLK(CLK), .D(_maxi_read_fsm), .Q(_d1__maxi_read_fsm), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __maxi_read_fsm_cond_3_0_1_reg ( .CLK(CLK), .D(_22722_), .Q(__maxi_read_fsm_cond_3_0_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_15_reg ( .CLK(CLK), .D(_22721_), .Q(axim_flag_15), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __maxi_read_fsm_cond_4_1_1_reg ( .CLK(CLK), .D(_22718_), .Q(__maxi_read_fsm_cond_4_1_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37986_ ( .CLK(CLK), .D(_22717_), .Q(_wdata_17), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _wvalid_18_reg ( .CLK(CLK), .D(_22715_), .Q(_wvalid_18), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __maxi_read_fsm_cond_3_2_1_reg ( .CLK(CLK), .D(_22711_), .Q(__maxi_read_fsm_cond_3_2_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37989_ ( .CLK(CLK), .D(_22710_), .Q(_wdata_30), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _wvalid_31_reg ( .CLK(CLK), .D(_22708_), .Q(_wvalid_31), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __maxi_read_fsm_cond_3_3_1_reg ( .CLK(CLK), .D(_22704_), .Q(__maxi_read_fsm_cond_3_3_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37992_ ( .CLK(CLK), .D(_22703_), .Q(_wdata_159), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _wvalid_160_reg ( .CLK(CLK), .D(_22701_), .Q(_wvalid_160), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __maxi_read_fsm_cond_3_4_1_reg ( .CLK(CLK), .D(_22697_), .Q(__maxi_read_fsm_cond_3_4_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37995_ ( .CLK(CLK), .D(_22696_), .Q(_wdata_216), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _wvalid_217_reg ( .CLK(CLK), .D(_22694_), .Q(_wvalid_217), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __maxi_read_fsm_cond_3_5_1_reg ( .CLK(CLK), .D(_22690_), .Q(__maxi_read_fsm_cond_3_5_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _37998_ ( .CLK(CLK), .D(_22689_), .Q(_wdata_273), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _wvalid_274_reg ( .CLK(CLK), .D(_22687_), .Q(_wvalid_274), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __maxi_read_fsm_cond_3_6_1_reg ( .CLK(CLK), .D(_22683_), .Q(__maxi_read_fsm_cond_3_6_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38001_ ( .CLK(CLK), .D(_22682_), .Q(_wdata_851), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _wvalid_852_reg ( .CLK(CLK), .D(_22680_), .Q(_wvalid_852), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __maxi_read_fsm_cond_3_7_1_reg ( .CLK(CLK), .D(_22676_), .Q(__maxi_read_fsm_cond_3_7_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38004_ ( .CLK(CLK), .D(_22675_), .Q(_wdata_962), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _wvalid_963_reg ( .CLK(CLK), .D(_22673_), .Q(_wvalid_963), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __maxi_read_fsm_cond_3_8_1_reg ( .CLK(CLK), .D(_22669_), .Q(__maxi_read_fsm_cond_3_8_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38007_ ( .CLK(CLK), .D(_22668_), .Q(_wdata_973), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _wvalid_974_reg ( .CLK(CLK), .D(_22666_), .Q(_wvalid_974), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __maxi_read_fsm_cond_3_9_1_reg ( .CLK(CLK), .D(_22662_), .Q(__maxi_read_fsm_cond_3_9_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38010_ ( .CLK(CLK), .D(_22848_), .Q(control_conv2d_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38011_ ( .CLK(CLK), .D(_22846_), .Q(conv2d_8_act_base_offset_row), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38012_ ( .CLK(CLK), .D(_22845_), .Q(conv2d_8_act_base_offset_bat), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38013_ ( .CLK(CLK), .D(_22844_), .Q(conv2d_8_filter_base_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38014_ ( .CLK(CLK), .D(_22843_), .Q(conv2d_8_out_base_offset_val), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38015_ ( .CLK(CLK), .D(_22842_), .Q(conv2d_8_out_base_offset_col), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38016_ ( .CLK(CLK), .D(_22841_), .Q(conv2d_8_out_base_offset_row), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38017_ ( .CLK(CLK), .D(_22839_), .Q(conv2d_8_out_base_offset_bat), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38018_ ( .CLK(CLK), .D(_22838_), .Q(conv2d_8_out_base_offset_och), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) conv2d_8_dma_flag_0_reg ( .CLK(CLK), .D(_22837_), .Q(conv2d_8_dma_flag_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) conv2d_8_dma_flag_1_reg ( .CLK(CLK), .D(_22836_), .Q(conv2d_8_dma_flag_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) conv2d_8_dma_flag_2_reg ( .CLK(CLK), .D(_22835_), .Q(conv2d_8_dma_flag_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38022_ ( .CLK(CLK), .D(_22834_), .Q(conv2d_8_sync_out_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38023_ ( .CLK(CLK), .D(_22833_), .Q(conv2d_8_next_out_write_size), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38024_ ( .CLK(CLK), .D(_22832_), .Q(conv2d_8_row_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38025_ ( .CLK(CLK), .D(_22831_), .Q(conv2d_8_bat_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38026_ ( .CLK(CLK), .D(_22830_), .Q(conv2d_8_och_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _38027_ ( .CLK(CLK), .D(_22829_), .Q(conv2d_8_row_select), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38028_ ( .CLK(CLK), .D(_22827_), .Q(conv2d_8_out_row_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38029_ ( .CLK(CLK), .D(_22825_), .Q(conv2d_8_out_ram_select), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38030_ ( .CLK(CLK), .D(_22824_), .Q(conv2d_8_prev_row_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38031_ ( .CLK(CLK), .D(_22823_), .Q(conv2d_8_prev_bat_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38032_ ( .CLK(CLK), .D(_22822_), .Q(conv2d_8_prev_och_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _38033_ ( .CLK(CLK), .D(_22821_), .Q(conv2d_8_prev_row_select), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38034_ ( .CLK(CLK), .D(_22820_), .Q(conv2d_8_act_page_comp_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38035_ ( .CLK(CLK), .D(_22817_), .Q(conv2d_8_act_page_comp_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38036_ ( .CLK(CLK), .D(_22814_), .Q(conv2d_8_act_page_comp_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38037_ ( .CLK(CLK), .D(_22811_), .Q(conv2d_8_act_page_dma_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38038_ ( .CLK(CLK), .D(_22808_), .Q(conv2d_8_act_page_dma_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38039_ ( .CLK(CLK), .D(_22805_), .Q(conv2d_8_act_page_dma_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38040_ ( .CLK(CLK), .D(_22802_), .Q(conv2d_8_filter_page_comp_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38041_ ( .CLK(CLK), .D(_22800_), .Q(conv2d_8_filter_page_dma_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) conv2d_8_out_page_reg ( .CLK(CLK), .D(_22798_), .Q(conv2d_8_out_page), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38043_ ( .CLK(CLK), .D(_22797_), .Q(conv2d_8_out_page_comp_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38044_ ( .CLK(CLK), .D(_22796_), .Q(conv2d_8_out_page_dma_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38045_ ( .CLK(CLK), .D(_22795_), .Q(conv2d_8_out_laddr_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) conv2d_8_skip_read_filter_reg ( .CLK(CLK), .D(_22794_), .Q(conv2d_8_skip_read_filter), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) conv2d_8_skip_read_act_reg ( .CLK(CLK), .D(_22793_), .Q(conv2d_8_skip_read_act), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) conv2d_8_skip_comp_reg ( .CLK(CLK), .D(_22792_), .Q(conv2d_8_skip_comp), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) conv2d_8_skip_write_out_reg  ( .CLK(CLK), .D(_03072_), .Q(conv2d_8_skip_write_out) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_9_reg ( .CLK(CLK), .D(_22790_), .Q(axim_flag_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38051_ ( .CLK(CLK), .D(control_conv2d_8), .Q(_d1_control_conv2d_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_conv2d_8_cond_3_0_1_reg ( .CLK(CLK), .D(_22787_), .Q(_control_conv2d_8_cond_3_0_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_16_reg ( .CLK(CLK), .D(_22786_), .Q(axim_flag_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_conv2d_8_cond_8_1_1_reg ( .CLK(CLK), .D(_22783_), .Q(_control_conv2d_8_cond_8_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) set_req_28_reg ( .CLK(CLK), .D(_22782_), .Q(set_req_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_conv2d_8_cond_14_2_1_reg ( .CLK(CLK), .D(_22779_), .Q(_control_conv2d_8_cond_14_2_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_29_reg ( .CLK(CLK), .D(_22778_), .Q(axim_flag_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_conv2d_8_cond_15_3_1_reg ( .CLK(CLK), .D(_22775_), .Q(_control_conv2d_8_cond_15_3_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) set_req_157_reg ( .CLK(CLK), .D(_22774_), .Q(set_req_157), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_conv2d_8_cond_23_4_1_reg ( .CLK(CLK), .D(_22771_), .Q(_control_conv2d_8_cond_23_4_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_158_reg ( .CLK(CLK), .D(_22770_), .Q(axim_flag_158), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_conv2d_8_cond_24_5_1_reg ( .CLK(CLK), .D(_22767_), .Q(_control_conv2d_8_cond_24_5_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) set_req_214_reg ( .CLK(CLK), .D(_22766_), .Q(set_req_214), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_conv2d_8_cond_30_6_1_reg ( .CLK(CLK), .D(_22763_), .Q(_control_conv2d_8_cond_30_6_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_215_reg ( .CLK(CLK), .D(_22762_), .Q(axim_flag_215), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_conv2d_8_cond_31_7_1_reg ( .CLK(CLK), .D(_22759_), .Q(_control_conv2d_8_cond_31_7_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) set_req_271_reg ( .CLK(CLK), .D(_22758_), .Q(set_req_271), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_conv2d_8_cond_37_8_1_reg ( .CLK(CLK), .D(_22755_), .Q(_control_conv2d_8_cond_37_8_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_272_reg ( .CLK(CLK), .D(_22754_), .Q(axim_flag_272), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_conv2d_8_cond_38_9_1_reg ( .CLK(CLK), .D(_22751_), .Q(_control_conv2d_8_cond_38_9_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) axim_flag_798_reg ( .CLK(CLK), .D(_22750_), .Q(axim_flag_798), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _control_conv2d_8_cond_48_10_1_reg ( .CLK(CLK), .D(_22747_), .Q(_control_conv2d_8_cond_48_10_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) conv2d_8_control_param_index_reg ( .CLK(CLK), .D(_22868_), .Q(conv2d_8_control_param_index), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) max_pool_serial_9_control_param_index_reg ( .CLK(CLK), .D(_22867_), .Q(max_pool_serial_9_control_param_index), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38075_ ( .CLK(CLK), .D(_22866_), .Q(main_fsm), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38076_ ( .CLK(CLK), .D(_22865_), .Q(conv2d_8_objaddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38077_ ( .CLK(CLK), .D(_22864_), .Q(conv2d_8_arg_objaddr_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38078_ ( .CLK(CLK), .D(_22863_), .Q(conv2d_8_arg_objaddr_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38079_ ( .CLK(CLK), .D(_22862_), .Q(conv2d_8_arg_objaddr_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38080_ ( .CLK(CLK), .D(_22861_), .Q(conv2d_8_arg_objaddr_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38081_ ( .CLK(CLK), .D(_22860_), .Q(max_pool_serial_9_objaddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38082_ ( .CLK(CLK), .D(_22859_), .Q(max_pool_serial_9_arg_objaddr_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38083_ ( .CLK(CLK), .D(_22858_), .Q(matmul_15_objaddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38084_ ( .CLK(CLK), .D(_22857_), .Q(matmul_15_arg_objaddr_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38085_ ( .CLK(CLK), .D(_22856_), .Q(matmul_15_arg_objaddr_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38086_ ( .CLK(CLK), .D(_22855_), .Q(matmul_15_arg_objaddr_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38087_ ( .CLK(CLK), .D(_22854_), .Q(matmul_15_arg_objaddr_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38088_ ( .CLK(CLK), .D(_22874_), .Q(_stream_matmul_15_fsm), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_start_reg ( .CLK(CLK), .D(_22873_), .Q(_stream_matmul_15_start), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_end_flag_reg ( .CLK(CLK), .D(_22871_), .Q(_stream_matmul_15_end_flag), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_term_sink_reg ( .CLK(CLK), .D(_22870_), .Q(_stream_matmul_15_term_sink), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_source_busy_reg ( .CLK(CLK), .D(_22869_), .Q(_stream_matmul_15_source_busy), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38093_ ( .CLK(CLK), .D(_23114_), .Q(_stream_matmul_15_constant_0_next_constant_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_constant_1_next_constant_data_reg ( .CLK(CLK), .D(_23113_), .Q(_stream_matmul_15_constant_1_next_constant_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_constant_2_next_constant_data_reg ( .CLK(CLK), .D(_23112_), .Q(_stream_matmul_15_constant_2_next_constant_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_constant_3_next_constant_data_reg ( .CLK(CLK), .D(_23111_), .Q(_stream_matmul_15_constant_3_next_constant_data), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_15_source_6_idle_reg  ( .CLK(CLK), .D(_02622_), .Q(_stream_matmul_15_source_6_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38098_ ( .CLK(CLK), .D(_23108_), .Q(_stream_matmul_15_source_6_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38099_ ( .CLK(CLK), .D(_23107_), .Q(_stream_matmul_15_source_6_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38100_ ( .CLK(CLK), .D(_23106_), .Q(_stream_matmul_15_source_6_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38101_ ( .CLK(CLK), .D(_23105_), .Q(_stream_matmul_15_source_6_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38102_ ( .CLK(CLK), .D(_23104_), .Q(_stream_matmul_15_source_6_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_source_6_source_ram_renable_reg ( .CLK(CLK), .D(_23103_), .Q(_stream_matmul_15_source_6_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_source_6_source_ram_rvalid_reg ( .CLK(CLK), .D(_23101_), .Q(_stream_matmul_15_source_6_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_15_source_8_idle_reg  ( .CLK(CLK), .D(_02631_), .Q(_stream_matmul_15_source_8_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38106_ ( .CLK(CLK), .D(_23098_), .Q(_stream_matmul_15_source_8_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38107_ ( .CLK(CLK), .D(_23097_), .Q(_stream_matmul_15_source_8_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38108_ ( .CLK(CLK), .D(_23096_), .Q(_stream_matmul_15_source_8_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38109_ ( .CLK(CLK), .D(_23095_), .Q(_stream_matmul_15_source_8_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38110_ ( .CLK(CLK), .D(_23094_), .Q(_stream_matmul_15_source_8_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_source_8_source_ram_renable_reg ( .CLK(CLK), .D(_23093_), .Q(_stream_matmul_15_source_8_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_source_8_source_ram_rvalid_reg ( .CLK(CLK), .D(_23091_), .Q(_stream_matmul_15_source_8_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_15_source_10_idle_reg  ( .CLK(CLK), .D(_02598_), .Q(_stream_matmul_15_source_10_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38114_ ( .CLK(CLK), .D(_23089_), .Q(_stream_matmul_15_source_10_source_empty_data), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_15_source_12_idle_reg  ( .CLK(CLK), .D(_02600_), .Q(_stream_matmul_15_source_12_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38116_ ( .CLK(CLK), .D(_23087_), .Q(_stream_matmul_15_source_12_source_empty_data), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_15_source_14_idle_reg  ( .CLK(CLK), .D(_02602_), .Q(_stream_matmul_15_source_14_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38118_ ( .CLK(CLK), .D(_23085_), .Q(_stream_matmul_15_source_14_source_empty_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_constant_15_next_constant_data_reg ( .CLK(CLK), .D(_23084_), .Q(_stream_matmul_15_constant_15_next_constant_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_constant_16_next_constant_data_reg ( .CLK(CLK), .D(_23083_), .Q(_stream_matmul_15_constant_16_next_constant_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _38121_ ( .CLK(CLK), .D(_23082_), .Q(_stream_matmul_15_constant_17_next_constant_data), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_15_source_19_idle_reg  ( .CLK(CLK), .D(_02604_), .Q(_stream_matmul_15_source_19_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38123_ ( .CLK(CLK), .D(_23079_), .Q(_stream_matmul_15_source_19_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38124_ ( .CLK(CLK), .D(_23078_), .Q(_stream_matmul_15_source_19_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38125_ ( .CLK(CLK), .D(_23077_), .Q(_stream_matmul_15_source_19_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38126_ ( .CLK(CLK), .D(_23076_), .Q(_stream_matmul_15_source_19_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38127_ ( .CLK(CLK), .D(_23075_), .Q(_stream_matmul_15_source_19_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_source_19_source_ram_renable_reg ( .CLK(CLK), .D(_23074_), .Q(_stream_matmul_15_source_19_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_source_19_source_ram_rvalid_reg ( .CLK(CLK), .D(_23072_), .Q(_stream_matmul_15_source_19_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_15_source_20_idle_reg  ( .CLK(CLK), .D(_02613_), .Q(_stream_matmul_15_source_20_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38131_ ( .CLK(CLK), .D(_23069_), .Q(_stream_matmul_15_source_20_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38132_ ( .CLK(CLK), .D(_23068_), .Q(_stream_matmul_15_source_20_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38133_ ( .CLK(CLK), .D(_23067_), .Q(_stream_matmul_15_source_20_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38134_ ( .CLK(CLK), .D(_23066_), .Q(_stream_matmul_15_source_20_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38135_ ( .CLK(CLK), .D(_23065_), .Q(_stream_matmul_15_source_20_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_source_20_source_ram_renable_reg ( .CLK(CLK), .D(_23064_), .Q(_stream_matmul_15_source_20_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_source_20_source_ram_rvalid_reg ( .CLK(CLK), .D(_23062_), .Q(_stream_matmul_15_source_20_source_ram_rvalid), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38138_ ( .CLK(CLK), .D(_23061_), .Q(_stream_matmul_15_sink_21_sink_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38139_ ( .CLK(CLK), .D(_23060_), .Q(_stream_matmul_15_sink_21_sink_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38140_ ( .CLK(CLK), .D(_23059_), .Q(_stream_matmul_15_sink_21_sink_size), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38141_ ( .CLK(CLK), .D(_23058_), .Q(_stream_matmul_15_sink_21_sink_stride), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38142_ ( .CLK(CLK), .D(_23057_), .Q(_stream_matmul_15_sink_21_sink_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38143_ ( .CLK(CLK), .D(_23055_), .Q(_stream_matmul_15_sink_21_sink_stride_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38144_ ( .CLK(CLK), .D(_23054_), .Q(_stream_matmul_15_sink_21_sink_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38145_ ( .CLK(CLK), .D(_23053_), .Q(_stream_matmul_15_sink_21_sink_waddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_matmul_15_sink_21_sink_wenable_reg ( .CLK(CLK), .D(_23051_), .Q(_stream_matmul_15_sink_21_sink_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38147_ ( .CLK(CLK), .D(_23050_), .Q(_stream_matmul_15_sink_21_sink_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38148_ ( .CLK(CLK), .D(__variable_wdata_792), .Q(_cond_data_797), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38149_ ( .CLK(CLK), .D(__variable_wdata_799), .Q(_cond_data_804), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38150_ ( .CLK(CLK), .D(__variable_wdata_806), .Q(_cond_data_811), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38151_ ( .CLK(CLK), .D(__variable_wdata_813), .Q(_cond_data_818), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38152_ ( .CLK(CLK), .D(__variable_wdata_820), .Q(_cond_data_825), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _eq_data_831_reg ( .CLK(CLK), .D(_05230_), .Q(_eq_data_831), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _eq_data_835_reg ( .CLK(CLK), .D(_05231_), .Q(_eq_data_835), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pointer_data_850_reg ( .CLK(CLK), .D(__variable_wdata_779), .Q(_pointer_data_850), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38156_ ( .CLK(CLK), .D(__variable_wdata_830), .Q(__delay_data_1378), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1382_reg ( .CLK(CLK), .D(__variable_wdata_826), .Q(__delay_data_1382), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38158_ ( .CLK(CLK), .D(__variable_wdata_844), .Q(__delay_data_1383), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1389_reg ( .CLK(CLK), .D(__variable_wdata_827), .Q(__delay_data_1389), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38160_ ( .CLK(CLK), .D(__variable_wdata_776), .Q(__delay_data_1404), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _38161_ ( .CLK(CLK), .D(__variable_wdata_828), .Q(__delay_data_1442), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38162_ ( .CLK(CLK), .D(_26632_), .Q(_cond_data_833), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38163_ ( .CLK(CLK), .D(_22240_), .Q(_plus_data_855), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38164_ ( .CLK(CLK), .D(_22241_), .Q(_plus_data_860), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38165_ ( .CLK(CLK), .D(_22242_), .Q(_plus_data_865), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1379_reg ( .CLK(CLK), .D(_eq_data_835), .Q(__delay_data_1379), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1380_reg ( .CLK(CLK), .D(_pointer_data_850), .Q(__delay_data_1380), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38168_ ( .CLK(CLK), .D(__delay_data_1383), .Q(__delay_data_1384), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38169_ ( .CLK(CLK), .D(__delay_data_1404), .Q(__delay_data_1405), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38170_ ( .CLK(CLK), .D(_cond_data_797), .Q(__delay_data_1420), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38171_ ( .CLK(CLK), .D(_cond_data_804), .Q(__delay_data_1443), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38172_ ( .CLK(CLK), .D(_26633_), .Q(_cond_data_837), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1381_reg ( .CLK(CLK), .D(__delay_data_1380), .Q(__delay_data_1381), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38174_ ( .CLK(CLK), .D(__delay_data_1384), .Q(__delay_data_1385), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38175_ ( .CLK(CLK), .D(_plus_data_855), .Q(__delay_data_1387), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38176_ ( .CLK(CLK), .D(_plus_data_860), .Q(__delay_data_1390), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38177_ ( .CLK(CLK), .D(__delay_data_1405), .Q(__delay_data_1406), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38178_ ( .CLK(CLK), .D(__delay_data_1420), .Q(__delay_data_1421), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38179_ ( .CLK(CLK), .D(__delay_data_1443), .Q(__delay_data_1444), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38180_ ( .CLK(CLK), .D(_plus_data_865), .Q(__delay_data_1466), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38181_ ( .CLK(CLK), .D(_26634_), .Q(_cond_data_853), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38182_ ( .CLK(CLK), .D(__delay_data_1385), .Q(__delay_data_1386), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38183_ ( .CLK(CLK), .D(__delay_data_1387), .Q(__delay_data_1388), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38184_ ( .CLK(CLK), .D(__delay_data_1390), .Q(__delay_data_1391), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38185_ ( .CLK(CLK), .D(__delay_data_1406), .Q(__delay_data_1407), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38186_ ( .CLK(CLK), .D(__delay_data_1421), .Q(__delay_data_1422), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38187_ ( .CLK(CLK), .D(__delay_data_1444), .Q(__delay_data_1445), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38188_ ( .CLK(CLK), .D(__delay_data_1466), .Q(__delay_data_1467), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38189_ ( .CLK(CLK), .D(__delay_data_1391), .Q(__delay_data_1392), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38190_ ( .CLK(CLK), .D(__delay_data_1407), .Q(__delay_data_1408), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38191_ ( .CLK(CLK), .D(__delay_data_1422), .Q(__delay_data_1423), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38192_ ( .CLK(CLK), .D(__delay_data_1445), .Q(__delay_data_1446), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38193_ ( .CLK(CLK), .D(__delay_data_1467), .Q(__delay_data_1468), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38194_ ( .CLK(CLK), .D(__delay_data_1392), .Q(__delay_data_1393), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38195_ ( .CLK(CLK), .D(__delay_data_1408), .Q(__delay_data_1409), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38196_ ( .CLK(CLK), .D(__delay_data_1423), .Q(__delay_data_1424), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38197_ ( .CLK(CLK), .D(__delay_data_1446), .Q(__delay_data_1447), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38198_ ( .CLK(CLK), .D(__delay_data_1468), .Q(__delay_data_1469), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38199_ ( .CLK(CLK), .D(__delay_data_1393), .Q(__delay_data_1394), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38200_ ( .CLK(CLK), .D(__delay_data_1409), .Q(__delay_data_1410), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38201_ ( .CLK(CLK), .D(__delay_data_1424), .Q(__delay_data_1425), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38202_ ( .CLK(CLK), .D(__delay_data_1447), .Q(__delay_data_1448), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38203_ ( .CLK(CLK), .D(__delay_data_1469), .Q(__delay_data_1470), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38204_ ( .CLK(CLK), .D(__delay_data_1394), .Q(__delay_data_1395), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38205_ ( .CLK(CLK), .D(__delay_data_1410), .Q(__delay_data_1411), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38206_ ( .CLK(CLK), .D(__delay_data_1425), .Q(__delay_data_1426), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38207_ ( .CLK(CLK), .D(__delay_data_1448), .Q(__delay_data_1449), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38208_ ( .CLK(CLK), .D(__delay_data_1470), .Q(__delay_data_1471), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38209_ ( .CLK(CLK), .D(__delay_data_1395), .Q(__delay_data_1396), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38210_ ( .CLK(CLK), .D(__delay_data_1411), .Q(__delay_data_1412), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38211_ ( .CLK(CLK), .D(__delay_data_1426), .Q(__delay_data_1427), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38212_ ( .CLK(CLK), .D(__delay_data_1449), .Q(__delay_data_1450), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38213_ ( .CLK(CLK), .D(__delay_data_1471), .Q(__delay_data_1472), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38214_ ( .CLK(CLK), .D(__delay_data_1396), .Q(__delay_data_1397), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38215_ ( .CLK(CLK), .D(__delay_data_1412), .Q(__delay_data_1413), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38216_ ( .CLK(CLK), .D(__delay_data_1427), .Q(__delay_data_1428), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38217_ ( .CLK(CLK), .D(__delay_data_1450), .Q(__delay_data_1451), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38218_ ( .CLK(CLK), .D(__delay_data_1472), .Q(__delay_data_1473), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38219_ ( .CLK(CLK), .D(__delay_data_1397), .Q(__delay_data_1398), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38220_ ( .CLK(CLK), .D(__delay_data_1413), .Q(__delay_data_1414), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38221_ ( .CLK(CLK), .D(__delay_data_1428), .Q(__delay_data_1429), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38222_ ( .CLK(CLK), .D(__delay_data_1451), .Q(__delay_data_1452), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38223_ ( .CLK(CLK), .D(__delay_data_1473), .Q(__delay_data_1474), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38224_ ( .CLK(CLK), .D(__delay_data_1398), .Q(__delay_data_1399), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38225_ ( .CLK(CLK), .D(__delay_data_1414), .Q(__delay_data_1415), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38226_ ( .CLK(CLK), .D(__delay_data_1429), .Q(__delay_data_1430), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38227_ ( .CLK(CLK), .D(__delay_data_1452), .Q(__delay_data_1453), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38228_ ( .CLK(CLK), .D(__delay_data_1474), .Q(__delay_data_1475), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38229_ ( .CLK(CLK), .D(__delay_data_1399), .Q(__delay_data_1400), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38230_ ( .CLK(CLK), .D(__delay_data_1415), .Q(__delay_data_1416), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38231_ ( .CLK(CLK), .D(__delay_data_1430), .Q(__delay_data_1431), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38232_ ( .CLK(CLK), .D(__delay_data_1453), .Q(__delay_data_1454), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38233_ ( .CLK(CLK), .D(__delay_data_1475), .Q(__delay_data_1476), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _38234_ ( .CLK(CLK), .D(_sra_data_66), .Q(__substreamoutput_data_856), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38235_ ( .CLK(CLK), .D(__delay_data_1400), .Q(__delay_data_1401), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38236_ ( .CLK(CLK), .D(__delay_data_1416), .Q(__delay_data_1417), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38237_ ( .CLK(CLK), .D(__delay_data_1431), .Q(__delay_data_1432), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38238_ ( .CLK(CLK), .D(__delay_data_1454), .Q(__delay_data_1455), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38239_ ( .CLK(CLK), .D(__delay_data_1476), .Q(__delay_data_1477), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38240_ ( .CLK(CLK), .D(__delay_data_1401), .Q(__delay_data_1402), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38241_ ( .CLK(CLK), .D(__delay_data_1417), .Q(__delay_data_1418), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38242_ ( .CLK(CLK), .D(__delay_data_1432), .Q(__delay_data_1433), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38243_ ( .CLK(CLK), .D(__delay_data_1455), .Q(__delay_data_1456), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38244_ ( .CLK(CLK), .D(__delay_data_1477), .Q(__delay_data_1478), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38245_ ( .CLK(CLK), .D(__variable_wdata_20), .Q(__substreamoutput_data_858), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38246_ ( .CLK(CLK), .D(__delay_data_1402), .Q(__delay_data_1403), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38247_ ( .CLK(CLK), .D(__delay_data_1418), .Q(__delay_data_1419), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38248_ ( .CLK(CLK), .D(__delay_data_1433), .Q(__delay_data_1434), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38249_ ( .CLK(CLK), .D(__delay_data_1456), .Q(__delay_data_1457), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38250_ ( .CLK(CLK), .D(__delay_data_1478), .Q(__delay_data_1479), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38251_ ( .CLK(CLK), .D(__delay_data_1434), .Q(__delay_data_1435), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38252_ ( .CLK(CLK), .D(__delay_data_1457), .Q(__delay_data_1458), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38253_ ( .CLK(CLK), .D(__delay_data_1479), .Q(__delay_data_1480), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38254_ ( .CLK(CLK), .D(__delay_data_1435), .Q(__delay_data_1436), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38255_ ( .CLK(CLK), .D(__delay_data_1458), .Q(__delay_data_1459), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38256_ ( .CLK(CLK), .D(__delay_data_1480), .Q(__delay_data_1481), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38257_ ( .CLK(CLK), .D(__delay_data_1436), .Q(__delay_data_1437), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38258_ ( .CLK(CLK), .D(__delay_data_1459), .Q(__delay_data_1460), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38259_ ( .CLK(CLK), .D(__delay_data_1481), .Q(__delay_data_1482), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38260_ ( .CLK(CLK), .D(__delay_data_1437), .Q(__delay_data_1438), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38261_ ( .CLK(CLK), .D(__delay_data_1460), .Q(__delay_data_1461), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38262_ ( .CLK(CLK), .D(__delay_data_1482), .Q(__delay_data_1483), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38263_ ( .CLK(CLK), .D(__delay_data_1438), .Q(__delay_data_1439), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38264_ ( .CLK(CLK), .D(__delay_data_1461), .Q(__delay_data_1462), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38265_ ( .CLK(CLK), .D(__delay_data_1483), .Q(__delay_data_1484), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38266_ ( .CLK(CLK), .D(__delay_data_1439), .Q(__delay_data_1440), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38267_ ( .CLK(CLK), .D(__delay_data_1462), .Q(__delay_data_1463), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38268_ ( .CLK(CLK), .D(__delay_data_1484), .Q(__delay_data_1485), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38269_ ( .CLK(CLK), .D(_sra_data_19), .Q(__substreamoutput_data_861), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __substreamoutput_data_862_reg ( .CLK(CLK), .D(__delay_data_738), .Q(__substreamoutput_data_862), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38271_ ( .CLK(CLK), .D(__delay_data_1440), .Q(__delay_data_1441), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38272_ ( .CLK(CLK), .D(__delay_data_1463), .Q(__delay_data_1464), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38273_ ( .CLK(CLK), .D(__delay_data_1485), .Q(__delay_data_1486), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38274_ ( .CLK(CLK), .D(_22243_), .Q(_plus_data_863), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38275_ ( .CLK(CLK), .D(__delay_data_1464), .Q(__delay_data_1465), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38276_ ( .CLK(CLK), .D(__delay_data_1486), .Q(__delay_data_1487), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1488_reg ( .CLK(CLK), .D(__substreamoutput_data_862), .Q(__delay_data_1488), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1489_reg ( .CLK(CLK), .D(__delay_data_1488), .Q(__delay_data_1489), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1490_reg ( .CLK(CLK), .D(__delay_data_1489), .Q(__delay_data_1490), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1491_reg ( .CLK(CLK), .D(__delay_data_1490), .Q(__delay_data_1491), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1492_reg ( .CLK(CLK), .D(__delay_data_1491), .Q(__delay_data_1492), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1493_reg ( .CLK(CLK), .D(__delay_data_1492), .Q(__delay_data_1493), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1494_reg ( .CLK(CLK), .D(__delay_data_1493), .Q(__delay_data_1494), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1495_reg ( .CLK(CLK), .D(__delay_data_1494), .Q(__delay_data_1495), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1496_reg ( .CLK(CLK), .D(__delay_data_1495), .Q(__delay_data_1496), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1497_reg ( .CLK(CLK), .D(__delay_data_1496), .Q(__delay_data_1497), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38287_ ( .CLK(CLK), .D(_cond_data_51), .Q(__substreamoutput_data_866), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1498_reg ( .CLK(CLK), .D(__delay_data_1497), .Q(__delay_data_1498), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38289_ ( .CLK(CLK), .D(_23049_), .Q(__variable_wdata_776), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __variable_wdata_777_reg ( .CLK(CLK), .D(_23048_), .Q(__variable_wdata_777), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __variable_wdata_778_reg ( .CLK(CLK), .D(_23047_), .Q(__variable_wdata_778), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __variable_wdata_779_reg ( .CLK(CLK), .D(_23046_), .Q(__variable_wdata_779), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38293_ ( .CLK(CLK), .D(_23045_), .Q(_source_stream_matmul_15_source_6_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38294_ ( .CLK(CLK), .D(_23042_), .Q(_source_stream_matmul_15_source_6_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38295_ ( .CLK(CLK), .D(_23039_), .Q(_source_stream_matmul_15_source_6_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38296_ ( .CLK(CLK), .D(_23036_), .Q(_source_stream_matmul_15_source_6_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38297_ ( .CLK(CLK), .D(_23033_), .Q(_source_stream_matmul_15_source_6_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38298_ ( .CLK(CLK), .D(_23032_), .Q(_source_stream_matmul_15_source_6_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38299_ ( .CLK(CLK), .D(_23031_), .Q(_source_stream_matmul_15_source_6_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38300_ ( .CLK(CLK), .D(_23030_), .Q(_source_stream_matmul_15_source_6_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38301_ ( .CLK(CLK), .D(_23029_), .Q(_source_stream_matmul_15_source_6_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38302_ ( .CLK(CLK), .D(_23028_), .Q(_source_stream_matmul_15_source_6_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38303_ ( .CLK(CLK), .D(_23027_), .Q(_source_stream_matmul_15_source_6_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38304_ ( .CLK(CLK), .D(_23026_), .Q(_source_stream_matmul_15_source_6_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38305_ ( .CLK(CLK), .D(_23025_), .Q(_source_stream_matmul_15_source_6_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38306_ ( .CLK(CLK), .D(_23022_), .Q(_source_stream_matmul_15_source_6_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38307_ ( .CLK(CLK), .D(_23019_), .Q(_source_stream_matmul_15_source_6_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38308_ ( .CLK(CLK), .D(_23016_), .Q(_source_stream_matmul_15_source_6_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38309_ ( .CLK(CLK), .D(_23013_), .Q(_source_stream_matmul_15_source_6_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38310_ ( .CLK(CLK), .D(_23012_), .Q(_source_stream_matmul_15_source_6_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38311_ ( .CLK(CLK), .D(_23011_), .Q(_source_stream_matmul_15_source_6_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38312_ ( .CLK(CLK), .D(_23010_), .Q(_source_stream_matmul_15_source_6_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38313_ ( .CLK(CLK), .D(_23009_), .Q(_source_stream_matmul_15_source_6_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38314_ ( .CLK(CLK), .D(_23008_), .Q(_source_stream_matmul_15_source_6_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38315_ ( .CLK(CLK), .D(_23007_), .Q(_source_stream_matmul_15_source_6_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38316_ ( .CLK(CLK), .D(_23006_), .Q(_source_stream_matmul_15_source_6_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38317_ ( .CLK(CLK), .D(_23005_), .Q(__variable_wdata_792), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38318_ ( .CLK(CLK), .D(_23004_), .Q(_source_stream_matmul_15_source_8_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38319_ ( .CLK(CLK), .D(_23001_), .Q(_source_stream_matmul_15_source_8_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38320_ ( .CLK(CLK), .D(_22998_), .Q(_source_stream_matmul_15_source_8_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38321_ ( .CLK(CLK), .D(_22995_), .Q(_source_stream_matmul_15_source_8_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38322_ ( .CLK(CLK), .D(_22992_), .Q(_source_stream_matmul_15_source_8_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38323_ ( .CLK(CLK), .D(_22991_), .Q(_source_stream_matmul_15_source_8_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38324_ ( .CLK(CLK), .D(_22990_), .Q(_source_stream_matmul_15_source_8_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38325_ ( .CLK(CLK), .D(_22989_), .Q(_source_stream_matmul_15_source_8_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38326_ ( .CLK(CLK), .D(_22988_), .Q(_source_stream_matmul_15_source_8_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38327_ ( .CLK(CLK), .D(_22987_), .Q(_source_stream_matmul_15_source_8_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38328_ ( .CLK(CLK), .D(_22986_), .Q(_source_stream_matmul_15_source_8_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38329_ ( .CLK(CLK), .D(_22985_), .Q(_source_stream_matmul_15_source_8_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38330_ ( .CLK(CLK), .D(_22984_), .Q(_source_stream_matmul_15_source_8_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38331_ ( .CLK(CLK), .D(_22981_), .Q(_source_stream_matmul_15_source_8_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38332_ ( .CLK(CLK), .D(_22978_), .Q(_source_stream_matmul_15_source_8_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38333_ ( .CLK(CLK), .D(_22975_), .Q(_source_stream_matmul_15_source_8_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38334_ ( .CLK(CLK), .D(_22972_), .Q(_source_stream_matmul_15_source_8_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38335_ ( .CLK(CLK), .D(_22971_), .Q(_source_stream_matmul_15_source_8_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38336_ ( .CLK(CLK), .D(_22970_), .Q(_source_stream_matmul_15_source_8_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38337_ ( .CLK(CLK), .D(_22969_), .Q(_source_stream_matmul_15_source_8_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38338_ ( .CLK(CLK), .D(_22968_), .Q(_source_stream_matmul_15_source_8_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38339_ ( .CLK(CLK), .D(_22967_), .Q(_source_stream_matmul_15_source_8_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38340_ ( .CLK(CLK), .D(_22966_), .Q(_source_stream_matmul_15_source_8_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38341_ ( .CLK(CLK), .D(_22965_), .Q(_source_stream_matmul_15_source_8_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38342_ ( .CLK(CLK), .D(_22964_), .Q(__variable_wdata_799), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38343_ ( .CLK(CLK), .D(_22963_), .Q(__variable_wdata_806), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38344_ ( .CLK(CLK), .D(_22962_), .Q(__variable_wdata_813), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38345_ ( .CLK(CLK), .D(_22961_), .Q(__variable_wdata_820), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __variable_wdata_826_reg ( .CLK(CLK), .D(_22960_), .Q(__variable_wdata_826), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __variable_wdata_827_reg ( .CLK(CLK), .D(_22959_), .Q(__variable_wdata_827), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _38348_ ( .CLK(CLK), .D(_22958_), .Q(__variable_wdata_828), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38349_ ( .CLK(CLK), .D(_22957_), .Q(_source_stream_matmul_15_source_19_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38350_ ( .CLK(CLK), .D(_22954_), .Q(_source_stream_matmul_15_source_19_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38351_ ( .CLK(CLK), .D(_22951_), .Q(_source_stream_matmul_15_source_19_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38352_ ( .CLK(CLK), .D(_22948_), .Q(_source_stream_matmul_15_source_19_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38353_ ( .CLK(CLK), .D(_22945_), .Q(_source_stream_matmul_15_source_19_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38354_ ( .CLK(CLK), .D(_22944_), .Q(_source_stream_matmul_15_source_19_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38355_ ( .CLK(CLK), .D(_22943_), .Q(_source_stream_matmul_15_source_19_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38356_ ( .CLK(CLK), .D(_22942_), .Q(_source_stream_matmul_15_source_19_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38357_ ( .CLK(CLK), .D(_22941_), .Q(_source_stream_matmul_15_source_19_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38358_ ( .CLK(CLK), .D(_22940_), .Q(_source_stream_matmul_15_source_19_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38359_ ( .CLK(CLK), .D(_22939_), .Q(_source_stream_matmul_15_source_19_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38360_ ( .CLK(CLK), .D(_22938_), .Q(_source_stream_matmul_15_source_19_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38361_ ( .CLK(CLK), .D(_22937_), .Q(_source_stream_matmul_15_source_19_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38362_ ( .CLK(CLK), .D(_22934_), .Q(_source_stream_matmul_15_source_19_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38363_ ( .CLK(CLK), .D(_22931_), .Q(_source_stream_matmul_15_source_19_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38364_ ( .CLK(CLK), .D(_22928_), .Q(_source_stream_matmul_15_source_19_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38365_ ( .CLK(CLK), .D(_22925_), .Q(_source_stream_matmul_15_source_19_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38366_ ( .CLK(CLK), .D(_22924_), .Q(_source_stream_matmul_15_source_19_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38367_ ( .CLK(CLK), .D(_22923_), .Q(_source_stream_matmul_15_source_19_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38368_ ( .CLK(CLK), .D(_22922_), .Q(_source_stream_matmul_15_source_19_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38369_ ( .CLK(CLK), .D(_22921_), .Q(_source_stream_matmul_15_source_19_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38370_ ( .CLK(CLK), .D(_22920_), .Q(_source_stream_matmul_15_source_19_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38371_ ( .CLK(CLK), .D(_22919_), .Q(_source_stream_matmul_15_source_19_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38372_ ( .CLK(CLK), .D(_22918_), .Q(_source_stream_matmul_15_source_19_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38373_ ( .CLK(CLK), .D(_22917_), .Q(__variable_wdata_830), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38374_ ( .CLK(CLK), .D(_22916_), .Q(_source_stream_matmul_15_source_20_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38375_ ( .CLK(CLK), .D(_22913_), .Q(_source_stream_matmul_15_source_20_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38376_ ( .CLK(CLK), .D(_22910_), .Q(_source_stream_matmul_15_source_20_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38377_ ( .CLK(CLK), .D(_22907_), .Q(_source_stream_matmul_15_source_20_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38378_ ( .CLK(CLK), .D(_22904_), .Q(_source_stream_matmul_15_source_20_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38379_ ( .CLK(CLK), .D(_22903_), .Q(_source_stream_matmul_15_source_20_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38380_ ( .CLK(CLK), .D(_22902_), .Q(_source_stream_matmul_15_source_20_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38381_ ( .CLK(CLK), .D(_22901_), .Q(_source_stream_matmul_15_source_20_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38382_ ( .CLK(CLK), .D(_22900_), .Q(_source_stream_matmul_15_source_20_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38383_ ( .CLK(CLK), .D(_22899_), .Q(_source_stream_matmul_15_source_20_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38384_ ( .CLK(CLK), .D(_22898_), .Q(_source_stream_matmul_15_source_20_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38385_ ( .CLK(CLK), .D(_22897_), .Q(_source_stream_matmul_15_source_20_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38386_ ( .CLK(CLK), .D(_22896_), .Q(_source_stream_matmul_15_source_20_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38387_ ( .CLK(CLK), .D(_22893_), .Q(_source_stream_matmul_15_source_20_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38388_ ( .CLK(CLK), .D(_22890_), .Q(_source_stream_matmul_15_source_20_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38389_ ( .CLK(CLK), .D(_22887_), .Q(_source_stream_matmul_15_source_20_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38390_ ( .CLK(CLK), .D(_22884_), .Q(_source_stream_matmul_15_source_20_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38391_ ( .CLK(CLK), .D(_22883_), .Q(_source_stream_matmul_15_source_20_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38392_ ( .CLK(CLK), .D(_22882_), .Q(_source_stream_matmul_15_source_20_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38393_ ( .CLK(CLK), .D(_22881_), .Q(_source_stream_matmul_15_source_20_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38394_ ( .CLK(CLK), .D(_22880_), .Q(_source_stream_matmul_15_source_20_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38395_ ( .CLK(CLK), .D(_22879_), .Q(_source_stream_matmul_15_source_20_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38396_ ( .CLK(CLK), .D(_22878_), .Q(_source_stream_matmul_15_source_20_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38397_ ( .CLK(CLK), .D(_22877_), .Q(_source_stream_matmul_15_source_20_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38398_ ( .CLK(CLK), .D(_22876_), .Q(__variable_wdata_844), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _set_flag_1034_reg ( .CLK(CLK), .D(_22875_), .Q(_set_flag_1034), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38400_ ( .CLK(CLK), .D(_22261_), .Q(__stream_matmul_15_sink_21_sink_offset_0_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38401_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_1), .Q(__stream_matmul_15_sink_21_sink_offset_0_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38402_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_2), .Q(__stream_matmul_15_sink_21_sink_offset_0_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38403_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_3), .Q(__stream_matmul_15_sink_21_sink_offset_0_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38404_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_4), .Q(__stream_matmul_15_sink_21_sink_offset_0_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38405_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_5), .Q(__stream_matmul_15_sink_21_sink_offset_0_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38406_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_6), .Q(__stream_matmul_15_sink_21_sink_offset_0_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38407_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_7), .Q(__stream_matmul_15_sink_21_sink_offset_0_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38408_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_8), .Q(__stream_matmul_15_sink_21_sink_offset_0_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38409_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_9), .Q(__stream_matmul_15_sink_21_sink_offset_0_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38410_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_10), .Q(__stream_matmul_15_sink_21_sink_offset_0_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38411_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_11), .Q(__stream_matmul_15_sink_21_sink_offset_0_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38412_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_12), .Q(__stream_matmul_15_sink_21_sink_offset_0_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38413_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_13), .Q(__stream_matmul_15_sink_21_sink_offset_0_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38414_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_14), .Q(__stream_matmul_15_sink_21_sink_offset_0_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38415_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_15), .Q(__stream_matmul_15_sink_21_sink_offset_0_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38416_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_16), .Q(__stream_matmul_15_sink_21_sink_offset_0_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38417_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_17), .Q(__stream_matmul_15_sink_21_sink_offset_0_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38418_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_18), .Q(__stream_matmul_15_sink_21_sink_offset_0_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38419_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_19), .Q(__stream_matmul_15_sink_21_sink_offset_0_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38420_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_20), .Q(__stream_matmul_15_sink_21_sink_offset_0_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38421_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_21), .Q(__stream_matmul_15_sink_21_sink_offset_0_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38422_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_22), .Q(__stream_matmul_15_sink_21_sink_offset_0_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38423_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_23), .Q(__stream_matmul_15_sink_21_sink_offset_0_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38424_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_24), .Q(__stream_matmul_15_sink_21_sink_offset_0_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38425_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_25), .Q(__stream_matmul_15_sink_21_sink_offset_0_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38426_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_26), .Q(__stream_matmul_15_sink_21_sink_offset_0_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38427_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_27), .Q(__stream_matmul_15_sink_21_sink_offset_0_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38428_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_28), .Q(__stream_matmul_15_sink_21_sink_offset_0_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38429_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_29), .Q(__stream_matmul_15_sink_21_sink_offset_0_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38430_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_30), .Q(__stream_matmul_15_sink_21_sink_offset_0_31), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38431_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_31), .Q(__stream_matmul_15_sink_21_sink_offset_0_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38432_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_32), .Q(__stream_matmul_15_sink_21_sink_offset_0_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38433_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_33), .Q(__stream_matmul_15_sink_21_sink_offset_0_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38434_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_34), .Q(__stream_matmul_15_sink_21_sink_offset_0_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38435_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_35), .Q(__stream_matmul_15_sink_21_sink_offset_0_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38436_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_offset_0_36), .Q(__stream_matmul_15_sink_21_sink_offset_0_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38437_ ( .CLK(CLK), .D({ 1'h0, matmul_15_next_stream_num_ops }), .Q(__stream_matmul_15_sink_21_sink_size_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38438_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_1), .Q(__stream_matmul_15_sink_21_sink_size_1_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38439_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_2), .Q(__stream_matmul_15_sink_21_sink_size_1_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38440_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_3), .Q(__stream_matmul_15_sink_21_sink_size_1_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38441_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_4), .Q(__stream_matmul_15_sink_21_sink_size_1_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38442_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_5), .Q(__stream_matmul_15_sink_21_sink_size_1_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38443_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_6), .Q(__stream_matmul_15_sink_21_sink_size_1_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38444_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_7), .Q(__stream_matmul_15_sink_21_sink_size_1_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38445_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_8), .Q(__stream_matmul_15_sink_21_sink_size_1_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38446_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_9), .Q(__stream_matmul_15_sink_21_sink_size_1_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38447_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_10), .Q(__stream_matmul_15_sink_21_sink_size_1_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38448_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_11), .Q(__stream_matmul_15_sink_21_sink_size_1_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38449_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_12), .Q(__stream_matmul_15_sink_21_sink_size_1_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38450_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_13), .Q(__stream_matmul_15_sink_21_sink_size_1_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38451_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_14), .Q(__stream_matmul_15_sink_21_sink_size_1_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38452_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_15), .Q(__stream_matmul_15_sink_21_sink_size_1_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38453_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_16), .Q(__stream_matmul_15_sink_21_sink_size_1_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38454_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_17), .Q(__stream_matmul_15_sink_21_sink_size_1_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38455_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_18), .Q(__stream_matmul_15_sink_21_sink_size_1_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38456_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_19), .Q(__stream_matmul_15_sink_21_sink_size_1_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38457_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_20), .Q(__stream_matmul_15_sink_21_sink_size_1_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38458_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_21), .Q(__stream_matmul_15_sink_21_sink_size_1_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38459_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_22), .Q(__stream_matmul_15_sink_21_sink_size_1_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38460_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_23), .Q(__stream_matmul_15_sink_21_sink_size_1_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38461_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_24), .Q(__stream_matmul_15_sink_21_sink_size_1_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38462_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_25), .Q(__stream_matmul_15_sink_21_sink_size_1_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38463_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_26), .Q(__stream_matmul_15_sink_21_sink_size_1_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38464_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_27), .Q(__stream_matmul_15_sink_21_sink_size_1_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38465_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_28), .Q(__stream_matmul_15_sink_21_sink_size_1_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38466_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_29), .Q(__stream_matmul_15_sink_21_sink_size_1_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38467_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_30), .Q(__stream_matmul_15_sink_21_sink_size_1_31), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38468_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_31), .Q(__stream_matmul_15_sink_21_sink_size_1_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38469_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_32), .Q(__stream_matmul_15_sink_21_sink_size_1_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38470_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_33), .Q(__stream_matmul_15_sink_21_sink_size_1_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38471_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_34), .Q(__stream_matmul_15_sink_21_sink_size_1_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38472_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_35), .Q(__stream_matmul_15_sink_21_sink_size_1_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38473_ ( .CLK(CLK), .D(__stream_matmul_15_sink_21_sink_size_1_36), .Q(__stream_matmul_15_sink_21_sink_size_1_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_1_reg ( .CLK(CLK), .D(_set_flag_1034), .Q(__set_flag_1034_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_2_reg ( .CLK(CLK), .D(__set_flag_1034_1), .Q(__set_flag_1034_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_3_reg ( .CLK(CLK), .D(__set_flag_1034_2), .Q(__set_flag_1034_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_4_reg ( .CLK(CLK), .D(__set_flag_1034_3), .Q(__set_flag_1034_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_5_reg ( .CLK(CLK), .D(__set_flag_1034_4), .Q(__set_flag_1034_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_6_reg ( .CLK(CLK), .D(__set_flag_1034_5), .Q(__set_flag_1034_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_7_reg ( .CLK(CLK), .D(__set_flag_1034_6), .Q(__set_flag_1034_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_8_reg ( .CLK(CLK), .D(__set_flag_1034_7), .Q(__set_flag_1034_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_9_reg ( .CLK(CLK), .D(__set_flag_1034_8), .Q(__set_flag_1034_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_10_reg ( .CLK(CLK), .D(__set_flag_1034_9), .Q(__set_flag_1034_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_11_reg ( .CLK(CLK), .D(__set_flag_1034_10), .Q(__set_flag_1034_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_12_reg ( .CLK(CLK), .D(__set_flag_1034_11), .Q(__set_flag_1034_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_13_reg ( .CLK(CLK), .D(__set_flag_1034_12), .Q(__set_flag_1034_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_14_reg ( .CLK(CLK), .D(__set_flag_1034_13), .Q(__set_flag_1034_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_15_reg ( .CLK(CLK), .D(__set_flag_1034_14), .Q(__set_flag_1034_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_16_reg ( .CLK(CLK), .D(__set_flag_1034_15), .Q(__set_flag_1034_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_17_reg ( .CLK(CLK), .D(__set_flag_1034_16), .Q(__set_flag_1034_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_18_reg ( .CLK(CLK), .D(__set_flag_1034_17), .Q(__set_flag_1034_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_19_reg ( .CLK(CLK), .D(__set_flag_1034_18), .Q(__set_flag_1034_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_20_reg ( .CLK(CLK), .D(__set_flag_1034_19), .Q(__set_flag_1034_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_21_reg ( .CLK(CLK), .D(__set_flag_1034_20), .Q(__set_flag_1034_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_22_reg ( .CLK(CLK), .D(__set_flag_1034_21), .Q(__set_flag_1034_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_23_reg ( .CLK(CLK), .D(__set_flag_1034_22), .Q(__set_flag_1034_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_24_reg ( .CLK(CLK), .D(__set_flag_1034_23), .Q(__set_flag_1034_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_25_reg ( .CLK(CLK), .D(__set_flag_1034_24), .Q(__set_flag_1034_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_26_reg ( .CLK(CLK), .D(__set_flag_1034_25), .Q(__set_flag_1034_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_27_reg ( .CLK(CLK), .D(__set_flag_1034_26), .Q(__set_flag_1034_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_28_reg ( .CLK(CLK), .D(__set_flag_1034_27), .Q(__set_flag_1034_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_29_reg ( .CLK(CLK), .D(__set_flag_1034_28), .Q(__set_flag_1034_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_30_reg ( .CLK(CLK), .D(__set_flag_1034_29), .Q(__set_flag_1034_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_31_reg ( .CLK(CLK), .D(__set_flag_1034_30), .Q(__set_flag_1034_31), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_32_reg ( .CLK(CLK), .D(__set_flag_1034_31), .Q(__set_flag_1034_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_33_reg ( .CLK(CLK), .D(__set_flag_1034_32), .Q(__set_flag_1034_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_34_reg ( .CLK(CLK), .D(__set_flag_1034_33), .Q(__set_flag_1034_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_35_reg ( .CLK(CLK), .D(__set_flag_1034_34), .Q(__set_flag_1034_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_36_reg ( .CLK(CLK), .D(__set_flag_1034_35), .Q(__set_flag_1034_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_1034_37_reg ( .CLK(CLK), .D(__set_flag_1034_36), .Q(__set_flag_1034_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_1_reg ( .CLK(CLK), .D(_stream_matmul_15_start), .Q(__stream_matmul_15_start_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_2_reg ( .CLK(CLK), .D(__stream_matmul_15_start_1), .Q(__stream_matmul_15_start_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_3_reg ( .CLK(CLK), .D(__stream_matmul_15_start_2), .Q(__stream_matmul_15_start_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_4_reg ( .CLK(CLK), .D(__stream_matmul_15_start_3), .Q(__stream_matmul_15_start_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_5_reg ( .CLK(CLK), .D(__stream_matmul_15_start_4), .Q(__stream_matmul_15_start_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_6_reg ( .CLK(CLK), .D(__stream_matmul_15_start_5), .Q(__stream_matmul_15_start_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_7_reg ( .CLK(CLK), .D(__stream_matmul_15_start_6), .Q(__stream_matmul_15_start_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_8_reg ( .CLK(CLK), .D(__stream_matmul_15_start_7), .Q(__stream_matmul_15_start_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_9_reg ( .CLK(CLK), .D(__stream_matmul_15_start_8), .Q(__stream_matmul_15_start_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_10_reg ( .CLK(CLK), .D(__stream_matmul_15_start_9), .Q(__stream_matmul_15_start_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_11_reg ( .CLK(CLK), .D(__stream_matmul_15_start_10), .Q(__stream_matmul_15_start_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_12_reg ( .CLK(CLK), .D(__stream_matmul_15_start_11), .Q(__stream_matmul_15_start_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_13_reg ( .CLK(CLK), .D(__stream_matmul_15_start_12), .Q(__stream_matmul_15_start_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_14_reg ( .CLK(CLK), .D(__stream_matmul_15_start_13), .Q(__stream_matmul_15_start_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_15_reg ( .CLK(CLK), .D(__stream_matmul_15_start_14), .Q(__stream_matmul_15_start_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_16_reg ( .CLK(CLK), .D(__stream_matmul_15_start_15), .Q(__stream_matmul_15_start_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_17_reg ( .CLK(CLK), .D(__stream_matmul_15_start_16), .Q(__stream_matmul_15_start_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_18_reg ( .CLK(CLK), .D(__stream_matmul_15_start_17), .Q(__stream_matmul_15_start_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_19_reg ( .CLK(CLK), .D(__stream_matmul_15_start_18), .Q(__stream_matmul_15_start_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_20_reg ( .CLK(CLK), .D(__stream_matmul_15_start_19), .Q(__stream_matmul_15_start_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_21_reg ( .CLK(CLK), .D(__stream_matmul_15_start_20), .Q(__stream_matmul_15_start_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_22_reg ( .CLK(CLK), .D(__stream_matmul_15_start_21), .Q(__stream_matmul_15_start_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_23_reg ( .CLK(CLK), .D(__stream_matmul_15_start_22), .Q(__stream_matmul_15_start_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_24_reg ( .CLK(CLK), .D(__stream_matmul_15_start_23), .Q(__stream_matmul_15_start_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_25_reg ( .CLK(CLK), .D(__stream_matmul_15_start_24), .Q(__stream_matmul_15_start_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_26_reg ( .CLK(CLK), .D(__stream_matmul_15_start_25), .Q(__stream_matmul_15_start_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_27_reg ( .CLK(CLK), .D(__stream_matmul_15_start_26), .Q(__stream_matmul_15_start_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_28_reg ( .CLK(CLK), .D(__stream_matmul_15_start_27), .Q(__stream_matmul_15_start_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_29_reg ( .CLK(CLK), .D(__stream_matmul_15_start_28), .Q(__stream_matmul_15_start_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_30_reg ( .CLK(CLK), .D(__stream_matmul_15_start_29), .Q(__stream_matmul_15_start_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_31_reg ( .CLK(CLK), .D(__stream_matmul_15_start_30), .Q(__stream_matmul_15_start_31), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_32_reg ( .CLK(CLK), .D(__stream_matmul_15_start_31), .Q(__stream_matmul_15_start_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_33_reg ( .CLK(CLK), .D(__stream_matmul_15_start_32), .Q(__stream_matmul_15_start_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_34_reg ( .CLK(CLK), .D(__stream_matmul_15_start_33), .Q(__stream_matmul_15_start_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_35_reg ( .CLK(CLK), .D(__stream_matmul_15_start_34), .Q(__stream_matmul_15_start_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_36_reg ( .CLK(CLK), .D(__stream_matmul_15_start_35), .Q(__stream_matmul_15_start_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_37_reg ( .CLK(CLK), .D(__stream_matmul_15_start_36), .Q(__stream_matmul_15_start_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_matmul_15_start_38_reg ( .CLK(CLK), .D(__stream_matmul_15_start_37), .Q(__stream_matmul_15_start_38), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_1_reg ( .CLK(CLK), .D(_tmp_1037), .Q(__tmp_1059_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_2_reg ( .CLK(CLK), .D(__tmp_1059_1), .Q(__tmp_1059_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_3_reg ( .CLK(CLK), .D(__tmp_1059_2), .Q(__tmp_1059_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_4_reg ( .CLK(CLK), .D(__tmp_1059_3), .Q(__tmp_1059_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_5_reg ( .CLK(CLK), .D(__tmp_1059_4), .Q(__tmp_1059_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_6_reg ( .CLK(CLK), .D(__tmp_1059_5), .Q(__tmp_1059_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_7_reg ( .CLK(CLK), .D(__tmp_1059_6), .Q(__tmp_1059_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_8_reg ( .CLK(CLK), .D(__tmp_1059_7), .Q(__tmp_1059_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_9_reg ( .CLK(CLK), .D(__tmp_1059_8), .Q(__tmp_1059_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_10_reg ( .CLK(CLK), .D(__tmp_1059_9), .Q(__tmp_1059_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_11_reg ( .CLK(CLK), .D(__tmp_1059_10), .Q(__tmp_1059_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_12_reg ( .CLK(CLK), .D(__tmp_1059_11), .Q(__tmp_1059_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_13_reg ( .CLK(CLK), .D(__tmp_1059_12), .Q(__tmp_1059_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_14_reg ( .CLK(CLK), .D(__tmp_1059_13), .Q(__tmp_1059_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_15_reg ( .CLK(CLK), .D(__tmp_1059_14), .Q(__tmp_1059_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_16_reg ( .CLK(CLK), .D(__tmp_1059_15), .Q(__tmp_1059_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_17_reg ( .CLK(CLK), .D(__tmp_1059_16), .Q(__tmp_1059_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_18_reg ( .CLK(CLK), .D(__tmp_1059_17), .Q(__tmp_1059_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_19_reg ( .CLK(CLK), .D(__tmp_1059_18), .Q(__tmp_1059_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_20_reg ( .CLK(CLK), .D(__tmp_1059_19), .Q(__tmp_1059_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_21_reg ( .CLK(CLK), .D(__tmp_1059_20), .Q(__tmp_1059_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_22_reg ( .CLK(CLK), .D(__tmp_1059_21), .Q(__tmp_1059_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_23_reg ( .CLK(CLK), .D(__tmp_1059_22), .Q(__tmp_1059_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_24_reg ( .CLK(CLK), .D(__tmp_1059_23), .Q(__tmp_1059_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_25_reg ( .CLK(CLK), .D(__tmp_1059_24), .Q(__tmp_1059_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_26_reg ( .CLK(CLK), .D(__tmp_1059_25), .Q(__tmp_1059_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_27_reg ( .CLK(CLK), .D(__tmp_1059_26), .Q(__tmp_1059_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1059_28_reg ( .CLK(CLK), .D(__tmp_1059_27), .Q(__tmp_1059_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1115_35_reg ( .CLK(CLK), .D(__tmp_1117_34), .Q(__tmp_1115_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1115_36_reg ( .CLK(CLK), .D(__tmp_1115_35), .Q(__tmp_1115_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1115_37_reg ( .CLK(CLK), .D(__tmp_1115_36), .Q(__tmp_1115_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1115_38_reg ( .CLK(CLK), .D(__tmp_1115_37), .Q(__tmp_1115_38), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_13_reg ( .CLK(CLK), .D(__tmp_1107_12), .Q(__tmp_1117_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_14_reg ( .CLK(CLK), .D(__tmp_1117_13), .Q(__tmp_1117_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_15_reg ( .CLK(CLK), .D(__tmp_1117_14), .Q(__tmp_1117_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_16_reg ( .CLK(CLK), .D(__tmp_1117_15), .Q(__tmp_1117_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_17_reg ( .CLK(CLK), .D(__tmp_1117_16), .Q(__tmp_1117_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_18_reg ( .CLK(CLK), .D(__tmp_1117_17), .Q(__tmp_1117_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_19_reg ( .CLK(CLK), .D(__tmp_1117_18), .Q(__tmp_1117_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_20_reg ( .CLK(CLK), .D(__tmp_1117_19), .Q(__tmp_1117_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_21_reg ( .CLK(CLK), .D(__tmp_1117_20), .Q(__tmp_1117_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_22_reg ( .CLK(CLK), .D(__tmp_1117_21), .Q(__tmp_1117_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_23_reg ( .CLK(CLK), .D(__tmp_1117_22), .Q(__tmp_1117_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_24_reg ( .CLK(CLK), .D(__tmp_1117_23), .Q(__tmp_1117_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_25_reg ( .CLK(CLK), .D(__tmp_1117_24), .Q(__tmp_1117_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_26_reg ( .CLK(CLK), .D(__tmp_1117_25), .Q(__tmp_1117_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_27_reg ( .CLK(CLK), .D(__tmp_1117_26), .Q(__tmp_1117_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_28_reg ( .CLK(CLK), .D(__tmp_1117_27), .Q(__tmp_1117_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_29_reg ( .CLK(CLK), .D(__tmp_1117_28), .Q(__tmp_1117_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_30_reg ( .CLK(CLK), .D(__tmp_1117_29), .Q(__tmp_1117_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_31_reg ( .CLK(CLK), .D(__tmp_1117_30), .Q(__tmp_1117_31), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_32_reg ( .CLK(CLK), .D(__tmp_1117_31), .Q(__tmp_1117_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_33_reg ( .CLK(CLK), .D(__tmp_1117_32), .Q(__tmp_1117_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1117_34_reg ( .CLK(CLK), .D(__tmp_1117_33), .Q(__tmp_1117_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38603_ ( .CLK(CLK), .D(_23122_), .Q(_stream_max_pool_serial_9_fsm), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_max_pool_serial_9_start_reg ( .CLK(CLK), .D(_23121_), .Q(_stream_max_pool_serial_9_start), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_max_pool_serial_9_end_flag_reg ( .CLK(CLK), .D(_23119_), .Q(_stream_max_pool_serial_9_end_flag), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_max_pool_serial_9_term_sink_reg ( .CLK(CLK), .D(_23118_), .Q(_stream_max_pool_serial_9_term_sink), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_max_pool_serial_9_source_busy_reg ( .CLK(CLK), .D(_23117_), .Q(_stream_max_pool_serial_9_source_busy), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_max_pool_serial_9_reduce_reset_reg  ( .CLK(CLK), .D(_02647_), .Q(_stream_max_pool_serial_9_reduce_reset) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38609_ ( .CLK(CLK), .D(_23194_), .Q(_stream_max_pool_serial_9_constant_0_next_constant_data), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_max_pool_serial_9_source_1_idle_reg  ( .CLK(CLK), .D(_02659_), .Q(_stream_max_pool_serial_9_source_1_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38611_ ( .CLK(CLK), .D(_23191_), .Q(_stream_max_pool_serial_9_source_1_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38612_ ( .CLK(CLK), .D(_23190_), .Q(_stream_max_pool_serial_9_source_1_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38613_ ( .CLK(CLK), .D(_23189_), .Q(_stream_max_pool_serial_9_source_1_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38614_ ( .CLK(CLK), .D(_23188_), .Q(_stream_max_pool_serial_9_source_1_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38615_ ( .CLK(CLK), .D(_23187_), .Q(_stream_max_pool_serial_9_source_1_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_max_pool_serial_9_source_1_source_ram_renable_reg ( .CLK(CLK), .D(_23186_), .Q(_stream_max_pool_serial_9_source_1_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_max_pool_serial_9_source_1_source_ram_rvalid_reg ( .CLK(CLK), .D(_23184_), .Q(_stream_max_pool_serial_9_source_1_source_ram_rvalid), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _38618_ ( .CLK(CLK), .D(_23183_), .Q(_stream_max_pool_serial_9_constant_2_next_constant_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38619_ ( .CLK(CLK), .D(_23182_), .Q(_stream_max_pool_serial_9_sink_3_sink_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38620_ ( .CLK(CLK), .D(_23181_), .Q(_stream_max_pool_serial_9_sink_3_sink_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38621_ ( .CLK(CLK), .D(_23180_), .Q(_stream_max_pool_serial_9_sink_3_sink_size), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38622_ ( .CLK(CLK), .D(_23179_), .Q(_stream_max_pool_serial_9_sink_3_sink_stride), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38623_ ( .CLK(CLK), .D(_23178_), .Q(_stream_max_pool_serial_9_sink_3_sink_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38624_ ( .CLK(CLK), .D(_23176_), .Q(_stream_max_pool_serial_9_sink_3_sink_stride_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38625_ ( .CLK(CLK), .D(_23175_), .Q(_stream_max_pool_serial_9_sink_3_sink_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38626_ ( .CLK(CLK), .D(_23174_), .Q(_stream_max_pool_serial_9_sink_3_sink_waddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_max_pool_serial_9_sink_3_sink_wenable_reg ( .CLK(CLK), .D(_23172_), .Q(_stream_max_pool_serial_9_sink_3_sink_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38628_ ( .CLK(CLK), .D(_23171_), .Q(_stream_max_pool_serial_9_sink_3_sink_wdata), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _38629_ ( .CLK(CLK), .D(_01468_), .Q(_counter_data_762) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _38630_ ( .CLK(CLK), .D(_23168_), .Q(_counter_count_762), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _38631_ ( .CLK(CLK), .D(__variable_wdata_759), .Q(__delay_data_1372), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38632_ ( .CLK(CLK), .D(__variable_wdata_758), .Q(__delay_data_1373), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38633_ ( .CLK(CLK), .D(__variable_wdata_757), .Q(__delay_data_1375), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pointer_data_764_reg ( .CLK(CLK), .D(_25911_[0]), .Q(_pointer_data_764), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38635_ ( .CLK(CLK), .D(__delay_data_1373), .Q(__delay_data_1374), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38636_ ( .CLK(CLK), .D(__delay_data_1375), .Q(__delay_data_1376), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38637_ ( .CLK(CLK), .D(_26631_), .Q(_cond_data_771), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38638_ ( .CLK(CLK), .D(__delay_data_1376), .Q(__delay_data_1377), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38639_ ( .CLK(CLK), .D(_reducecustom_data_191), .Q(__substreamoutput_data_773), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __substreamoutput_data_774_reg ( .CLK(CLK), .D(_pulse_data_193), .Q(__substreamoutput_data_774), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38641_ ( .CLK(CLK), .D(_23167_), .Q(__variable_wdata_757), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _38642_ ( .CLK(CLK), .D(_23166_), .Q(__variable_wdata_759), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38643_ ( .CLK(CLK), .D(_23165_), .Q(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38644_ ( .CLK(CLK), .D(_23162_), .Q(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38645_ ( .CLK(CLK), .D(_23159_), .Q(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38646_ ( .CLK(CLK), .D(_23156_), .Q(_source_stream_max_pool_serial_9_source_1_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38647_ ( .CLK(CLK), .D(_23153_), .Q(_source_stream_max_pool_serial_9_source_1_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38648_ ( .CLK(CLK), .D(_23152_), .Q(_source_stream_max_pool_serial_9_source_1_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38649_ ( .CLK(CLK), .D(_23151_), .Q(_source_stream_max_pool_serial_9_source_1_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38650_ ( .CLK(CLK), .D(_23150_), .Q(_source_stream_max_pool_serial_9_source_1_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38651_ ( .CLK(CLK), .D(_23149_), .Q(_source_stream_max_pool_serial_9_source_1_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38652_ ( .CLK(CLK), .D(_23148_), .Q(_source_stream_max_pool_serial_9_source_1_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38653_ ( .CLK(CLK), .D(_23147_), .Q(_source_stream_max_pool_serial_9_source_1_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38654_ ( .CLK(CLK), .D(_23146_), .Q(_source_stream_max_pool_serial_9_source_1_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38655_ ( .CLK(CLK), .D(_23145_), .Q(_source_stream_max_pool_serial_9_source_1_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38656_ ( .CLK(CLK), .D(_23142_), .Q(_source_stream_max_pool_serial_9_source_1_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38657_ ( .CLK(CLK), .D(_23139_), .Q(_source_stream_max_pool_serial_9_source_1_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38658_ ( .CLK(CLK), .D(_23136_), .Q(_source_stream_max_pool_serial_9_source_1_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38659_ ( .CLK(CLK), .D(_23133_), .Q(_source_stream_max_pool_serial_9_source_1_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38660_ ( .CLK(CLK), .D(_23132_), .Q(_source_stream_max_pool_serial_9_source_1_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38661_ ( .CLK(CLK), .D(_23131_), .Q(_source_stream_max_pool_serial_9_source_1_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38662_ ( .CLK(CLK), .D(_23130_), .Q(_source_stream_max_pool_serial_9_source_1_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38663_ ( .CLK(CLK), .D(_23129_), .Q(_source_stream_max_pool_serial_9_source_1_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38664_ ( .CLK(CLK), .D(_23128_), .Q(_source_stream_max_pool_serial_9_source_1_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38665_ ( .CLK(CLK), .D(_23127_), .Q(_source_stream_max_pool_serial_9_source_1_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38666_ ( .CLK(CLK), .D(_23126_), .Q(_source_stream_max_pool_serial_9_source_1_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38667_ ( .CLK(CLK), .D(_23125_), .Q(__variable_wdata_758), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _set_flag_874_reg ( .CLK(CLK), .D(_23124_), .Q(_set_flag_874), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38669_ ( .CLK(CLK), .D(_22238_), .Q(__stream_max_pool_serial_9_sink_3_sink_offset_0_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38670_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_offset_0_1), .Q(__stream_max_pool_serial_9_sink_3_sink_offset_0_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38671_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_offset_0_2), .Q(__stream_max_pool_serial_9_sink_3_sink_offset_0_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38672_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_offset_0_3), .Q(__stream_max_pool_serial_9_sink_3_sink_offset_0_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38673_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_offset_0_4), .Q(__stream_max_pool_serial_9_sink_3_sink_offset_0_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38674_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_offset_0_5), .Q(__stream_max_pool_serial_9_sink_3_sink_offset_0_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38675_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_offset_0_6), .Q(__stream_max_pool_serial_9_sink_3_sink_offset_0_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38676_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_offset_0_7), .Q(__stream_max_pool_serial_9_sink_3_sink_offset_0_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38677_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_offset_0_8), .Q(__stream_max_pool_serial_9_sink_3_sink_offset_0_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38678_ ( .CLK(CLK), .D({ 28'h0000000, cparam_max_pool_serial_9_inc_out_laddr }), .Q(__stream_max_pool_serial_9_sink_3_sink_size_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38679_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_size_1_1), .Q(__stream_max_pool_serial_9_sink_3_sink_size_1_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38680_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_size_1_2), .Q(__stream_max_pool_serial_9_sink_3_sink_size_1_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38681_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_size_1_3), .Q(__stream_max_pool_serial_9_sink_3_sink_size_1_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38682_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_size_1_4), .Q(__stream_max_pool_serial_9_sink_3_sink_size_1_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38683_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_size_1_5), .Q(__stream_max_pool_serial_9_sink_3_sink_size_1_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38684_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_size_1_6), .Q(__stream_max_pool_serial_9_sink_3_sink_size_1_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38685_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_size_1_7), .Q(__stream_max_pool_serial_9_sink_3_sink_size_1_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38686_ ( .CLK(CLK), .D(__stream_max_pool_serial_9_sink_3_sink_size_1_8), .Q(__stream_max_pool_serial_9_sink_3_sink_size_1_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_874_1_reg ( .CLK(CLK), .D(_set_flag_874), .Q(__set_flag_874_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_874_2_reg ( .CLK(CLK), .D(__set_flag_874_1), .Q(__set_flag_874_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_874_3_reg ( .CLK(CLK), .D(__set_flag_874_2), .Q(__set_flag_874_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_874_4_reg ( .CLK(CLK), .D(__set_flag_874_3), .Q(__set_flag_874_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_874_5_reg ( .CLK(CLK), .D(__set_flag_874_4), .Q(__set_flag_874_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_874_6_reg ( .CLK(CLK), .D(__set_flag_874_5), .Q(__set_flag_874_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_874_7_reg ( .CLK(CLK), .D(__set_flag_874_6), .Q(__set_flag_874_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_874_8_reg ( .CLK(CLK), .D(__set_flag_874_7), .Q(__set_flag_874_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_874_9_reg ( .CLK(CLK), .D(__set_flag_874_8), .Q(__set_flag_874_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_max_pool_serial_9_start_1_reg ( .CLK(CLK), .D(_stream_max_pool_serial_9_start), .Q(__stream_max_pool_serial_9_start_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_max_pool_serial_9_start_2_reg ( .CLK(CLK), .D(__stream_max_pool_serial_9_start_1), .Q(__stream_max_pool_serial_9_start_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_max_pool_serial_9_start_3_reg ( .CLK(CLK), .D(__stream_max_pool_serial_9_start_2), .Q(__stream_max_pool_serial_9_start_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_max_pool_serial_9_start_4_reg ( .CLK(CLK), .D(__stream_max_pool_serial_9_start_3), .Q(__stream_max_pool_serial_9_start_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_max_pool_serial_9_start_5_reg ( .CLK(CLK), .D(__stream_max_pool_serial_9_start_4), .Q(__stream_max_pool_serial_9_start_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_max_pool_serial_9_start_6_reg ( .CLK(CLK), .D(__stream_max_pool_serial_9_start_5), .Q(__stream_max_pool_serial_9_start_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_max_pool_serial_9_start_7_reg ( .CLK(CLK), .D(__stream_max_pool_serial_9_start_6), .Q(__stream_max_pool_serial_9_start_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_max_pool_serial_9_start_8_reg ( .CLK(CLK), .D(__stream_max_pool_serial_9_start_7), .Q(__stream_max_pool_serial_9_start_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_max_pool_serial_9_start_9_reg ( .CLK(CLK), .D(__stream_max_pool_serial_9_start_8), .Q(__stream_max_pool_serial_9_start_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_max_pool_serial_9_start_10_reg ( .CLK(CLK), .D(__stream_max_pool_serial_9_start_9), .Q(__stream_max_pool_serial_9_start_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _set_flag_876_reg ( .CLK(CLK), .D(_23123_), .Q(_set_flag_876), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_880_8_reg ( .CLK(CLK), .D(__tmp_884_7), .Q(__tmp_880_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_880_9_reg ( .CLK(CLK), .D(__tmp_880_8), .Q(__tmp_880_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_884_1_reg ( .CLK(CLK), .D(_tmp_878), .Q(__tmp_884_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_884_2_reg ( .CLK(CLK), .D(__tmp_884_1), .Q(__tmp_884_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_884_3_reg ( .CLK(CLK), .D(__tmp_884_2), .Q(__tmp_884_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_884_4_reg ( .CLK(CLK), .D(__tmp_884_3), .Q(__tmp_884_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_884_5_reg ( .CLK(CLK), .D(__tmp_884_4), .Q(__tmp_884_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_884_6_reg ( .CLK(CLK), .D(__tmp_884_5), .Q(__tmp_884_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_884_7_reg ( .CLK(CLK), .D(__tmp_884_6), .Q(__tmp_884_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_906_7_reg ( .CLK(CLK), .D(__tmp_908_6), .Q(__tmp_906_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_906_8_reg ( .CLK(CLK), .D(__tmp_906_7), .Q(__tmp_906_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_906_9_reg ( .CLK(CLK), .D(__tmp_906_8), .Q(__tmp_906_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_906_10_reg ( .CLK(CLK), .D(__tmp_906_9), .Q(__tmp_906_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_908_1_reg ( .CLK(CLK), .D(_tmp_894), .Q(__tmp_908_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_908_2_reg ( .CLK(CLK), .D(__tmp_908_1), .Q(__tmp_908_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_908_3_reg ( .CLK(CLK), .D(__tmp_908_2), .Q(__tmp_908_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_908_4_reg ( .CLK(CLK), .D(__tmp_908_3), .Q(__tmp_908_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_908_5_reg ( .CLK(CLK), .D(__tmp_908_4), .Q(__tmp_908_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_908_6_reg ( .CLK(CLK), .D(__tmp_908_5), .Q(__tmp_908_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38726_ ( .CLK(CLK), .D(_23200_), .Q(_stream_conv2d_8_fsm), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_start_reg ( .CLK(CLK), .D(_23199_), .Q(_stream_conv2d_8_start), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_end_flag_reg ( .CLK(CLK), .D(_23197_), .Q(_stream_conv2d_8_end_flag), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_term_sink_reg ( .CLK(CLK), .D(_23196_), .Q(_stream_conv2d_8_term_sink), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_busy_reg ( .CLK(CLK), .D(_23195_), .Q(_stream_conv2d_8_source_busy), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _38731_ ( .CLK(CLK), .D(_24256_), .Q(_stream_conv2d_8_constant_0_next_constant_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _38732_ ( .CLK(CLK), .D(_24255_), .Q(_stream_conv2d_8_constant_1_next_constant_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _38733_ ( .CLK(CLK), .D(_24254_), .Q(_stream_conv2d_8_constant_2_next_constant_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _38734_ ( .CLK(CLK), .D(_24253_), .Q(_stream_conv2d_8_constant_3_next_constant_data), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_6_idle_reg  ( .CLK(CLK), .D(_02557_), .Q(_stream_conv2d_8_source_6_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38736_ ( .CLK(CLK), .D(_24250_), .Q(_stream_conv2d_8_source_6_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38737_ ( .CLK(CLK), .D(_24249_), .Q(_stream_conv2d_8_source_6_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38738_ ( .CLK(CLK), .D(_24248_), .Q(_stream_conv2d_8_source_6_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38739_ ( .CLK(CLK), .D(_24247_), .Q(_stream_conv2d_8_source_6_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38740_ ( .CLK(CLK), .D(_24246_), .Q(_stream_conv2d_8_source_6_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_6_source_ram_renable_reg ( .CLK(CLK), .D(_24245_), .Q(_stream_conv2d_8_source_6_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_6_source_ram_rvalid_reg ( .CLK(CLK), .D(_24243_), .Q(_stream_conv2d_8_source_6_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_8_idle_reg  ( .CLK(CLK), .D(_02566_), .Q(_stream_conv2d_8_source_8_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38744_ ( .CLK(CLK), .D(_24240_), .Q(_stream_conv2d_8_source_8_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38745_ ( .CLK(CLK), .D(_24239_), .Q(_stream_conv2d_8_source_8_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38746_ ( .CLK(CLK), .D(_24238_), .Q(_stream_conv2d_8_source_8_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38747_ ( .CLK(CLK), .D(_24237_), .Q(_stream_conv2d_8_source_8_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38748_ ( .CLK(CLK), .D(_24236_), .Q(_stream_conv2d_8_source_8_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_8_source_ram_renable_reg ( .CLK(CLK), .D(_24235_), .Q(_stream_conv2d_8_source_8_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_8_source_ram_rvalid_reg ( .CLK(CLK), .D(_24233_), .Q(_stream_conv2d_8_source_8_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_10_idle_reg  ( .CLK(CLK), .D(_02389_), .Q(_stream_conv2d_8_source_10_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38752_ ( .CLK(CLK), .D(_24231_), .Q(_stream_conv2d_8_source_10_source_empty_data), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_12_idle_reg  ( .CLK(CLK), .D(_02391_), .Q(_stream_conv2d_8_source_12_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38754_ ( .CLK(CLK), .D(_24229_), .Q(_stream_conv2d_8_source_12_source_empty_data), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_14_idle_reg  ( .CLK(CLK), .D(_02393_), .Q(_stream_conv2d_8_source_14_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38756_ ( .CLK(CLK), .D(_24227_), .Q(_stream_conv2d_8_source_14_source_empty_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_constant_15_next_constant_data_reg ( .CLK(CLK), .D(_24226_), .Q(_stream_conv2d_8_constant_15_next_constant_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_constant_16_next_constant_data_reg ( .CLK(CLK), .D(_24225_), .Q(_stream_conv2d_8_constant_16_next_constant_data), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _38759_ ( .CLK(CLK), .D(_24224_), .Q(_stream_conv2d_8_constant_17_next_constant_data), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_19_idle_reg  ( .CLK(CLK), .D(_02395_), .Q(_stream_conv2d_8_source_19_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38761_ ( .CLK(CLK), .D(_24221_), .Q(_stream_conv2d_8_source_19_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38762_ ( .CLK(CLK), .D(_24220_), .Q(_stream_conv2d_8_source_19_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38763_ ( .CLK(CLK), .D(_24219_), .Q(_stream_conv2d_8_source_19_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38764_ ( .CLK(CLK), .D(_24218_), .Q(_stream_conv2d_8_source_19_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38765_ ( .CLK(CLK), .D(_24217_), .Q(_stream_conv2d_8_source_19_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_19_source_ram_renable_reg ( .CLK(CLK), .D(_24216_), .Q(_stream_conv2d_8_source_19_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_19_source_ram_rvalid_reg ( .CLK(CLK), .D(_24214_), .Q(_stream_conv2d_8_source_19_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_20_idle_reg  ( .CLK(CLK), .D(_02404_), .Q(_stream_conv2d_8_source_20_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38769_ ( .CLK(CLK), .D(_24211_), .Q(_stream_conv2d_8_source_20_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38770_ ( .CLK(CLK), .D(_24210_), .Q(_stream_conv2d_8_source_20_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38771_ ( .CLK(CLK), .D(_24209_), .Q(_stream_conv2d_8_source_20_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38772_ ( .CLK(CLK), .D(_24208_), .Q(_stream_conv2d_8_source_20_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38773_ ( .CLK(CLK), .D(_24207_), .Q(_stream_conv2d_8_source_20_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_20_source_ram_renable_reg ( .CLK(CLK), .D(_24206_), .Q(_stream_conv2d_8_source_20_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_20_source_ram_rvalid_reg ( .CLK(CLK), .D(_24204_), .Q(_stream_conv2d_8_source_20_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_21_idle_reg  ( .CLK(CLK), .D(_02413_), .Q(_stream_conv2d_8_source_21_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38777_ ( .CLK(CLK), .D(_24201_), .Q(_stream_conv2d_8_source_21_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38778_ ( .CLK(CLK), .D(_24200_), .Q(_stream_conv2d_8_source_21_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38779_ ( .CLK(CLK), .D(_24199_), .Q(_stream_conv2d_8_source_21_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38780_ ( .CLK(CLK), .D(_24198_), .Q(_stream_conv2d_8_source_21_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38781_ ( .CLK(CLK), .D(_24197_), .Q(_stream_conv2d_8_source_21_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_21_source_ram_renable_reg ( .CLK(CLK), .D(_24196_), .Q(_stream_conv2d_8_source_21_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_21_source_ram_rvalid_reg ( .CLK(CLK), .D(_24194_), .Q(_stream_conv2d_8_source_21_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_22_idle_reg  ( .CLK(CLK), .D(_02422_), .Q(_stream_conv2d_8_source_22_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38785_ ( .CLK(CLK), .D(_24191_), .Q(_stream_conv2d_8_source_22_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38786_ ( .CLK(CLK), .D(_24190_), .Q(_stream_conv2d_8_source_22_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38787_ ( .CLK(CLK), .D(_24189_), .Q(_stream_conv2d_8_source_22_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38788_ ( .CLK(CLK), .D(_24188_), .Q(_stream_conv2d_8_source_22_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38789_ ( .CLK(CLK), .D(_24187_), .Q(_stream_conv2d_8_source_22_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_22_source_ram_renable_reg ( .CLK(CLK), .D(_24186_), .Q(_stream_conv2d_8_source_22_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_22_source_ram_rvalid_reg ( .CLK(CLK), .D(_24184_), .Q(_stream_conv2d_8_source_22_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_23_idle_reg  ( .CLK(CLK), .D(_02431_), .Q(_stream_conv2d_8_source_23_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38793_ ( .CLK(CLK), .D(_24181_), .Q(_stream_conv2d_8_source_23_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38794_ ( .CLK(CLK), .D(_24180_), .Q(_stream_conv2d_8_source_23_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38795_ ( .CLK(CLK), .D(_24179_), .Q(_stream_conv2d_8_source_23_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38796_ ( .CLK(CLK), .D(_24178_), .Q(_stream_conv2d_8_source_23_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38797_ ( .CLK(CLK), .D(_24177_), .Q(_stream_conv2d_8_source_23_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_23_source_ram_renable_reg ( .CLK(CLK), .D(_24176_), .Q(_stream_conv2d_8_source_23_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_23_source_ram_rvalid_reg ( .CLK(CLK), .D(_24174_), .Q(_stream_conv2d_8_source_23_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_24_idle_reg  ( .CLK(CLK), .D(_02440_), .Q(_stream_conv2d_8_source_24_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38801_ ( .CLK(CLK), .D(_24171_), .Q(_stream_conv2d_8_source_24_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38802_ ( .CLK(CLK), .D(_24170_), .Q(_stream_conv2d_8_source_24_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38803_ ( .CLK(CLK), .D(_24169_), .Q(_stream_conv2d_8_source_24_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38804_ ( .CLK(CLK), .D(_24168_), .Q(_stream_conv2d_8_source_24_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38805_ ( .CLK(CLK), .D(_24167_), .Q(_stream_conv2d_8_source_24_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_24_source_ram_renable_reg ( .CLK(CLK), .D(_24166_), .Q(_stream_conv2d_8_source_24_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_24_source_ram_rvalid_reg ( .CLK(CLK), .D(_24164_), .Q(_stream_conv2d_8_source_24_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_25_idle_reg  ( .CLK(CLK), .D(_02449_), .Q(_stream_conv2d_8_source_25_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38809_ ( .CLK(CLK), .D(_24161_), .Q(_stream_conv2d_8_source_25_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38810_ ( .CLK(CLK), .D(_24160_), .Q(_stream_conv2d_8_source_25_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38811_ ( .CLK(CLK), .D(_24159_), .Q(_stream_conv2d_8_source_25_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38812_ ( .CLK(CLK), .D(_24158_), .Q(_stream_conv2d_8_source_25_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38813_ ( .CLK(CLK), .D(_24157_), .Q(_stream_conv2d_8_source_25_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_25_source_ram_renable_reg ( .CLK(CLK), .D(_24156_), .Q(_stream_conv2d_8_source_25_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_25_source_ram_rvalid_reg ( .CLK(CLK), .D(_24154_), .Q(_stream_conv2d_8_source_25_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_26_idle_reg  ( .CLK(CLK), .D(_02458_), .Q(_stream_conv2d_8_source_26_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38817_ ( .CLK(CLK), .D(_24151_), .Q(_stream_conv2d_8_source_26_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38818_ ( .CLK(CLK), .D(_24150_), .Q(_stream_conv2d_8_source_26_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38819_ ( .CLK(CLK), .D(_24149_), .Q(_stream_conv2d_8_source_26_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38820_ ( .CLK(CLK), .D(_24148_), .Q(_stream_conv2d_8_source_26_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38821_ ( .CLK(CLK), .D(_24147_), .Q(_stream_conv2d_8_source_26_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_26_source_ram_renable_reg ( .CLK(CLK), .D(_24146_), .Q(_stream_conv2d_8_source_26_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_26_source_ram_rvalid_reg ( .CLK(CLK), .D(_24144_), .Q(_stream_conv2d_8_source_26_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_27_idle_reg  ( .CLK(CLK), .D(_02467_), .Q(_stream_conv2d_8_source_27_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38825_ ( .CLK(CLK), .D(_24141_), .Q(_stream_conv2d_8_source_27_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38826_ ( .CLK(CLK), .D(_24140_), .Q(_stream_conv2d_8_source_27_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38827_ ( .CLK(CLK), .D(_24139_), .Q(_stream_conv2d_8_source_27_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38828_ ( .CLK(CLK), .D(_24138_), .Q(_stream_conv2d_8_source_27_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38829_ ( .CLK(CLK), .D(_24137_), .Q(_stream_conv2d_8_source_27_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_27_source_ram_renable_reg ( .CLK(CLK), .D(_24136_), .Q(_stream_conv2d_8_source_27_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_27_source_ram_rvalid_reg ( .CLK(CLK), .D(_24134_), .Q(_stream_conv2d_8_source_27_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_28_idle_reg  ( .CLK(CLK), .D(_02476_), .Q(_stream_conv2d_8_source_28_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38833_ ( .CLK(CLK), .D(_24131_), .Q(_stream_conv2d_8_source_28_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38834_ ( .CLK(CLK), .D(_24130_), .Q(_stream_conv2d_8_source_28_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38835_ ( .CLK(CLK), .D(_24129_), .Q(_stream_conv2d_8_source_28_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38836_ ( .CLK(CLK), .D(_24128_), .Q(_stream_conv2d_8_source_28_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38837_ ( .CLK(CLK), .D(_24127_), .Q(_stream_conv2d_8_source_28_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_28_source_ram_renable_reg ( .CLK(CLK), .D(_24126_), .Q(_stream_conv2d_8_source_28_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_28_source_ram_rvalid_reg ( .CLK(CLK), .D(_24124_), .Q(_stream_conv2d_8_source_28_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_29_idle_reg  ( .CLK(CLK), .D(_02485_), .Q(_stream_conv2d_8_source_29_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38841_ ( .CLK(CLK), .D(_24121_), .Q(_stream_conv2d_8_source_29_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38842_ ( .CLK(CLK), .D(_24120_), .Q(_stream_conv2d_8_source_29_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38843_ ( .CLK(CLK), .D(_24119_), .Q(_stream_conv2d_8_source_29_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38844_ ( .CLK(CLK), .D(_24118_), .Q(_stream_conv2d_8_source_29_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38845_ ( .CLK(CLK), .D(_24117_), .Q(_stream_conv2d_8_source_29_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_29_source_ram_renable_reg ( .CLK(CLK), .D(_24116_), .Q(_stream_conv2d_8_source_29_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_29_source_ram_rvalid_reg ( .CLK(CLK), .D(_24114_), .Q(_stream_conv2d_8_source_29_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_30_idle_reg  ( .CLK(CLK), .D(_02494_), .Q(_stream_conv2d_8_source_30_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38849_ ( .CLK(CLK), .D(_24111_), .Q(_stream_conv2d_8_source_30_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38850_ ( .CLK(CLK), .D(_24110_), .Q(_stream_conv2d_8_source_30_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38851_ ( .CLK(CLK), .D(_24109_), .Q(_stream_conv2d_8_source_30_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38852_ ( .CLK(CLK), .D(_24108_), .Q(_stream_conv2d_8_source_30_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38853_ ( .CLK(CLK), .D(_24107_), .Q(_stream_conv2d_8_source_30_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_30_source_ram_renable_reg ( .CLK(CLK), .D(_24106_), .Q(_stream_conv2d_8_source_30_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_30_source_ram_rvalid_reg ( .CLK(CLK), .D(_24104_), .Q(_stream_conv2d_8_source_30_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_31_idle_reg  ( .CLK(CLK), .D(_02503_), .Q(_stream_conv2d_8_source_31_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38857_ ( .CLK(CLK), .D(_24101_), .Q(_stream_conv2d_8_source_31_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38858_ ( .CLK(CLK), .D(_24100_), .Q(_stream_conv2d_8_source_31_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38859_ ( .CLK(CLK), .D(_24099_), .Q(_stream_conv2d_8_source_31_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38860_ ( .CLK(CLK), .D(_24098_), .Q(_stream_conv2d_8_source_31_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38861_ ( .CLK(CLK), .D(_24097_), .Q(_stream_conv2d_8_source_31_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_31_source_ram_renable_reg ( .CLK(CLK), .D(_24096_), .Q(_stream_conv2d_8_source_31_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_31_source_ram_rvalid_reg ( .CLK(CLK), .D(_24094_), .Q(_stream_conv2d_8_source_31_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_32_idle_reg  ( .CLK(CLK), .D(_02512_), .Q(_stream_conv2d_8_source_32_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38865_ ( .CLK(CLK), .D(_24091_), .Q(_stream_conv2d_8_source_32_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38866_ ( .CLK(CLK), .D(_24090_), .Q(_stream_conv2d_8_source_32_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38867_ ( .CLK(CLK), .D(_24089_), .Q(_stream_conv2d_8_source_32_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38868_ ( .CLK(CLK), .D(_24088_), .Q(_stream_conv2d_8_source_32_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38869_ ( .CLK(CLK), .D(_24087_), .Q(_stream_conv2d_8_source_32_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_32_source_ram_renable_reg ( .CLK(CLK), .D(_24086_), .Q(_stream_conv2d_8_source_32_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_32_source_ram_rvalid_reg ( .CLK(CLK), .D(_24084_), .Q(_stream_conv2d_8_source_32_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_33_idle_reg  ( .CLK(CLK), .D(_02521_), .Q(_stream_conv2d_8_source_33_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38873_ ( .CLK(CLK), .D(_24081_), .Q(_stream_conv2d_8_source_33_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38874_ ( .CLK(CLK), .D(_24080_), .Q(_stream_conv2d_8_source_33_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38875_ ( .CLK(CLK), .D(_24079_), .Q(_stream_conv2d_8_source_33_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38876_ ( .CLK(CLK), .D(_24078_), .Q(_stream_conv2d_8_source_33_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38877_ ( .CLK(CLK), .D(_24077_), .Q(_stream_conv2d_8_source_33_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_33_source_ram_renable_reg ( .CLK(CLK), .D(_24076_), .Q(_stream_conv2d_8_source_33_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_33_source_ram_rvalid_reg ( .CLK(CLK), .D(_24074_), .Q(_stream_conv2d_8_source_33_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_34_idle_reg  ( .CLK(CLK), .D(_02530_), .Q(_stream_conv2d_8_source_34_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38881_ ( .CLK(CLK), .D(_24071_), .Q(_stream_conv2d_8_source_34_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38882_ ( .CLK(CLK), .D(_24070_), .Q(_stream_conv2d_8_source_34_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38883_ ( .CLK(CLK), .D(_24069_), .Q(_stream_conv2d_8_source_34_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38884_ ( .CLK(CLK), .D(_24068_), .Q(_stream_conv2d_8_source_34_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38885_ ( .CLK(CLK), .D(_24067_), .Q(_stream_conv2d_8_source_34_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_34_source_ram_renable_reg ( .CLK(CLK), .D(_24066_), .Q(_stream_conv2d_8_source_34_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_34_source_ram_rvalid_reg ( .CLK(CLK), .D(_24064_), .Q(_stream_conv2d_8_source_34_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_35_idle_reg  ( .CLK(CLK), .D(_02539_), .Q(_stream_conv2d_8_source_35_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38889_ ( .CLK(CLK), .D(_24061_), .Q(_stream_conv2d_8_source_35_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38890_ ( .CLK(CLK), .D(_24060_), .Q(_stream_conv2d_8_source_35_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38891_ ( .CLK(CLK), .D(_24059_), .Q(_stream_conv2d_8_source_35_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38892_ ( .CLK(CLK), .D(_24058_), .Q(_stream_conv2d_8_source_35_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38893_ ( .CLK(CLK), .D(_24057_), .Q(_stream_conv2d_8_source_35_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_35_source_ram_renable_reg ( .CLK(CLK), .D(_24056_), .Q(_stream_conv2d_8_source_35_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_35_source_ram_rvalid_reg ( .CLK(CLK), .D(_24054_), .Q(_stream_conv2d_8_source_35_source_ram_rvalid), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_8_source_36_idle_reg  ( .CLK(CLK), .D(_02548_), .Q(_stream_conv2d_8_source_36_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38897_ ( .CLK(CLK), .D(_24051_), .Q(_stream_conv2d_8_source_36_source_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38898_ ( .CLK(CLK), .D(_24050_), .Q(_stream_conv2d_8_source_36_source_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38899_ ( .CLK(CLK), .D(_24049_), .Q(_stream_conv2d_8_source_36_source_offset_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38900_ ( .CLK(CLK), .D(_24048_), .Q(_stream_conv2d_8_source_36_source_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38901_ ( .CLK(CLK), .D(_24047_), .Q(_stream_conv2d_8_source_36_source_ram_raddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_36_source_ram_renable_reg ( .CLK(CLK), .D(_24046_), .Q(_stream_conv2d_8_source_36_source_ram_renable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_source_36_source_ram_rvalid_reg ( .CLK(CLK), .D(_24044_), .Q(_stream_conv2d_8_source_36_source_ram_rvalid), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(3), .SRST_POLARITY(1'h1), .SRST_VALUE(3'h0) ) _38904_ ( .CLK(CLK), .D(_24043_), .Q(_stream_conv2d_8_sink_37_sink_mode), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38905_ ( .CLK(CLK), .D(_24042_), .Q(_stream_conv2d_8_sink_37_sink_offset), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38906_ ( .CLK(CLK), .D(_24041_), .Q(_stream_conv2d_8_sink_37_sink_size), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38907_ ( .CLK(CLK), .D(_24040_), .Q(_stream_conv2d_8_sink_37_sink_stride), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _38908_ ( .CLK(CLK), .D(_24039_), .Q(_stream_conv2d_8_sink_37_sink_count), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38909_ ( .CLK(CLK), .D(_24037_), .Q(_stream_conv2d_8_sink_37_sink_stride_buf), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38910_ ( .CLK(CLK), .D(_24036_), .Q(_stream_conv2d_8_sink_37_sink_ram_sel), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38911_ ( .CLK(CLK), .D(_24035_), .Q(_stream_conv2d_8_sink_37_sink_waddr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _stream_conv2d_8_sink_37_sink_wenable_reg ( .CLK(CLK), .D(_24033_), .Q(_stream_conv2d_8_sink_37_sink_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38913_ ( .CLK(CLK), .D(_24032_), .Q(_stream_conv2d_8_sink_37_sink_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _38914_ ( .CLK(CLK), .D(__variable_wdata_210), .Q(_cond_data_215), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38915_ ( .CLK(CLK), .D(__variable_wdata_217), .Q(_cond_data_222), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38916_ ( .CLK(CLK), .D(__variable_wdata_224), .Q(_cond_data_229), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38917_ ( .CLK(CLK), .D(__variable_wdata_231), .Q(_cond_data_236), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38918_ ( .CLK(CLK), .D(__variable_wdata_238), .Q(_cond_data_243), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _eq_data_337_reg ( .CLK(CLK), .D(_05224_), .Q(_eq_data_337), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _eq_data_341_reg ( .CLK(CLK), .D(_05225_), .Q(_eq_data_341), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _eq_data_344_reg ( .CLK(CLK), .D(_05226_), .Q(_eq_data_344), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _eq_data_427_reg ( .CLK(CLK), .D(_05227_), .Q(_eq_data_427), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _eq_data_431_reg ( .CLK(CLK), .D(_05228_), .Q(_eq_data_431), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _eq_data_434_reg ( .CLK(CLK), .D(_05229_), .Q(_eq_data_434), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pointer_data_536_reg ( .CLK(CLK), .D(__variable_wdata_197[0]), .Q(_pointer_data_536), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pointer_data_538_reg ( .CLK(CLK), .D(__variable_wdata_197[1]), .Q(_pointer_data_538), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pointer_data_540_reg ( .CLK(CLK), .D(__variable_wdata_197[2]), .Q(_pointer_data_540), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pointer_data_542_reg ( .CLK(CLK), .D(__variable_wdata_197[3]), .Q(_pointer_data_542), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pointer_data_544_reg ( .CLK(CLK), .D(__variable_wdata_197[4]), .Q(_pointer_data_544), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pointer_data_546_reg ( .CLK(CLK), .D(__variable_wdata_197[5]), .Q(_pointer_data_546), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pointer_data_548_reg ( .CLK(CLK), .D(__variable_wdata_197[6]), .Q(_pointer_data_548), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pointer_data_550_reg ( .CLK(CLK), .D(__variable_wdata_197[7]), .Q(_pointer_data_550), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pointer_data_552_reg ( .CLK(CLK), .D(__variable_wdata_197[8]), .Q(_pointer_data_552), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38934_ ( .CLK(CLK), .D(__variable_wdata_250), .Q(__delay_data_868), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38935_ ( .CLK(CLK), .D(__variable_wdata_249), .Q(__delay_data_870), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38936_ ( .CLK(CLK), .D(__variable_wdata_248), .Q(__delay_data_874), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38937_ ( .CLK(CLK), .D(__variable_wdata_253), .Q(__delay_data_877), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38938_ ( .CLK(CLK), .D(__variable_wdata_252), .Q(__delay_data_879), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38939_ ( .CLK(CLK), .D(__variable_wdata_251), .Q(__delay_data_883), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38940_ ( .CLK(CLK), .D(__variable_wdata_256), .Q(__delay_data_886), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38941_ ( .CLK(CLK), .D(__variable_wdata_255), .Q(__delay_data_888), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38942_ ( .CLK(CLK), .D(__variable_wdata_254), .Q(__delay_data_892), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_916_reg ( .CLK(CLK), .D(__variable_wdata_244), .Q(__delay_data_916), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38944_ ( .CLK(CLK), .D(__variable_wdata_482), .Q(__delay_data_917), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38945_ ( .CLK(CLK), .D(__variable_wdata_483), .Q(__delay_data_967), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38946_ ( .CLK(CLK), .D(__variable_wdata_484), .Q(__delay_data_1014), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38947_ ( .CLK(CLK), .D(__variable_wdata_485), .Q(__delay_data_1048), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38948_ ( .CLK(CLK), .D(__variable_wdata_486), .Q(__delay_data_1082), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38949_ ( .CLK(CLK), .D(__variable_wdata_487), .Q(__delay_data_1116), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38950_ ( .CLK(CLK), .D(__variable_wdata_488), .Q(__delay_data_1149), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38951_ ( .CLK(CLK), .D(__variable_wdata_489), .Q(__delay_data_1182), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38952_ ( .CLK(CLK), .D(__variable_wdata_490), .Q(__delay_data_1215), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1229_reg ( .CLK(CLK), .D(__variable_wdata_245), .Q(__delay_data_1229), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _38954_ ( .CLK(CLK), .D(__variable_wdata_194), .Q(__delay_data_1250), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _38955_ ( .CLK(CLK), .D(__variable_wdata_246), .Q(__delay_data_1300), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38956_ ( .CLK(CLK), .D(_26564_), .Q(_cond_data_259), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38957_ ( .CLK(CLK), .D(_26565_), .Q(_cond_data_269), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38958_ ( .CLK(CLK), .D(_26566_), .Q(_cond_data_279), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38959_ ( .CLK(CLK), .D(_26567_), .Q(_cond_data_289), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38960_ ( .CLK(CLK), .D(_26568_), .Q(_cond_data_299), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38961_ ( .CLK(CLK), .D(_26569_), .Q(_cond_data_309), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38962_ ( .CLK(CLK), .D(_26570_), .Q(_cond_data_319), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38963_ ( .CLK(CLK), .D(_26571_), .Q(_cond_data_329), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38964_ ( .CLK(CLK), .D(_26572_), .Q(_cond_data_339), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38965_ ( .CLK(CLK), .D(_22136_), .Q(_plus_data_723), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38966_ ( .CLK(CLK), .D(_22137_), .Q(_plus_data_739), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38967_ ( .CLK(CLK), .D(_22138_), .Q(_plus_data_750), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_869_reg ( .CLK(CLK), .D(_eq_data_341), .Q(__delay_data_869), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38969_ ( .CLK(CLK), .D(__delay_data_870), .Q(__delay_data_871), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38970_ ( .CLK(CLK), .D(__delay_data_874), .Q(__delay_data_875), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38971_ ( .CLK(CLK), .D(__delay_data_879), .Q(__delay_data_880), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38972_ ( .CLK(CLK), .D(__delay_data_883), .Q(__delay_data_884), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38973_ ( .CLK(CLK), .D(__delay_data_888), .Q(__delay_data_889), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38974_ ( .CLK(CLK), .D(__delay_data_892), .Q(__delay_data_893), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_910_reg ( .CLK(CLK), .D(_pointer_data_536), .Q(__delay_data_910), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38976_ ( .CLK(CLK), .D(__delay_data_917), .Q(__delay_data_918), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38977_ ( .CLK(CLK), .D(__delay_data_868), .Q(__delay_data_932), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38978_ ( .CLK(CLK), .D(__delay_data_877), .Q(__delay_data_937), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38979_ ( .CLK(CLK), .D(__delay_data_886), .Q(__delay_data_942), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_961_reg ( .CLK(CLK), .D(_pointer_data_538), .Q(__delay_data_961), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38981_ ( .CLK(CLK), .D(__delay_data_967), .Q(__delay_data_968), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_990_reg ( .CLK(CLK), .D(_eq_data_344), .Q(__delay_data_990), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1008_reg ( .CLK(CLK), .D(_pointer_data_540), .Q(__delay_data_1008), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38984_ ( .CLK(CLK), .D(__delay_data_1014), .Q(__delay_data_1015), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1042_reg ( .CLK(CLK), .D(_pointer_data_542), .Q(__delay_data_1042), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38986_ ( .CLK(CLK), .D(__delay_data_1048), .Q(__delay_data_1049), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1076_reg ( .CLK(CLK), .D(_pointer_data_544), .Q(__delay_data_1076), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38988_ ( .CLK(CLK), .D(__delay_data_1082), .Q(__delay_data_1083), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1110_reg ( .CLK(CLK), .D(_pointer_data_546), .Q(__delay_data_1110), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38990_ ( .CLK(CLK), .D(__delay_data_1116), .Q(__delay_data_1117), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1143_reg ( .CLK(CLK), .D(_pointer_data_548), .Q(__delay_data_1143), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38992_ ( .CLK(CLK), .D(__delay_data_1149), .Q(__delay_data_1150), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1176_reg ( .CLK(CLK), .D(_pointer_data_550), .Q(__delay_data_1176), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38994_ ( .CLK(CLK), .D(__delay_data_1182), .Q(__delay_data_1183), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1196_reg ( .CLK(CLK), .D(_eq_data_427), .Q(__delay_data_1196), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1199_reg ( .CLK(CLK), .D(_eq_data_431), .Q(__delay_data_1199), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1203_reg ( .CLK(CLK), .D(_eq_data_434), .Q(__delay_data_1203), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1209_reg ( .CLK(CLK), .D(_pointer_data_552), .Q(__delay_data_1209), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _38999_ ( .CLK(CLK), .D(__delay_data_1215), .Q(__delay_data_1216), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39000_ ( .CLK(CLK), .D(__delay_data_1250), .Q(__delay_data_1251), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39001_ ( .CLK(CLK), .D(_cond_data_215), .Q(__delay_data_1272), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39002_ ( .CLK(CLK), .D(_cond_data_222), .Q(__delay_data_1301), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39003_ ( .CLK(CLK), .D(_26573_), .Q(_cond_data_263), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39004_ ( .CLK(CLK), .D(_26574_), .Q(_cond_data_273), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39005_ ( .CLK(CLK), .D(_26575_), .Q(_cond_data_283), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39006_ ( .CLK(CLK), .D(_26576_), .Q(_cond_data_293), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39007_ ( .CLK(CLK), .D(_26577_), .Q(_cond_data_303), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39008_ ( .CLK(CLK), .D(_26578_), .Q(_cond_data_313), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39009_ ( .CLK(CLK), .D(_26579_), .Q(_cond_data_323), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39010_ ( .CLK(CLK), .D(_26580_), .Q(_cond_data_333), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39011_ ( .CLK(CLK), .D(_26581_), .Q(_cond_data_343), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39012_ ( .CLK(CLK), .D(__delay_data_875), .Q(__delay_data_876), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39013_ ( .CLK(CLK), .D(__delay_data_884), .Q(__delay_data_885), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39014_ ( .CLK(CLK), .D(__delay_data_893), .Q(__delay_data_894), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_911_reg ( .CLK(CLK), .D(__delay_data_910), .Q(__delay_data_911), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39016_ ( .CLK(CLK), .D(__delay_data_918), .Q(__delay_data_919), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39017_ ( .CLK(CLK), .D(__delay_data_871), .Q(__delay_data_935), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39018_ ( .CLK(CLK), .D(__delay_data_880), .Q(__delay_data_940), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39019_ ( .CLK(CLK), .D(__delay_data_889), .Q(__delay_data_945), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_962_reg ( .CLK(CLK), .D(__delay_data_961), .Q(__delay_data_962), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39021_ ( .CLK(CLK), .D(__delay_data_968), .Q(__delay_data_969), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39022_ ( .CLK(CLK), .D(__delay_data_932), .Q(__delay_data_984), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39023_ ( .CLK(CLK), .D(__delay_data_937), .Q(__delay_data_988), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_991_reg ( .CLK(CLK), .D(__delay_data_990), .Q(__delay_data_991), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39025_ ( .CLK(CLK), .D(__delay_data_942), .Q(__delay_data_992), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1009_reg ( .CLK(CLK), .D(__delay_data_1008), .Q(__delay_data_1009), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39027_ ( .CLK(CLK), .D(__delay_data_1015), .Q(__delay_data_1016), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1043_reg ( .CLK(CLK), .D(__delay_data_1042), .Q(__delay_data_1043), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39029_ ( .CLK(CLK), .D(__delay_data_1049), .Q(__delay_data_1050), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1077_reg ( .CLK(CLK), .D(__delay_data_1076), .Q(__delay_data_1077), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39031_ ( .CLK(CLK), .D(__delay_data_1083), .Q(__delay_data_1084), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1111_reg ( .CLK(CLK), .D(__delay_data_1110), .Q(__delay_data_1111), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39033_ ( .CLK(CLK), .D(__delay_data_1117), .Q(__delay_data_1118), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1144_reg ( .CLK(CLK), .D(__delay_data_1143), .Q(__delay_data_1144), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39035_ ( .CLK(CLK), .D(__delay_data_1150), .Q(__delay_data_1151), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1177_reg ( .CLK(CLK), .D(__delay_data_1176), .Q(__delay_data_1177), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39037_ ( .CLK(CLK), .D(__delay_data_1183), .Q(__delay_data_1184), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1197_reg ( .CLK(CLK), .D(__delay_data_1196), .Q(__delay_data_1197), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1200_reg ( .CLK(CLK), .D(__delay_data_1199), .Q(__delay_data_1200), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1204_reg ( .CLK(CLK), .D(__delay_data_1203), .Q(__delay_data_1204), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1210_reg ( .CLK(CLK), .D(__delay_data_1209), .Q(__delay_data_1210), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39042_ ( .CLK(CLK), .D(__delay_data_1216), .Q(__delay_data_1217), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39043_ ( .CLK(CLK), .D(_plus_data_723), .Q(__delay_data_1223), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39044_ ( .CLK(CLK), .D(_plus_data_739), .Q(__delay_data_1230), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39045_ ( .CLK(CLK), .D(__delay_data_1251), .Q(__delay_data_1252), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39046_ ( .CLK(CLK), .D(__delay_data_1272), .Q(__delay_data_1273), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39047_ ( .CLK(CLK), .D(__delay_data_1301), .Q(__delay_data_1302), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39048_ ( .CLK(CLK), .D(_plus_data_750), .Q(__delay_data_1330), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39049_ ( .CLK(CLK), .D(_26582_), .Q(_cond_data_266), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39050_ ( .CLK(CLK), .D(_26583_), .Q(_cond_data_276), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39051_ ( .CLK(CLK), .D(_26584_), .Q(_cond_data_286), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39052_ ( .CLK(CLK), .D(_26585_), .Q(_cond_data_296), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39053_ ( .CLK(CLK), .D(_26586_), .Q(_cond_data_306), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39054_ ( .CLK(CLK), .D(_26587_), .Q(_cond_data_316), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39055_ ( .CLK(CLK), .D(_26588_), .Q(_cond_data_326), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39056_ ( .CLK(CLK), .D(_26589_), .Q(_cond_data_336), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39057_ ( .CLK(CLK), .D(_26590_), .Q(_cond_data_346), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_912_reg ( .CLK(CLK), .D(__delay_data_911), .Q(__delay_data_912), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39059_ ( .CLK(CLK), .D(__delay_data_919), .Q(__delay_data_920), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_963_reg ( .CLK(CLK), .D(__delay_data_962), .Q(__delay_data_963), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39061_ ( .CLK(CLK), .D(__delay_data_969), .Q(__delay_data_970), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1010_reg ( .CLK(CLK), .D(__delay_data_1009), .Q(__delay_data_1010), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39063_ ( .CLK(CLK), .D(__delay_data_1016), .Q(__delay_data_1017), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1044_reg ( .CLK(CLK), .D(__delay_data_1043), .Q(__delay_data_1044), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39065_ ( .CLK(CLK), .D(__delay_data_1050), .Q(__delay_data_1051), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1078_reg ( .CLK(CLK), .D(__delay_data_1077), .Q(__delay_data_1078), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39067_ ( .CLK(CLK), .D(__delay_data_1084), .Q(__delay_data_1085), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1112_reg ( .CLK(CLK), .D(__delay_data_1111), .Q(__delay_data_1112), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39069_ ( .CLK(CLK), .D(__delay_data_1118), .Q(__delay_data_1119), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1145_reg ( .CLK(CLK), .D(__delay_data_1144), .Q(__delay_data_1145), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39071_ ( .CLK(CLK), .D(__delay_data_1151), .Q(__delay_data_1152), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1178_reg ( .CLK(CLK), .D(__delay_data_1177), .Q(__delay_data_1178), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39073_ ( .CLK(CLK), .D(__delay_data_1184), .Q(__delay_data_1185), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1198_reg ( .CLK(CLK), .D(__delay_data_1197), .Q(__delay_data_1198), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1201_reg ( .CLK(CLK), .D(__delay_data_1200), .Q(__delay_data_1201), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1205_reg ( .CLK(CLK), .D(__delay_data_1204), .Q(__delay_data_1205), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1211_reg ( .CLK(CLK), .D(__delay_data_1210), .Q(__delay_data_1211), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39078_ ( .CLK(CLK), .D(__delay_data_1217), .Q(__delay_data_1218), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39079_ ( .CLK(CLK), .D(__delay_data_1223), .Q(__delay_data_1224), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39080_ ( .CLK(CLK), .D(__delay_data_1230), .Q(__delay_data_1231), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39081_ ( .CLK(CLK), .D(__delay_data_1252), .Q(__delay_data_1253), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39082_ ( .CLK(CLK), .D(__delay_data_1273), .Q(__delay_data_1274), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39083_ ( .CLK(CLK), .D(__delay_data_1302), .Q(__delay_data_1303), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39084_ ( .CLK(CLK), .D(__delay_data_1330), .Q(__delay_data_1331), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39085_ ( .CLK(CLK), .D(_26591_), .Q(_cond_data_349), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39086_ ( .CLK(CLK), .D(_26592_), .Q(_cond_data_359), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39087_ ( .CLK(CLK), .D(_26593_), .Q(_cond_data_369), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39088_ ( .CLK(CLK), .D(_26594_), .Q(_cond_data_379), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39089_ ( .CLK(CLK), .D(_26595_), .Q(_cond_data_389), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39090_ ( .CLK(CLK), .D(_26596_), .Q(_cond_data_399), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39091_ ( .CLK(CLK), .D(_26597_), .Q(_cond_data_409), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39092_ ( .CLK(CLK), .D(_26598_), .Q(_cond_data_419), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39093_ ( .CLK(CLK), .D(_26599_), .Q(_cond_data_429), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39094_ ( .CLK(CLK), .D(_cond_data_296), .Q(__delay_data_902), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39095_ ( .CLK(CLK), .D(_cond_data_266), .Q(__delay_data_908), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_913_reg ( .CLK(CLK), .D(__delay_data_912), .Q(__delay_data_913), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39097_ ( .CLK(CLK), .D(__delay_data_920), .Q(__delay_data_921), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39098_ ( .CLK(CLK), .D(_cond_data_306), .Q(__delay_data_953), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39099_ ( .CLK(CLK), .D(_cond_data_276), .Q(__delay_data_959), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_964_reg ( .CLK(CLK), .D(__delay_data_963), .Q(__delay_data_964), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39101_ ( .CLK(CLK), .D(__delay_data_970), .Q(__delay_data_971), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39102_ ( .CLK(CLK), .D(_cond_data_316), .Q(__delay_data_1000), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39103_ ( .CLK(CLK), .D(_cond_data_286), .Q(__delay_data_1006), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1011_reg ( .CLK(CLK), .D(__delay_data_1010), .Q(__delay_data_1011), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39105_ ( .CLK(CLK), .D(__delay_data_1017), .Q(__delay_data_1018), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39106_ ( .CLK(CLK), .D(_cond_data_326), .Q(__delay_data_1035), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1045_reg ( .CLK(CLK), .D(__delay_data_1044), .Q(__delay_data_1045), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39108_ ( .CLK(CLK), .D(__delay_data_1051), .Q(__delay_data_1052), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39109_ ( .CLK(CLK), .D(_cond_data_336), .Q(__delay_data_1069), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1079_reg ( .CLK(CLK), .D(__delay_data_1078), .Q(__delay_data_1079), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39111_ ( .CLK(CLK), .D(__delay_data_1085), .Q(__delay_data_1086), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39112_ ( .CLK(CLK), .D(_cond_data_346), .Q(__delay_data_1103), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1113_reg ( .CLK(CLK), .D(__delay_data_1112), .Q(__delay_data_1113), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39114_ ( .CLK(CLK), .D(__delay_data_1119), .Q(__delay_data_1120), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1146_reg ( .CLK(CLK), .D(__delay_data_1145), .Q(__delay_data_1146), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39116_ ( .CLK(CLK), .D(__delay_data_1152), .Q(__delay_data_1153), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1179_reg ( .CLK(CLK), .D(__delay_data_1178), .Q(__delay_data_1179), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39118_ ( .CLK(CLK), .D(__delay_data_1185), .Q(__delay_data_1186), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1202_reg ( .CLK(CLK), .D(__delay_data_1201), .Q(__delay_data_1202), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1206_reg ( .CLK(CLK), .D(__delay_data_1205), .Q(__delay_data_1206), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1212_reg ( .CLK(CLK), .D(__delay_data_1211), .Q(__delay_data_1212), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39122_ ( .CLK(CLK), .D(__delay_data_1218), .Q(__delay_data_1219), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39123_ ( .CLK(CLK), .D(__delay_data_1224), .Q(__delay_data_1225), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39124_ ( .CLK(CLK), .D(__delay_data_1231), .Q(__delay_data_1232), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39125_ ( .CLK(CLK), .D(__delay_data_1253), .Q(__delay_data_1254), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39126_ ( .CLK(CLK), .D(__delay_data_1274), .Q(__delay_data_1275), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39127_ ( .CLK(CLK), .D(__delay_data_1303), .Q(__delay_data_1304), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39128_ ( .CLK(CLK), .D(__delay_data_1331), .Q(__delay_data_1332), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39129_ ( .CLK(CLK), .D(_26600_), .Q(_cond_data_353), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39130_ ( .CLK(CLK), .D(_26601_), .Q(_cond_data_363), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39131_ ( .CLK(CLK), .D(_26602_), .Q(_cond_data_373), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39132_ ( .CLK(CLK), .D(_26603_), .Q(_cond_data_383), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39133_ ( .CLK(CLK), .D(_26604_), .Q(_cond_data_393), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39134_ ( .CLK(CLK), .D(_26605_), .Q(_cond_data_403), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39135_ ( .CLK(CLK), .D(_26606_), .Q(_cond_data_413), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39136_ ( .CLK(CLK), .D(_26607_), .Q(_cond_data_423), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39137_ ( .CLK(CLK), .D(_26608_), .Q(_cond_data_433), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39138_ ( .CLK(CLK), .D(__delay_data_908), .Q(__delay_data_909), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_914_reg ( .CLK(CLK), .D(__delay_data_913), .Q(__delay_data_914), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39140_ ( .CLK(CLK), .D(__delay_data_921), .Q(__delay_data_922), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39141_ ( .CLK(CLK), .D(__delay_data_959), .Q(__delay_data_960), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_965_reg ( .CLK(CLK), .D(__delay_data_964), .Q(__delay_data_965), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39143_ ( .CLK(CLK), .D(__delay_data_971), .Q(__delay_data_972), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39144_ ( .CLK(CLK), .D(__delay_data_1006), .Q(__delay_data_1007), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1012_reg ( .CLK(CLK), .D(__delay_data_1011), .Q(__delay_data_1012), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39146_ ( .CLK(CLK), .D(__delay_data_1018), .Q(__delay_data_1019), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39147_ ( .CLK(CLK), .D(__delay_data_902), .Q(__delay_data_1041), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1046_reg ( .CLK(CLK), .D(__delay_data_1045), .Q(__delay_data_1046), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39149_ ( .CLK(CLK), .D(__delay_data_1052), .Q(__delay_data_1053), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39150_ ( .CLK(CLK), .D(__delay_data_953), .Q(__delay_data_1075), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1080_reg ( .CLK(CLK), .D(__delay_data_1079), .Q(__delay_data_1080), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39152_ ( .CLK(CLK), .D(__delay_data_1086), .Q(__delay_data_1087), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39153_ ( .CLK(CLK), .D(__delay_data_1000), .Q(__delay_data_1109), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1114_reg ( .CLK(CLK), .D(__delay_data_1113), .Q(__delay_data_1114), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39155_ ( .CLK(CLK), .D(__delay_data_1120), .Q(__delay_data_1121), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39156_ ( .CLK(CLK), .D(__delay_data_1035), .Q(__delay_data_1142), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1147_reg ( .CLK(CLK), .D(__delay_data_1146), .Q(__delay_data_1147), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39158_ ( .CLK(CLK), .D(__delay_data_1153), .Q(__delay_data_1154), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39159_ ( .CLK(CLK), .D(__delay_data_1069), .Q(__delay_data_1175), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1180_reg ( .CLK(CLK), .D(__delay_data_1179), .Q(__delay_data_1180), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39161_ ( .CLK(CLK), .D(__delay_data_1186), .Q(__delay_data_1187), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1207_reg ( .CLK(CLK), .D(__delay_data_1206), .Q(__delay_data_1207), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39163_ ( .CLK(CLK), .D(__delay_data_1103), .Q(__delay_data_1208), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1213_reg ( .CLK(CLK), .D(__delay_data_1212), .Q(__delay_data_1213), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39165_ ( .CLK(CLK), .D(__delay_data_1219), .Q(__delay_data_1220), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39166_ ( .CLK(CLK), .D(__delay_data_1225), .Q(__delay_data_1226), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39167_ ( .CLK(CLK), .D(__delay_data_1232), .Q(__delay_data_1233), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39168_ ( .CLK(CLK), .D(__delay_data_1254), .Q(__delay_data_1255), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39169_ ( .CLK(CLK), .D(__delay_data_1275), .Q(__delay_data_1276), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39170_ ( .CLK(CLK), .D(__delay_data_1304), .Q(__delay_data_1305), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39171_ ( .CLK(CLK), .D(__delay_data_1332), .Q(__delay_data_1333), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39172_ ( .CLK(CLK), .D(_26609_), .Q(_cond_data_356), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39173_ ( .CLK(CLK), .D(_26610_), .Q(_cond_data_366), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39174_ ( .CLK(CLK), .D(_26611_), .Q(_cond_data_376), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39175_ ( .CLK(CLK), .D(_26612_), .Q(_cond_data_386), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39176_ ( .CLK(CLK), .D(_26613_), .Q(_cond_data_396), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39177_ ( .CLK(CLK), .D(_26614_), .Q(_cond_data_406), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39178_ ( .CLK(CLK), .D(_26615_), .Q(_cond_data_416), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39179_ ( .CLK(CLK), .D(_26616_), .Q(_cond_data_426), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39180_ ( .CLK(CLK), .D(_26617_), .Q(_cond_data_436), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_915_reg ( .CLK(CLK), .D(__delay_data_914), .Q(__delay_data_915), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39182_ ( .CLK(CLK), .D(__delay_data_922), .Q(__delay_data_923), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_966_reg ( .CLK(CLK), .D(__delay_data_965), .Q(__delay_data_966), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39184_ ( .CLK(CLK), .D(__delay_data_972), .Q(__delay_data_973), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1013_reg ( .CLK(CLK), .D(__delay_data_1012), .Q(__delay_data_1013), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39186_ ( .CLK(CLK), .D(__delay_data_1019), .Q(__delay_data_1020), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1047_reg ( .CLK(CLK), .D(__delay_data_1046), .Q(__delay_data_1047), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39188_ ( .CLK(CLK), .D(__delay_data_1053), .Q(__delay_data_1054), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1081_reg ( .CLK(CLK), .D(__delay_data_1080), .Q(__delay_data_1081), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39190_ ( .CLK(CLK), .D(__delay_data_1087), .Q(__delay_data_1088), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1115_reg ( .CLK(CLK), .D(__delay_data_1114), .Q(__delay_data_1115), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39192_ ( .CLK(CLK), .D(__delay_data_1121), .Q(__delay_data_1122), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1148_reg ( .CLK(CLK), .D(__delay_data_1147), .Q(__delay_data_1148), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39194_ ( .CLK(CLK), .D(__delay_data_1154), .Q(__delay_data_1155), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1181_reg ( .CLK(CLK), .D(__delay_data_1180), .Q(__delay_data_1181), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39196_ ( .CLK(CLK), .D(__delay_data_1187), .Q(__delay_data_1188), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1214_reg ( .CLK(CLK), .D(__delay_data_1213), .Q(__delay_data_1214), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39198_ ( .CLK(CLK), .D(__delay_data_1220), .Q(__delay_data_1221), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39199_ ( .CLK(CLK), .D(__delay_data_1226), .Q(__delay_data_1227), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39200_ ( .CLK(CLK), .D(__delay_data_1233), .Q(__delay_data_1234), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39201_ ( .CLK(CLK), .D(__delay_data_1255), .Q(__delay_data_1256), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39202_ ( .CLK(CLK), .D(__delay_data_1276), .Q(__delay_data_1277), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39203_ ( .CLK(CLK), .D(__delay_data_1305), .Q(__delay_data_1306), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39204_ ( .CLK(CLK), .D(__delay_data_1333), .Q(__delay_data_1334), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39205_ ( .CLK(CLK), .D(_26618_), .Q(_cond_data_555), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39206_ ( .CLK(CLK), .D(_26619_), .Q(_cond_data_557), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39207_ ( .CLK(CLK), .D(_26620_), .Q(_cond_data_559), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39208_ ( .CLK(CLK), .D(_26621_), .Q(_cond_data_561), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39209_ ( .CLK(CLK), .D(_26622_), .Q(_cond_data_563), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39210_ ( .CLK(CLK), .D(_26623_), .Q(_cond_data_565), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39211_ ( .CLK(CLK), .D(_26624_), .Q(_cond_data_567), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39212_ ( .CLK(CLK), .D(_26625_), .Q(_cond_data_569), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39213_ ( .CLK(CLK), .D(_26626_), .Q(_cond_data_571), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39214_ ( .CLK(CLK), .D(__delay_data_923), .Q(__delay_data_924), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39215_ ( .CLK(CLK), .D(__delay_data_973), .Q(__delay_data_974), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39216_ ( .CLK(CLK), .D(__delay_data_1020), .Q(__delay_data_1021), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39217_ ( .CLK(CLK), .D(__delay_data_1054), .Q(__delay_data_1055), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39218_ ( .CLK(CLK), .D(__delay_data_1088), .Q(__delay_data_1089), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39219_ ( .CLK(CLK), .D(__delay_data_1122), .Q(__delay_data_1123), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39220_ ( .CLK(CLK), .D(__delay_data_1155), .Q(__delay_data_1156), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39221_ ( .CLK(CLK), .D(__delay_data_1188), .Q(__delay_data_1189), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39222_ ( .CLK(CLK), .D(__delay_data_1221), .Q(__delay_data_1222), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39223_ ( .CLK(CLK), .D(__delay_data_1227), .Q(__delay_data_1228), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39224_ ( .CLK(CLK), .D(__delay_data_1234), .Q(__delay_data_1235), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39225_ ( .CLK(CLK), .D(__delay_data_1256), .Q(__delay_data_1257), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39226_ ( .CLK(CLK), .D(__delay_data_1277), .Q(__delay_data_1278), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39227_ ( .CLK(CLK), .D(__delay_data_1306), .Q(__delay_data_1307), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39228_ ( .CLK(CLK), .D(__delay_data_1334), .Q(__delay_data_1335), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39229_ ( .CLK(CLK), .D(__delay_data_1235), .Q(__delay_data_1236), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39230_ ( .CLK(CLK), .D(__delay_data_1257), .Q(__delay_data_1258), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39231_ ( .CLK(CLK), .D(__delay_data_1278), .Q(__delay_data_1279), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39232_ ( .CLK(CLK), .D(__delay_data_1307), .Q(__delay_data_1308), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39233_ ( .CLK(CLK), .D(__delay_data_1335), .Q(__delay_data_1336), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39234_ ( .CLK(CLK), .D(__delay_data_1236), .Q(__delay_data_1237), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39235_ ( .CLK(CLK), .D(__delay_data_1258), .Q(__delay_data_1259), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39236_ ( .CLK(CLK), .D(__delay_data_1279), .Q(__delay_data_1280), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39237_ ( .CLK(CLK), .D(__delay_data_1308), .Q(__delay_data_1309), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39238_ ( .CLK(CLK), .D(__delay_data_1336), .Q(__delay_data_1337), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39239_ ( .CLK(CLK), .D(__delay_data_1237), .Q(__delay_data_1238), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39240_ ( .CLK(CLK), .D(__delay_data_1259), .Q(__delay_data_1260), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39241_ ( .CLK(CLK), .D(__delay_data_1280), .Q(__delay_data_1281), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39242_ ( .CLK(CLK), .D(__delay_data_1309), .Q(__delay_data_1310), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39243_ ( .CLK(CLK), .D(__delay_data_1337), .Q(__delay_data_1338), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39244_ ( .CLK(CLK), .D(__delay_data_1238), .Q(__delay_data_1239), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39245_ ( .CLK(CLK), .D(__delay_data_1260), .Q(__delay_data_1261), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39246_ ( .CLK(CLK), .D(__delay_data_1281), .Q(__delay_data_1282), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39247_ ( .CLK(CLK), .D(__delay_data_1310), .Q(__delay_data_1311), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39248_ ( .CLK(CLK), .D(__delay_data_1338), .Q(__delay_data_1339), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39249_ ( .CLK(CLK), .D(__delay_data_1239), .Q(__delay_data_1240), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39250_ ( .CLK(CLK), .D(__delay_data_1261), .Q(__delay_data_1262), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39251_ ( .CLK(CLK), .D(__delay_data_1282), .Q(__delay_data_1283), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39252_ ( .CLK(CLK), .D(__delay_data_1311), .Q(__delay_data_1312), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39253_ ( .CLK(CLK), .D(__delay_data_1339), .Q(__delay_data_1340), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39254_ ( .CLK(CLK), .D(__delay_data_1240), .Q(__delay_data_1241), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39255_ ( .CLK(CLK), .D(__delay_data_1262), .Q(__delay_data_1263), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39256_ ( .CLK(CLK), .D(__delay_data_1283), .Q(__delay_data_1284), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39257_ ( .CLK(CLK), .D(__delay_data_1312), .Q(__delay_data_1313), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39258_ ( .CLK(CLK), .D(__delay_data_1340), .Q(__delay_data_1341), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39259_ ( .CLK(CLK), .D(__delay_data_1241), .Q(__delay_data_1242), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39260_ ( .CLK(CLK), .D(__delay_data_1263), .Q(__delay_data_1264), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39261_ ( .CLK(CLK), .D(__delay_data_1284), .Q(__delay_data_1285), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39262_ ( .CLK(CLK), .D(__delay_data_1313), .Q(__delay_data_1314), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39263_ ( .CLK(CLK), .D(__delay_data_1341), .Q(__delay_data_1342), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39264_ ( .CLK(CLK), .D(__delay_data_1242), .Q(__delay_data_1243), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39265_ ( .CLK(CLK), .D(__delay_data_1264), .Q(__delay_data_1265), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39266_ ( .CLK(CLK), .D(__delay_data_1285), .Q(__delay_data_1286), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39267_ ( .CLK(CLK), .D(__delay_data_1314), .Q(__delay_data_1315), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39268_ ( .CLK(CLK), .D(__delay_data_1342), .Q(__delay_data_1343), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39269_ ( .CLK(CLK), .D(__delay_data_1243), .Q(__delay_data_1244), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39270_ ( .CLK(CLK), .D(__delay_data_1265), .Q(__delay_data_1266), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39271_ ( .CLK(CLK), .D(__delay_data_1286), .Q(__delay_data_1287), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39272_ ( .CLK(CLK), .D(__delay_data_1315), .Q(__delay_data_1316), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39273_ ( .CLK(CLK), .D(__delay_data_1343), .Q(__delay_data_1344), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _39274_ ( .CLK(CLK), .D(_sra_data_81), .Q(__substreamoutput_data_605), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _39275_ ( .CLK(CLK), .D(_sra_data_96), .Q(__substreamoutput_data_622), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _39276_ ( .CLK(CLK), .D(_sra_data_111), .Q(__substreamoutput_data_639), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _39277_ ( .CLK(CLK), .D(_sra_data_126), .Q(__substreamoutput_data_656), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _39278_ ( .CLK(CLK), .D(_sra_data_141), .Q(__substreamoutput_data_673), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _39279_ ( .CLK(CLK), .D(_sra_data_156), .Q(__substreamoutput_data_690), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _39280_ ( .CLK(CLK), .D(_sra_data_171), .Q(__substreamoutput_data_707), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _39281_ ( .CLK(CLK), .D(_sra_data_186), .Q(__substreamoutput_data_724), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39282_ ( .CLK(CLK), .D(__delay_data_1244), .Q(__delay_data_1245), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39283_ ( .CLK(CLK), .D(__delay_data_1266), .Q(__delay_data_1267), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39284_ ( .CLK(CLK), .D(__delay_data_1287), .Q(__delay_data_1288), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39285_ ( .CLK(CLK), .D(__delay_data_1316), .Q(__delay_data_1317), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39286_ ( .CLK(CLK), .D(__delay_data_1344), .Q(__delay_data_1345), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39287_ ( .CLK(CLK), .D(__delay_data_1245), .Q(__delay_data_1246), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39288_ ( .CLK(CLK), .D(__delay_data_1267), .Q(__delay_data_1268), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39289_ ( .CLK(CLK), .D(__delay_data_1288), .Q(__delay_data_1289), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39290_ ( .CLK(CLK), .D(__delay_data_1317), .Q(__delay_data_1318), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39291_ ( .CLK(CLK), .D(__delay_data_1345), .Q(__delay_data_1346), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39292_ ( .CLK(CLK), .D(__delay_data_1246), .Q(__delay_data_1247), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39293_ ( .CLK(CLK), .D(__delay_data_1268), .Q(__delay_data_1269), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39294_ ( .CLK(CLK), .D(__delay_data_1289), .Q(__delay_data_1290), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39295_ ( .CLK(CLK), .D(__delay_data_1318), .Q(__delay_data_1319), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39296_ ( .CLK(CLK), .D(__delay_data_1346), .Q(__delay_data_1347), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39297_ ( .CLK(CLK), .D(__delay_data_1247), .Q(__delay_data_1248), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39298_ ( .CLK(CLK), .D(__delay_data_1269), .Q(__delay_data_1270), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39299_ ( .CLK(CLK), .D(__delay_data_1290), .Q(__delay_data_1291), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39300_ ( .CLK(CLK), .D(__delay_data_1319), .Q(__delay_data_1320), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39301_ ( .CLK(CLK), .D(__delay_data_1347), .Q(__delay_data_1348), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39302_ ( .CLK(CLK), .D(__plusn_data_35), .Q(__substreamoutput_data_726), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39303_ ( .CLK(CLK), .D(__delay_data_1248), .Q(__delay_data_1249), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39304_ ( .CLK(CLK), .D(__delay_data_1270), .Q(__delay_data_1271), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39305_ ( .CLK(CLK), .D(__delay_data_1291), .Q(__delay_data_1292), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39306_ ( .CLK(CLK), .D(__delay_data_1320), .Q(__delay_data_1321), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39307_ ( .CLK(CLK), .D(__delay_data_1348), .Q(__delay_data_1349), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39308_ ( .CLK(CLK), .D(__delay_data_1292), .Q(__delay_data_1293), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39309_ ( .CLK(CLK), .D(__delay_data_1321), .Q(__delay_data_1322), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39310_ ( .CLK(CLK), .D(__delay_data_1349), .Q(__delay_data_1350), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39311_ ( .CLK(CLK), .D(__delay_data_1293), .Q(__delay_data_1294), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39312_ ( .CLK(CLK), .D(__delay_data_1322), .Q(__delay_data_1323), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39313_ ( .CLK(CLK), .D(__delay_data_1350), .Q(__delay_data_1351), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39314_ ( .CLK(CLK), .D(__delay_data_1294), .Q(__delay_data_1295), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39315_ ( .CLK(CLK), .D(__delay_data_1323), .Q(__delay_data_1324), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39316_ ( .CLK(CLK), .D(__delay_data_1351), .Q(__delay_data_1352), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39317_ ( .CLK(CLK), .D(__delay_data_1295), .Q(__delay_data_1296), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39318_ ( .CLK(CLK), .D(__delay_data_1324), .Q(__delay_data_1325), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39319_ ( .CLK(CLK), .D(__delay_data_1352), .Q(__delay_data_1353), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39320_ ( .CLK(CLK), .D(__delay_data_1296), .Q(__delay_data_1297), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39321_ ( .CLK(CLK), .D(__delay_data_1325), .Q(__delay_data_1326), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39322_ ( .CLK(CLK), .D(__delay_data_1353), .Q(__delay_data_1354), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39323_ ( .CLK(CLK), .D(__delay_data_1297), .Q(__delay_data_1298), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39324_ ( .CLK(CLK), .D(__delay_data_1326), .Q(__delay_data_1327), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39325_ ( .CLK(CLK), .D(__delay_data_1354), .Q(__delay_data_1355), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39326_ ( .CLK(CLK), .D(__delay_data_1298), .Q(__delay_data_1299), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39327_ ( .CLK(CLK), .D(__delay_data_1327), .Q(__delay_data_1328), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39328_ ( .CLK(CLK), .D(__delay_data_1355), .Q(__delay_data_1356), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39329_ ( .CLK(CLK), .D(_22139_), .Q(_plus_data_742), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39330_ ( .CLK(CLK), .D(__delay_data_1328), .Q(__delay_data_1329), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39331_ ( .CLK(CLK), .D(__delay_data_1356), .Q(__delay_data_1357), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greaterthan_data_753_reg ( .CLK(CLK), .D(_05261_), .Q(_greaterthan_data_753), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39333_ ( .CLK(CLK), .D(__substreamoutput_data_866), .Q(__delay_data_1358), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1370_reg ( .CLK(CLK), .D(__delay_data_1498), .Q(__delay_data_1370), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39335_ ( .CLK(CLK), .D(_26627_), .Q(_cond_data_755), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_1371_reg ( .CLK(CLK), .D(__delay_data_1370), .Q(__delay_data_1371), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(5), .SRST_POLARITY(1'h1), .SRST_VALUE(5'h00) ) _39337_ ( .CLK(CLK), .D(_24031_), .Q(__variable_wdata_194), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _39338_ ( .CLK(CLK), .D(_24030_), .Q(__variable_wdata_195), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _39339_ ( .CLK(CLK), .D(_24029_), .Q(__variable_wdata_196), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _39340_ ( .CLK(CLK), .D(_24028_), .Q(__variable_wdata_197), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39341_ ( .CLK(CLK), .D(_24027_), .Q(_source_stream_conv2d_8_source_6_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39342_ ( .CLK(CLK), .D(_24024_), .Q(_source_stream_conv2d_8_source_6_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39343_ ( .CLK(CLK), .D(_24021_), .Q(_source_stream_conv2d_8_source_6_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39344_ ( .CLK(CLK), .D(_24018_), .Q(_source_stream_conv2d_8_source_6_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39345_ ( .CLK(CLK), .D(_24015_), .Q(_source_stream_conv2d_8_source_6_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39346_ ( .CLK(CLK), .D(_24014_), .Q(_source_stream_conv2d_8_source_6_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39347_ ( .CLK(CLK), .D(_24013_), .Q(_source_stream_conv2d_8_source_6_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39348_ ( .CLK(CLK), .D(_24012_), .Q(_source_stream_conv2d_8_source_6_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39349_ ( .CLK(CLK), .D(_24011_), .Q(_source_stream_conv2d_8_source_6_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39350_ ( .CLK(CLK), .D(_24010_), .Q(_source_stream_conv2d_8_source_6_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39351_ ( .CLK(CLK), .D(_24009_), .Q(_source_stream_conv2d_8_source_6_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39352_ ( .CLK(CLK), .D(_24008_), .Q(_source_stream_conv2d_8_source_6_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39353_ ( .CLK(CLK), .D(_24007_), .Q(_source_stream_conv2d_8_source_6_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39354_ ( .CLK(CLK), .D(_24004_), .Q(_source_stream_conv2d_8_source_6_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39355_ ( .CLK(CLK), .D(_24001_), .Q(_source_stream_conv2d_8_source_6_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39356_ ( .CLK(CLK), .D(_23998_), .Q(_source_stream_conv2d_8_source_6_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39357_ ( .CLK(CLK), .D(_23995_), .Q(_source_stream_conv2d_8_source_6_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39358_ ( .CLK(CLK), .D(_23994_), .Q(_source_stream_conv2d_8_source_6_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39359_ ( .CLK(CLK), .D(_23993_), .Q(_source_stream_conv2d_8_source_6_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39360_ ( .CLK(CLK), .D(_23992_), .Q(_source_stream_conv2d_8_source_6_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39361_ ( .CLK(CLK), .D(_23991_), .Q(_source_stream_conv2d_8_source_6_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39362_ ( .CLK(CLK), .D(_23990_), .Q(_source_stream_conv2d_8_source_6_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39363_ ( .CLK(CLK), .D(_23989_), .Q(_source_stream_conv2d_8_source_6_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39364_ ( .CLK(CLK), .D(_23988_), .Q(_source_stream_conv2d_8_source_6_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39365_ ( .CLK(CLK), .D(_23987_), .Q(__variable_wdata_210), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39366_ ( .CLK(CLK), .D(_23986_), .Q(_source_stream_conv2d_8_source_8_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39367_ ( .CLK(CLK), .D(_23983_), .Q(_source_stream_conv2d_8_source_8_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39368_ ( .CLK(CLK), .D(_23980_), .Q(_source_stream_conv2d_8_source_8_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39369_ ( .CLK(CLK), .D(_23977_), .Q(_source_stream_conv2d_8_source_8_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39370_ ( .CLK(CLK), .D(_23974_), .Q(_source_stream_conv2d_8_source_8_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39371_ ( .CLK(CLK), .D(_23973_), .Q(_source_stream_conv2d_8_source_8_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39372_ ( .CLK(CLK), .D(_23972_), .Q(_source_stream_conv2d_8_source_8_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39373_ ( .CLK(CLK), .D(_23971_), .Q(_source_stream_conv2d_8_source_8_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39374_ ( .CLK(CLK), .D(_23970_), .Q(_source_stream_conv2d_8_source_8_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39375_ ( .CLK(CLK), .D(_23969_), .Q(_source_stream_conv2d_8_source_8_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39376_ ( .CLK(CLK), .D(_23968_), .Q(_source_stream_conv2d_8_source_8_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39377_ ( .CLK(CLK), .D(_23967_), .Q(_source_stream_conv2d_8_source_8_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39378_ ( .CLK(CLK), .D(_23966_), .Q(_source_stream_conv2d_8_source_8_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39379_ ( .CLK(CLK), .D(_23963_), .Q(_source_stream_conv2d_8_source_8_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39380_ ( .CLK(CLK), .D(_23960_), .Q(_source_stream_conv2d_8_source_8_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39381_ ( .CLK(CLK), .D(_23957_), .Q(_source_stream_conv2d_8_source_8_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39382_ ( .CLK(CLK), .D(_23954_), .Q(_source_stream_conv2d_8_source_8_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39383_ ( .CLK(CLK), .D(_23953_), .Q(_source_stream_conv2d_8_source_8_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39384_ ( .CLK(CLK), .D(_23952_), .Q(_source_stream_conv2d_8_source_8_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39385_ ( .CLK(CLK), .D(_23951_), .Q(_source_stream_conv2d_8_source_8_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39386_ ( .CLK(CLK), .D(_23950_), .Q(_source_stream_conv2d_8_source_8_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39387_ ( .CLK(CLK), .D(_23949_), .Q(_source_stream_conv2d_8_source_8_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39388_ ( .CLK(CLK), .D(_23948_), .Q(_source_stream_conv2d_8_source_8_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39389_ ( .CLK(CLK), .D(_23947_), .Q(_source_stream_conv2d_8_source_8_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39390_ ( .CLK(CLK), .D(_23946_), .Q(__variable_wdata_217), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39391_ ( .CLK(CLK), .D(_23945_), .Q(__variable_wdata_224), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39392_ ( .CLK(CLK), .D(_23944_), .Q(__variable_wdata_231), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39393_ ( .CLK(CLK), .D(_23943_), .Q(__variable_wdata_238), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __variable_wdata_244_reg ( .CLK(CLK), .D(_23942_), .Q(__variable_wdata_244), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __variable_wdata_245_reg ( .CLK(CLK), .D(_23941_), .Q(__variable_wdata_245), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _39396_ ( .CLK(CLK), .D(_23940_), .Q(__variable_wdata_246), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39397_ ( .CLK(CLK), .D(_23939_), .Q(_source_stream_conv2d_8_source_19_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39398_ ( .CLK(CLK), .D(_23936_), .Q(_source_stream_conv2d_8_source_19_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39399_ ( .CLK(CLK), .D(_23933_), .Q(_source_stream_conv2d_8_source_19_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39400_ ( .CLK(CLK), .D(_23930_), .Q(_source_stream_conv2d_8_source_19_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39401_ ( .CLK(CLK), .D(_23927_), .Q(_source_stream_conv2d_8_source_19_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39402_ ( .CLK(CLK), .D(_23926_), .Q(_source_stream_conv2d_8_source_19_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39403_ ( .CLK(CLK), .D(_23925_), .Q(_source_stream_conv2d_8_source_19_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39404_ ( .CLK(CLK), .D(_23924_), .Q(_source_stream_conv2d_8_source_19_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39405_ ( .CLK(CLK), .D(_23923_), .Q(_source_stream_conv2d_8_source_19_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39406_ ( .CLK(CLK), .D(_23922_), .Q(_source_stream_conv2d_8_source_19_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39407_ ( .CLK(CLK), .D(_23921_), .Q(_source_stream_conv2d_8_source_19_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39408_ ( .CLK(CLK), .D(_23920_), .Q(_source_stream_conv2d_8_source_19_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39409_ ( .CLK(CLK), .D(_23919_), .Q(_source_stream_conv2d_8_source_19_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39410_ ( .CLK(CLK), .D(_23916_), .Q(_source_stream_conv2d_8_source_19_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39411_ ( .CLK(CLK), .D(_23913_), .Q(_source_stream_conv2d_8_source_19_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39412_ ( .CLK(CLK), .D(_23910_), .Q(_source_stream_conv2d_8_source_19_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39413_ ( .CLK(CLK), .D(_23907_), .Q(_source_stream_conv2d_8_source_19_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39414_ ( .CLK(CLK), .D(_23906_), .Q(_source_stream_conv2d_8_source_19_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39415_ ( .CLK(CLK), .D(_23905_), .Q(_source_stream_conv2d_8_source_19_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39416_ ( .CLK(CLK), .D(_23904_), .Q(_source_stream_conv2d_8_source_19_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39417_ ( .CLK(CLK), .D(_23903_), .Q(_source_stream_conv2d_8_source_19_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39418_ ( .CLK(CLK), .D(_23902_), .Q(_source_stream_conv2d_8_source_19_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39419_ ( .CLK(CLK), .D(_23901_), .Q(_source_stream_conv2d_8_source_19_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39420_ ( .CLK(CLK), .D(_23900_), .Q(_source_stream_conv2d_8_source_19_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39421_ ( .CLK(CLK), .D(_23899_), .Q(__variable_wdata_248), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39422_ ( .CLK(CLK), .D(_23898_), .Q(_source_stream_conv2d_8_source_20_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39423_ ( .CLK(CLK), .D(_23895_), .Q(_source_stream_conv2d_8_source_20_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39424_ ( .CLK(CLK), .D(_23892_), .Q(_source_stream_conv2d_8_source_20_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39425_ ( .CLK(CLK), .D(_23889_), .Q(_source_stream_conv2d_8_source_20_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39426_ ( .CLK(CLK), .D(_23886_), .Q(_source_stream_conv2d_8_source_20_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39427_ ( .CLK(CLK), .D(_23885_), .Q(_source_stream_conv2d_8_source_20_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39428_ ( .CLK(CLK), .D(_23884_), .Q(_source_stream_conv2d_8_source_20_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39429_ ( .CLK(CLK), .D(_23883_), .Q(_source_stream_conv2d_8_source_20_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39430_ ( .CLK(CLK), .D(_23882_), .Q(_source_stream_conv2d_8_source_20_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39431_ ( .CLK(CLK), .D(_23881_), .Q(_source_stream_conv2d_8_source_20_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39432_ ( .CLK(CLK), .D(_23880_), .Q(_source_stream_conv2d_8_source_20_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39433_ ( .CLK(CLK), .D(_23879_), .Q(_source_stream_conv2d_8_source_20_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39434_ ( .CLK(CLK), .D(_23878_), .Q(_source_stream_conv2d_8_source_20_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39435_ ( .CLK(CLK), .D(_23875_), .Q(_source_stream_conv2d_8_source_20_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39436_ ( .CLK(CLK), .D(_23872_), .Q(_source_stream_conv2d_8_source_20_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39437_ ( .CLK(CLK), .D(_23869_), .Q(_source_stream_conv2d_8_source_20_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39438_ ( .CLK(CLK), .D(_23866_), .Q(_source_stream_conv2d_8_source_20_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39439_ ( .CLK(CLK), .D(_23865_), .Q(_source_stream_conv2d_8_source_20_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39440_ ( .CLK(CLK), .D(_23864_), .Q(_source_stream_conv2d_8_source_20_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39441_ ( .CLK(CLK), .D(_23863_), .Q(_source_stream_conv2d_8_source_20_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39442_ ( .CLK(CLK), .D(_23862_), .Q(_source_stream_conv2d_8_source_20_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39443_ ( .CLK(CLK), .D(_23861_), .Q(_source_stream_conv2d_8_source_20_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39444_ ( .CLK(CLK), .D(_23860_), .Q(_source_stream_conv2d_8_source_20_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39445_ ( .CLK(CLK), .D(_23859_), .Q(_source_stream_conv2d_8_source_20_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39446_ ( .CLK(CLK), .D(_23858_), .Q(__variable_wdata_249), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39447_ ( .CLK(CLK), .D(_23857_), .Q(_source_stream_conv2d_8_source_21_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39448_ ( .CLK(CLK), .D(_23854_), .Q(_source_stream_conv2d_8_source_21_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39449_ ( .CLK(CLK), .D(_23851_), .Q(_source_stream_conv2d_8_source_21_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39450_ ( .CLK(CLK), .D(_23848_), .Q(_source_stream_conv2d_8_source_21_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39451_ ( .CLK(CLK), .D(_23845_), .Q(_source_stream_conv2d_8_source_21_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39452_ ( .CLK(CLK), .D(_23844_), .Q(_source_stream_conv2d_8_source_21_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39453_ ( .CLK(CLK), .D(_23843_), .Q(_source_stream_conv2d_8_source_21_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39454_ ( .CLK(CLK), .D(_23842_), .Q(_source_stream_conv2d_8_source_21_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39455_ ( .CLK(CLK), .D(_23841_), .Q(_source_stream_conv2d_8_source_21_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39456_ ( .CLK(CLK), .D(_23840_), .Q(_source_stream_conv2d_8_source_21_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39457_ ( .CLK(CLK), .D(_23839_), .Q(_source_stream_conv2d_8_source_21_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39458_ ( .CLK(CLK), .D(_23838_), .Q(_source_stream_conv2d_8_source_21_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39459_ ( .CLK(CLK), .D(_23837_), .Q(_source_stream_conv2d_8_source_21_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39460_ ( .CLK(CLK), .D(_23834_), .Q(_source_stream_conv2d_8_source_21_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39461_ ( .CLK(CLK), .D(_23831_), .Q(_source_stream_conv2d_8_source_21_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39462_ ( .CLK(CLK), .D(_23828_), .Q(_source_stream_conv2d_8_source_21_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39463_ ( .CLK(CLK), .D(_23825_), .Q(_source_stream_conv2d_8_source_21_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39464_ ( .CLK(CLK), .D(_23824_), .Q(_source_stream_conv2d_8_source_21_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39465_ ( .CLK(CLK), .D(_23823_), .Q(_source_stream_conv2d_8_source_21_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39466_ ( .CLK(CLK), .D(_23822_), .Q(_source_stream_conv2d_8_source_21_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39467_ ( .CLK(CLK), .D(_23821_), .Q(_source_stream_conv2d_8_source_21_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39468_ ( .CLK(CLK), .D(_23820_), .Q(_source_stream_conv2d_8_source_21_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39469_ ( .CLK(CLK), .D(_23819_), .Q(_source_stream_conv2d_8_source_21_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39470_ ( .CLK(CLK), .D(_23818_), .Q(_source_stream_conv2d_8_source_21_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39471_ ( .CLK(CLK), .D(_23817_), .Q(__variable_wdata_250), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39472_ ( .CLK(CLK), .D(_23816_), .Q(_source_stream_conv2d_8_source_22_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39473_ ( .CLK(CLK), .D(_23813_), .Q(_source_stream_conv2d_8_source_22_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39474_ ( .CLK(CLK), .D(_23810_), .Q(_source_stream_conv2d_8_source_22_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39475_ ( .CLK(CLK), .D(_23807_), .Q(_source_stream_conv2d_8_source_22_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39476_ ( .CLK(CLK), .D(_23804_), .Q(_source_stream_conv2d_8_source_22_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39477_ ( .CLK(CLK), .D(_23803_), .Q(_source_stream_conv2d_8_source_22_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39478_ ( .CLK(CLK), .D(_23802_), .Q(_source_stream_conv2d_8_source_22_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39479_ ( .CLK(CLK), .D(_23801_), .Q(_source_stream_conv2d_8_source_22_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39480_ ( .CLK(CLK), .D(_23800_), .Q(_source_stream_conv2d_8_source_22_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39481_ ( .CLK(CLK), .D(_23799_), .Q(_source_stream_conv2d_8_source_22_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39482_ ( .CLK(CLK), .D(_23798_), .Q(_source_stream_conv2d_8_source_22_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39483_ ( .CLK(CLK), .D(_23797_), .Q(_source_stream_conv2d_8_source_22_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39484_ ( .CLK(CLK), .D(_23796_), .Q(_source_stream_conv2d_8_source_22_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39485_ ( .CLK(CLK), .D(_23793_), .Q(_source_stream_conv2d_8_source_22_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39486_ ( .CLK(CLK), .D(_23790_), .Q(_source_stream_conv2d_8_source_22_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39487_ ( .CLK(CLK), .D(_23787_), .Q(_source_stream_conv2d_8_source_22_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39488_ ( .CLK(CLK), .D(_23784_), .Q(_source_stream_conv2d_8_source_22_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39489_ ( .CLK(CLK), .D(_23783_), .Q(_source_stream_conv2d_8_source_22_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39490_ ( .CLK(CLK), .D(_23782_), .Q(_source_stream_conv2d_8_source_22_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39491_ ( .CLK(CLK), .D(_23781_), .Q(_source_stream_conv2d_8_source_22_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39492_ ( .CLK(CLK), .D(_23780_), .Q(_source_stream_conv2d_8_source_22_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39493_ ( .CLK(CLK), .D(_23779_), .Q(_source_stream_conv2d_8_source_22_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39494_ ( .CLK(CLK), .D(_23778_), .Q(_source_stream_conv2d_8_source_22_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39495_ ( .CLK(CLK), .D(_23777_), .Q(_source_stream_conv2d_8_source_22_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39496_ ( .CLK(CLK), .D(_23776_), .Q(__variable_wdata_251), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39497_ ( .CLK(CLK), .D(_23775_), .Q(_source_stream_conv2d_8_source_23_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39498_ ( .CLK(CLK), .D(_23772_), .Q(_source_stream_conv2d_8_source_23_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39499_ ( .CLK(CLK), .D(_23769_), .Q(_source_stream_conv2d_8_source_23_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39500_ ( .CLK(CLK), .D(_23766_), .Q(_source_stream_conv2d_8_source_23_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39501_ ( .CLK(CLK), .D(_23763_), .Q(_source_stream_conv2d_8_source_23_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39502_ ( .CLK(CLK), .D(_23762_), .Q(_source_stream_conv2d_8_source_23_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39503_ ( .CLK(CLK), .D(_23761_), .Q(_source_stream_conv2d_8_source_23_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39504_ ( .CLK(CLK), .D(_23760_), .Q(_source_stream_conv2d_8_source_23_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39505_ ( .CLK(CLK), .D(_23759_), .Q(_source_stream_conv2d_8_source_23_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39506_ ( .CLK(CLK), .D(_23758_), .Q(_source_stream_conv2d_8_source_23_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39507_ ( .CLK(CLK), .D(_23757_), .Q(_source_stream_conv2d_8_source_23_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39508_ ( .CLK(CLK), .D(_23756_), .Q(_source_stream_conv2d_8_source_23_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39509_ ( .CLK(CLK), .D(_23755_), .Q(_source_stream_conv2d_8_source_23_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39510_ ( .CLK(CLK), .D(_23752_), .Q(_source_stream_conv2d_8_source_23_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39511_ ( .CLK(CLK), .D(_23749_), .Q(_source_stream_conv2d_8_source_23_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39512_ ( .CLK(CLK), .D(_23746_), .Q(_source_stream_conv2d_8_source_23_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39513_ ( .CLK(CLK), .D(_23743_), .Q(_source_stream_conv2d_8_source_23_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39514_ ( .CLK(CLK), .D(_23742_), .Q(_source_stream_conv2d_8_source_23_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39515_ ( .CLK(CLK), .D(_23741_), .Q(_source_stream_conv2d_8_source_23_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39516_ ( .CLK(CLK), .D(_23740_), .Q(_source_stream_conv2d_8_source_23_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39517_ ( .CLK(CLK), .D(_23739_), .Q(_source_stream_conv2d_8_source_23_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39518_ ( .CLK(CLK), .D(_23738_), .Q(_source_stream_conv2d_8_source_23_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39519_ ( .CLK(CLK), .D(_23737_), .Q(_source_stream_conv2d_8_source_23_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39520_ ( .CLK(CLK), .D(_23736_), .Q(_source_stream_conv2d_8_source_23_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39521_ ( .CLK(CLK), .D(_23735_), .Q(__variable_wdata_252), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39522_ ( .CLK(CLK), .D(_23734_), .Q(_source_stream_conv2d_8_source_24_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39523_ ( .CLK(CLK), .D(_23731_), .Q(_source_stream_conv2d_8_source_24_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39524_ ( .CLK(CLK), .D(_23728_), .Q(_source_stream_conv2d_8_source_24_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39525_ ( .CLK(CLK), .D(_23725_), .Q(_source_stream_conv2d_8_source_24_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39526_ ( .CLK(CLK), .D(_23722_), .Q(_source_stream_conv2d_8_source_24_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39527_ ( .CLK(CLK), .D(_23721_), .Q(_source_stream_conv2d_8_source_24_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39528_ ( .CLK(CLK), .D(_23720_), .Q(_source_stream_conv2d_8_source_24_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39529_ ( .CLK(CLK), .D(_23719_), .Q(_source_stream_conv2d_8_source_24_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39530_ ( .CLK(CLK), .D(_23718_), .Q(_source_stream_conv2d_8_source_24_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39531_ ( .CLK(CLK), .D(_23717_), .Q(_source_stream_conv2d_8_source_24_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39532_ ( .CLK(CLK), .D(_23716_), .Q(_source_stream_conv2d_8_source_24_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39533_ ( .CLK(CLK), .D(_23715_), .Q(_source_stream_conv2d_8_source_24_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39534_ ( .CLK(CLK), .D(_23714_), .Q(_source_stream_conv2d_8_source_24_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39535_ ( .CLK(CLK), .D(_23711_), .Q(_source_stream_conv2d_8_source_24_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39536_ ( .CLK(CLK), .D(_23708_), .Q(_source_stream_conv2d_8_source_24_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39537_ ( .CLK(CLK), .D(_23705_), .Q(_source_stream_conv2d_8_source_24_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39538_ ( .CLK(CLK), .D(_23702_), .Q(_source_stream_conv2d_8_source_24_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39539_ ( .CLK(CLK), .D(_23701_), .Q(_source_stream_conv2d_8_source_24_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39540_ ( .CLK(CLK), .D(_23700_), .Q(_source_stream_conv2d_8_source_24_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39541_ ( .CLK(CLK), .D(_23699_), .Q(_source_stream_conv2d_8_source_24_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39542_ ( .CLK(CLK), .D(_23698_), .Q(_source_stream_conv2d_8_source_24_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39543_ ( .CLK(CLK), .D(_23697_), .Q(_source_stream_conv2d_8_source_24_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39544_ ( .CLK(CLK), .D(_23696_), .Q(_source_stream_conv2d_8_source_24_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39545_ ( .CLK(CLK), .D(_23695_), .Q(_source_stream_conv2d_8_source_24_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39546_ ( .CLK(CLK), .D(_23694_), .Q(__variable_wdata_253), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39547_ ( .CLK(CLK), .D(_23693_), .Q(_source_stream_conv2d_8_source_25_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39548_ ( .CLK(CLK), .D(_23690_), .Q(_source_stream_conv2d_8_source_25_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39549_ ( .CLK(CLK), .D(_23687_), .Q(_source_stream_conv2d_8_source_25_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39550_ ( .CLK(CLK), .D(_23684_), .Q(_source_stream_conv2d_8_source_25_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39551_ ( .CLK(CLK), .D(_23681_), .Q(_source_stream_conv2d_8_source_25_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39552_ ( .CLK(CLK), .D(_23680_), .Q(_source_stream_conv2d_8_source_25_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39553_ ( .CLK(CLK), .D(_23679_), .Q(_source_stream_conv2d_8_source_25_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39554_ ( .CLK(CLK), .D(_23678_), .Q(_source_stream_conv2d_8_source_25_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39555_ ( .CLK(CLK), .D(_23677_), .Q(_source_stream_conv2d_8_source_25_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39556_ ( .CLK(CLK), .D(_23676_), .Q(_source_stream_conv2d_8_source_25_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39557_ ( .CLK(CLK), .D(_23675_), .Q(_source_stream_conv2d_8_source_25_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39558_ ( .CLK(CLK), .D(_23674_), .Q(_source_stream_conv2d_8_source_25_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39559_ ( .CLK(CLK), .D(_23673_), .Q(_source_stream_conv2d_8_source_25_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39560_ ( .CLK(CLK), .D(_23670_), .Q(_source_stream_conv2d_8_source_25_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39561_ ( .CLK(CLK), .D(_23667_), .Q(_source_stream_conv2d_8_source_25_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39562_ ( .CLK(CLK), .D(_23664_), .Q(_source_stream_conv2d_8_source_25_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39563_ ( .CLK(CLK), .D(_23661_), .Q(_source_stream_conv2d_8_source_25_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39564_ ( .CLK(CLK), .D(_23660_), .Q(_source_stream_conv2d_8_source_25_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39565_ ( .CLK(CLK), .D(_23659_), .Q(_source_stream_conv2d_8_source_25_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39566_ ( .CLK(CLK), .D(_23658_), .Q(_source_stream_conv2d_8_source_25_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39567_ ( .CLK(CLK), .D(_23657_), .Q(_source_stream_conv2d_8_source_25_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39568_ ( .CLK(CLK), .D(_23656_), .Q(_source_stream_conv2d_8_source_25_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39569_ ( .CLK(CLK), .D(_23655_), .Q(_source_stream_conv2d_8_source_25_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39570_ ( .CLK(CLK), .D(_23654_), .Q(_source_stream_conv2d_8_source_25_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39571_ ( .CLK(CLK), .D(_23653_), .Q(__variable_wdata_254), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39572_ ( .CLK(CLK), .D(_23652_), .Q(_source_stream_conv2d_8_source_26_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39573_ ( .CLK(CLK), .D(_23649_), .Q(_source_stream_conv2d_8_source_26_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39574_ ( .CLK(CLK), .D(_23646_), .Q(_source_stream_conv2d_8_source_26_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39575_ ( .CLK(CLK), .D(_23643_), .Q(_source_stream_conv2d_8_source_26_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39576_ ( .CLK(CLK), .D(_23640_), .Q(_source_stream_conv2d_8_source_26_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39577_ ( .CLK(CLK), .D(_23639_), .Q(_source_stream_conv2d_8_source_26_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39578_ ( .CLK(CLK), .D(_23638_), .Q(_source_stream_conv2d_8_source_26_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39579_ ( .CLK(CLK), .D(_23637_), .Q(_source_stream_conv2d_8_source_26_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39580_ ( .CLK(CLK), .D(_23636_), .Q(_source_stream_conv2d_8_source_26_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39581_ ( .CLK(CLK), .D(_23635_), .Q(_source_stream_conv2d_8_source_26_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39582_ ( .CLK(CLK), .D(_23634_), .Q(_source_stream_conv2d_8_source_26_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39583_ ( .CLK(CLK), .D(_23633_), .Q(_source_stream_conv2d_8_source_26_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39584_ ( .CLK(CLK), .D(_23632_), .Q(_source_stream_conv2d_8_source_26_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39585_ ( .CLK(CLK), .D(_23629_), .Q(_source_stream_conv2d_8_source_26_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39586_ ( .CLK(CLK), .D(_23626_), .Q(_source_stream_conv2d_8_source_26_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39587_ ( .CLK(CLK), .D(_23623_), .Q(_source_stream_conv2d_8_source_26_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39588_ ( .CLK(CLK), .D(_23620_), .Q(_source_stream_conv2d_8_source_26_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39589_ ( .CLK(CLK), .D(_23619_), .Q(_source_stream_conv2d_8_source_26_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39590_ ( .CLK(CLK), .D(_23618_), .Q(_source_stream_conv2d_8_source_26_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39591_ ( .CLK(CLK), .D(_23617_), .Q(_source_stream_conv2d_8_source_26_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39592_ ( .CLK(CLK), .D(_23616_), .Q(_source_stream_conv2d_8_source_26_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39593_ ( .CLK(CLK), .D(_23615_), .Q(_source_stream_conv2d_8_source_26_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39594_ ( .CLK(CLK), .D(_23614_), .Q(_source_stream_conv2d_8_source_26_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39595_ ( .CLK(CLK), .D(_23613_), .Q(_source_stream_conv2d_8_source_26_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39596_ ( .CLK(CLK), .D(_23612_), .Q(__variable_wdata_255), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39597_ ( .CLK(CLK), .D(_23611_), .Q(_source_stream_conv2d_8_source_27_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39598_ ( .CLK(CLK), .D(_23608_), .Q(_source_stream_conv2d_8_source_27_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39599_ ( .CLK(CLK), .D(_23605_), .Q(_source_stream_conv2d_8_source_27_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39600_ ( .CLK(CLK), .D(_23602_), .Q(_source_stream_conv2d_8_source_27_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39601_ ( .CLK(CLK), .D(_23599_), .Q(_source_stream_conv2d_8_source_27_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39602_ ( .CLK(CLK), .D(_23598_), .Q(_source_stream_conv2d_8_source_27_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39603_ ( .CLK(CLK), .D(_23597_), .Q(_source_stream_conv2d_8_source_27_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39604_ ( .CLK(CLK), .D(_23596_), .Q(_source_stream_conv2d_8_source_27_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39605_ ( .CLK(CLK), .D(_23595_), .Q(_source_stream_conv2d_8_source_27_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39606_ ( .CLK(CLK), .D(_23594_), .Q(_source_stream_conv2d_8_source_27_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39607_ ( .CLK(CLK), .D(_23593_), .Q(_source_stream_conv2d_8_source_27_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39608_ ( .CLK(CLK), .D(_23592_), .Q(_source_stream_conv2d_8_source_27_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39609_ ( .CLK(CLK), .D(_23591_), .Q(_source_stream_conv2d_8_source_27_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39610_ ( .CLK(CLK), .D(_23588_), .Q(_source_stream_conv2d_8_source_27_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39611_ ( .CLK(CLK), .D(_23585_), .Q(_source_stream_conv2d_8_source_27_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39612_ ( .CLK(CLK), .D(_23582_), .Q(_source_stream_conv2d_8_source_27_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39613_ ( .CLK(CLK), .D(_23579_), .Q(_source_stream_conv2d_8_source_27_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39614_ ( .CLK(CLK), .D(_23578_), .Q(_source_stream_conv2d_8_source_27_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39615_ ( .CLK(CLK), .D(_23577_), .Q(_source_stream_conv2d_8_source_27_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39616_ ( .CLK(CLK), .D(_23576_), .Q(_source_stream_conv2d_8_source_27_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39617_ ( .CLK(CLK), .D(_23575_), .Q(_source_stream_conv2d_8_source_27_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39618_ ( .CLK(CLK), .D(_23574_), .Q(_source_stream_conv2d_8_source_27_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39619_ ( .CLK(CLK), .D(_23573_), .Q(_source_stream_conv2d_8_source_27_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39620_ ( .CLK(CLK), .D(_23572_), .Q(_source_stream_conv2d_8_source_27_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39621_ ( .CLK(CLK), .D(_23571_), .Q(__variable_wdata_256), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39622_ ( .CLK(CLK), .D(_23570_), .Q(_source_stream_conv2d_8_source_28_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39623_ ( .CLK(CLK), .D(_23567_), .Q(_source_stream_conv2d_8_source_28_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39624_ ( .CLK(CLK), .D(_23564_), .Q(_source_stream_conv2d_8_source_28_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39625_ ( .CLK(CLK), .D(_23561_), .Q(_source_stream_conv2d_8_source_28_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39626_ ( .CLK(CLK), .D(_23558_), .Q(_source_stream_conv2d_8_source_28_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39627_ ( .CLK(CLK), .D(_23557_), .Q(_source_stream_conv2d_8_source_28_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39628_ ( .CLK(CLK), .D(_23556_), .Q(_source_stream_conv2d_8_source_28_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39629_ ( .CLK(CLK), .D(_23555_), .Q(_source_stream_conv2d_8_source_28_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39630_ ( .CLK(CLK), .D(_23554_), .Q(_source_stream_conv2d_8_source_28_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39631_ ( .CLK(CLK), .D(_23553_), .Q(_source_stream_conv2d_8_source_28_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39632_ ( .CLK(CLK), .D(_23552_), .Q(_source_stream_conv2d_8_source_28_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39633_ ( .CLK(CLK), .D(_23551_), .Q(_source_stream_conv2d_8_source_28_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39634_ ( .CLK(CLK), .D(_23550_), .Q(_source_stream_conv2d_8_source_28_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39635_ ( .CLK(CLK), .D(_23547_), .Q(_source_stream_conv2d_8_source_28_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39636_ ( .CLK(CLK), .D(_23544_), .Q(_source_stream_conv2d_8_source_28_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39637_ ( .CLK(CLK), .D(_23541_), .Q(_source_stream_conv2d_8_source_28_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39638_ ( .CLK(CLK), .D(_23538_), .Q(_source_stream_conv2d_8_source_28_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39639_ ( .CLK(CLK), .D(_23537_), .Q(_source_stream_conv2d_8_source_28_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39640_ ( .CLK(CLK), .D(_23536_), .Q(_source_stream_conv2d_8_source_28_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39641_ ( .CLK(CLK), .D(_23535_), .Q(_source_stream_conv2d_8_source_28_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39642_ ( .CLK(CLK), .D(_23534_), .Q(_source_stream_conv2d_8_source_28_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39643_ ( .CLK(CLK), .D(_23533_), .Q(_source_stream_conv2d_8_source_28_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39644_ ( .CLK(CLK), .D(_23532_), .Q(_source_stream_conv2d_8_source_28_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39645_ ( .CLK(CLK), .D(_23531_), .Q(_source_stream_conv2d_8_source_28_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39646_ ( .CLK(CLK), .D(_23530_), .Q(__variable_wdata_482), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39647_ ( .CLK(CLK), .D(_23529_), .Q(_source_stream_conv2d_8_source_29_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39648_ ( .CLK(CLK), .D(_23526_), .Q(_source_stream_conv2d_8_source_29_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39649_ ( .CLK(CLK), .D(_23523_), .Q(_source_stream_conv2d_8_source_29_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39650_ ( .CLK(CLK), .D(_23520_), .Q(_source_stream_conv2d_8_source_29_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39651_ ( .CLK(CLK), .D(_23517_), .Q(_source_stream_conv2d_8_source_29_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39652_ ( .CLK(CLK), .D(_23516_), .Q(_source_stream_conv2d_8_source_29_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39653_ ( .CLK(CLK), .D(_23515_), .Q(_source_stream_conv2d_8_source_29_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39654_ ( .CLK(CLK), .D(_23514_), .Q(_source_stream_conv2d_8_source_29_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39655_ ( .CLK(CLK), .D(_23513_), .Q(_source_stream_conv2d_8_source_29_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39656_ ( .CLK(CLK), .D(_23512_), .Q(_source_stream_conv2d_8_source_29_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39657_ ( .CLK(CLK), .D(_23511_), .Q(_source_stream_conv2d_8_source_29_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39658_ ( .CLK(CLK), .D(_23510_), .Q(_source_stream_conv2d_8_source_29_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39659_ ( .CLK(CLK), .D(_23509_), .Q(_source_stream_conv2d_8_source_29_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39660_ ( .CLK(CLK), .D(_23506_), .Q(_source_stream_conv2d_8_source_29_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39661_ ( .CLK(CLK), .D(_23503_), .Q(_source_stream_conv2d_8_source_29_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39662_ ( .CLK(CLK), .D(_23500_), .Q(_source_stream_conv2d_8_source_29_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39663_ ( .CLK(CLK), .D(_23497_), .Q(_source_stream_conv2d_8_source_29_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39664_ ( .CLK(CLK), .D(_23496_), .Q(_source_stream_conv2d_8_source_29_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39665_ ( .CLK(CLK), .D(_23495_), .Q(_source_stream_conv2d_8_source_29_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39666_ ( .CLK(CLK), .D(_23494_), .Q(_source_stream_conv2d_8_source_29_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39667_ ( .CLK(CLK), .D(_23493_), .Q(_source_stream_conv2d_8_source_29_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39668_ ( .CLK(CLK), .D(_23492_), .Q(_source_stream_conv2d_8_source_29_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39669_ ( .CLK(CLK), .D(_23491_), .Q(_source_stream_conv2d_8_source_29_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39670_ ( .CLK(CLK), .D(_23490_), .Q(_source_stream_conv2d_8_source_29_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39671_ ( .CLK(CLK), .D(_23489_), .Q(__variable_wdata_483), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39672_ ( .CLK(CLK), .D(_23488_), .Q(_source_stream_conv2d_8_source_30_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39673_ ( .CLK(CLK), .D(_23485_), .Q(_source_stream_conv2d_8_source_30_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39674_ ( .CLK(CLK), .D(_23482_), .Q(_source_stream_conv2d_8_source_30_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39675_ ( .CLK(CLK), .D(_23479_), .Q(_source_stream_conv2d_8_source_30_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39676_ ( .CLK(CLK), .D(_23476_), .Q(_source_stream_conv2d_8_source_30_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39677_ ( .CLK(CLK), .D(_23475_), .Q(_source_stream_conv2d_8_source_30_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39678_ ( .CLK(CLK), .D(_23474_), .Q(_source_stream_conv2d_8_source_30_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39679_ ( .CLK(CLK), .D(_23473_), .Q(_source_stream_conv2d_8_source_30_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39680_ ( .CLK(CLK), .D(_23472_), .Q(_source_stream_conv2d_8_source_30_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39681_ ( .CLK(CLK), .D(_23471_), .Q(_source_stream_conv2d_8_source_30_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39682_ ( .CLK(CLK), .D(_23470_), .Q(_source_stream_conv2d_8_source_30_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39683_ ( .CLK(CLK), .D(_23469_), .Q(_source_stream_conv2d_8_source_30_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39684_ ( .CLK(CLK), .D(_23468_), .Q(_source_stream_conv2d_8_source_30_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39685_ ( .CLK(CLK), .D(_23465_), .Q(_source_stream_conv2d_8_source_30_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39686_ ( .CLK(CLK), .D(_23462_), .Q(_source_stream_conv2d_8_source_30_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39687_ ( .CLK(CLK), .D(_23459_), .Q(_source_stream_conv2d_8_source_30_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39688_ ( .CLK(CLK), .D(_23456_), .Q(_source_stream_conv2d_8_source_30_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39689_ ( .CLK(CLK), .D(_23455_), .Q(_source_stream_conv2d_8_source_30_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39690_ ( .CLK(CLK), .D(_23454_), .Q(_source_stream_conv2d_8_source_30_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39691_ ( .CLK(CLK), .D(_23453_), .Q(_source_stream_conv2d_8_source_30_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39692_ ( .CLK(CLK), .D(_23452_), .Q(_source_stream_conv2d_8_source_30_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39693_ ( .CLK(CLK), .D(_23451_), .Q(_source_stream_conv2d_8_source_30_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39694_ ( .CLK(CLK), .D(_23450_), .Q(_source_stream_conv2d_8_source_30_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39695_ ( .CLK(CLK), .D(_23449_), .Q(_source_stream_conv2d_8_source_30_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39696_ ( .CLK(CLK), .D(_23448_), .Q(__variable_wdata_484), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39697_ ( .CLK(CLK), .D(_23447_), .Q(_source_stream_conv2d_8_source_31_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39698_ ( .CLK(CLK), .D(_23444_), .Q(_source_stream_conv2d_8_source_31_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39699_ ( .CLK(CLK), .D(_23441_), .Q(_source_stream_conv2d_8_source_31_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39700_ ( .CLK(CLK), .D(_23438_), .Q(_source_stream_conv2d_8_source_31_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39701_ ( .CLK(CLK), .D(_23435_), .Q(_source_stream_conv2d_8_source_31_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39702_ ( .CLK(CLK), .D(_23434_), .Q(_source_stream_conv2d_8_source_31_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39703_ ( .CLK(CLK), .D(_23433_), .Q(_source_stream_conv2d_8_source_31_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39704_ ( .CLK(CLK), .D(_23432_), .Q(_source_stream_conv2d_8_source_31_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39705_ ( .CLK(CLK), .D(_23431_), .Q(_source_stream_conv2d_8_source_31_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39706_ ( .CLK(CLK), .D(_23430_), .Q(_source_stream_conv2d_8_source_31_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39707_ ( .CLK(CLK), .D(_23429_), .Q(_source_stream_conv2d_8_source_31_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39708_ ( .CLK(CLK), .D(_23428_), .Q(_source_stream_conv2d_8_source_31_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39709_ ( .CLK(CLK), .D(_23427_), .Q(_source_stream_conv2d_8_source_31_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39710_ ( .CLK(CLK), .D(_23424_), .Q(_source_stream_conv2d_8_source_31_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39711_ ( .CLK(CLK), .D(_23421_), .Q(_source_stream_conv2d_8_source_31_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39712_ ( .CLK(CLK), .D(_23418_), .Q(_source_stream_conv2d_8_source_31_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39713_ ( .CLK(CLK), .D(_23415_), .Q(_source_stream_conv2d_8_source_31_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39714_ ( .CLK(CLK), .D(_23414_), .Q(_source_stream_conv2d_8_source_31_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39715_ ( .CLK(CLK), .D(_23413_), .Q(_source_stream_conv2d_8_source_31_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39716_ ( .CLK(CLK), .D(_23412_), .Q(_source_stream_conv2d_8_source_31_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39717_ ( .CLK(CLK), .D(_23411_), .Q(_source_stream_conv2d_8_source_31_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39718_ ( .CLK(CLK), .D(_23410_), .Q(_source_stream_conv2d_8_source_31_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39719_ ( .CLK(CLK), .D(_23409_), .Q(_source_stream_conv2d_8_source_31_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39720_ ( .CLK(CLK), .D(_23408_), .Q(_source_stream_conv2d_8_source_31_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39721_ ( .CLK(CLK), .D(_23407_), .Q(__variable_wdata_485), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39722_ ( .CLK(CLK), .D(_23406_), .Q(_source_stream_conv2d_8_source_32_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39723_ ( .CLK(CLK), .D(_23403_), .Q(_source_stream_conv2d_8_source_32_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39724_ ( .CLK(CLK), .D(_23400_), .Q(_source_stream_conv2d_8_source_32_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39725_ ( .CLK(CLK), .D(_23397_), .Q(_source_stream_conv2d_8_source_32_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39726_ ( .CLK(CLK), .D(_23394_), .Q(_source_stream_conv2d_8_source_32_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39727_ ( .CLK(CLK), .D(_23393_), .Q(_source_stream_conv2d_8_source_32_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39728_ ( .CLK(CLK), .D(_23392_), .Q(_source_stream_conv2d_8_source_32_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39729_ ( .CLK(CLK), .D(_23391_), .Q(_source_stream_conv2d_8_source_32_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39730_ ( .CLK(CLK), .D(_23390_), .Q(_source_stream_conv2d_8_source_32_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39731_ ( .CLK(CLK), .D(_23389_), .Q(_source_stream_conv2d_8_source_32_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39732_ ( .CLK(CLK), .D(_23388_), .Q(_source_stream_conv2d_8_source_32_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39733_ ( .CLK(CLK), .D(_23387_), .Q(_source_stream_conv2d_8_source_32_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39734_ ( .CLK(CLK), .D(_23386_), .Q(_source_stream_conv2d_8_source_32_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39735_ ( .CLK(CLK), .D(_23383_), .Q(_source_stream_conv2d_8_source_32_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39736_ ( .CLK(CLK), .D(_23380_), .Q(_source_stream_conv2d_8_source_32_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39737_ ( .CLK(CLK), .D(_23377_), .Q(_source_stream_conv2d_8_source_32_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39738_ ( .CLK(CLK), .D(_23374_), .Q(_source_stream_conv2d_8_source_32_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39739_ ( .CLK(CLK), .D(_23373_), .Q(_source_stream_conv2d_8_source_32_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39740_ ( .CLK(CLK), .D(_23372_), .Q(_source_stream_conv2d_8_source_32_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39741_ ( .CLK(CLK), .D(_23371_), .Q(_source_stream_conv2d_8_source_32_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39742_ ( .CLK(CLK), .D(_23370_), .Q(_source_stream_conv2d_8_source_32_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39743_ ( .CLK(CLK), .D(_23369_), .Q(_source_stream_conv2d_8_source_32_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39744_ ( .CLK(CLK), .D(_23368_), .Q(_source_stream_conv2d_8_source_32_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39745_ ( .CLK(CLK), .D(_23367_), .Q(_source_stream_conv2d_8_source_32_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39746_ ( .CLK(CLK), .D(_23366_), .Q(__variable_wdata_486), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39747_ ( .CLK(CLK), .D(_23365_), .Q(_source_stream_conv2d_8_source_33_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39748_ ( .CLK(CLK), .D(_23362_), .Q(_source_stream_conv2d_8_source_33_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39749_ ( .CLK(CLK), .D(_23359_), .Q(_source_stream_conv2d_8_source_33_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39750_ ( .CLK(CLK), .D(_23356_), .Q(_source_stream_conv2d_8_source_33_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39751_ ( .CLK(CLK), .D(_23353_), .Q(_source_stream_conv2d_8_source_33_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39752_ ( .CLK(CLK), .D(_23352_), .Q(_source_stream_conv2d_8_source_33_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39753_ ( .CLK(CLK), .D(_23351_), .Q(_source_stream_conv2d_8_source_33_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39754_ ( .CLK(CLK), .D(_23350_), .Q(_source_stream_conv2d_8_source_33_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39755_ ( .CLK(CLK), .D(_23349_), .Q(_source_stream_conv2d_8_source_33_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39756_ ( .CLK(CLK), .D(_23348_), .Q(_source_stream_conv2d_8_source_33_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39757_ ( .CLK(CLK), .D(_23347_), .Q(_source_stream_conv2d_8_source_33_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39758_ ( .CLK(CLK), .D(_23346_), .Q(_source_stream_conv2d_8_source_33_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39759_ ( .CLK(CLK), .D(_23345_), .Q(_source_stream_conv2d_8_source_33_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39760_ ( .CLK(CLK), .D(_23342_), .Q(_source_stream_conv2d_8_source_33_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39761_ ( .CLK(CLK), .D(_23339_), .Q(_source_stream_conv2d_8_source_33_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39762_ ( .CLK(CLK), .D(_23336_), .Q(_source_stream_conv2d_8_source_33_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39763_ ( .CLK(CLK), .D(_23333_), .Q(_source_stream_conv2d_8_source_33_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39764_ ( .CLK(CLK), .D(_23332_), .Q(_source_stream_conv2d_8_source_33_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39765_ ( .CLK(CLK), .D(_23331_), .Q(_source_stream_conv2d_8_source_33_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39766_ ( .CLK(CLK), .D(_23330_), .Q(_source_stream_conv2d_8_source_33_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39767_ ( .CLK(CLK), .D(_23329_), .Q(_source_stream_conv2d_8_source_33_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39768_ ( .CLK(CLK), .D(_23328_), .Q(_source_stream_conv2d_8_source_33_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39769_ ( .CLK(CLK), .D(_23327_), .Q(_source_stream_conv2d_8_source_33_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39770_ ( .CLK(CLK), .D(_23326_), .Q(_source_stream_conv2d_8_source_33_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39771_ ( .CLK(CLK), .D(_23325_), .Q(__variable_wdata_487), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39772_ ( .CLK(CLK), .D(_23324_), .Q(_source_stream_conv2d_8_source_34_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39773_ ( .CLK(CLK), .D(_23321_), .Q(_source_stream_conv2d_8_source_34_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39774_ ( .CLK(CLK), .D(_23318_), .Q(_source_stream_conv2d_8_source_34_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39775_ ( .CLK(CLK), .D(_23315_), .Q(_source_stream_conv2d_8_source_34_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39776_ ( .CLK(CLK), .D(_23312_), .Q(_source_stream_conv2d_8_source_34_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39777_ ( .CLK(CLK), .D(_23311_), .Q(_source_stream_conv2d_8_source_34_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39778_ ( .CLK(CLK), .D(_23310_), .Q(_source_stream_conv2d_8_source_34_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39779_ ( .CLK(CLK), .D(_23309_), .Q(_source_stream_conv2d_8_source_34_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39780_ ( .CLK(CLK), .D(_23308_), .Q(_source_stream_conv2d_8_source_34_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39781_ ( .CLK(CLK), .D(_23307_), .Q(_source_stream_conv2d_8_source_34_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39782_ ( .CLK(CLK), .D(_23306_), .Q(_source_stream_conv2d_8_source_34_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39783_ ( .CLK(CLK), .D(_23305_), .Q(_source_stream_conv2d_8_source_34_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39784_ ( .CLK(CLK), .D(_23304_), .Q(_source_stream_conv2d_8_source_34_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39785_ ( .CLK(CLK), .D(_23301_), .Q(_source_stream_conv2d_8_source_34_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39786_ ( .CLK(CLK), .D(_23298_), .Q(_source_stream_conv2d_8_source_34_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39787_ ( .CLK(CLK), .D(_23295_), .Q(_source_stream_conv2d_8_source_34_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39788_ ( .CLK(CLK), .D(_23292_), .Q(_source_stream_conv2d_8_source_34_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39789_ ( .CLK(CLK), .D(_23291_), .Q(_source_stream_conv2d_8_source_34_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39790_ ( .CLK(CLK), .D(_23290_), .Q(_source_stream_conv2d_8_source_34_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39791_ ( .CLK(CLK), .D(_23289_), .Q(_source_stream_conv2d_8_source_34_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39792_ ( .CLK(CLK), .D(_23288_), .Q(_source_stream_conv2d_8_source_34_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39793_ ( .CLK(CLK), .D(_23287_), .Q(_source_stream_conv2d_8_source_34_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39794_ ( .CLK(CLK), .D(_23286_), .Q(_source_stream_conv2d_8_source_34_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39795_ ( .CLK(CLK), .D(_23285_), .Q(_source_stream_conv2d_8_source_34_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39796_ ( .CLK(CLK), .D(_23284_), .Q(__variable_wdata_488), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39797_ ( .CLK(CLK), .D(_23283_), .Q(_source_stream_conv2d_8_source_35_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39798_ ( .CLK(CLK), .D(_23280_), .Q(_source_stream_conv2d_8_source_35_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39799_ ( .CLK(CLK), .D(_23277_), .Q(_source_stream_conv2d_8_source_35_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39800_ ( .CLK(CLK), .D(_23274_), .Q(_source_stream_conv2d_8_source_35_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39801_ ( .CLK(CLK), .D(_23271_), .Q(_source_stream_conv2d_8_source_35_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39802_ ( .CLK(CLK), .D(_23270_), .Q(_source_stream_conv2d_8_source_35_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39803_ ( .CLK(CLK), .D(_23269_), .Q(_source_stream_conv2d_8_source_35_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39804_ ( .CLK(CLK), .D(_23268_), .Q(_source_stream_conv2d_8_source_35_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39805_ ( .CLK(CLK), .D(_23267_), .Q(_source_stream_conv2d_8_source_35_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39806_ ( .CLK(CLK), .D(_23266_), .Q(_source_stream_conv2d_8_source_35_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39807_ ( .CLK(CLK), .D(_23265_), .Q(_source_stream_conv2d_8_source_35_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39808_ ( .CLK(CLK), .D(_23264_), .Q(_source_stream_conv2d_8_source_35_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39809_ ( .CLK(CLK), .D(_23263_), .Q(_source_stream_conv2d_8_source_35_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39810_ ( .CLK(CLK), .D(_23260_), .Q(_source_stream_conv2d_8_source_35_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39811_ ( .CLK(CLK), .D(_23257_), .Q(_source_stream_conv2d_8_source_35_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39812_ ( .CLK(CLK), .D(_23254_), .Q(_source_stream_conv2d_8_source_35_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39813_ ( .CLK(CLK), .D(_23251_), .Q(_source_stream_conv2d_8_source_35_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39814_ ( .CLK(CLK), .D(_23250_), .Q(_source_stream_conv2d_8_source_35_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39815_ ( .CLK(CLK), .D(_23249_), .Q(_source_stream_conv2d_8_source_35_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39816_ ( .CLK(CLK), .D(_23248_), .Q(_source_stream_conv2d_8_source_35_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39817_ ( .CLK(CLK), .D(_23247_), .Q(_source_stream_conv2d_8_source_35_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39818_ ( .CLK(CLK), .D(_23246_), .Q(_source_stream_conv2d_8_source_35_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39819_ ( .CLK(CLK), .D(_23245_), .Q(_source_stream_conv2d_8_source_35_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39820_ ( .CLK(CLK), .D(_23244_), .Q(_source_stream_conv2d_8_source_35_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39821_ ( .CLK(CLK), .D(_23243_), .Q(__variable_wdata_489), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39822_ ( .CLK(CLK), .D(_23242_), .Q(_source_stream_conv2d_8_source_36_pat_cur_offset_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39823_ ( .CLK(CLK), .D(_23239_), .Q(_source_stream_conv2d_8_source_36_pat_cur_offset_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39824_ ( .CLK(CLK), .D(_23236_), .Q(_source_stream_conv2d_8_source_36_pat_cur_offset_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39825_ ( .CLK(CLK), .D(_23233_), .Q(_source_stream_conv2d_8_source_36_pat_cur_offset_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39826_ ( .CLK(CLK), .D(_23230_), .Q(_source_stream_conv2d_8_source_36_pat_size_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39827_ ( .CLK(CLK), .D(_23229_), .Q(_source_stream_conv2d_8_source_36_pat_size_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39828_ ( .CLK(CLK), .D(_23228_), .Q(_source_stream_conv2d_8_source_36_pat_size_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39829_ ( .CLK(CLK), .D(_23227_), .Q(_source_stream_conv2d_8_source_36_pat_size_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39830_ ( .CLK(CLK), .D(_23226_), .Q(_source_stream_conv2d_8_source_36_pat_stride_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39831_ ( .CLK(CLK), .D(_23225_), .Q(_source_stream_conv2d_8_source_36_pat_stride_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39832_ ( .CLK(CLK), .D(_23224_), .Q(_source_stream_conv2d_8_source_36_pat_stride_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39833_ ( .CLK(CLK), .D(_23223_), .Q(_source_stream_conv2d_8_source_36_pat_stride_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39834_ ( .CLK(CLK), .D(_23222_), .Q(_source_stream_conv2d_8_source_36_pat_count_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39835_ ( .CLK(CLK), .D(_23219_), .Q(_source_stream_conv2d_8_source_36_pat_count_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39836_ ( .CLK(CLK), .D(_23216_), .Q(_source_stream_conv2d_8_source_36_pat_count_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39837_ ( .CLK(CLK), .D(_23213_), .Q(_source_stream_conv2d_8_source_36_pat_count_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39838_ ( .CLK(CLK), .D(_23210_), .Q(_source_stream_conv2d_8_source_36_pat_size_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39839_ ( .CLK(CLK), .D(_23209_), .Q(_source_stream_conv2d_8_source_36_pat_size_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39840_ ( .CLK(CLK), .D(_23208_), .Q(_source_stream_conv2d_8_source_36_pat_size_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39841_ ( .CLK(CLK), .D(_23207_), .Q(_source_stream_conv2d_8_source_36_pat_size_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39842_ ( .CLK(CLK), .D(_23206_), .Q(_source_stream_conv2d_8_source_36_pat_stride_buf_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39843_ ( .CLK(CLK), .D(_23205_), .Q(_source_stream_conv2d_8_source_36_pat_stride_buf_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39844_ ( .CLK(CLK), .D(_23204_), .Q(_source_stream_conv2d_8_source_36_pat_stride_buf_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39845_ ( .CLK(CLK), .D(_23203_), .Q(_source_stream_conv2d_8_source_36_pat_stride_buf_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _39846_ ( .CLK(CLK), .D(_23202_), .Q(__variable_wdata_490), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _set_flag_538_reg ( .CLK(CLK), .D(_23201_), .Q(_set_flag_538), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39848_ ( .CLK(CLK), .D(_22229_), .Q(__stream_conv2d_8_sink_37_sink_offset_0_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39849_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_1), .Q(__stream_conv2d_8_sink_37_sink_offset_0_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39850_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_2), .Q(__stream_conv2d_8_sink_37_sink_offset_0_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39851_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_3), .Q(__stream_conv2d_8_sink_37_sink_offset_0_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39852_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_4), .Q(__stream_conv2d_8_sink_37_sink_offset_0_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39853_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_5), .Q(__stream_conv2d_8_sink_37_sink_offset_0_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39854_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_6), .Q(__stream_conv2d_8_sink_37_sink_offset_0_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39855_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_7), .Q(__stream_conv2d_8_sink_37_sink_offset_0_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39856_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_8), .Q(__stream_conv2d_8_sink_37_sink_offset_0_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39857_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_9), .Q(__stream_conv2d_8_sink_37_sink_offset_0_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39858_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_10), .Q(__stream_conv2d_8_sink_37_sink_offset_0_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39859_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_11), .Q(__stream_conv2d_8_sink_37_sink_offset_0_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39860_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_12), .Q(__stream_conv2d_8_sink_37_sink_offset_0_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39861_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_13), .Q(__stream_conv2d_8_sink_37_sink_offset_0_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39862_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_14), .Q(__stream_conv2d_8_sink_37_sink_offset_0_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39863_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_15), .Q(__stream_conv2d_8_sink_37_sink_offset_0_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39864_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_16), .Q(__stream_conv2d_8_sink_37_sink_offset_0_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39865_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_17), .Q(__stream_conv2d_8_sink_37_sink_offset_0_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39866_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_18), .Q(__stream_conv2d_8_sink_37_sink_offset_0_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39867_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_19), .Q(__stream_conv2d_8_sink_37_sink_offset_0_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39868_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_20), .Q(__stream_conv2d_8_sink_37_sink_offset_0_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39869_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_21), .Q(__stream_conv2d_8_sink_37_sink_offset_0_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39870_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_22), .Q(__stream_conv2d_8_sink_37_sink_offset_0_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39871_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_23), .Q(__stream_conv2d_8_sink_37_sink_offset_0_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39872_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_24), .Q(__stream_conv2d_8_sink_37_sink_offset_0_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39873_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_25), .Q(__stream_conv2d_8_sink_37_sink_offset_0_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39874_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_26), .Q(__stream_conv2d_8_sink_37_sink_offset_0_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39875_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_27), .Q(__stream_conv2d_8_sink_37_sink_offset_0_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39876_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_28), .Q(__stream_conv2d_8_sink_37_sink_offset_0_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39877_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_29), .Q(__stream_conv2d_8_sink_37_sink_offset_0_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39878_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_30), .Q(__stream_conv2d_8_sink_37_sink_offset_0_31), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39879_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_31), .Q(__stream_conv2d_8_sink_37_sink_offset_0_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39880_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_32), .Q(__stream_conv2d_8_sink_37_sink_offset_0_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39881_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_33), .Q(__stream_conv2d_8_sink_37_sink_offset_0_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39882_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_34), .Q(__stream_conv2d_8_sink_37_sink_offset_0_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39883_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_35), .Q(__stream_conv2d_8_sink_37_sink_offset_0_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39884_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_36), .Q(__stream_conv2d_8_sink_37_sink_offset_0_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39885_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_37), .Q(__stream_conv2d_8_sink_37_sink_offset_0_38), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39886_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_38), .Q(__stream_conv2d_8_sink_37_sink_offset_0_39), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39887_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_39), .Q(__stream_conv2d_8_sink_37_sink_offset_0_40), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39888_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_40), .Q(__stream_conv2d_8_sink_37_sink_offset_0_41), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39889_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_41), .Q(__stream_conv2d_8_sink_37_sink_offset_0_42), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39890_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_42), .Q(__stream_conv2d_8_sink_37_sink_offset_0_43), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39891_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_43), .Q(__stream_conv2d_8_sink_37_sink_offset_0_44), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _39892_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_offset_0_44), .Q(__stream_conv2d_8_sink_37_sink_offset_0_45), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39893_ ( .CLK(CLK), .D({ 1'h0, conv2d_8_next_stream_num_ops }), .Q(__stream_conv2d_8_sink_37_sink_size_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39894_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_1), .Q(__stream_conv2d_8_sink_37_sink_size_1_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39895_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_2), .Q(__stream_conv2d_8_sink_37_sink_size_1_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39896_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_3), .Q(__stream_conv2d_8_sink_37_sink_size_1_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39897_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_4), .Q(__stream_conv2d_8_sink_37_sink_size_1_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39898_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_5), .Q(__stream_conv2d_8_sink_37_sink_size_1_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39899_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_6), .Q(__stream_conv2d_8_sink_37_sink_size_1_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39900_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_7), .Q(__stream_conv2d_8_sink_37_sink_size_1_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39901_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_8), .Q(__stream_conv2d_8_sink_37_sink_size_1_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39902_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_9), .Q(__stream_conv2d_8_sink_37_sink_size_1_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39903_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_10), .Q(__stream_conv2d_8_sink_37_sink_size_1_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39904_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_11), .Q(__stream_conv2d_8_sink_37_sink_size_1_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39905_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_12), .Q(__stream_conv2d_8_sink_37_sink_size_1_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39906_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_13), .Q(__stream_conv2d_8_sink_37_sink_size_1_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39907_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_14), .Q(__stream_conv2d_8_sink_37_sink_size_1_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39908_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_15), .Q(__stream_conv2d_8_sink_37_sink_size_1_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39909_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_16), .Q(__stream_conv2d_8_sink_37_sink_size_1_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39910_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_17), .Q(__stream_conv2d_8_sink_37_sink_size_1_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39911_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_18), .Q(__stream_conv2d_8_sink_37_sink_size_1_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39912_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_19), .Q(__stream_conv2d_8_sink_37_sink_size_1_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39913_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_20), .Q(__stream_conv2d_8_sink_37_sink_size_1_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39914_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_21), .Q(__stream_conv2d_8_sink_37_sink_size_1_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39915_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_22), .Q(__stream_conv2d_8_sink_37_sink_size_1_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39916_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_23), .Q(__stream_conv2d_8_sink_37_sink_size_1_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39917_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_24), .Q(__stream_conv2d_8_sink_37_sink_size_1_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39918_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_25), .Q(__stream_conv2d_8_sink_37_sink_size_1_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39919_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_26), .Q(__stream_conv2d_8_sink_37_sink_size_1_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39920_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_27), .Q(__stream_conv2d_8_sink_37_sink_size_1_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39921_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_28), .Q(__stream_conv2d_8_sink_37_sink_size_1_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39922_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_29), .Q(__stream_conv2d_8_sink_37_sink_size_1_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39923_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_30), .Q(__stream_conv2d_8_sink_37_sink_size_1_31), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39924_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_31), .Q(__stream_conv2d_8_sink_37_sink_size_1_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39925_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_32), .Q(__stream_conv2d_8_sink_37_sink_size_1_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39926_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_33), .Q(__stream_conv2d_8_sink_37_sink_size_1_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39927_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_34), .Q(__stream_conv2d_8_sink_37_sink_size_1_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39928_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_35), .Q(__stream_conv2d_8_sink_37_sink_size_1_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39929_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_36), .Q(__stream_conv2d_8_sink_37_sink_size_1_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39930_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_37), .Q(__stream_conv2d_8_sink_37_sink_size_1_38), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39931_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_38), .Q(__stream_conv2d_8_sink_37_sink_size_1_39), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39932_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_39), .Q(__stream_conv2d_8_sink_37_sink_size_1_40), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39933_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_40), .Q(__stream_conv2d_8_sink_37_sink_size_1_41), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39934_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_41), .Q(__stream_conv2d_8_sink_37_sink_size_1_42), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39935_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_42), .Q(__stream_conv2d_8_sink_37_sink_size_1_43), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39936_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_43), .Q(__stream_conv2d_8_sink_37_sink_size_1_44), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _39937_ ( .CLK(CLK), .D(__stream_conv2d_8_sink_37_sink_size_1_44), .Q(__stream_conv2d_8_sink_37_sink_size_1_45), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_1_reg ( .CLK(CLK), .D(_set_flag_538), .Q(__set_flag_538_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_2_reg ( .CLK(CLK), .D(__set_flag_538_1), .Q(__set_flag_538_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_3_reg ( .CLK(CLK), .D(__set_flag_538_2), .Q(__set_flag_538_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_4_reg ( .CLK(CLK), .D(__set_flag_538_3), .Q(__set_flag_538_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_5_reg ( .CLK(CLK), .D(__set_flag_538_4), .Q(__set_flag_538_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_6_reg ( .CLK(CLK), .D(__set_flag_538_5), .Q(__set_flag_538_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_7_reg ( .CLK(CLK), .D(__set_flag_538_6), .Q(__set_flag_538_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_8_reg ( .CLK(CLK), .D(__set_flag_538_7), .Q(__set_flag_538_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_9_reg ( .CLK(CLK), .D(__set_flag_538_8), .Q(__set_flag_538_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_10_reg ( .CLK(CLK), .D(__set_flag_538_9), .Q(__set_flag_538_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_11_reg ( .CLK(CLK), .D(__set_flag_538_10), .Q(__set_flag_538_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_12_reg ( .CLK(CLK), .D(__set_flag_538_11), .Q(__set_flag_538_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_13_reg ( .CLK(CLK), .D(__set_flag_538_12), .Q(__set_flag_538_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_14_reg ( .CLK(CLK), .D(__set_flag_538_13), .Q(__set_flag_538_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_15_reg ( .CLK(CLK), .D(__set_flag_538_14), .Q(__set_flag_538_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_16_reg ( .CLK(CLK), .D(__set_flag_538_15), .Q(__set_flag_538_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_17_reg ( .CLK(CLK), .D(__set_flag_538_16), .Q(__set_flag_538_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_18_reg ( .CLK(CLK), .D(__set_flag_538_17), .Q(__set_flag_538_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_19_reg ( .CLK(CLK), .D(__set_flag_538_18), .Q(__set_flag_538_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_20_reg ( .CLK(CLK), .D(__set_flag_538_19), .Q(__set_flag_538_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_21_reg ( .CLK(CLK), .D(__set_flag_538_20), .Q(__set_flag_538_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_22_reg ( .CLK(CLK), .D(__set_flag_538_21), .Q(__set_flag_538_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_23_reg ( .CLK(CLK), .D(__set_flag_538_22), .Q(__set_flag_538_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_24_reg ( .CLK(CLK), .D(__set_flag_538_23), .Q(__set_flag_538_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_25_reg ( .CLK(CLK), .D(__set_flag_538_24), .Q(__set_flag_538_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_26_reg ( .CLK(CLK), .D(__set_flag_538_25), .Q(__set_flag_538_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_27_reg ( .CLK(CLK), .D(__set_flag_538_26), .Q(__set_flag_538_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_28_reg ( .CLK(CLK), .D(__set_flag_538_27), .Q(__set_flag_538_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_29_reg ( .CLK(CLK), .D(__set_flag_538_28), .Q(__set_flag_538_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_30_reg ( .CLK(CLK), .D(__set_flag_538_29), .Q(__set_flag_538_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_31_reg ( .CLK(CLK), .D(__set_flag_538_30), .Q(__set_flag_538_31), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_32_reg ( .CLK(CLK), .D(__set_flag_538_31), .Q(__set_flag_538_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_33_reg ( .CLK(CLK), .D(__set_flag_538_32), .Q(__set_flag_538_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_34_reg ( .CLK(CLK), .D(__set_flag_538_33), .Q(__set_flag_538_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_35_reg ( .CLK(CLK), .D(__set_flag_538_34), .Q(__set_flag_538_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_36_reg ( .CLK(CLK), .D(__set_flag_538_35), .Q(__set_flag_538_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_37_reg ( .CLK(CLK), .D(__set_flag_538_36), .Q(__set_flag_538_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_38_reg ( .CLK(CLK), .D(__set_flag_538_37), .Q(__set_flag_538_38), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_39_reg ( .CLK(CLK), .D(__set_flag_538_38), .Q(__set_flag_538_39), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_40_reg ( .CLK(CLK), .D(__set_flag_538_39), .Q(__set_flag_538_40), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_41_reg ( .CLK(CLK), .D(__set_flag_538_40), .Q(__set_flag_538_41), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_42_reg ( .CLK(CLK), .D(__set_flag_538_41), .Q(__set_flag_538_42), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_43_reg ( .CLK(CLK), .D(__set_flag_538_42), .Q(__set_flag_538_43), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_44_reg ( .CLK(CLK), .D(__set_flag_538_43), .Q(__set_flag_538_44), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __set_flag_538_45_reg ( .CLK(CLK), .D(__set_flag_538_44), .Q(__set_flag_538_45), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_1_reg ( .CLK(CLK), .D(_stream_conv2d_8_start), .Q(__stream_conv2d_8_start_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_2_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_1), .Q(__stream_conv2d_8_start_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_3_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_2), .Q(__stream_conv2d_8_start_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_4_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_3), .Q(__stream_conv2d_8_start_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_5_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_4), .Q(__stream_conv2d_8_start_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_6_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_5), .Q(__stream_conv2d_8_start_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_7_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_6), .Q(__stream_conv2d_8_start_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_8_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_7), .Q(__stream_conv2d_8_start_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_9_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_8), .Q(__stream_conv2d_8_start_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_10_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_9), .Q(__stream_conv2d_8_start_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_11_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_10), .Q(__stream_conv2d_8_start_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_12_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_11), .Q(__stream_conv2d_8_start_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_13_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_12), .Q(__stream_conv2d_8_start_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_14_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_13), .Q(__stream_conv2d_8_start_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_15_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_14), .Q(__stream_conv2d_8_start_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_16_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_15), .Q(__stream_conv2d_8_start_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_17_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_16), .Q(__stream_conv2d_8_start_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_18_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_17), .Q(__stream_conv2d_8_start_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_19_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_18), .Q(__stream_conv2d_8_start_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_20_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_19), .Q(__stream_conv2d_8_start_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_21_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_20), .Q(__stream_conv2d_8_start_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_22_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_21), .Q(__stream_conv2d_8_start_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_23_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_22), .Q(__stream_conv2d_8_start_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_24_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_23), .Q(__stream_conv2d_8_start_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_25_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_24), .Q(__stream_conv2d_8_start_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_26_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_25), .Q(__stream_conv2d_8_start_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_27_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_26), .Q(__stream_conv2d_8_start_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_28_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_27), .Q(__stream_conv2d_8_start_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_29_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_28), .Q(__stream_conv2d_8_start_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_30_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_29), .Q(__stream_conv2d_8_start_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_31_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_30), .Q(__stream_conv2d_8_start_31), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_32_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_31), .Q(__stream_conv2d_8_start_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_33_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_32), .Q(__stream_conv2d_8_start_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_34_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_33), .Q(__stream_conv2d_8_start_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_35_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_34), .Q(__stream_conv2d_8_start_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_36_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_35), .Q(__stream_conv2d_8_start_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_37_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_36), .Q(__stream_conv2d_8_start_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_38_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_37), .Q(__stream_conv2d_8_start_38), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_39_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_38), .Q(__stream_conv2d_8_start_39), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_40_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_39), .Q(__stream_conv2d_8_start_40), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_41_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_40), .Q(__stream_conv2d_8_start_41), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_42_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_41), .Q(__stream_conv2d_8_start_42), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_43_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_42), .Q(__stream_conv2d_8_start_43), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_44_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_43), .Q(__stream_conv2d_8_start_44), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_45_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_44), .Q(__stream_conv2d_8_start_45), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __stream_conv2d_8_start_46_reg ( .CLK(CLK), .D(__stream_conv2d_8_start_45), .Q(__stream_conv2d_8_start_46), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_1_reg ( .CLK(CLK), .D(_tmp_541), .Q(__tmp_627_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_2_reg ( .CLK(CLK), .D(__tmp_627_1), .Q(__tmp_627_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_3_reg ( .CLK(CLK), .D(__tmp_627_2), .Q(__tmp_627_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_4_reg ( .CLK(CLK), .D(__tmp_627_3), .Q(__tmp_627_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_5_reg ( .CLK(CLK), .D(__tmp_627_4), .Q(__tmp_627_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_6_reg ( .CLK(CLK), .D(__tmp_627_5), .Q(__tmp_627_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_7_reg ( .CLK(CLK), .D(__tmp_627_6), .Q(__tmp_627_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_8_reg ( .CLK(CLK), .D(__tmp_627_7), .Q(__tmp_627_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_9_reg ( .CLK(CLK), .D(__tmp_627_8), .Q(__tmp_627_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_10_reg ( .CLK(CLK), .D(__tmp_627_9), .Q(__tmp_627_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_11_reg ( .CLK(CLK), .D(__tmp_627_10), .Q(__tmp_627_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_12_reg ( .CLK(CLK), .D(__tmp_627_11), .Q(__tmp_627_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_13_reg ( .CLK(CLK), .D(__tmp_627_12), .Q(__tmp_627_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_14_reg ( .CLK(CLK), .D(__tmp_627_13), .Q(__tmp_627_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_15_reg ( .CLK(CLK), .D(__tmp_627_14), .Q(__tmp_627_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_16_reg ( .CLK(CLK), .D(__tmp_627_15), .Q(__tmp_627_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_17_reg ( .CLK(CLK), .D(__tmp_627_16), .Q(__tmp_627_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_18_reg ( .CLK(CLK), .D(__tmp_627_17), .Q(__tmp_627_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_19_reg ( .CLK(CLK), .D(__tmp_627_18), .Q(__tmp_627_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_20_reg ( .CLK(CLK), .D(__tmp_627_19), .Q(__tmp_627_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_21_reg ( .CLK(CLK), .D(__tmp_627_20), .Q(__tmp_627_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_22_reg ( .CLK(CLK), .D(__tmp_627_21), .Q(__tmp_627_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_23_reg ( .CLK(CLK), .D(__tmp_627_22), .Q(__tmp_627_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_24_reg ( .CLK(CLK), .D(__tmp_627_23), .Q(__tmp_627_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_25_reg ( .CLK(CLK), .D(__tmp_627_24), .Q(__tmp_627_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_26_reg ( .CLK(CLK), .D(__tmp_627_25), .Q(__tmp_627_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_27_reg ( .CLK(CLK), .D(__tmp_627_26), .Q(__tmp_627_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_28_reg ( .CLK(CLK), .D(__tmp_627_27), .Q(__tmp_627_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_29_reg ( .CLK(CLK), .D(__tmp_627_28), .Q(__tmp_627_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_30_reg ( .CLK(CLK), .D(__tmp_627_29), .Q(__tmp_627_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_31_reg ( .CLK(CLK), .D(__tmp_627_30), .Q(__tmp_627_31), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_32_reg ( .CLK(CLK), .D(__tmp_627_31), .Q(__tmp_627_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_33_reg ( .CLK(CLK), .D(__tmp_627_32), .Q(__tmp_627_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_627_34_reg ( .CLK(CLK), .D(__tmp_627_33), .Q(__tmp_627_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_795_43_reg ( .CLK(CLK), .D(__tmp_797_42), .Q(__tmp_795_43), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_795_44_reg ( .CLK(CLK), .D(__tmp_795_43), .Q(__tmp_795_44), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_795_45_reg ( .CLK(CLK), .D(__tmp_795_44), .Q(__tmp_795_45), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_795_46_reg ( .CLK(CLK), .D(__tmp_795_45), .Q(__tmp_795_46), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_13_reg ( .CLK(CLK), .D(__tmp_787_12), .Q(__tmp_797_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_14_reg ( .CLK(CLK), .D(__tmp_797_13), .Q(__tmp_797_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_15_reg ( .CLK(CLK), .D(__tmp_797_14), .Q(__tmp_797_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_16_reg ( .CLK(CLK), .D(__tmp_797_15), .Q(__tmp_797_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_17_reg ( .CLK(CLK), .D(__tmp_797_16), .Q(__tmp_797_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_18_reg ( .CLK(CLK), .D(__tmp_797_17), .Q(__tmp_797_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_19_reg ( .CLK(CLK), .D(__tmp_797_18), .Q(__tmp_797_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_20_reg ( .CLK(CLK), .D(__tmp_797_19), .Q(__tmp_797_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_21_reg ( .CLK(CLK), .D(__tmp_797_20), .Q(__tmp_797_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_22_reg ( .CLK(CLK), .D(__tmp_797_21), .Q(__tmp_797_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_23_reg ( .CLK(CLK), .D(__tmp_797_22), .Q(__tmp_797_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_24_reg ( .CLK(CLK), .D(__tmp_797_23), .Q(__tmp_797_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_25_reg ( .CLK(CLK), .D(__tmp_797_24), .Q(__tmp_797_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_26_reg ( .CLK(CLK), .D(__tmp_797_25), .Q(__tmp_797_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_27_reg ( .CLK(CLK), .D(__tmp_797_26), .Q(__tmp_797_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_28_reg ( .CLK(CLK), .D(__tmp_797_27), .Q(__tmp_797_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_29_reg ( .CLK(CLK), .D(__tmp_797_28), .Q(__tmp_797_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_30_reg ( .CLK(CLK), .D(__tmp_797_29), .Q(__tmp_797_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_31_reg ( .CLK(CLK), .D(__tmp_797_30), .Q(__tmp_797_31), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_32_reg ( .CLK(CLK), .D(__tmp_797_31), .Q(__tmp_797_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_33_reg ( .CLK(CLK), .D(__tmp_797_32), .Q(__tmp_797_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_34_reg ( .CLK(CLK), .D(__tmp_797_33), .Q(__tmp_797_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_35_reg ( .CLK(CLK), .D(__tmp_797_34), .Q(__tmp_797_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_36_reg ( .CLK(CLK), .D(__tmp_797_35), .Q(__tmp_797_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_37_reg ( .CLK(CLK), .D(__tmp_797_36), .Q(__tmp_797_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_38_reg ( .CLK(CLK), .D(__tmp_797_37), .Q(__tmp_797_38), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_39_reg ( .CLK(CLK), .D(__tmp_797_38), .Q(__tmp_797_39), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_40_reg ( .CLK(CLK), .D(__tmp_797_39), .Q(__tmp_797_40), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_41_reg ( .CLK(CLK), .D(__tmp_797_40), .Q(__tmp_797_41), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_797_42_reg ( .CLK(CLK), .D(__tmp_797_41), .Q(__tmp_797_42), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __reduce_max_13_reduce_reset_reg  ( .CLK(CLK), .D(_00620_), .Q(__reduce_max_13_reduce_reset) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream__reduce_max_13_x_data_cond_772_42_reg ( .CLK(CLK), .D(_24260_), .Q(_substream__reduce_max_13_x_data_cond_772_42), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream__reduce_max_13_size_data_cond_772_43_reg ( .CLK(CLK), .D(_24258_), .Q(_substream__reduce_max_13_size_data_cond_772_43), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _40100_ ( .CLK(CLK), .D(_01714_), .Q(_reducecustom_data_191) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40101_ ( .CLK(CLK), .D(_24266_), .Q(_reducecustom_count_191), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pulse_data_193_reg ( .CLK(CLK), .D(_05237_), .Q(_pulse_data_193), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40103_ ( .CLK(CLK), .D(_24265_), .Q(_pulse_count_193), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40104_ ( .CLK(CLK), .D(_24264_), .Q(__variable_wdata_187), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40105_ ( .CLK(CLK), .D(_24263_), .Q(__variable_wdata_188), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_12_x_data_cond_708_24_reg ( .CLK(CLK), .D(_24274_), .Q(_substream_mul_12_x_data_cond_708_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_12_y_data_cond_708_25_reg ( .CLK(CLK), .D(_24272_), .Q(_substream_mul_12_y_data_cond_708_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_12_rshift_data_cond_708_26_reg ( .CLK(CLK), .D(_24270_), .Q(_substream_mul_12_rshift_data_cond_708_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greaterthan_data_175_reg ( .CLK(CLK), .D(_05259_), .Q(_greaterthan_data_175), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40110_ ( .CLK(CLK), .D(_26015_), .Q(_minus_data_177), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40111_ ( .CLK(CLK), .D(__variable_wdata_172), .Q(__delay_data_710), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40112_ ( .CLK(CLK), .D(__variable_wdata_173), .Q(__delay_data_713), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40113_ ( .CLK(CLK), .D(__variable_wdata_174), .Q(__delay_data_716), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(18), .SRST_POLARITY(1'h1), .SRST_VALUE(18'h00000) ) _40114_ ( .CLK(CLK), .D(_25921_), .Q(_sll_data_179), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_709_reg ( .CLK(CLK), .D(_greaterthan_data_175), .Q(__delay_data_709), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40116_ ( .CLK(CLK), .D(__delay_data_710), .Q(__delay_data_711), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40117_ ( .CLK(CLK), .D(__delay_data_713), .Q(__delay_data_714), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40118_ ( .CLK(CLK), .D(__delay_data_716), .Q(__delay_data_717), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40119_ ( .CLK(CLK), .D(_26538_[15:0]), .Q(_cond_data_183), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40120_ ( .CLK(CLK), .D(__delay_data_711), .Q(__delay_data_712), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40121_ ( .CLK(CLK), .D(__delay_data_714), .Q(__delay_data_715), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40122_ ( .CLK(CLK), .D(__delay_data_717), .Q(__delay_data_718), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40123_ ( .CLK(CLK), .D(\__muladd_madd_185.madd._pipe_madd1 ), .Q(__muladd_madd_odata_reg_185), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40124_ ( .CLK(CLK), .D(__delay_data_718), .Q(__delay_data_719), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40125_ ( .CLK(CLK), .D(__delay_data_719), .Q(__delay_data_720), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40126_ ( .CLK(CLK), .D(__delay_data_720), .Q(__delay_data_721), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40127_ ( .CLK(CLK), .D(__delay_data_721), .Q(__delay_data_722), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40128_ ( .CLK(CLK), .D(_25934_), .Q(_sra_data_186), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40129_ ( .CLK(CLK), .D(_24277_), .Q(__variable_wdata_172), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40130_ ( .CLK(CLK), .D(_24276_), .Q(__variable_wdata_173), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40131_ ( .CLK(CLK), .D(_24275_), .Q(__variable_wdata_174), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_11_x_data_cond_691_21_reg ( .CLK(CLK), .D(_24283_), .Q(_substream_mul_11_x_data_cond_691_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_11_y_data_cond_691_22_reg ( .CLK(CLK), .D(_24281_), .Q(_substream_mul_11_y_data_cond_691_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_11_rshift_data_cond_691_23_reg ( .CLK(CLK), .D(_24279_), .Q(_substream_mul_11_rshift_data_cond_691_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greaterthan_data_160_reg ( .CLK(CLK), .D(_05258_), .Q(_greaterthan_data_160), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40136_ ( .CLK(CLK), .D(_26014_), .Q(_minus_data_162), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40137_ ( .CLK(CLK), .D(__variable_wdata_157), .Q(__delay_data_693), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40138_ ( .CLK(CLK), .D(__variable_wdata_158), .Q(__delay_data_696), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40139_ ( .CLK(CLK), .D(__variable_wdata_159), .Q(__delay_data_699), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(18), .SRST_POLARITY(1'h1), .SRST_VALUE(18'h00000) ) _40140_ ( .CLK(CLK), .D(_25920_), .Q(_sll_data_164), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_692_reg ( .CLK(CLK), .D(_greaterthan_data_160), .Q(__delay_data_692), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40142_ ( .CLK(CLK), .D(__delay_data_693), .Q(__delay_data_694), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40143_ ( .CLK(CLK), .D(__delay_data_696), .Q(__delay_data_697), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40144_ ( .CLK(CLK), .D(__delay_data_699), .Q(__delay_data_700), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40145_ ( .CLK(CLK), .D(_26537_[15:0]), .Q(_cond_data_168), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40146_ ( .CLK(CLK), .D(__delay_data_694), .Q(__delay_data_695), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40147_ ( .CLK(CLK), .D(__delay_data_697), .Q(__delay_data_698), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40148_ ( .CLK(CLK), .D(__delay_data_700), .Q(__delay_data_701), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40149_ ( .CLK(CLK), .D(\__muladd_madd_170.madd._pipe_madd1 ), .Q(__muladd_madd_odata_reg_170), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40150_ ( .CLK(CLK), .D(__delay_data_701), .Q(__delay_data_702), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40151_ ( .CLK(CLK), .D(__delay_data_702), .Q(__delay_data_703), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40152_ ( .CLK(CLK), .D(__delay_data_703), .Q(__delay_data_704), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40153_ ( .CLK(CLK), .D(__delay_data_704), .Q(__delay_data_705), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40154_ ( .CLK(CLK), .D(_25933_), .Q(_sra_data_171), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40155_ ( .CLK(CLK), .D(_24286_), .Q(__variable_wdata_157), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40156_ ( .CLK(CLK), .D(_24285_), .Q(__variable_wdata_158), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40157_ ( .CLK(CLK), .D(_24284_), .Q(__variable_wdata_159), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_10_x_data_cond_674_18_reg ( .CLK(CLK), .D(_24292_), .Q(_substream_mul_10_x_data_cond_674_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_10_y_data_cond_674_19_reg ( .CLK(CLK), .D(_24290_), .Q(_substream_mul_10_y_data_cond_674_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_10_rshift_data_cond_674_20_reg ( .CLK(CLK), .D(_24288_), .Q(_substream_mul_10_rshift_data_cond_674_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greaterthan_data_145_reg ( .CLK(CLK), .D(_05257_), .Q(_greaterthan_data_145), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40162_ ( .CLK(CLK), .D(_26013_), .Q(_minus_data_147), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40163_ ( .CLK(CLK), .D(__variable_wdata_142), .Q(__delay_data_676), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40164_ ( .CLK(CLK), .D(__variable_wdata_143), .Q(__delay_data_679), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40165_ ( .CLK(CLK), .D(__variable_wdata_144), .Q(__delay_data_682), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(18), .SRST_POLARITY(1'h1), .SRST_VALUE(18'h00000) ) _40166_ ( .CLK(CLK), .D(_25919_), .Q(_sll_data_149), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_675_reg ( .CLK(CLK), .D(_greaterthan_data_145), .Q(__delay_data_675), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40168_ ( .CLK(CLK), .D(__delay_data_676), .Q(__delay_data_677), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40169_ ( .CLK(CLK), .D(__delay_data_679), .Q(__delay_data_680), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40170_ ( .CLK(CLK), .D(__delay_data_682), .Q(__delay_data_683), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40171_ ( .CLK(CLK), .D(_26536_[15:0]), .Q(_cond_data_153), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40172_ ( .CLK(CLK), .D(__delay_data_677), .Q(__delay_data_678), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40173_ ( .CLK(CLK), .D(__delay_data_680), .Q(__delay_data_681), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40174_ ( .CLK(CLK), .D(__delay_data_683), .Q(__delay_data_684), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40175_ ( .CLK(CLK), .D(\__muladd_madd_155.madd._pipe_madd1 ), .Q(__muladd_madd_odata_reg_155), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40176_ ( .CLK(CLK), .D(__delay_data_684), .Q(__delay_data_685), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40177_ ( .CLK(CLK), .D(__delay_data_685), .Q(__delay_data_686), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40178_ ( .CLK(CLK), .D(__delay_data_686), .Q(__delay_data_687), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40179_ ( .CLK(CLK), .D(__delay_data_687), .Q(__delay_data_688), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40180_ ( .CLK(CLK), .D(_25932_), .Q(_sra_data_156), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40181_ ( .CLK(CLK), .D(_24295_), .Q(__variable_wdata_142), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40182_ ( .CLK(CLK), .D(_24294_), .Q(__variable_wdata_143), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40183_ ( .CLK(CLK), .D(_24293_), .Q(__variable_wdata_144), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_9_x_data_cond_657_15_reg ( .CLK(CLK), .D(_24301_), .Q(_substream_mul_9_x_data_cond_657_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_9_y_data_cond_657_16_reg ( .CLK(CLK), .D(_24299_), .Q(_substream_mul_9_y_data_cond_657_16), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_9_rshift_data_cond_657_17_reg ( .CLK(CLK), .D(_24297_), .Q(_substream_mul_9_rshift_data_cond_657_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greaterthan_data_130_reg ( .CLK(CLK), .D(_05256_), .Q(_greaterthan_data_130), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40188_ ( .CLK(CLK), .D(_26012_), .Q(_minus_data_132), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40189_ ( .CLK(CLK), .D(__variable_wdata_127), .Q(__delay_data_659), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40190_ ( .CLK(CLK), .D(__variable_wdata_128), .Q(__delay_data_662), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40191_ ( .CLK(CLK), .D(__variable_wdata_129), .Q(__delay_data_665), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(18), .SRST_POLARITY(1'h1), .SRST_VALUE(18'h00000) ) _40192_ ( .CLK(CLK), .D(_25918_), .Q(_sll_data_134), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_658_reg ( .CLK(CLK), .D(_greaterthan_data_130), .Q(__delay_data_658), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40194_ ( .CLK(CLK), .D(__delay_data_659), .Q(__delay_data_660), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40195_ ( .CLK(CLK), .D(__delay_data_662), .Q(__delay_data_663), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40196_ ( .CLK(CLK), .D(__delay_data_665), .Q(__delay_data_666), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40197_ ( .CLK(CLK), .D(_26535_[15:0]), .Q(_cond_data_138), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40198_ ( .CLK(CLK), .D(__delay_data_660), .Q(__delay_data_661), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40199_ ( .CLK(CLK), .D(__delay_data_663), .Q(__delay_data_664), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40200_ ( .CLK(CLK), .D(__delay_data_666), .Q(__delay_data_667), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40201_ ( .CLK(CLK), .D(\__muladd_madd_140.madd._pipe_madd1 ), .Q(__muladd_madd_odata_reg_140), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40202_ ( .CLK(CLK), .D(__delay_data_667), .Q(__delay_data_668), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40203_ ( .CLK(CLK), .D(__delay_data_668), .Q(__delay_data_669), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40204_ ( .CLK(CLK), .D(__delay_data_669), .Q(__delay_data_670), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40205_ ( .CLK(CLK), .D(__delay_data_670), .Q(__delay_data_671), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40206_ ( .CLK(CLK), .D(_25931_), .Q(_sra_data_141), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40207_ ( .CLK(CLK), .D(_24304_), .Q(__variable_wdata_127), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40208_ ( .CLK(CLK), .D(_24303_), .Q(__variable_wdata_128), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40209_ ( .CLK(CLK), .D(_24302_), .Q(__variable_wdata_129), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_8_x_data_cond_640_12_reg ( .CLK(CLK), .D(_24310_), .Q(_substream_mul_8_x_data_cond_640_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_8_y_data_cond_640_13_reg ( .CLK(CLK), .D(_24308_), .Q(_substream_mul_8_y_data_cond_640_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_8_rshift_data_cond_640_14_reg ( .CLK(CLK), .D(_24306_), .Q(_substream_mul_8_rshift_data_cond_640_14), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greaterthan_data_115_reg ( .CLK(CLK), .D(_05255_), .Q(_greaterthan_data_115), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40214_ ( .CLK(CLK), .D(_26011_), .Q(_minus_data_117), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40215_ ( .CLK(CLK), .D(__variable_wdata_112), .Q(__delay_data_642), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40216_ ( .CLK(CLK), .D(__variable_wdata_113), .Q(__delay_data_645), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40217_ ( .CLK(CLK), .D(__variable_wdata_114), .Q(__delay_data_648), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(18), .SRST_POLARITY(1'h1), .SRST_VALUE(18'h00000) ) _40218_ ( .CLK(CLK), .D(_25917_), .Q(_sll_data_119), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_641_reg ( .CLK(CLK), .D(_greaterthan_data_115), .Q(__delay_data_641), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40220_ ( .CLK(CLK), .D(__delay_data_642), .Q(__delay_data_643), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40221_ ( .CLK(CLK), .D(__delay_data_645), .Q(__delay_data_646), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40222_ ( .CLK(CLK), .D(__delay_data_648), .Q(__delay_data_649), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40223_ ( .CLK(CLK), .D(_26534_[15:0]), .Q(_cond_data_123), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40224_ ( .CLK(CLK), .D(__delay_data_643), .Q(__delay_data_644), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40225_ ( .CLK(CLK), .D(__delay_data_646), .Q(__delay_data_647), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40226_ ( .CLK(CLK), .D(__delay_data_649), .Q(__delay_data_650), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40227_ ( .CLK(CLK), .D(\__muladd_madd_125.madd._pipe_madd1 ), .Q(__muladd_madd_odata_reg_125), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40228_ ( .CLK(CLK), .D(__delay_data_650), .Q(__delay_data_651), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40229_ ( .CLK(CLK), .D(__delay_data_651), .Q(__delay_data_652), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40230_ ( .CLK(CLK), .D(__delay_data_652), .Q(__delay_data_653), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40231_ ( .CLK(CLK), .D(__delay_data_653), .Q(__delay_data_654), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40232_ ( .CLK(CLK), .D(_25930_), .Q(_sra_data_126), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40233_ ( .CLK(CLK), .D(_24313_), .Q(__variable_wdata_112), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40234_ ( .CLK(CLK), .D(_24312_), .Q(__variable_wdata_113), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40235_ ( .CLK(CLK), .D(_24311_), .Q(__variable_wdata_114), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_7_x_data_cond_623_9_reg ( .CLK(CLK), .D(_24319_), .Q(_substream_mul_7_x_data_cond_623_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_7_y_data_cond_623_10_reg ( .CLK(CLK), .D(_24317_), .Q(_substream_mul_7_y_data_cond_623_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_7_rshift_data_cond_623_11_reg ( .CLK(CLK), .D(_24315_), .Q(_substream_mul_7_rshift_data_cond_623_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greaterthan_data_100_reg ( .CLK(CLK), .D(_05254_), .Q(_greaterthan_data_100), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40240_ ( .CLK(CLK), .D(_26010_), .Q(_minus_data_102), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40241_ ( .CLK(CLK), .D(__variable_wdata_97), .Q(__delay_data_625), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40242_ ( .CLK(CLK), .D(__variable_wdata_98), .Q(__delay_data_628), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40243_ ( .CLK(CLK), .D(__variable_wdata_99), .Q(__delay_data_631), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(18), .SRST_POLARITY(1'h1), .SRST_VALUE(18'h00000) ) _40244_ ( .CLK(CLK), .D(_25916_), .Q(_sll_data_104), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_624_reg ( .CLK(CLK), .D(_greaterthan_data_100), .Q(__delay_data_624), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40246_ ( .CLK(CLK), .D(__delay_data_625), .Q(__delay_data_626), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40247_ ( .CLK(CLK), .D(__delay_data_628), .Q(__delay_data_629), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40248_ ( .CLK(CLK), .D(__delay_data_631), .Q(__delay_data_632), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40249_ ( .CLK(CLK), .D(_26533_[15:0]), .Q(_cond_data_108), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40250_ ( .CLK(CLK), .D(__delay_data_626), .Q(__delay_data_627), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40251_ ( .CLK(CLK), .D(__delay_data_629), .Q(__delay_data_630), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40252_ ( .CLK(CLK), .D(__delay_data_632), .Q(__delay_data_633), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40253_ ( .CLK(CLK), .D(\__muladd_madd_110.madd._pipe_madd1 ), .Q(__muladd_madd_odata_reg_110), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40254_ ( .CLK(CLK), .D(__delay_data_633), .Q(__delay_data_634), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40255_ ( .CLK(CLK), .D(__delay_data_634), .Q(__delay_data_635), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40256_ ( .CLK(CLK), .D(__delay_data_635), .Q(__delay_data_636), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40257_ ( .CLK(CLK), .D(__delay_data_636), .Q(__delay_data_637), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40258_ ( .CLK(CLK), .D(_25929_), .Q(_sra_data_111), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40259_ ( .CLK(CLK), .D(_24322_), .Q(__variable_wdata_97), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40260_ ( .CLK(CLK), .D(_24321_), .Q(__variable_wdata_98), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40261_ ( .CLK(CLK), .D(_24320_), .Q(__variable_wdata_99), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_6_x_data_cond_606_6_reg ( .CLK(CLK), .D(_24328_), .Q(_substream_mul_6_x_data_cond_606_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_6_y_data_cond_606_7_reg ( .CLK(CLK), .D(_24326_), .Q(_substream_mul_6_y_data_cond_606_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_6_rshift_data_cond_606_8_reg ( .CLK(CLK), .D(_24324_), .Q(_substream_mul_6_rshift_data_cond_606_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greaterthan_data_85_reg ( .CLK(CLK), .D(_05253_), .Q(_greaterthan_data_85), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40266_ ( .CLK(CLK), .D(_26009_), .Q(_minus_data_87), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40267_ ( .CLK(CLK), .D(__variable_wdata_82), .Q(__delay_data_608), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40268_ ( .CLK(CLK), .D(__variable_wdata_83), .Q(__delay_data_611), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40269_ ( .CLK(CLK), .D(__variable_wdata_84), .Q(__delay_data_614), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(18), .SRST_POLARITY(1'h1), .SRST_VALUE(18'h00000) ) _40270_ ( .CLK(CLK), .D(_25915_), .Q(_sll_data_89), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_607_reg ( .CLK(CLK), .D(_greaterthan_data_85), .Q(__delay_data_607), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40272_ ( .CLK(CLK), .D(__delay_data_608), .Q(__delay_data_609), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40273_ ( .CLK(CLK), .D(__delay_data_611), .Q(__delay_data_612), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40274_ ( .CLK(CLK), .D(__delay_data_614), .Q(__delay_data_615), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40275_ ( .CLK(CLK), .D(_26532_[15:0]), .Q(_cond_data_93), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40276_ ( .CLK(CLK), .D(__delay_data_609), .Q(__delay_data_610), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40277_ ( .CLK(CLK), .D(__delay_data_612), .Q(__delay_data_613), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40278_ ( .CLK(CLK), .D(__delay_data_615), .Q(__delay_data_616), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40279_ ( .CLK(CLK), .D(\__muladd_madd_95.madd._pipe_madd1 ), .Q(__muladd_madd_odata_reg_95), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40280_ ( .CLK(CLK), .D(__delay_data_616), .Q(__delay_data_617), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40281_ ( .CLK(CLK), .D(__delay_data_617), .Q(__delay_data_618), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40282_ ( .CLK(CLK), .D(__delay_data_618), .Q(__delay_data_619), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40283_ ( .CLK(CLK), .D(__delay_data_619), .Q(__delay_data_620), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40284_ ( .CLK(CLK), .D(_25928_), .Q(_sra_data_96), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40285_ ( .CLK(CLK), .D(_24331_), .Q(__variable_wdata_82), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40286_ ( .CLK(CLK), .D(_24330_), .Q(__variable_wdata_83), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40287_ ( .CLK(CLK), .D(_24329_), .Q(__variable_wdata_84), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_5_x_data_cond_589_3_reg ( .CLK(CLK), .D(_24337_), .Q(_substream_mul_5_x_data_cond_589_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_5_y_data_cond_589_4_reg ( .CLK(CLK), .D(_24335_), .Q(_substream_mul_5_y_data_cond_589_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_5_rshift_data_cond_589_5_reg ( .CLK(CLK), .D(_24333_), .Q(_substream_mul_5_rshift_data_cond_589_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greaterthan_data_70_reg ( .CLK(CLK), .D(_05252_), .Q(_greaterthan_data_70), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40292_ ( .CLK(CLK), .D(_26008_), .Q(_minus_data_72), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40293_ ( .CLK(CLK), .D(__variable_wdata_67), .Q(__delay_data_591), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40294_ ( .CLK(CLK), .D(__variable_wdata_68), .Q(__delay_data_594), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40295_ ( .CLK(CLK), .D(__variable_wdata_69), .Q(__delay_data_597), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(18), .SRST_POLARITY(1'h1), .SRST_VALUE(18'h00000) ) _40296_ ( .CLK(CLK), .D(_25914_), .Q(_sll_data_74), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_590_reg ( .CLK(CLK), .D(_greaterthan_data_70), .Q(__delay_data_590), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40298_ ( .CLK(CLK), .D(__delay_data_591), .Q(__delay_data_592), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40299_ ( .CLK(CLK), .D(__delay_data_594), .Q(__delay_data_595), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40300_ ( .CLK(CLK), .D(__delay_data_597), .Q(__delay_data_598), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40301_ ( .CLK(CLK), .D(_26531_[15:0]), .Q(_cond_data_78), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40302_ ( .CLK(CLK), .D(__delay_data_592), .Q(__delay_data_593), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40303_ ( .CLK(CLK), .D(__delay_data_595), .Q(__delay_data_596), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40304_ ( .CLK(CLK), .D(__delay_data_598), .Q(__delay_data_599), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40305_ ( .CLK(CLK), .D(\__muladd_madd_80.madd._pipe_madd1 ), .Q(__muladd_madd_odata_reg_80), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40306_ ( .CLK(CLK), .D(__delay_data_599), .Q(__delay_data_600), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40307_ ( .CLK(CLK), .D(__delay_data_600), .Q(__delay_data_601), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40308_ ( .CLK(CLK), .D(__delay_data_601), .Q(__delay_data_602), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40309_ ( .CLK(CLK), .D(__delay_data_602), .Q(__delay_data_603), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40310_ ( .CLK(CLK), .D(_25927_), .Q(_sra_data_81), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40311_ ( .CLK(CLK), .D(_24340_), .Q(__variable_wdata_67), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40312_ ( .CLK(CLK), .D(_24339_), .Q(__variable_wdata_68), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40313_ ( .CLK(CLK), .D(_24338_), .Q(__variable_wdata_69), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_4_x_data_cond_572_0_reg ( .CLK(CLK), .D(_24352_), .Q(_substream_mul_4_x_data_cond_572_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_4_y_data_cond_572_1_reg ( .CLK(CLK), .D(_24350_), .Q(_substream_mul_4_y_data_cond_572_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_4_rshift_data_cond_572_2_reg ( .CLK(CLK), .D(_24348_), .Q(_substream_mul_4_rshift_data_cond_572_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_4_x_data_cond_854_44_reg ( .CLK(CLK), .D(_24346_), .Q(_substream_mul_4_x_data_cond_854_44), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_4_y_data_cond_854_45_reg ( .CLK(CLK), .D(_24344_), .Q(_substream_mul_4_y_data_cond_854_45), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_4_rshift_data_cond_854_46_reg ( .CLK(CLK), .D(_24342_), .Q(_substream_mul_4_rshift_data_cond_854_46), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greaterthan_data_55_reg ( .CLK(CLK), .D(_05251_), .Q(_greaterthan_data_55), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40321_ ( .CLK(CLK), .D(_26007_), .Q(_minus_data_57), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40322_ ( .CLK(CLK), .D(__variable_wdata_52), .Q(__delay_data_574), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40323_ ( .CLK(CLK), .D(__variable_wdata_53), .Q(__delay_data_577), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40324_ ( .CLK(CLK), .D(__variable_wdata_54), .Q(__delay_data_580), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(18), .SRST_POLARITY(1'h1), .SRST_VALUE(18'h00000) ) _40325_ ( .CLK(CLK), .D(_25913_), .Q(_sll_data_59), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_573_reg ( .CLK(CLK), .D(_greaterthan_data_55), .Q(__delay_data_573), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40327_ ( .CLK(CLK), .D(__delay_data_574), .Q(__delay_data_575), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40328_ ( .CLK(CLK), .D(__delay_data_577), .Q(__delay_data_578), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40329_ ( .CLK(CLK), .D(__delay_data_580), .Q(__delay_data_581), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40330_ ( .CLK(CLK), .D(_26530_[15:0]), .Q(_cond_data_63), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40331_ ( .CLK(CLK), .D(__delay_data_575), .Q(__delay_data_576), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40332_ ( .CLK(CLK), .D(__delay_data_578), .Q(__delay_data_579), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40333_ ( .CLK(CLK), .D(__delay_data_581), .Q(__delay_data_582), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40334_ ( .CLK(CLK), .D(\__muladd_madd_65.madd._pipe_madd1 ), .Q(__muladd_madd_odata_reg_65), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40335_ ( .CLK(CLK), .D(__delay_data_582), .Q(__delay_data_583), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40336_ ( .CLK(CLK), .D(__delay_data_583), .Q(__delay_data_584), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40337_ ( .CLK(CLK), .D(__delay_data_584), .Q(__delay_data_585), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40338_ ( .CLK(CLK), .D(__delay_data_585), .Q(__delay_data_586), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(16), .SRST_POLARITY(1'h1), .SRST_VALUE(16'h0000) ) _40339_ ( .CLK(CLK), .D(_25926_), .Q(_sra_data_66), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40340_ ( .CLK(CLK), .D(_24358_), .Q(__variable_wdata_52), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40341_ ( .CLK(CLK), .D(_24356_), .Q(__variable_wdata_53), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40342_ ( .CLK(CLK), .D(_24354_), .Q(__variable_wdata_54), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_rshift_clip_3_x_data_cond_743_39_reg ( .CLK(CLK), .D(_24370_), .Q(_substream_mul_rshift_clip_3_x_data_cond_743_39), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_rshift_clip_3_y_data_cond_743_40_reg ( .CLK(CLK), .D(_24368_), .Q(_substream_mul_rshift_clip_3_y_data_cond_743_40), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_rshift_clip_3_rshift_data_cond_743_41_reg ( .CLK(CLK), .D(_24366_), .Q(_substream_mul_rshift_clip_3_rshift_data_cond_743_41), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_rshift_clip_3_x_data_cond_864_51_reg ( .CLK(CLK), .D(_24364_), .Q(_substream_mul_rshift_clip_3_x_data_cond_864_51), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_rshift_clip_3_y_data_cond_864_52_reg ( .CLK(CLK), .D(_24362_), .Q(_substream_mul_rshift_clip_3_y_data_cond_864_52), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_mul_rshift_clip_3_rshift_data_cond_864_53_reg ( .CLK(CLK), .D(_24360_), .Q(_substream_mul_rshift_clip_3_rshift_data_cond_864_53), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(40), .SRST_POLARITY(1'h1), .SRST_VALUE(40'h0000000000) ) _40349_ ( .CLK(CLK), .D(\_times_mul_39.mult._pipe_mul1 ), .Q(_times_mul_odata_reg_39), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(6), .SRST_POLARITY(1'h1), .SRST_VALUE(6'h00) ) _40350_ ( .CLK(CLK), .D(__variable_wdata_38), .Q(__delay_data_744), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(6), .SRST_POLARITY(1'h1), .SRST_VALUE(6'h00) ) _40351_ ( .CLK(CLK), .D(__delay_data_744), .Q(__delay_data_745), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(6), .SRST_POLARITY(1'h1), .SRST_VALUE(6'h00) ) _40352_ ( .CLK(CLK), .D(__delay_data_745), .Q(__delay_data_746), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(6), .SRST_POLARITY(1'h1), .SRST_VALUE(6'h00) ) _40353_ ( .CLK(CLK), .D(__delay_data_746), .Q(__delay_data_747), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(40), .SRST_POLARITY(1'h1), .SRST_VALUE(40'h0000000000) ) _40354_ ( .CLK(CLK), .D(_25925_), .Q(_sra_data_40), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greaterthan_data_41_reg ( .CLK(CLK), .D(_05250_), .Q(_greaterthan_data_41), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _lessthan_data_45_reg ( .CLK(CLK), .D(_05872_), .Q(_lessthan_data_45), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greatereq_data_49_reg ( .CLK(CLK), .D(_05235_), .Q(_greatereq_data_49), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(40), .SRST_POLARITY(1'h1), .SRST_VALUE(40'h0000000000) ) _40358_ ( .CLK(CLK), .D(_sra_data_40), .Q(__delay_data_748), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(40), .SRST_POLARITY(1'h1), .SRST_VALUE(40'h0000000000) ) _40359_ ( .CLK(CLK), .D(_26514_), .Q(_cond_data_43), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(40), .SRST_POLARITY(1'h1), .SRST_VALUE(40'h0000000000) ) _40360_ ( .CLK(CLK), .D(_26515_), .Q(_cond_data_47), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_749_reg ( .CLK(CLK), .D(_greatereq_data_49), .Q(__delay_data_749), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40362_ ( .CLK(CLK), .D(_26516_[7:0]), .Q(_cond_data_51), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40363_ ( .CLK(CLK), .D(_24376_), .Q(__variable_wdata_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40364_ ( .CLK(CLK), .D(_24374_), .Q(__variable_wdata_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(6), .SRST_POLARITY(1'h1), .SRST_VALUE(6'h00) ) _40365_ ( .CLK(CLK), .D(_24372_), .Q(__variable_wdata_38), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_787_10_reg ( .CLK(CLK), .D(__tmp_775_9), .Q(__tmp_787_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_787_11_reg ( .CLK(CLK), .D(__tmp_787_10), .Q(__tmp_787_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_787_12_reg ( .CLK(CLK), .D(__tmp_787_11), .Q(__tmp_787_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1107_10_reg ( .CLK(CLK), .D(__tmp_1095_9), .Q(__tmp_1107_10), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1107_11_reg ( .CLK(CLK), .D(__tmp_1107_10), .Q(__tmp_1107_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1107_12_reg ( .CLK(CLK), .D(__tmp_1107_11), .Q(__tmp_1107_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_add_tree_2_var0_data_cond_725_27_reg ( .CLK(CLK), .D(_24394_), .Q(_substream_add_tree_2_var0_data_cond_725_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_add_tree_2_var1_data_cond_725_28_reg ( .CLK(CLK), .D(_24392_), .Q(_substream_add_tree_2_var1_data_cond_725_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_add_tree_2_var2_data_cond_725_29_reg ( .CLK(CLK), .D(_24390_), .Q(_substream_add_tree_2_var2_data_cond_725_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_add_tree_2_var3_data_cond_725_30_reg ( .CLK(CLK), .D(_24388_), .Q(_substream_add_tree_2_var3_data_cond_725_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_add_tree_2_var4_data_cond_725_31_reg ( .CLK(CLK), .D(_24386_), .Q(_substream_add_tree_2_var4_data_cond_725_31), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_add_tree_2_var5_data_cond_725_32_reg ( .CLK(CLK), .D(_24384_), .Q(_substream_add_tree_2_var5_data_cond_725_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_add_tree_2_var6_data_cond_725_33_reg ( .CLK(CLK), .D(_24382_), .Q(_substream_add_tree_2_var6_data_cond_725_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_add_tree_2_var7_data_cond_725_34_reg ( .CLK(CLK), .D(_24380_), .Q(_substream_add_tree_2_var7_data_cond_725_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_add_tree_2_var8_data_cond_725_35_reg ( .CLK(CLK), .D(_24378_), .Q(_substream_add_tree_2_var8_data_cond_725_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40381_ ( .CLK(CLK), .D(_22127_), .Q(__plusn_data_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40382_ ( .CLK(CLK), .D(_22129_), .Q(__plusn_data_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40383_ ( .CLK(CLK), .D(_22131_), .Q(__plusn_data_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40384_ ( .CLK(CLK), .D(_22133_), .Q(__plusn_data_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40385_ ( .CLK(CLK), .D(_24403_), .Q(__variable_wdata_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40386_ ( .CLK(CLK), .D(_24402_), .Q(__variable_wdata_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40387_ ( .CLK(CLK), .D(_24401_), .Q(__variable_wdata_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40388_ ( .CLK(CLK), .D(_24400_), .Q(__variable_wdata_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40389_ ( .CLK(CLK), .D(_24399_), .Q(__variable_wdata_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40390_ ( .CLK(CLK), .D(_24398_), .Q(__variable_wdata_27), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40391_ ( .CLK(CLK), .D(_24397_), .Q(__variable_wdata_28), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40392_ ( .CLK(CLK), .D(_24396_), .Q(__variable_wdata_29), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40393_ ( .CLK(CLK), .D(_24395_), .Q(__variable_wdata_30), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_add_tree_1_var0_data_cond_857_47_reg ( .CLK(CLK), .D(_24405_), .Q(_substream_add_tree_1_var0_data_cond_857_47), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40395_ ( .CLK(CLK), .D(_24406_), .Q(__variable_wdata_20), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _acc_0_reduce_reset_reg  ( .CLK(CLK), .D(_01356_), .Q(_acc_0_reduce_reset) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_acc_0_x_data_cond_727_36_reg ( .CLK(CLK), .D(_24418_), .Q(_substream_acc_0_x_data_cond_727_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_acc_0_rshift_data_cond_727_37_reg ( .CLK(CLK), .D(_24416_), .Q(_substream_acc_0_rshift_data_cond_727_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_acc_0_size_data_cond_727_38_reg ( .CLK(CLK), .D(_24414_), .Q(_substream_acc_0_size_data_cond_727_38), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_acc_0_x_data_cond_859_48_reg ( .CLK(CLK), .D(_24412_), .Q(_substream_acc_0_x_data_cond_859_48), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_acc_0_rshift_data_cond_859_49_reg ( .CLK(CLK), .D(_24410_), .Q(_substream_acc_0_rshift_data_cond_859_49), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _substream_acc_0_size_data_cond_859_50_reg ( .CLK(CLK), .D(_24408_), .Q(_substream_acc_0_size_data_cond_859_50), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _greaterthan_data_3_reg ( .CLK(CLK), .D(_05249_), .Q(_greaterthan_data_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(6), .SRST_POLARITY(1'h1), .SRST_VALUE(6'h00) ) _40404_ ( .CLK(CLK), .D(_26006_), .Q(_minus_data_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40405_ ( .CLK(CLK), .D(_24432_), .Q(_reduceadd_data_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _40406_ ( .CLK(CLK), .D(_24430_), .Q(_reduceadd_count_15), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _pulse_data_17_reg ( .CLK(CLK), .D(_05234_), .Q(_pulse_data_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _40408_ ( .CLK(CLK), .D(_24429_), .Q(_pulse_count_17), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(6), .SRST_POLARITY(1'h1), .SRST_VALUE(6'h00) ) _40409_ ( .CLK(CLK), .D(__variable_wdata_1), .Q(__delay_data_731), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(66), .SRST_POLARITY(1'h1), .SRST_VALUE(66'h00000000000000000) ) _40410_ ( .CLK(CLK), .D(_25912_), .Q(_sll_data_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_728_reg ( .CLK(CLK), .D(_greaterthan_data_3), .Q(__delay_data_728), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40412_ ( .CLK(CLK), .D(_reduceadd_data_15), .Q(__delay_data_729), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(6), .SRST_POLARITY(1'h1), .SRST_VALUE(6'h00) ) _40413_ ( .CLK(CLK), .D(__delay_data_731), .Q(__delay_data_732), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_735_reg ( .CLK(CLK), .D(_pulse_data_17), .Q(__delay_data_735), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40415_ ( .CLK(CLK), .D(_26513_[31:0]), .Q(_cond_data_11), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40416_ ( .CLK(CLK), .D(__delay_data_729), .Q(__delay_data_730), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(6), .SRST_POLARITY(1'h1), .SRST_VALUE(6'h00) ) _40417_ ( .CLK(CLK), .D(__delay_data_732), .Q(__delay_data_733), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_736_reg ( .CLK(CLK), .D(__delay_data_735), .Q(__delay_data_736), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40419_ ( .CLK(CLK), .D(_22125_), .Q(_plus_data_18), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(6), .SRST_POLARITY(1'h1), .SRST_VALUE(6'h00) ) _40420_ ( .CLK(CLK), .D(__delay_data_733), .Q(__delay_data_734), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_737_reg ( .CLK(CLK), .D(__delay_data_736), .Q(__delay_data_737), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40422_ ( .CLK(CLK), .D(_25924_), .Q(_sra_data_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __delay_data_738_reg ( .CLK(CLK), .D(__delay_data_737), .Q(__delay_data_738), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40424_ ( .CLK(CLK), .D(_24428_), .Q(__variable_wdata_0), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(6), .SRST_POLARITY(1'h1), .SRST_VALUE(6'h00) ) _40425_ ( .CLK(CLK), .D(_24426_), .Q(__variable_wdata_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40426_ ( .CLK(CLK), .D(_24424_), .Q(__variable_wdata_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_775_1_reg ( .CLK(CLK), .D(_tmp_771), .Q(__tmp_775_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_775_2_reg ( .CLK(CLK), .D(__tmp_775_1), .Q(__tmp_775_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_775_3_reg ( .CLK(CLK), .D(__tmp_775_2), .Q(__tmp_775_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_775_4_reg ( .CLK(CLK), .D(__tmp_775_3), .Q(__tmp_775_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_775_5_reg ( .CLK(CLK), .D(__tmp_775_4), .Q(__tmp_775_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_775_6_reg ( .CLK(CLK), .D(__tmp_775_5), .Q(__tmp_775_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_775_7_reg ( .CLK(CLK), .D(__tmp_775_6), .Q(__tmp_775_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_775_8_reg ( .CLK(CLK), .D(__tmp_775_7), .Q(__tmp_775_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_775_9_reg ( .CLK(CLK), .D(__tmp_775_8), .Q(__tmp_775_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1095_1_reg ( .CLK(CLK), .D(_tmp_1091), .Q(__tmp_1095_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1095_2_reg ( .CLK(CLK), .D(__tmp_1095_1), .Q(__tmp_1095_2), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1095_3_reg ( .CLK(CLK), .D(__tmp_1095_2), .Q(__tmp_1095_3), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1095_4_reg ( .CLK(CLK), .D(__tmp_1095_3), .Q(__tmp_1095_4), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1095_5_reg ( .CLK(CLK), .D(__tmp_1095_4), .Q(__tmp_1095_5), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1095_6_reg ( .CLK(CLK), .D(__tmp_1095_5), .Q(__tmp_1095_6), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1095_7_reg ( .CLK(CLK), .D(__tmp_1095_6), .Q(__tmp_1095_7), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1095_8_reg ( .CLK(CLK), .D(__tmp_1095_7), .Q(__tmp_1095_8), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1095_9_reg ( .CLK(CLK), .D(__tmp_1095_8), .Q(__tmp_1095_9), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(7), .SRST_POLARITY(1'h1), .SRST_VALUE(7'h00) ) _40445_ ( .CLK(CLK), .D(_24443_), .Q(ram_w32_l128_id0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(7), .SRST_POLARITY(1'h1), .SRST_VALUE(7'h00) ) _40446_ ( .CLK(CLK), .D(_24441_), .Q(ram_w32_l128_id0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40447_ ( .CLK(CLK), .D(_24439_), .Q(ram_w32_l128_id0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w32_l128_id0_1_wenable_reg ( .CLK(CLK), .D(_24438_), .Q(ram_w32_l128_id0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40449_ ( .CLK(CLK), .D(_24436_), .Q(_tmp_12), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_13_reg ( .CLK(CLK), .D(_24434_), .Q(_tmp_13), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w32_l128_id0_cond_2_1_reg ( .CLK(CLK), .D(_tmp_336), .Q(_ram_w32_l128_id0_cond_2_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w32_l128_id0_cond_4_1_reg ( .CLK(CLK), .D(_tmp_992), .Q(_ram_w32_l128_id0_cond_4_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40453_ ( .CLK(CLK), .D(_24464_), .Q(ram_w8_l2048_id19_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40454_ ( .CLK(CLK), .D(_24463_), .Q(ram_w8_l2048_id19_3_0_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id19_3_0_wenable_reg ( .CLK(CLK), .D(_24462_), .Q(ram_w8_l2048_id19_3_0_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40456_ ( .CLK(CLK), .D(_24460_), .Q(ram_w8_l2048_id19_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id19_3_cond_0_1_reg ( .CLK(CLK), .D(_05665_), .Q(_ram_w8_l2048_id19_3_cond_0_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_835_reg ( .CLK(CLK), .D(_24458_), .Q(_tmp_835), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_840_1_reg ( .CLK(CLK), .D(_tmp_840), .Q(__tmp_840_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40460_ ( .CLK(CLK), .D(_tmp_841), .Q(__tmp_841_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_842_reg ( .CLK(CLK), .D(_24456_), .Q(_tmp_842), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_843_reg ( .CLK(CLK), .D(_24453_), .Q(_tmp_843), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_844_reg ( .CLK(CLK), .D(_24451_), .Q(_tmp_844), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_845_reg ( .CLK(CLK), .D(_24447_), .Q(_tmp_845), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40465_ ( .CLK(CLK), .D(_24445_), .Q(_tmp_846), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40466_ ( .CLK(CLK), .D(_24485_), .Q(ram_w8_l2048_id19_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40467_ ( .CLK(CLK), .D(_24484_), .Q(ram_w8_l2048_id19_2_0_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id19_2_0_wenable_reg ( .CLK(CLK), .D(_24483_), .Q(ram_w8_l2048_id19_2_0_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40469_ ( .CLK(CLK), .D(_24481_), .Q(ram_w8_l2048_id19_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id19_2_cond_0_1_reg ( .CLK(CLK), .D(_05659_), .Q(_ram_w8_l2048_id19_2_cond_0_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_823_reg ( .CLK(CLK), .D(_24479_), .Q(_tmp_823), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_828_1_reg ( .CLK(CLK), .D(_tmp_828), .Q(__tmp_828_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40473_ ( .CLK(CLK), .D(_tmp_829), .Q(__tmp_829_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_830_reg ( .CLK(CLK), .D(_24477_), .Q(_tmp_830), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_831_reg ( .CLK(CLK), .D(_24474_), .Q(_tmp_831), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_832_reg ( .CLK(CLK), .D(_24472_), .Q(_tmp_832), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_833_reg ( .CLK(CLK), .D(_24468_), .Q(_tmp_833), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40478_ ( .CLK(CLK), .D(_24466_), .Q(_tmp_834), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40479_ ( .CLK(CLK), .D(_24506_), .Q(ram_w8_l2048_id19_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40480_ ( .CLK(CLK), .D(_24505_), .Q(ram_w8_l2048_id19_1_0_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id19_1_0_wenable_reg ( .CLK(CLK), .D(_24504_), .Q(ram_w8_l2048_id19_1_0_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40482_ ( .CLK(CLK), .D(_24502_), .Q(ram_w8_l2048_id19_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id19_1_cond_0_1_reg ( .CLK(CLK), .D(_05653_), .Q(_ram_w8_l2048_id19_1_cond_0_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_811_reg ( .CLK(CLK), .D(_24500_), .Q(_tmp_811), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_816_1_reg ( .CLK(CLK), .D(_tmp_816), .Q(__tmp_816_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40486_ ( .CLK(CLK), .D(_tmp_817), .Q(__tmp_817_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_818_reg ( .CLK(CLK), .D(_24498_), .Q(_tmp_818), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_819_reg ( .CLK(CLK), .D(_24495_), .Q(_tmp_819), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_820_reg ( .CLK(CLK), .D(_24493_), .Q(_tmp_820), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_821_reg ( .CLK(CLK), .D(_24489_), .Q(_tmp_821), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40491_ ( .CLK(CLK), .D(_24487_), .Q(_tmp_822), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40492_ ( .CLK(CLK), .D(_24509_), .Q(_dataflow_cat_data_74), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_cat_valid_74_reg ( .CLK(CLK), .D(_24508_), .Q(_dataflow_cat_valid_74), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40494_ ( .CLK(CLK), .D(_24530_), .Q(ram_w8_l2048_id19_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40495_ ( .CLK(CLK), .D(_24529_), .Q(ram_w8_l2048_id19_0_0_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id19_0_0_wenable_reg ( .CLK(CLK), .D(_24528_), .Q(ram_w8_l2048_id19_0_0_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40497_ ( .CLK(CLK), .D(_24526_), .Q(ram_w8_l2048_id19_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id19_0_cond_0_1_reg ( .CLK(CLK), .D(_05644_), .Q(_ram_w8_l2048_id19_0_cond_0_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_799_reg ( .CLK(CLK), .D(_24524_), .Q(_tmp_799), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_804_1_reg ( .CLK(CLK), .D(_tmp_804), .Q(__tmp_804_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40501_ ( .CLK(CLK), .D(_tmp_805), .Q(__tmp_805_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_806_reg ( .CLK(CLK), .D(_24522_), .Q(_tmp_806), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_807_reg ( .CLK(CLK), .D(_24519_), .Q(_tmp_807), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_808_reg ( .CLK(CLK), .D(_24517_), .Q(_tmp_808), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_809_reg ( .CLK(CLK), .D(_24513_), .Q(_tmp_809), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40506_ ( .CLK(CLK), .D(_24511_), .Q(_tmp_810), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40507_ ( .CLK(CLK), .D(_24535_), .Q(ram_w8_l2048_id18_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40508_ ( .CLK(CLK), .D(_24534_), .Q(ram_w8_l2048_id18_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40509_ ( .CLK(CLK), .D(_24533_), .Q(ram_w8_l2048_id18_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id18_3_1_wenable_reg ( .CLK(CLK), .D(_24532_), .Q(ram_w8_l2048_id18_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40511_ ( .CLK(CLK), .D(_24540_), .Q(ram_w8_l2048_id18_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40512_ ( .CLK(CLK), .D(_24539_), .Q(ram_w8_l2048_id18_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40513_ ( .CLK(CLK), .D(_24538_), .Q(ram_w8_l2048_id18_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id18_2_1_wenable_reg ( .CLK(CLK), .D(_24537_), .Q(ram_w8_l2048_id18_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40515_ ( .CLK(CLK), .D(_24545_), .Q(ram_w8_l2048_id18_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40516_ ( .CLK(CLK), .D(_24544_), .Q(ram_w8_l2048_id18_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40517_ ( .CLK(CLK), .D(_24543_), .Q(ram_w8_l2048_id18_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id18_1_1_wenable_reg ( .CLK(CLK), .D(_24542_), .Q(ram_w8_l2048_id18_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40519_ ( .CLK(CLK), .D(_24550_), .Q(ram_w8_l2048_id18_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40520_ ( .CLK(CLK), .D(_24549_), .Q(ram_w8_l2048_id18_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40521_ ( .CLK(CLK), .D(_24548_), .Q(ram_w8_l2048_id18_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id18_0_1_wenable_reg ( .CLK(CLK), .D(_24547_), .Q(ram_w8_l2048_id18_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id18_0_cond_2_1_reg ( .CLK(CLK), .D(_tmp_447), .Q(_ram_w8_l2048_id18_0_cond_2_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40524_ ( .CLK(CLK), .D(_24555_), .Q(ram_w8_l2048_id17_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40525_ ( .CLK(CLK), .D(_24554_), .Q(ram_w8_l2048_id17_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40526_ ( .CLK(CLK), .D(_24553_), .Q(ram_w8_l2048_id17_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id17_3_1_wenable_reg ( .CLK(CLK), .D(_24552_), .Q(ram_w8_l2048_id17_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40528_ ( .CLK(CLK), .D(_24560_), .Q(ram_w8_l2048_id17_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40529_ ( .CLK(CLK), .D(_24559_), .Q(ram_w8_l2048_id17_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40530_ ( .CLK(CLK), .D(_24558_), .Q(ram_w8_l2048_id17_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id17_2_1_wenable_reg ( .CLK(CLK), .D(_24557_), .Q(ram_w8_l2048_id17_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40532_ ( .CLK(CLK), .D(_24565_), .Q(ram_w8_l2048_id17_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40533_ ( .CLK(CLK), .D(_24564_), .Q(ram_w8_l2048_id17_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40534_ ( .CLK(CLK), .D(_24563_), .Q(ram_w8_l2048_id17_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id17_1_1_wenable_reg ( .CLK(CLK), .D(_24562_), .Q(ram_w8_l2048_id17_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40536_ ( .CLK(CLK), .D(_24570_), .Q(ram_w8_l2048_id17_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40537_ ( .CLK(CLK), .D(_24569_), .Q(ram_w8_l2048_id17_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40538_ ( .CLK(CLK), .D(_24568_), .Q(ram_w8_l2048_id17_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id17_0_1_wenable_reg ( .CLK(CLK), .D(_24567_), .Q(ram_w8_l2048_id17_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id17_0_cond_2_1_reg ( .CLK(CLK), .D(_tmp_437), .Q(_ram_w8_l2048_id17_0_cond_2_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40541_ ( .CLK(CLK), .D(_24591_), .Q(ram_w8_l2048_id16_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40542_ ( .CLK(CLK), .D(_24590_), .Q(ram_w8_l2048_id16_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40543_ ( .CLK(CLK), .D(_24589_), .Q(ram_w8_l2048_id16_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id16_3_1_wenable_reg ( .CLK(CLK), .D(_24588_), .Q(ram_w8_l2048_id16_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40545_ ( .CLK(CLK), .D(_24586_), .Q(_tmp_314), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40546_ ( .CLK(CLK), .D(_24583_), .Q(_tmp_315), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_316_reg ( .CLK(CLK), .D(_24581_), .Q(_tmp_316), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40548_ ( .CLK(CLK), .D(_24579_), .Q(_tmp_317), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40549_ ( .CLK(CLK), .D(_24577_), .Q(_tmp_318), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40550_ ( .CLK(CLK), .D(_24575_), .Q(_tmp_319), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _40551_ ( .CLK(CLK), .D(_24573_), .Q(_tmp_326), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40552_ ( .CLK(CLK), .D(_24612_), .Q(ram_w8_l2048_id16_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40553_ ( .CLK(CLK), .D(_24611_), .Q(ram_w8_l2048_id16_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40554_ ( .CLK(CLK), .D(_24610_), .Q(ram_w8_l2048_id16_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id16_2_1_wenable_reg ( .CLK(CLK), .D(_24609_), .Q(ram_w8_l2048_id16_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40556_ ( .CLK(CLK), .D(_24607_), .Q(_tmp_301), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40557_ ( .CLK(CLK), .D(_24604_), .Q(_tmp_302), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_303_reg ( .CLK(CLK), .D(_24602_), .Q(_tmp_303), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40559_ ( .CLK(CLK), .D(_24600_), .Q(_tmp_304), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40560_ ( .CLK(CLK), .D(_24598_), .Q(_tmp_305), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40561_ ( .CLK(CLK), .D(_24596_), .Q(_tmp_306), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _40562_ ( .CLK(CLK), .D(_24594_), .Q(_tmp_313), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40563_ ( .CLK(CLK), .D(_24633_), .Q(ram_w8_l2048_id16_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40564_ ( .CLK(CLK), .D(_24632_), .Q(ram_w8_l2048_id16_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40565_ ( .CLK(CLK), .D(_24631_), .Q(ram_w8_l2048_id16_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id16_1_1_wenable_reg ( .CLK(CLK), .D(_24630_), .Q(ram_w8_l2048_id16_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40567_ ( .CLK(CLK), .D(_24628_), .Q(_tmp_288), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40568_ ( .CLK(CLK), .D(_24625_), .Q(_tmp_289), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_290_reg ( .CLK(CLK), .D(_24623_), .Q(_tmp_290), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40570_ ( .CLK(CLK), .D(_24621_), .Q(_tmp_291), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40571_ ( .CLK(CLK), .D(_24619_), .Q(_tmp_292), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40572_ ( .CLK(CLK), .D(_24617_), .Q(_tmp_293), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _40573_ ( .CLK(CLK), .D(_24615_), .Q(_tmp_300), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40574_ ( .CLK(CLK), .D(_24654_), .Q(ram_w8_l2048_id16_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40575_ ( .CLK(CLK), .D(_24653_), .Q(ram_w8_l2048_id16_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40576_ ( .CLK(CLK), .D(_24652_), .Q(ram_w8_l2048_id16_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id16_0_1_wenable_reg ( .CLK(CLK), .D(_24651_), .Q(ram_w8_l2048_id16_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40578_ ( .CLK(CLK), .D(_24649_), .Q(_tmp_275), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40579_ ( .CLK(CLK), .D(_24646_), .Q(_tmp_276), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_277_reg ( .CLK(CLK), .D(_24644_), .Q(_tmp_277), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40581_ ( .CLK(CLK), .D(_24642_), .Q(_tmp_278), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40582_ ( .CLK(CLK), .D(_24640_), .Q(_tmp_279), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40583_ ( .CLK(CLK), .D(_24638_), .Q(_tmp_280), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _40584_ ( .CLK(CLK), .D(_24636_), .Q(_tmp_287), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id16_0_cond_3_1_reg ( .CLK(CLK), .D(_tmp_427), .Q(_ram_w8_l2048_id16_0_cond_3_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40586_ ( .CLK(CLK), .D(_24659_), .Q(ram_w8_l2048_id15_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40587_ ( .CLK(CLK), .D(_24658_), .Q(ram_w8_l2048_id15_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40588_ ( .CLK(CLK), .D(_24657_), .Q(ram_w8_l2048_id15_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id15_3_1_wenable_reg ( .CLK(CLK), .D(_24656_), .Q(ram_w8_l2048_id15_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40590_ ( .CLK(CLK), .D(_24664_), .Q(ram_w8_l2048_id15_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40591_ ( .CLK(CLK), .D(_24663_), .Q(ram_w8_l2048_id15_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40592_ ( .CLK(CLK), .D(_24662_), .Q(ram_w8_l2048_id15_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id15_2_1_wenable_reg ( .CLK(CLK), .D(_24661_), .Q(ram_w8_l2048_id15_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40594_ ( .CLK(CLK), .D(_24669_), .Q(ram_w8_l2048_id15_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40595_ ( .CLK(CLK), .D(_24668_), .Q(ram_w8_l2048_id15_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40596_ ( .CLK(CLK), .D(_24667_), .Q(ram_w8_l2048_id15_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id15_1_1_wenable_reg ( .CLK(CLK), .D(_24666_), .Q(ram_w8_l2048_id15_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40598_ ( .CLK(CLK), .D(_24674_), .Q(ram_w8_l2048_id15_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40599_ ( .CLK(CLK), .D(_24673_), .Q(ram_w8_l2048_id15_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40600_ ( .CLK(CLK), .D(_24672_), .Q(ram_w8_l2048_id15_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id15_0_1_wenable_reg ( .CLK(CLK), .D(_24671_), .Q(ram_w8_l2048_id15_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id15_0_cond_2_1_reg ( .CLK(CLK), .D(_tmp_417), .Q(_ram_w8_l2048_id15_0_cond_2_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40603_ ( .CLK(CLK), .D(_24679_), .Q(ram_w8_l2048_id14_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40604_ ( .CLK(CLK), .D(_24678_), .Q(ram_w8_l2048_id14_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40605_ ( .CLK(CLK), .D(_24677_), .Q(ram_w8_l2048_id14_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id14_3_1_wenable_reg ( .CLK(CLK), .D(_24676_), .Q(ram_w8_l2048_id14_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40607_ ( .CLK(CLK), .D(_24684_), .Q(ram_w8_l2048_id14_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40608_ ( .CLK(CLK), .D(_24683_), .Q(ram_w8_l2048_id14_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40609_ ( .CLK(CLK), .D(_24682_), .Q(ram_w8_l2048_id14_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id14_2_1_wenable_reg ( .CLK(CLK), .D(_24681_), .Q(ram_w8_l2048_id14_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40611_ ( .CLK(CLK), .D(_24689_), .Q(ram_w8_l2048_id14_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40612_ ( .CLK(CLK), .D(_24688_), .Q(ram_w8_l2048_id14_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40613_ ( .CLK(CLK), .D(_24687_), .Q(ram_w8_l2048_id14_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id14_1_1_wenable_reg ( .CLK(CLK), .D(_24686_), .Q(ram_w8_l2048_id14_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40615_ ( .CLK(CLK), .D(_24694_), .Q(ram_w8_l2048_id14_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40616_ ( .CLK(CLK), .D(_24693_), .Q(ram_w8_l2048_id14_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40617_ ( .CLK(CLK), .D(_24692_), .Q(ram_w8_l2048_id14_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id14_0_1_wenable_reg ( .CLK(CLK), .D(_24691_), .Q(ram_w8_l2048_id14_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id14_0_cond_2_1_reg ( .CLK(CLK), .D(_tmp_407), .Q(_ram_w8_l2048_id14_0_cond_2_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40620_ ( .CLK(CLK), .D(_24715_), .Q(ram_w8_l2048_id13_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40621_ ( .CLK(CLK), .D(_24714_), .Q(ram_w8_l2048_id13_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40622_ ( .CLK(CLK), .D(_24713_), .Q(ram_w8_l2048_id13_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id13_3_1_wenable_reg ( .CLK(CLK), .D(_24712_), .Q(ram_w8_l2048_id13_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40624_ ( .CLK(CLK), .D(_24710_), .Q(_tmp_257), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40625_ ( .CLK(CLK), .D(_24707_), .Q(_tmp_258), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_259_reg ( .CLK(CLK), .D(_24705_), .Q(_tmp_259), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40627_ ( .CLK(CLK), .D(_24703_), .Q(_tmp_260), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40628_ ( .CLK(CLK), .D(_24701_), .Q(_tmp_261), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40629_ ( .CLK(CLK), .D(_24699_), .Q(_tmp_262), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _40630_ ( .CLK(CLK), .D(_24697_), .Q(_tmp_269), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40631_ ( .CLK(CLK), .D(_24736_), .Q(ram_w8_l2048_id13_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40632_ ( .CLK(CLK), .D(_24735_), .Q(ram_w8_l2048_id13_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40633_ ( .CLK(CLK), .D(_24734_), .Q(ram_w8_l2048_id13_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id13_2_1_wenable_reg ( .CLK(CLK), .D(_24733_), .Q(ram_w8_l2048_id13_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40635_ ( .CLK(CLK), .D(_24731_), .Q(_tmp_244), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40636_ ( .CLK(CLK), .D(_24728_), .Q(_tmp_245), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_246_reg ( .CLK(CLK), .D(_24726_), .Q(_tmp_246), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40638_ ( .CLK(CLK), .D(_24724_), .Q(_tmp_247), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40639_ ( .CLK(CLK), .D(_24722_), .Q(_tmp_248), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40640_ ( .CLK(CLK), .D(_24720_), .Q(_tmp_249), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _40641_ ( .CLK(CLK), .D(_24718_), .Q(_tmp_256), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40642_ ( .CLK(CLK), .D(_24757_), .Q(ram_w8_l2048_id13_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40643_ ( .CLK(CLK), .D(_24756_), .Q(ram_w8_l2048_id13_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40644_ ( .CLK(CLK), .D(_24755_), .Q(ram_w8_l2048_id13_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id13_1_1_wenable_reg ( .CLK(CLK), .D(_24754_), .Q(ram_w8_l2048_id13_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40646_ ( .CLK(CLK), .D(_24752_), .Q(_tmp_231), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40647_ ( .CLK(CLK), .D(_24749_), .Q(_tmp_232), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_233_reg ( .CLK(CLK), .D(_24747_), .Q(_tmp_233), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40649_ ( .CLK(CLK), .D(_24745_), .Q(_tmp_234), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40650_ ( .CLK(CLK), .D(_24743_), .Q(_tmp_235), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40651_ ( .CLK(CLK), .D(_24741_), .Q(_tmp_236), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _40652_ ( .CLK(CLK), .D(_24739_), .Q(_tmp_243), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40653_ ( .CLK(CLK), .D(_24778_), .Q(ram_w8_l2048_id13_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40654_ ( .CLK(CLK), .D(_24777_), .Q(ram_w8_l2048_id13_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40655_ ( .CLK(CLK), .D(_24776_), .Q(ram_w8_l2048_id13_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id13_0_1_wenable_reg ( .CLK(CLK), .D(_24775_), .Q(ram_w8_l2048_id13_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40657_ ( .CLK(CLK), .D(_24773_), .Q(_tmp_218), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40658_ ( .CLK(CLK), .D(_24770_), .Q(_tmp_219), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_220_reg ( .CLK(CLK), .D(_24768_), .Q(_tmp_220), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40660_ ( .CLK(CLK), .D(_24766_), .Q(_tmp_221), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40661_ ( .CLK(CLK), .D(_24764_), .Q(_tmp_222), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40662_ ( .CLK(CLK), .D(_24762_), .Q(_tmp_223), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _40663_ ( .CLK(CLK), .D(_24760_), .Q(_tmp_230), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id13_0_cond_3_1_reg ( .CLK(CLK), .D(_tmp_397), .Q(_ram_w8_l2048_id13_0_cond_3_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40665_ ( .CLK(CLK), .D(_24783_), .Q(ram_w8_l2048_id12_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40666_ ( .CLK(CLK), .D(_24782_), .Q(ram_w8_l2048_id12_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40667_ ( .CLK(CLK), .D(_24781_), .Q(ram_w8_l2048_id12_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id12_3_1_wenable_reg ( .CLK(CLK), .D(_24780_), .Q(ram_w8_l2048_id12_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40669_ ( .CLK(CLK), .D(_24788_), .Q(ram_w8_l2048_id12_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40670_ ( .CLK(CLK), .D(_24787_), .Q(ram_w8_l2048_id12_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40671_ ( .CLK(CLK), .D(_24786_), .Q(ram_w8_l2048_id12_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id12_2_1_wenable_reg ( .CLK(CLK), .D(_24785_), .Q(ram_w8_l2048_id12_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40673_ ( .CLK(CLK), .D(_24793_), .Q(ram_w8_l2048_id12_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40674_ ( .CLK(CLK), .D(_24792_), .Q(ram_w8_l2048_id12_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40675_ ( .CLK(CLK), .D(_24791_), .Q(ram_w8_l2048_id12_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id12_1_1_wenable_reg ( .CLK(CLK), .D(_24790_), .Q(ram_w8_l2048_id12_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40677_ ( .CLK(CLK), .D(_24798_), .Q(ram_w8_l2048_id12_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40678_ ( .CLK(CLK), .D(_24797_), .Q(ram_w8_l2048_id12_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40679_ ( .CLK(CLK), .D(_24796_), .Q(ram_w8_l2048_id12_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id12_0_1_wenable_reg ( .CLK(CLK), .D(_24795_), .Q(ram_w8_l2048_id12_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id12_0_cond_2_1_reg ( .CLK(CLK), .D(_tmp_387), .Q(_ram_w8_l2048_id12_0_cond_2_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40682_ ( .CLK(CLK), .D(_24803_), .Q(ram_w8_l2048_id11_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40683_ ( .CLK(CLK), .D(_24802_), .Q(ram_w8_l2048_id11_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40684_ ( .CLK(CLK), .D(_24801_), .Q(ram_w8_l2048_id11_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id11_3_1_wenable_reg ( .CLK(CLK), .D(_24800_), .Q(ram_w8_l2048_id11_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40686_ ( .CLK(CLK), .D(_24808_), .Q(ram_w8_l2048_id11_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40687_ ( .CLK(CLK), .D(_24807_), .Q(ram_w8_l2048_id11_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40688_ ( .CLK(CLK), .D(_24806_), .Q(ram_w8_l2048_id11_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id11_2_1_wenable_reg ( .CLK(CLK), .D(_24805_), .Q(ram_w8_l2048_id11_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40690_ ( .CLK(CLK), .D(_24813_), .Q(ram_w8_l2048_id11_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40691_ ( .CLK(CLK), .D(_24812_), .Q(ram_w8_l2048_id11_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40692_ ( .CLK(CLK), .D(_24811_), .Q(ram_w8_l2048_id11_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id11_1_1_wenable_reg ( .CLK(CLK), .D(_24810_), .Q(ram_w8_l2048_id11_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40694_ ( .CLK(CLK), .D(_24818_), .Q(ram_w8_l2048_id11_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40695_ ( .CLK(CLK), .D(_24817_), .Q(ram_w8_l2048_id11_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40696_ ( .CLK(CLK), .D(_24816_), .Q(ram_w8_l2048_id11_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id11_0_1_wenable_reg ( .CLK(CLK), .D(_24815_), .Q(ram_w8_l2048_id11_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id11_0_cond_2_1_reg ( .CLK(CLK), .D(_tmp_377), .Q(_ram_w8_l2048_id11_0_cond_2_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40699_ ( .CLK(CLK), .D(_24839_), .Q(ram_w8_l2048_id10_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40700_ ( .CLK(CLK), .D(_24838_), .Q(ram_w8_l2048_id10_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40701_ ( .CLK(CLK), .D(_24837_), .Q(ram_w8_l2048_id10_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id10_3_1_wenable_reg ( .CLK(CLK), .D(_24836_), .Q(ram_w8_l2048_id10_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40703_ ( .CLK(CLK), .D(_24834_), .Q(_tmp_200), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40704_ ( .CLK(CLK), .D(_24831_), .Q(_tmp_201), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_202_reg ( .CLK(CLK), .D(_24829_), .Q(_tmp_202), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40706_ ( .CLK(CLK), .D(_24827_), .Q(_tmp_203), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40707_ ( .CLK(CLK), .D(_24825_), .Q(_tmp_204), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40708_ ( .CLK(CLK), .D(_24823_), .Q(_tmp_205), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _40709_ ( .CLK(CLK), .D(_24821_), .Q(_tmp_212), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40710_ ( .CLK(CLK), .D(_24860_), .Q(ram_w8_l2048_id10_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40711_ ( .CLK(CLK), .D(_24859_), .Q(ram_w8_l2048_id10_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40712_ ( .CLK(CLK), .D(_24858_), .Q(ram_w8_l2048_id10_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id10_2_1_wenable_reg ( .CLK(CLK), .D(_24857_), .Q(ram_w8_l2048_id10_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40714_ ( .CLK(CLK), .D(_24855_), .Q(_tmp_187), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40715_ ( .CLK(CLK), .D(_24852_), .Q(_tmp_188), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_189_reg ( .CLK(CLK), .D(_24850_), .Q(_tmp_189), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40717_ ( .CLK(CLK), .D(_24848_), .Q(_tmp_190), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40718_ ( .CLK(CLK), .D(_24846_), .Q(_tmp_191), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40719_ ( .CLK(CLK), .D(_24844_), .Q(_tmp_192), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _40720_ ( .CLK(CLK), .D(_24842_), .Q(_tmp_199), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40721_ ( .CLK(CLK), .D(_24881_), .Q(ram_w8_l2048_id10_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40722_ ( .CLK(CLK), .D(_24880_), .Q(ram_w8_l2048_id10_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40723_ ( .CLK(CLK), .D(_24879_), .Q(ram_w8_l2048_id10_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id10_1_1_wenable_reg ( .CLK(CLK), .D(_24878_), .Q(ram_w8_l2048_id10_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40725_ ( .CLK(CLK), .D(_24876_), .Q(_tmp_174), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40726_ ( .CLK(CLK), .D(_24873_), .Q(_tmp_175), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_176_reg ( .CLK(CLK), .D(_24871_), .Q(_tmp_176), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40728_ ( .CLK(CLK), .D(_24869_), .Q(_tmp_177), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40729_ ( .CLK(CLK), .D(_24867_), .Q(_tmp_178), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40730_ ( .CLK(CLK), .D(_24865_), .Q(_tmp_179), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _40731_ ( .CLK(CLK), .D(_24863_), .Q(_tmp_186), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40732_ ( .CLK(CLK), .D(_24902_), .Q(ram_w8_l2048_id10_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40733_ ( .CLK(CLK), .D(_24901_), .Q(ram_w8_l2048_id10_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40734_ ( .CLK(CLK), .D(_24900_), .Q(ram_w8_l2048_id10_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id10_0_1_wenable_reg ( .CLK(CLK), .D(_24899_), .Q(ram_w8_l2048_id10_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40736_ ( .CLK(CLK), .D(_24897_), .Q(_tmp_161), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40737_ ( .CLK(CLK), .D(_24894_), .Q(_tmp_162), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_163_reg ( .CLK(CLK), .D(_24892_), .Q(_tmp_163), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40739_ ( .CLK(CLK), .D(_24890_), .Q(_tmp_164), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40740_ ( .CLK(CLK), .D(_24888_), .Q(_tmp_165), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40741_ ( .CLK(CLK), .D(_24886_), .Q(_tmp_166), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(2), .SRST_POLARITY(1'h1), .SRST_VALUE(2'h0) ) _40742_ ( .CLK(CLK), .D(_24884_), .Q(_tmp_173), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id10_0_cond_3_1_reg ( .CLK(CLK), .D(_tmp_367), .Q(_ram_w8_l2048_id10_0_cond_3_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40744_ ( .CLK(CLK), .D(_24907_), .Q(ram_w8_l2048_id9_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40745_ ( .CLK(CLK), .D(_24906_), .Q(ram_w8_l2048_id9_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40746_ ( .CLK(CLK), .D(_24905_), .Q(ram_w8_l2048_id9_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id9_3_1_wenable_reg ( .CLK(CLK), .D(_24904_), .Q(ram_w8_l2048_id9_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40748_ ( .CLK(CLK), .D(_24912_), .Q(ram_w8_l2048_id9_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40749_ ( .CLK(CLK), .D(_24911_), .Q(ram_w8_l2048_id9_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40750_ ( .CLK(CLK), .D(_24910_), .Q(ram_w8_l2048_id9_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id9_2_1_wenable_reg ( .CLK(CLK), .D(_24909_), .Q(ram_w8_l2048_id9_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id9_2_cond_0_1_reg ( .CLK(CLK), .D(1'h1), .Q(_ram_w8_l2048_id9_2_cond_0_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40753_ ( .CLK(CLK), .D(_24917_), .Q(ram_w8_l2048_id9_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40754_ ( .CLK(CLK), .D(_24916_), .Q(ram_w8_l2048_id9_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40755_ ( .CLK(CLK), .D(_24915_), .Q(ram_w8_l2048_id9_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id9_1_1_wenable_reg ( .CLK(CLK), .D(_24914_), .Q(ram_w8_l2048_id9_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40757_ ( .CLK(CLK), .D(_24922_), .Q(ram_w8_l2048_id9_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40758_ ( .CLK(CLK), .D(_24921_), .Q(ram_w8_l2048_id9_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40759_ ( .CLK(CLK), .D(_24920_), .Q(ram_w8_l2048_id9_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id9_0_1_wenable_reg ( .CLK(CLK), .D(_24919_), .Q(ram_w8_l2048_id9_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id9_0_cond_1_1_reg ( .CLK(CLK), .D(_tmp_537), .Q(_ram_w8_l2048_id9_0_cond_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40762_ ( .CLK(CLK), .D(_24927_), .Q(ram_w8_l2048_id8_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40763_ ( .CLK(CLK), .D(_24926_), .Q(ram_w8_l2048_id8_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40764_ ( .CLK(CLK), .D(_24925_), .Q(ram_w8_l2048_id8_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id8_3_1_wenable_reg ( .CLK(CLK), .D(_24924_), .Q(ram_w8_l2048_id8_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id8_3_cond_1_1_reg ( .CLK(CLK), .D(_tmp_527), .Q(_ram_w8_l2048_id8_3_cond_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40767_ ( .CLK(CLK), .D(_24932_), .Q(ram_w8_l2048_id8_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40768_ ( .CLK(CLK), .D(_24931_), .Q(ram_w8_l2048_id8_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40769_ ( .CLK(CLK), .D(_24930_), .Q(ram_w8_l2048_id8_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id8_2_1_wenable_reg ( .CLK(CLK), .D(_24929_), .Q(ram_w8_l2048_id8_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40771_ ( .CLK(CLK), .D(_24937_), .Q(ram_w8_l2048_id8_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40772_ ( .CLK(CLK), .D(_24936_), .Q(ram_w8_l2048_id8_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40773_ ( .CLK(CLK), .D(_24935_), .Q(ram_w8_l2048_id8_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id8_1_1_wenable_reg ( .CLK(CLK), .D(_24934_), .Q(ram_w8_l2048_id8_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40775_ ( .CLK(CLK), .D(_24942_), .Q(ram_w8_l2048_id8_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40776_ ( .CLK(CLK), .D(_24941_), .Q(ram_w8_l2048_id8_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40777_ ( .CLK(CLK), .D(_24940_), .Q(ram_w8_l2048_id8_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id8_0_1_wenable_reg ( .CLK(CLK), .D(_24939_), .Q(ram_w8_l2048_id8_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40779_ ( .CLK(CLK), .D(_24947_), .Q(ram_w8_l2048_id7_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40780_ ( .CLK(CLK), .D(_24946_), .Q(ram_w8_l2048_id7_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40781_ ( .CLK(CLK), .D(_24945_), .Q(ram_w8_l2048_id7_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id7_3_1_wenable_reg ( .CLK(CLK), .D(_24944_), .Q(ram_w8_l2048_id7_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id7_3_cond_1_1_reg ( .CLK(CLK), .D(_tmp_517), .Q(_ram_w8_l2048_id7_3_cond_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40784_ ( .CLK(CLK), .D(_24952_), .Q(ram_w8_l2048_id7_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40785_ ( .CLK(CLK), .D(_24951_), .Q(ram_w8_l2048_id7_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40786_ ( .CLK(CLK), .D(_24950_), .Q(ram_w8_l2048_id7_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id7_2_1_wenable_reg ( .CLK(CLK), .D(_24949_), .Q(ram_w8_l2048_id7_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40788_ ( .CLK(CLK), .D(_24957_), .Q(ram_w8_l2048_id7_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40789_ ( .CLK(CLK), .D(_24956_), .Q(ram_w8_l2048_id7_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40790_ ( .CLK(CLK), .D(_24955_), .Q(ram_w8_l2048_id7_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id7_1_1_wenable_reg ( .CLK(CLK), .D(_24954_), .Q(ram_w8_l2048_id7_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40792_ ( .CLK(CLK), .D(_24962_), .Q(ram_w8_l2048_id7_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40793_ ( .CLK(CLK), .D(_24961_), .Q(ram_w8_l2048_id7_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40794_ ( .CLK(CLK), .D(_24960_), .Q(ram_w8_l2048_id7_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id7_0_1_wenable_reg ( .CLK(CLK), .D(_24959_), .Q(ram_w8_l2048_id7_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40796_ ( .CLK(CLK), .D(_24967_), .Q(ram_w8_l2048_id6_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40797_ ( .CLK(CLK), .D(_24966_), .Q(ram_w8_l2048_id6_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40798_ ( .CLK(CLK), .D(_24965_), .Q(ram_w8_l2048_id6_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id6_3_1_wenable_reg ( .CLK(CLK), .D(_24964_), .Q(ram_w8_l2048_id6_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id6_3_cond_1_1_reg ( .CLK(CLK), .D(_tmp_507), .Q(_ram_w8_l2048_id6_3_cond_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40801_ ( .CLK(CLK), .D(_24972_), .Q(ram_w8_l2048_id6_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40802_ ( .CLK(CLK), .D(_24971_), .Q(ram_w8_l2048_id6_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40803_ ( .CLK(CLK), .D(_24970_), .Q(ram_w8_l2048_id6_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id6_2_1_wenable_reg ( .CLK(CLK), .D(_24969_), .Q(ram_w8_l2048_id6_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40805_ ( .CLK(CLK), .D(_24977_), .Q(ram_w8_l2048_id6_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40806_ ( .CLK(CLK), .D(_24976_), .Q(ram_w8_l2048_id6_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40807_ ( .CLK(CLK), .D(_24975_), .Q(ram_w8_l2048_id6_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id6_1_1_wenable_reg ( .CLK(CLK), .D(_24974_), .Q(ram_w8_l2048_id6_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40809_ ( .CLK(CLK), .D(_24982_), .Q(ram_w8_l2048_id6_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40810_ ( .CLK(CLK), .D(_24981_), .Q(ram_w8_l2048_id6_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40811_ ( .CLK(CLK), .D(_24980_), .Q(ram_w8_l2048_id6_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id6_0_1_wenable_reg ( .CLK(CLK), .D(_24979_), .Q(ram_w8_l2048_id6_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40813_ ( .CLK(CLK), .D(_24987_), .Q(ram_w8_l2048_id5_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40814_ ( .CLK(CLK), .D(_24986_), .Q(ram_w8_l2048_id5_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40815_ ( .CLK(CLK), .D(_24985_), .Q(ram_w8_l2048_id5_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id5_3_1_wenable_reg ( .CLK(CLK), .D(_24984_), .Q(ram_w8_l2048_id5_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id5_3_cond_1_1_reg ( .CLK(CLK), .D(_tmp_497), .Q(_ram_w8_l2048_id5_3_cond_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40818_ ( .CLK(CLK), .D(_24992_), .Q(ram_w8_l2048_id5_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40819_ ( .CLK(CLK), .D(_24991_), .Q(ram_w8_l2048_id5_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40820_ ( .CLK(CLK), .D(_24990_), .Q(ram_w8_l2048_id5_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id5_2_1_wenable_reg ( .CLK(CLK), .D(_24989_), .Q(ram_w8_l2048_id5_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40822_ ( .CLK(CLK), .D(_24997_), .Q(ram_w8_l2048_id5_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40823_ ( .CLK(CLK), .D(_24996_), .Q(ram_w8_l2048_id5_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40824_ ( .CLK(CLK), .D(_24995_), .Q(ram_w8_l2048_id5_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id5_1_1_wenable_reg ( .CLK(CLK), .D(_24994_), .Q(ram_w8_l2048_id5_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40826_ ( .CLK(CLK), .D(_25002_), .Q(ram_w8_l2048_id5_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40827_ ( .CLK(CLK), .D(_25001_), .Q(ram_w8_l2048_id5_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40828_ ( .CLK(CLK), .D(_25000_), .Q(ram_w8_l2048_id5_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id5_0_1_wenable_reg ( .CLK(CLK), .D(_24999_), .Q(ram_w8_l2048_id5_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40830_ ( .CLK(CLK), .D(_25007_), .Q(ram_w8_l2048_id4_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40831_ ( .CLK(CLK), .D(_25006_), .Q(ram_w8_l2048_id4_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40832_ ( .CLK(CLK), .D(_25005_), .Q(ram_w8_l2048_id4_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id4_3_1_wenable_reg ( .CLK(CLK), .D(_25004_), .Q(ram_w8_l2048_id4_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id4_3_cond_1_1_reg ( .CLK(CLK), .D(_tmp_487), .Q(_ram_w8_l2048_id4_3_cond_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40835_ ( .CLK(CLK), .D(_25012_), .Q(ram_w8_l2048_id4_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40836_ ( .CLK(CLK), .D(_25011_), .Q(ram_w8_l2048_id4_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40837_ ( .CLK(CLK), .D(_25010_), .Q(ram_w8_l2048_id4_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id4_2_1_wenable_reg ( .CLK(CLK), .D(_25009_), .Q(ram_w8_l2048_id4_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40839_ ( .CLK(CLK), .D(_25017_), .Q(ram_w8_l2048_id4_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40840_ ( .CLK(CLK), .D(_25016_), .Q(ram_w8_l2048_id4_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40841_ ( .CLK(CLK), .D(_25015_), .Q(ram_w8_l2048_id4_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id4_1_1_wenable_reg ( .CLK(CLK), .D(_25014_), .Q(ram_w8_l2048_id4_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40843_ ( .CLK(CLK), .D(_25022_), .Q(ram_w8_l2048_id4_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40844_ ( .CLK(CLK), .D(_25021_), .Q(ram_w8_l2048_id4_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40845_ ( .CLK(CLK), .D(_25020_), .Q(ram_w8_l2048_id4_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id4_0_1_wenable_reg ( .CLK(CLK), .D(_25019_), .Q(ram_w8_l2048_id4_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40847_ ( .CLK(CLK), .D(_25027_), .Q(ram_w8_l2048_id3_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40848_ ( .CLK(CLK), .D(_25026_), .Q(ram_w8_l2048_id3_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40849_ ( .CLK(CLK), .D(_25025_), .Q(ram_w8_l2048_id3_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id3_3_1_wenable_reg ( .CLK(CLK), .D(_25024_), .Q(ram_w8_l2048_id3_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id3_3_cond_1_1_reg ( .CLK(CLK), .D(_tmp_477), .Q(_ram_w8_l2048_id3_3_cond_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40852_ ( .CLK(CLK), .D(_25032_), .Q(ram_w8_l2048_id3_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40853_ ( .CLK(CLK), .D(_25031_), .Q(ram_w8_l2048_id3_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40854_ ( .CLK(CLK), .D(_25030_), .Q(ram_w8_l2048_id3_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id3_2_1_wenable_reg ( .CLK(CLK), .D(_25029_), .Q(ram_w8_l2048_id3_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40856_ ( .CLK(CLK), .D(_25037_), .Q(ram_w8_l2048_id3_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40857_ ( .CLK(CLK), .D(_25036_), .Q(ram_w8_l2048_id3_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40858_ ( .CLK(CLK), .D(_25035_), .Q(ram_w8_l2048_id3_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id3_1_1_wenable_reg ( .CLK(CLK), .D(_25034_), .Q(ram_w8_l2048_id3_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40860_ ( .CLK(CLK), .D(_25042_), .Q(ram_w8_l2048_id3_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40861_ ( .CLK(CLK), .D(_25041_), .Q(ram_w8_l2048_id3_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40862_ ( .CLK(CLK), .D(_25040_), .Q(ram_w8_l2048_id3_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id3_0_1_wenable_reg ( .CLK(CLK), .D(_25039_), .Q(ram_w8_l2048_id3_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40864_ ( .CLK(CLK), .D(_25056_), .Q(ram_w8_l2048_id2_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40865_ ( .CLK(CLK), .D(_25054_), .Q(ram_w8_l2048_id2_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40866_ ( .CLK(CLK), .D(_25051_), .Q(ram_w8_l2048_id2_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id2_3_1_wenable_reg ( .CLK(CLK), .D(_25049_), .Q(ram_w8_l2048_id2_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id2_3_cond_1_1_reg ( .CLK(CLK), .D(_tmp_467), .Q(_ram_w8_l2048_id2_3_cond_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40869_ ( .CLK(CLK), .D(_25046_), .Q(_tmp_981), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_982_reg ( .CLK(CLK), .D(_25044_), .Q(_tmp_982), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id2_3_cond_4_1_reg ( .CLK(CLK), .D(_tmp_1023), .Q(_ram_w8_l2048_id2_3_cond_4_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40872_ ( .CLK(CLK), .D(_25070_), .Q(ram_w8_l2048_id2_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40873_ ( .CLK(CLK), .D(_25068_), .Q(ram_w8_l2048_id2_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40874_ ( .CLK(CLK), .D(_25065_), .Q(ram_w8_l2048_id2_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id2_2_1_wenable_reg ( .CLK(CLK), .D(_25063_), .Q(ram_w8_l2048_id2_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40876_ ( .CLK(CLK), .D(_25060_), .Q(_tmp_979), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_980_reg ( .CLK(CLK), .D(_25058_), .Q(_tmp_980), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40878_ ( .CLK(CLK), .D(_25084_), .Q(ram_w8_l2048_id2_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40879_ ( .CLK(CLK), .D(_25082_), .Q(ram_w8_l2048_id2_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40880_ ( .CLK(CLK), .D(_25079_), .Q(ram_w8_l2048_id2_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id2_1_1_wenable_reg ( .CLK(CLK), .D(_25077_), .Q(ram_w8_l2048_id2_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40882_ ( .CLK(CLK), .D(_25074_), .Q(_tmp_977), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_978_reg ( .CLK(CLK), .D(_25072_), .Q(_tmp_978), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40884_ ( .CLK(CLK), .D(_25098_), .Q(ram_w8_l2048_id2_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40885_ ( .CLK(CLK), .D(_25096_), .Q(ram_w8_l2048_id2_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40886_ ( .CLK(CLK), .D(_25093_), .Q(ram_w8_l2048_id2_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id2_0_1_wenable_reg ( .CLK(CLK), .D(_25091_), .Q(ram_w8_l2048_id2_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40888_ ( .CLK(CLK), .D(_25088_), .Q(_tmp_975), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_976_reg ( .CLK(CLK), .D(_25086_), .Q(_tmp_976), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40890_ ( .CLK(CLK), .D(_25161_), .Q(ram_w8_l2048_id1_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40891_ ( .CLK(CLK), .D(_25158_), .Q(ram_w8_l2048_id1_3_0_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id1_3_0_wenable_reg ( .CLK(CLK), .D(_25157_), .Q(ram_w8_l2048_id1_3_0_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40893_ ( .CLK(CLK), .D(_25155_), .Q(ram_w8_l2048_id1_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40894_ ( .CLK(CLK), .D(_25150_), .Q(ram_w8_l2048_id1_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id1_3_1_wenable_reg ( .CLK(CLK), .D(_25148_), .Q(ram_w8_l2048_id1_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40896_ ( .CLK(CLK), .D(_25145_), .Q(_tmp_125), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40897_ ( .CLK(CLK), .D(_25142_), .Q(_tmp_126), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_127_reg ( .CLK(CLK), .D(_25140_), .Q(_tmp_127), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40899_ ( .CLK(CLK), .D(_25138_), .Q(_tmp_128), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40900_ ( .CLK(CLK), .D(_25136_), .Q(_tmp_129), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40901_ ( .CLK(CLK), .D(_25134_), .Q(_tmp_130), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40902_ ( .CLK(CLK), .D(_25132_), .Q(_tmp_131), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40903_ ( .CLK(CLK), .D(_25130_), .Q(_tmp_132), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40904_ ( .CLK(CLK), .D(_25128_), .Q(_tmp_133), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40905_ ( .CLK(CLK), .D(_25126_), .Q(_tmp_134), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40906_ ( .CLK(CLK), .D(_25124_), .Q(_tmp_135), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40907_ ( .CLK(CLK), .D(_25122_), .Q(_tmp_136), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40908_ ( .CLK(CLK), .D(_25120_), .Q(_tmp_155), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id1_3_cond_2_1_reg ( .CLK(CLK), .D(_tmp_457), .Q(_ram_w8_l2048_id1_3_cond_2_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40910_ ( .CLK(CLK), .D(_25117_), .Q(_tmp_859), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_860_reg ( .CLK(CLK), .D(_25115_), .Q(_tmp_860), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id1_3_cond_5_1_reg ( .CLK(CLK), .D(_tmp_873), .Q(_ram_w8_l2048_id1_3_cond_5_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id1_3_cond_7_1_reg ( .CLK(CLK), .D(_05542_), .Q(_ram_w8_l2048_id1_3_cond_7_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1155_reg ( .CLK(CLK), .D(_25113_), .Q(_tmp_1155), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1160_1_reg ( .CLK(CLK), .D(_tmp_1160), .Q(__tmp_1160_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40916_ ( .CLK(CLK), .D(_tmp_1161), .Q(__tmp_1161_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1162_reg ( .CLK(CLK), .D(_25111_), .Q(_tmp_1162), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1163_reg ( .CLK(CLK), .D(_25108_), .Q(_tmp_1163), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1164_reg ( .CLK(CLK), .D(_25106_), .Q(_tmp_1164), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1165_reg ( .CLK(CLK), .D(_25102_), .Q(_tmp_1165), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40921_ ( .CLK(CLK), .D(_25100_), .Q(_tmp_1166), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40922_ ( .CLK(CLK), .D(_25224_), .Q(ram_w8_l2048_id1_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40923_ ( .CLK(CLK), .D(_25221_), .Q(ram_w8_l2048_id1_2_0_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id1_2_0_wenable_reg ( .CLK(CLK), .D(_25220_), .Q(ram_w8_l2048_id1_2_0_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40925_ ( .CLK(CLK), .D(_25218_), .Q(ram_w8_l2048_id1_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40926_ ( .CLK(CLK), .D(_25213_), .Q(ram_w8_l2048_id1_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id1_2_1_wenable_reg ( .CLK(CLK), .D(_25211_), .Q(ram_w8_l2048_id1_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40928_ ( .CLK(CLK), .D(_25208_), .Q(_tmp_94), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40929_ ( .CLK(CLK), .D(_25205_), .Q(_tmp_95), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_96_reg ( .CLK(CLK), .D(_25203_), .Q(_tmp_96), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40931_ ( .CLK(CLK), .D(_25201_), .Q(_tmp_97), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40932_ ( .CLK(CLK), .D(_25199_), .Q(_tmp_98), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40933_ ( .CLK(CLK), .D(_25197_), .Q(_tmp_99), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40934_ ( .CLK(CLK), .D(_25195_), .Q(_tmp_100), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40935_ ( .CLK(CLK), .D(_25193_), .Q(_tmp_101), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40936_ ( .CLK(CLK), .D(_25191_), .Q(_tmp_102), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40937_ ( .CLK(CLK), .D(_25189_), .Q(_tmp_103), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40938_ ( .CLK(CLK), .D(_25187_), .Q(_tmp_104), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40939_ ( .CLK(CLK), .D(_25185_), .Q(_tmp_105), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40940_ ( .CLK(CLK), .D(_25183_), .Q(_tmp_124), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40941_ ( .CLK(CLK), .D(_25180_), .Q(_tmp_857), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_858_reg ( .CLK(CLK), .D(_25178_), .Q(_tmp_858), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id1_2_cond_7_1_reg ( .CLK(CLK), .D(_05521_), .Q(_ram_w8_l2048_id1_2_cond_7_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1143_reg ( .CLK(CLK), .D(_25176_), .Q(_tmp_1143), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1148_1_reg ( .CLK(CLK), .D(_tmp_1148), .Q(__tmp_1148_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40946_ ( .CLK(CLK), .D(_tmp_1149), .Q(__tmp_1149_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1150_reg ( .CLK(CLK), .D(_25174_), .Q(_tmp_1150), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1151_reg ( .CLK(CLK), .D(_25171_), .Q(_tmp_1151), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1152_reg ( .CLK(CLK), .D(_25169_), .Q(_tmp_1152), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1153_reg ( .CLK(CLK), .D(_25165_), .Q(_tmp_1153), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40951_ ( .CLK(CLK), .D(_25163_), .Q(_tmp_1154), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40952_ ( .CLK(CLK), .D(_25287_), .Q(ram_w8_l2048_id1_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40953_ ( .CLK(CLK), .D(_25284_), .Q(ram_w8_l2048_id1_1_0_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id1_1_0_wenable_reg ( .CLK(CLK), .D(_25283_), .Q(ram_w8_l2048_id1_1_0_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40955_ ( .CLK(CLK), .D(_25281_), .Q(ram_w8_l2048_id1_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40956_ ( .CLK(CLK), .D(_25276_), .Q(ram_w8_l2048_id1_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id1_1_1_wenable_reg ( .CLK(CLK), .D(_25274_), .Q(ram_w8_l2048_id1_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40958_ ( .CLK(CLK), .D(_25271_), .Q(_tmp_63), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40959_ ( .CLK(CLK), .D(_25268_), .Q(_tmp_64), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_65_reg ( .CLK(CLK), .D(_25266_), .Q(_tmp_65), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40961_ ( .CLK(CLK), .D(_25264_), .Q(_tmp_66), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40962_ ( .CLK(CLK), .D(_25262_), .Q(_tmp_67), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40963_ ( .CLK(CLK), .D(_25260_), .Q(_tmp_68), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40964_ ( .CLK(CLK), .D(_25258_), .Q(_tmp_69), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40965_ ( .CLK(CLK), .D(_25256_), .Q(_tmp_70), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40966_ ( .CLK(CLK), .D(_25254_), .Q(_tmp_71), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40967_ ( .CLK(CLK), .D(_25252_), .Q(_tmp_72), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40968_ ( .CLK(CLK), .D(_25250_), .Q(_tmp_73), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40969_ ( .CLK(CLK), .D(_25248_), .Q(_tmp_74), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _40970_ ( .CLK(CLK), .D(_25246_), .Q(_tmp_93), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40971_ ( .CLK(CLK), .D(_25243_), .Q(_tmp_855), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_856_reg ( .CLK(CLK), .D(_25241_), .Q(_tmp_856), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id1_1_cond_7_1_reg ( .CLK(CLK), .D(_05500_), .Q(_ram_w8_l2048_id1_1_cond_7_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1131_reg ( .CLK(CLK), .D(_25239_), .Q(_tmp_1131), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1136_1_reg ( .CLK(CLK), .D(_tmp_1136), .Q(__tmp_1136_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40976_ ( .CLK(CLK), .D(_tmp_1137), .Q(__tmp_1137_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1138_reg ( .CLK(CLK), .D(_25237_), .Q(_tmp_1138), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1139_reg ( .CLK(CLK), .D(_25234_), .Q(_tmp_1139), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1140_reg ( .CLK(CLK), .D(_25232_), .Q(_tmp_1140), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1141_reg ( .CLK(CLK), .D(_25228_), .Q(_tmp_1141), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40981_ ( .CLK(CLK), .D(_25226_), .Q(_tmp_1142), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _40982_ ( .CLK(CLK), .D(_25290_), .Q(_dataflow_cat_data_131), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_cat_valid_131_reg ( .CLK(CLK), .D(_25289_), .Q(_dataflow_cat_valid_131), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40984_ ( .CLK(CLK), .D(_25353_), .Q(ram_w8_l2048_id1_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40985_ ( .CLK(CLK), .D(_25350_), .Q(ram_w8_l2048_id1_0_0_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id1_0_0_wenable_reg ( .CLK(CLK), .D(_25349_), .Q(ram_w8_l2048_id1_0_0_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40987_ ( .CLK(CLK), .D(_25347_), .Q(ram_w8_l2048_id1_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _40988_ ( .CLK(CLK), .D(_25342_), .Q(ram_w8_l2048_id1_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id1_0_1_wenable_reg ( .CLK(CLK), .D(_25340_), .Q(ram_w8_l2048_id1_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _40990_ ( .CLK(CLK), .D(_25337_), .Q(_tmp_32), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _40991_ ( .CLK(CLK), .D(_25334_), .Q(_tmp_33), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_34_reg ( .CLK(CLK), .D(_25332_), .Q(_tmp_34), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40993_ ( .CLK(CLK), .D(_25330_), .Q(_tmp_35), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40994_ ( .CLK(CLK), .D(_25328_), .Q(_tmp_36), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40995_ ( .CLK(CLK), .D(_25326_), .Q(_tmp_37), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40996_ ( .CLK(CLK), .D(_25324_), .Q(_tmp_38), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40997_ ( .CLK(CLK), .D(_25322_), .Q(_tmp_39), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40998_ ( .CLK(CLK), .D(_25320_), .Q(_tmp_40), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _40999_ ( .CLK(CLK), .D(_25318_), .Q(_tmp_41), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _41000_ ( .CLK(CLK), .D(_25316_), .Q(_tmp_42), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _41001_ ( .CLK(CLK), .D(_25314_), .Q(_tmp_43), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _41002_ ( .CLK(CLK), .D(_25312_), .Q(_tmp_62), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41003_ ( .CLK(CLK), .D(_25309_), .Q(_tmp_853), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_854_reg ( .CLK(CLK), .D(_25307_), .Q(_tmp_854), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id1_0_cond_7_1_reg ( .CLK(CLK), .D(_05476_), .Q(_ram_w8_l2048_id1_0_cond_7_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1119_reg ( .CLK(CLK), .D(_25305_), .Q(_tmp_1119), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_1124_1_reg ( .CLK(CLK), .D(_tmp_1124), .Q(__tmp_1124_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41008_ ( .CLK(CLK), .D(_tmp_1125), .Q(__tmp_1125_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1126_reg ( .CLK(CLK), .D(_25303_), .Q(_tmp_1126), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1127_reg ( .CLK(CLK), .D(_25300_), .Q(_tmp_1127), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1128_reg ( .CLK(CLK), .D(_25298_), .Q(_tmp_1128), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1129_reg ( .CLK(CLK), .D(_25294_), .Q(_tmp_1129), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41013_ ( .CLK(CLK), .D(_25292_), .Q(_tmp_1130), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _41014_ ( .CLK(CLK), .D(_25385_), .Q(ram_w8_l2048_id0_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41015_ ( .CLK(CLK), .D(_25382_), .Q(ram_w8_l2048_id0_3_0_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id0_3_0_wenable_reg ( .CLK(CLK), .D(_25381_), .Q(ram_w8_l2048_id0_3_0_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _41017_ ( .CLK(CLK), .D(_25379_), .Q(ram_w8_l2048_id0_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41018_ ( .CLK(CLK), .D(_25375_), .Q(ram_w8_l2048_id0_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id0_3_1_wenable_reg ( .CLK(CLK), .D(_25374_), .Q(ram_w8_l2048_id0_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41020_ ( .CLK(CLK), .D(_25372_), .Q(_tmp_25), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_26_reg ( .CLK(CLK), .D(_25370_), .Q(_tmp_26), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id0_3_cond_1_1_reg ( .CLK(CLK), .D(_tmp_347), .Q(_ram_w8_l2048_id0_3_cond_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id0_3_cond_3_1_reg ( .CLK(CLK), .D(_05453_), .Q(_ram_w8_l2048_id0_3_cond_3_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_946_reg ( .CLK(CLK), .D(_25368_), .Q(_tmp_946), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_951_1_reg ( .CLK(CLK), .D(_tmp_951), .Q(__tmp_951_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41026_ ( .CLK(CLK), .D(_tmp_952), .Q(__tmp_952_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_953_reg ( .CLK(CLK), .D(_25366_), .Q(_tmp_953), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_954_reg ( .CLK(CLK), .D(_25363_), .Q(_tmp_954), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_955_reg ( .CLK(CLK), .D(_25361_), .Q(_tmp_955), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_956_reg ( .CLK(CLK), .D(_25357_), .Q(_tmp_956), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41031_ ( .CLK(CLK), .D(_25355_), .Q(_tmp_957), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id0_3_cond_4_1_reg ( .CLK(CLK), .D(_tmp_1003), .Q(_ram_w8_l2048_id0_3_cond_4_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _41033_ ( .CLK(CLK), .D(_25417_), .Q(ram_w8_l2048_id0_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41034_ ( .CLK(CLK), .D(_25414_), .Q(ram_w8_l2048_id0_2_0_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id0_2_0_wenable_reg ( .CLK(CLK), .D(_25413_), .Q(ram_w8_l2048_id0_2_0_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _41036_ ( .CLK(CLK), .D(_25411_), .Q(ram_w8_l2048_id0_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41037_ ( .CLK(CLK), .D(_25407_), .Q(ram_w8_l2048_id0_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id0_2_1_wenable_reg ( .CLK(CLK), .D(_25406_), .Q(ram_w8_l2048_id0_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41039_ ( .CLK(CLK), .D(_25404_), .Q(_tmp_23), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_24_reg ( .CLK(CLK), .D(_25402_), .Q(_tmp_24), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id0_2_cond_3_1_reg ( .CLK(CLK), .D(_05445_), .Q(_ram_w8_l2048_id0_2_cond_3_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_934_reg ( .CLK(CLK), .D(_25400_), .Q(_tmp_934), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_939_1_reg ( .CLK(CLK), .D(_tmp_939), .Q(__tmp_939_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41044_ ( .CLK(CLK), .D(_tmp_940), .Q(__tmp_940_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_941_reg ( .CLK(CLK), .D(_25398_), .Q(_tmp_941), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_942_reg ( .CLK(CLK), .D(_25395_), .Q(_tmp_942), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_943_reg ( .CLK(CLK), .D(_25393_), .Q(_tmp_943), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_944_reg ( .CLK(CLK), .D(_25389_), .Q(_tmp_944), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41049_ ( .CLK(CLK), .D(_25387_), .Q(_tmp_945), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _41050_ ( .CLK(CLK), .D(_25449_), .Q(ram_w8_l2048_id0_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41051_ ( .CLK(CLK), .D(_25446_), .Q(ram_w8_l2048_id0_1_0_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id0_1_0_wenable_reg ( .CLK(CLK), .D(_25445_), .Q(ram_w8_l2048_id0_1_0_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _41053_ ( .CLK(CLK), .D(_25443_), .Q(ram_w8_l2048_id0_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41054_ ( .CLK(CLK), .D(_25439_), .Q(ram_w8_l2048_id0_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id0_1_1_wenable_reg ( .CLK(CLK), .D(_25438_), .Q(ram_w8_l2048_id0_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41056_ ( .CLK(CLK), .D(_25436_), .Q(_tmp_21), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_22_reg ( .CLK(CLK), .D(_25434_), .Q(_tmp_22), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id0_1_cond_3_1_reg ( .CLK(CLK), .D(_05437_), .Q(_ram_w8_l2048_id0_1_cond_3_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_922_reg ( .CLK(CLK), .D(_25432_), .Q(_tmp_922), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_927_1_reg ( .CLK(CLK), .D(_tmp_927), .Q(__tmp_927_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41061_ ( .CLK(CLK), .D(_tmp_928), .Q(__tmp_928_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_929_reg ( .CLK(CLK), .D(_25430_), .Q(_tmp_929), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_930_reg ( .CLK(CLK), .D(_25427_), .Q(_tmp_930), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_931_reg ( .CLK(CLK), .D(_25425_), .Q(_tmp_931), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_932_reg ( .CLK(CLK), .D(_25421_), .Q(_tmp_932), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41066_ ( .CLK(CLK), .D(_25419_), .Q(_tmp_933), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41067_ ( .CLK(CLK), .D(_25452_), .Q(_dataflow_cat_data_96), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_cat_valid_96_reg ( .CLK(CLK), .D(_25451_), .Q(_dataflow_cat_valid_96), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _41069_ ( .CLK(CLK), .D(_25484_), .Q(ram_w8_l2048_id0_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41070_ ( .CLK(CLK), .D(_25481_), .Q(ram_w8_l2048_id0_0_0_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id0_0_0_wenable_reg ( .CLK(CLK), .D(_25480_), .Q(ram_w8_l2048_id0_0_0_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _41072_ ( .CLK(CLK), .D(_25478_), .Q(ram_w8_l2048_id0_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41073_ ( .CLK(CLK), .D(_25474_), .Q(ram_w8_l2048_id0_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l2048_id0_0_1_wenable_reg ( .CLK(CLK), .D(_25473_), .Q(ram_w8_l2048_id0_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41075_ ( .CLK(CLK), .D(_25471_), .Q(_tmp_19), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_20_reg ( .CLK(CLK), .D(_25469_), .Q(_tmp_20), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l2048_id0_0_cond_3_1_reg ( .CLK(CLK), .D(_05426_), .Q(_ram_w8_l2048_id0_0_cond_3_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_910_reg ( .CLK(CLK), .D(_25467_), .Q(_tmp_910), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) __tmp_915_1_reg ( .CLK(CLK), .D(_tmp_915), .Q(__tmp_915_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41080_ ( .CLK(CLK), .D(_tmp_916), .Q(__tmp_916_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_917_reg ( .CLK(CLK), .D(_25465_), .Q(_tmp_917), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_918_reg ( .CLK(CLK), .D(_25462_), .Q(_tmp_918), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_919_reg ( .CLK(CLK), .D(_25460_), .Q(_tmp_919), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_920_reg ( .CLK(CLK), .D(_25456_), .Q(_tmp_920), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41085_ ( .CLK(CLK), .D(_25454_), .Q(_tmp_921), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _41086_ ( .CLK(CLK), .D(_25494_), .Q(ram_w8_l4096_id0_3_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _41087_ ( .CLK(CLK), .D(_25493_), .Q(ram_w8_l4096_id0_3_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41088_ ( .CLK(CLK), .D(_25491_), .Q(ram_w8_l4096_id0_3_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l4096_id0_3_1_wenable_reg ( .CLK(CLK), .D(_25490_), .Q(ram_w8_l4096_id0_3_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41090_ ( .CLK(CLK), .D(_25488_), .Q(_tmp_970), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_971_reg ( .CLK(CLK), .D(_25486_), .Q(_tmp_971), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _ram_w8_l4096_id0_3_cond_1_1_reg ( .CLK(CLK), .D(_tmp_1033), .Q(_ram_w8_l4096_id0_3_cond_1_1), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _41093_ ( .CLK(CLK), .D(_25504_), .Q(ram_w8_l4096_id0_2_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _41094_ ( .CLK(CLK), .D(_25503_), .Q(ram_w8_l4096_id0_2_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41095_ ( .CLK(CLK), .D(_25501_), .Q(ram_w8_l4096_id0_2_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l4096_id0_2_1_wenable_reg ( .CLK(CLK), .D(_25500_), .Q(ram_w8_l4096_id0_2_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41097_ ( .CLK(CLK), .D(_25498_), .Q(_tmp_968), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_969_reg ( .CLK(CLK), .D(_25496_), .Q(_tmp_969), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _41099_ ( .CLK(CLK), .D(_25514_), .Q(ram_w8_l4096_id0_1_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _41100_ ( .CLK(CLK), .D(_25513_), .Q(ram_w8_l4096_id0_1_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41101_ ( .CLK(CLK), .D(_25511_), .Q(ram_w8_l4096_id0_1_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l4096_id0_1_1_wenable_reg ( .CLK(CLK), .D(_25510_), .Q(ram_w8_l4096_id0_1_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41103_ ( .CLK(CLK), .D(_25508_), .Q(_tmp_966), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_967_reg ( .CLK(CLK), .D(_25506_), .Q(_tmp_967), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _41105_ ( .CLK(CLK), .D(_25524_), .Q(ram_w8_l4096_id0_0_0_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(10), .SRST_POLARITY(1'h1), .SRST_VALUE(10'h000) ) _41106_ ( .CLK(CLK), .D(_25523_), .Q(ram_w8_l4096_id0_0_1_addr), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41107_ ( .CLK(CLK), .D(_25521_), .Q(ram_w8_l4096_id0_0_1_wdata), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) ram_w8_l4096_id0_0_1_wenable_reg ( .CLK(CLK), .D(_25520_), .Q(ram_w8_l4096_id0_0_1_wenable), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(34), .SRST_POLARITY(1'h1), .SRST_VALUE(34'h000000000) ) _41109_ ( .CLK(CLK), .D(_25518_), .Q(_tmp_964), .SRST(RST) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_965_reg ( .CLK(CLK), .D(_25516_), .Q(_tmp_965), .SRST(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) RST_reg  ( .CLK(CLK), .D(_00000_), .Q(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _rst_logic_1_reg  ( .CLK(CLK), .D(rst_logic), .Q(_rst_logic_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _rst_logic_2_reg  ( .CLK(CLK), .D(_rst_logic_1), .Q(_rst_logic_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41114_ ( .CLK(CLK), .D(_25527_), .Q(_saxi_register_fsm), .SRST(_RESETN_inv_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _41115_ ( .CLK(CLK), .D(_02883_), .Q(_tmp_5) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) saxi_bvalid_reg ( .CLK(CLK), .D(_25590_), .Q(saxi_bvalid), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41117_ ( .CLK(CLK), .D(_25588_), .Q(saxi_rdata), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) saxi_rvalid_reg ( .CLK(CLK), .D(_25587_), .Q(saxi_rvalid), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41119_ ( .CLK(CLK), .D(_25584_), .Q(_saxi_register_0), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41120_ ( .CLK(CLK), .D(_25582_), .Q(_saxi_register_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41121_ ( .CLK(CLK), .D(_25580_), .Q(_saxi_register_2), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41122_ ( .CLK(CLK), .D(_25578_), .Q(_saxi_register_3), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41123_ ( .CLK(CLK), .D(_25576_), .Q(_saxi_register_4), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41124_ ( .CLK(CLK), .D(_25573_), .Q(_saxi_register_5), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41125_ ( .CLK(CLK), .D(_25568_), .Q(_saxi_register_6), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41126_ ( .CLK(CLK), .D(_25565_), .Q(_saxi_register_7), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41127_ ( .CLK(CLK), .D(_25562_), .Q(_saxi_register_8), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41128_ ( .CLK(CLK), .D(_25560_), .Q(_saxi_register_9), .SRST(_RESETN_inv_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41129_ ( .CLK(CLK), .D(_01730_), .Q(_saxi_register_10) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41130_ ( .CLK(CLK), .D(_25556_), .Q(_saxi_register_11), .SRST(_RESETN_inv_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41131_ ( .CLK(CLK), .D(_01732_), .Q(_saxi_register_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41132_ ( .CLK(CLK), .D(_01733_), .Q(_saxi_register_13) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_0_reg ( .CLK(CLK), .D(_25550_), .Q(_saxi_flag_0), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_1_reg ( .CLK(CLK), .D(_25549_), .Q(_saxi_flag_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_2_reg ( .CLK(CLK), .D(_25548_), .Q(_saxi_flag_2), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_3_reg ( .CLK(CLK), .D(_25547_), .Q(_saxi_flag_3), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_4_reg ( .CLK(CLK), .D(_25546_), .Q(_saxi_flag_4), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_5_reg ( .CLK(CLK), .D(_25544_), .Q(_saxi_flag_5), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_6_reg ( .CLK(CLK), .D(_25541_), .Q(_saxi_flag_6), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_7_reg ( .CLK(CLK), .D(_25540_), .Q(_saxi_flag_7), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_8_reg ( .CLK(CLK), .D(_25539_), .Q(_saxi_flag_8), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_9_reg ( .CLK(CLK), .D(_25538_), .Q(_saxi_flag_9), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_10_reg ( .CLK(CLK), .D(_25537_), .Q(_saxi_flag_10), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_11_reg ( .CLK(CLK), .D(_25536_), .Q(_saxi_flag_11), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_12_reg ( .CLK(CLK), .D(_25535_), .Q(_saxi_flag_12), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_flag_13_reg ( .CLK(CLK), .D(_25534_), .Q(_saxi_flag_13), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(6), .SRST_POLARITY(1'h1), .SRST_VALUE(6'h00) ) _41147_ ( .CLK(CLK), .D(_25533_), .Q(_tmp_0), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1_reg ( .CLK(CLK), .D(_25531_), .Q(_tmp_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_2_reg ( .CLK(CLK), .D(_25530_), .Q(_tmp_2), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_3_reg ( .CLK(CLK), .D(saxi_awvalid), .Q(_tmp_3), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_4_reg ( .CLK(CLK), .D(saxi_arvalid), .Q(_tmp_4), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _saxi_cond_0_1_reg ( .CLK(CLK), .D(1'h1), .Q(_saxi_cond_0_1), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41153_ ( .CLK(CLK), .D(_25689_), .Q(_dataflow_slice_data_4), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_4_reg ( .CLK(CLK), .D(_25688_), .Q(_dataflow_slice_valid_4), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41155_ ( .CLK(CLK), .D(_25686_), .Q(_dataflow_slice_data_7), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_7_reg ( .CLK(CLK), .D(_25685_), .Q(_dataflow_slice_valid_7), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41157_ ( .CLK(CLK), .D(_25683_), .Q(_dataflow_slice_data_10), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_10_reg ( .CLK(CLK), .D(_25682_), .Q(_dataflow_slice_valid_10), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41159_ ( .CLK(CLK), .D(_25680_), .Q(_dataflow_slice_data_13), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_13_reg ( .CLK(CLK), .D(_25679_), .Q(_dataflow_slice_valid_13), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41161_ ( .CLK(CLK), .D(_25677_), .Q(_dataflow_slice_data_17), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_17_reg ( .CLK(CLK), .D(_25676_), .Q(_dataflow_slice_valid_17), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41163_ ( .CLK(CLK), .D(_25674_), .Q(_dataflow_slice_data_20), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_20_reg ( .CLK(CLK), .D(_25673_), .Q(_dataflow_slice_valid_20), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41165_ ( .CLK(CLK), .D(_25671_), .Q(_dataflow_slice_data_23), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_23_reg ( .CLK(CLK), .D(_25670_), .Q(_dataflow_slice_valid_23), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41167_ ( .CLK(CLK), .D(_25668_), .Q(_dataflow_slice_data_26), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_26_reg ( .CLK(CLK), .D(_25667_), .Q(_dataflow_slice_valid_26), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41169_ ( .CLK(CLK), .D(_25665_), .Q(_dataflow_slice_data_30), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_30_reg ( .CLK(CLK), .D(_25664_), .Q(_dataflow_slice_valid_30), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41171_ ( .CLK(CLK), .D(_25662_), .Q(_dataflow_slice_data_33), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_33_reg ( .CLK(CLK), .D(_25661_), .Q(_dataflow_slice_valid_33), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41173_ ( .CLK(CLK), .D(_25659_), .Q(_dataflow_slice_data_36), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_36_reg ( .CLK(CLK), .D(_25658_), .Q(_dataflow_slice_valid_36), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41175_ ( .CLK(CLK), .D(_25656_), .Q(_dataflow_slice_data_39), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_39_reg ( .CLK(CLK), .D(_25655_), .Q(_dataflow_slice_valid_39), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41177_ ( .CLK(CLK), .D(_25653_), .Q(_dataflow_slice_data_43), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_43_reg ( .CLK(CLK), .D(_25652_), .Q(_dataflow_slice_valid_43), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41179_ ( .CLK(CLK), .D(_25650_), .Q(_dataflow_slice_data_46), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_46_reg ( .CLK(CLK), .D(_25649_), .Q(_dataflow_slice_valid_46), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41181_ ( .CLK(CLK), .D(_25647_), .Q(_dataflow_slice_data_49), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_49_reg ( .CLK(CLK), .D(_25646_), .Q(_dataflow_slice_valid_49), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41183_ ( .CLK(CLK), .D(_25644_), .Q(_dataflow_slice_data_52), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_52_reg ( .CLK(CLK), .D(_25643_), .Q(_dataflow_slice_valid_52), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41185_ ( .CLK(CLK), .D(_25641_), .Q(_dataflow_slice_data_56), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_56_reg ( .CLK(CLK), .D(_25640_), .Q(_dataflow_slice_valid_56), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41187_ ( .CLK(CLK), .D(_25638_), .Q(_dataflow_slice_data_59), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_59_reg ( .CLK(CLK), .D(_25637_), .Q(_dataflow_slice_valid_59), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41189_ ( .CLK(CLK), .D(_25635_), .Q(_dataflow_slice_data_62), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_62_reg ( .CLK(CLK), .D(_25634_), .Q(_dataflow_slice_valid_62), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41191_ ( .CLK(CLK), .D(_25632_), .Q(_dataflow_slice_data_65), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_65_reg ( .CLK(CLK), .D(_25631_), .Q(_dataflow_slice_valid_65), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41193_ ( .CLK(CLK), .D(_25629_), .Q(_dataflow_slice_data_78), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_78_reg ( .CLK(CLK), .D(_25628_), .Q(_dataflow_slice_valid_78), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41195_ ( .CLK(CLK), .D(_25626_), .Q(_dataflow_slice_data_81), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_81_reg ( .CLK(CLK), .D(_25625_), .Q(_dataflow_slice_valid_81), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41197_ ( .CLK(CLK), .D(_25623_), .Q(_dataflow_slice_data_84), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_84_reg ( .CLK(CLK), .D(_25622_), .Q(_dataflow_slice_valid_84), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41199_ ( .CLK(CLK), .D(_25620_), .Q(_dataflow_slice_data_87), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_87_reg ( .CLK(CLK), .D(_25619_), .Q(_dataflow_slice_valid_87), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41201_ ( .CLK(CLK), .D(_25617_), .Q(_dataflow_slice_data_100), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_100_reg ( .CLK(CLK), .D(_25616_), .Q(_dataflow_slice_valid_100), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41203_ ( .CLK(CLK), .D(_25614_), .Q(_dataflow_slice_data_103), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_103_reg ( .CLK(CLK), .D(_25613_), .Q(_dataflow_slice_valid_103), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41205_ ( .CLK(CLK), .D(_25611_), .Q(_dataflow_slice_data_106), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_106_reg ( .CLK(CLK), .D(_25610_), .Q(_dataflow_slice_valid_106), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41207_ ( .CLK(CLK), .D(_25608_), .Q(_dataflow_slice_data_109), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_109_reg ( .CLK(CLK), .D(_25607_), .Q(_dataflow_slice_valid_109), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41209_ ( .CLK(CLK), .D(_25605_), .Q(_dataflow_slice_data_113), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_113_reg ( .CLK(CLK), .D(_25604_), .Q(_dataflow_slice_valid_113), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41211_ ( .CLK(CLK), .D(_25602_), .Q(_dataflow_slice_data_116), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_116_reg ( .CLK(CLK), .D(_25601_), .Q(_dataflow_slice_valid_116), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41213_ ( .CLK(CLK), .D(_25599_), .Q(_dataflow_slice_data_119), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_119_reg ( .CLK(CLK), .D(_25598_), .Q(_dataflow_slice_valid_119), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41215_ ( .CLK(CLK), .D(_25596_), .Q(_dataflow_slice_data_122), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow_slice_valid_122_reg ( .CLK(CLK), .D(_25595_), .Q(_dataflow_slice_valid_122), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41217_ ( .CLK(CLK), .D(_25593_), .Q(_dataflow__delay_data_132), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _dataflow__delay_valid_132_reg ( .CLK(CLK), .D(_25592_), .Q(_dataflow__delay_valid_132), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41219_ ( .CLK(CLK), .D(_25910_), .Q(maxi_awaddr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41220_ ( .CLK(CLK), .D(_25909_), .Q(maxi_awlen), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) maxi_awvalid_reg ( .CLK(CLK), .D(_25908_), .Q(maxi_awvalid), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41222_ ( .CLK(CLK), .D(_25904_), .Q(maxi_wdata), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(4), .SRST_POLARITY(1'h1), .SRST_VALUE(4'h0) ) _41223_ ( .CLK(CLK), .D(_25901_), .Q(maxi_wstrb), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) maxi_wlast_reg ( .CLK(CLK), .D(_25898_), .Q(maxi_wlast), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) maxi_wvalid_reg ( .CLK(CLK), .D(_25890_), .Q(maxi_wvalid), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41226_ ( .CLK(CLK), .D(_25885_), .Q(maxi_araddr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41227_ ( .CLK(CLK), .D(_25884_), .Q(maxi_arlen), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) maxi_arvalid_reg ( .CLK(CLK), .D(_25883_), .Q(maxi_arvalid), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_read_start_reg ( .CLK(CLK), .D(_25880_), .Q(_maxi_read_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41230_ ( .CLK(CLK), .D(_25871_), .Q(_maxi_read_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41231_ ( .CLK(CLK), .D(_25862_), .Q(_maxi_read_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41232_ ( .CLK(CLK), .D(_25853_), .Q(_maxi_read_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41233_ ( .CLK(CLK), .D(_25844_), .Q(_maxi_read_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41234_ ( .CLK(CLK), .D(_25835_), .Q(_maxi_read_local_stride), .SRST(_RESETN_inv_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_read_idle_reg  ( .CLK(CLK), .D(_01646_), .Q(_maxi_read_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_write_start_reg ( .CLK(CLK), .D(_25816_), .Q(_maxi_write_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41237_ ( .CLK(CLK), .D(_25813_), .Q(_maxi_write_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41238_ ( .CLK(CLK), .D(_25810_), .Q(_maxi_write_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41239_ ( .CLK(CLK), .D(_25807_), .Q(_maxi_write_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41240_ ( .CLK(CLK), .D(_25804_), .Q(_maxi_write_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41241_ ( .CLK(CLK), .D(_25801_), .Q(_maxi_write_local_stride), .SRST(_RESETN_inv_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_write_idle_reg  ( .CLK(CLK), .D(_01657_), .Q(_maxi_write_idle) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41243_ ( .CLK(CLK), .D(_saxi_register_9), .Q(_maxi_global_base_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_ram_w32_l128_id0_1_read_start_reg ( .CLK(CLK), .D(_25794_), .Q(_maxi_ram_w32_l128_id0_1_read_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41245_ ( .CLK(CLK), .D(_25792_), .Q(_maxi_ram_w32_l128_id0_1_read_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41246_ ( .CLK(CLK), .D(_25790_), .Q(_maxi_ram_w32_l128_id0_1_read_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41247_ ( .CLK(CLK), .D(_25788_), .Q(_maxi_ram_w32_l128_id0_1_read_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41248_ ( .CLK(CLK), .D(_25786_), .Q(_maxi_ram_w32_l128_id0_1_read_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41249_ ( .CLK(CLK), .D(_25784_), .Q(_maxi_ram_w32_l128_id0_1_read_local_stride), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _41250_ ( .CLK(CLK), .D(_25782_), .Q(_tmp_14), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_ram_w8_l2048_id0_1_read_start_reg ( .CLK(CLK), .D(_25780_), .Q(_maxi_ram_w8_l2048_id0_1_read_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41252_ ( .CLK(CLK), .D(_25778_), .Q(_maxi_ram_w8_l2048_id0_1_read_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41253_ ( .CLK(CLK), .D(_25776_), .Q(_maxi_ram_w8_l2048_id0_1_read_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41254_ ( .CLK(CLK), .D(_25774_), .Q(_maxi_ram_w8_l2048_id0_1_read_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41255_ ( .CLK(CLK), .D(_25772_), .Q(_maxi_ram_w8_l2048_id0_1_read_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41256_ ( .CLK(CLK), .D(_25770_), .Q(_maxi_ram_w8_l2048_id0_1_read_local_stride), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_start_reg ( .CLK(CLK), .D(_25768_), .Q(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41258_ ( .CLK(CLK), .D(_25767_), .Q(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41259_ ( .CLK(CLK), .D(_25766_), .Q(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41260_ ( .CLK(CLK), .D(_25765_), .Q(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41261_ ( .CLK(CLK), .D(_25764_), .Q(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41262_ ( .CLK(CLK), .D(_25763_), .Q(_maxi_ram_w8_l2048_id1_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_ram_w8_l2048_id8_ram_w8_l2048_id9_1_read_local_stride), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_start_reg ( .CLK(CLK), .D(_25762_), .Q(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41264_ ( .CLK(CLK), .D(_25761_), .Q(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41265_ ( .CLK(CLK), .D(_25760_), .Q(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41266_ ( .CLK(CLK), .D(_25759_), .Q(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41267_ ( .CLK(CLK), .D(_25758_), .Q(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41268_ ( .CLK(CLK), .D(_25757_), .Q(_maxi_ram_w8_l2048_id10_ram_w8_l2048_id11_ram_w8_l2048_id12_1_read_local_stride), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_start_reg ( .CLK(CLK), .D(_25756_), .Q(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41270_ ( .CLK(CLK), .D(_25755_), .Q(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41271_ ( .CLK(CLK), .D(_25754_), .Q(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41272_ ( .CLK(CLK), .D(_25753_), .Q(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41273_ ( .CLK(CLK), .D(_25752_), .Q(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41274_ ( .CLK(CLK), .D(_25751_), .Q(_maxi_ram_w8_l2048_id13_ram_w8_l2048_id14_ram_w8_l2048_id15_1_read_local_stride), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_start_reg ( .CLK(CLK), .D(_25750_), .Q(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41276_ ( .CLK(CLK), .D(_25749_), .Q(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41277_ ( .CLK(CLK), .D(_25748_), .Q(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41278_ ( .CLK(CLK), .D(_25747_), .Q(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41279_ ( .CLK(CLK), .D(_25746_), .Q(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41280_ ( .CLK(CLK), .D(_25745_), .Q(_maxi_ram_w8_l2048_id16_ram_w8_l2048_id17_ram_w8_l2048_id18_1_read_local_stride), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_ram_w8_l2048_id19_1_write_start_reg ( .CLK(CLK), .D(_25744_), .Q(_maxi_ram_w8_l2048_id19_1_write_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41282_ ( .CLK(CLK), .D(_25743_), .Q(_maxi_ram_w8_l2048_id19_1_write_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41283_ ( .CLK(CLK), .D(_25742_), .Q(_maxi_ram_w8_l2048_id19_1_write_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41284_ ( .CLK(CLK), .D(_25741_), .Q(_maxi_ram_w8_l2048_id19_1_write_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41285_ ( .CLK(CLK), .D(_25740_), .Q(_maxi_ram_w8_l2048_id19_1_write_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41286_ ( .CLK(CLK), .D(_25739_), .Q(_maxi_ram_w8_l2048_id19_1_write_local_stride), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(9), .SRST_POLARITY(1'h1), .SRST_VALUE(9'h000) ) _41287_ ( .CLK(CLK), .D(_25738_), .Q(_tmp_847), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_848_reg ( .CLK(CLK), .D(_25734_), .Q(_tmp_848), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_ram_w8_l2048_id1_1_read_start_reg ( .CLK(CLK), .D(_25731_), .Q(_maxi_ram_w8_l2048_id1_1_read_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41290_ ( .CLK(CLK), .D(_25729_), .Q(_maxi_ram_w8_l2048_id1_1_read_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41291_ ( .CLK(CLK), .D(_25727_), .Q(_maxi_ram_w8_l2048_id1_1_read_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41292_ ( .CLK(CLK), .D(_25725_), .Q(_maxi_ram_w8_l2048_id1_1_read_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41293_ ( .CLK(CLK), .D(_25723_), .Q(_maxi_ram_w8_l2048_id1_1_read_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41294_ ( .CLK(CLK), .D(_25721_), .Q(_maxi_ram_w8_l2048_id1_1_read_local_stride), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_ram_w8_l2048_id0_1_write_start_reg ( .CLK(CLK), .D(_25719_), .Q(_maxi_ram_w8_l2048_id0_1_write_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41296_ ( .CLK(CLK), .D(_25718_), .Q(_maxi_ram_w8_l2048_id0_1_write_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41297_ ( .CLK(CLK), .D(_25717_), .Q(_maxi_ram_w8_l2048_id0_1_write_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41298_ ( .CLK(CLK), .D(_25716_), .Q(_maxi_ram_w8_l2048_id0_1_write_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41299_ ( .CLK(CLK), .D(_25715_), .Q(_maxi_ram_w8_l2048_id0_1_write_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41300_ ( .CLK(CLK), .D(_25714_), .Q(_maxi_ram_w8_l2048_id0_1_write_local_stride), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_958_reg ( .CLK(CLK), .D(_25713_), .Q(_tmp_958), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_ram_w8_l4096_id0_1_read_start_reg ( .CLK(CLK), .D(_25710_), .Q(_maxi_ram_w8_l4096_id0_1_read_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41303_ ( .CLK(CLK), .D(_25709_), .Q(_maxi_ram_w8_l4096_id0_1_read_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41304_ ( .CLK(CLK), .D(_25708_), .Q(_maxi_ram_w8_l4096_id0_1_read_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41305_ ( .CLK(CLK), .D(_25707_), .Q(_maxi_ram_w8_l4096_id0_1_read_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41306_ ( .CLK(CLK), .D(_25706_), .Q(_maxi_ram_w8_l4096_id0_1_read_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41307_ ( .CLK(CLK), .D(_25705_), .Q(_maxi_ram_w8_l4096_id0_1_read_local_stride), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_ram_w8_l2048_id2_1_read_start_reg ( .CLK(CLK), .D(_25704_), .Q(_maxi_ram_w8_l2048_id2_1_read_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41309_ ( .CLK(CLK), .D(_25703_), .Q(_maxi_ram_w8_l2048_id2_1_read_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41310_ ( .CLK(CLK), .D(_25702_), .Q(_maxi_ram_w8_l2048_id2_1_read_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41311_ ( .CLK(CLK), .D(_25701_), .Q(_maxi_ram_w8_l2048_id2_1_read_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41312_ ( .CLK(CLK), .D(_25700_), .Q(_maxi_ram_w8_l2048_id2_1_read_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41313_ ( .CLK(CLK), .D(_25699_), .Q(_maxi_ram_w8_l2048_id2_1_read_local_stride), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _maxi_ram_w8_l2048_id1_1_write_start_reg ( .CLK(CLK), .D(_25698_), .Q(_maxi_ram_w8_l2048_id1_1_write_start), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(8), .SRST_POLARITY(1'h1), .SRST_VALUE(8'h00) ) _41315_ ( .CLK(CLK), .D(_25697_), .Q(_maxi_ram_w8_l2048_id1_1_write_op_sel), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41316_ ( .CLK(CLK), .D(_25696_), .Q(_maxi_ram_w8_l2048_id1_1_write_local_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41317_ ( .CLK(CLK), .D(_25695_), .Q(_maxi_ram_w8_l2048_id1_1_write_global_addr), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(33), .SRST_POLARITY(1'h1), .SRST_VALUE(33'h000000000) ) _41318_ ( .CLK(CLK), .D(_25694_), .Q(_maxi_ram_w8_l2048_id1_1_write_size), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(32), .SRST_POLARITY(1'h1), .SRST_VALUE(0) ) _41319_ ( .CLK(CLK), .D(_25693_), .Q(_maxi_ram_w8_l2048_id1_1_write_local_stride), .SRST(_RESETN_inv_2) );
  \$sdff #( .CLK_POLARITY(1'h1), .WIDTH(1), .SRST_POLARITY(1'h1), .SRST_VALUE(1'h0) ) _tmp_1167_reg ( .CLK(CLK), .D(_25692_), .Q(_tmp_1167), .SRST(_RESETN_inv_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _RESETN_inv_1_reg  ( .CLK(CLK), .D(RESETN_inv), .Q(_RESETN_inv_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _RESETN_inv_2_reg  ( .CLK(CLK), .D(_RESETN_inv_1), .Q(_RESETN_inv_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49075_ ( .CLK(CLK), .D(_cond_data_108), .Q(\__muladd_madd_110.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49076_ ( .CLK(CLK), .D(__delay_data_630), .Q(\__muladd_madd_110.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49077_ ( .CLK(CLK), .D(\__muladd_madd_110.madd._madd ), .Q(\__muladd_madd_110.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49078_ ( .CLK(CLK), .D(__delay_data_627), .Q(\__muladd_madd_110.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49079_ ( .CLK(CLK), .D(\__muladd_madd_110.madd._pipe_madd0 ), .Q(\__muladd_madd_110.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49082_ ( .CLK(CLK), .D(_cond_data_123), .Q(\__muladd_madd_125.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49083_ ( .CLK(CLK), .D(__delay_data_647), .Q(\__muladd_madd_125.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49084_ ( .CLK(CLK), .D(\__muladd_madd_125.madd._madd ), .Q(\__muladd_madd_125.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49085_ ( .CLK(CLK), .D(__delay_data_644), .Q(\__muladd_madd_125.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49086_ ( .CLK(CLK), .D(\__muladd_madd_125.madd._pipe_madd0 ), .Q(\__muladd_madd_125.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49089_ ( .CLK(CLK), .D(_cond_data_138), .Q(\__muladd_madd_140.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49090_ ( .CLK(CLK), .D(__delay_data_664), .Q(\__muladd_madd_140.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49091_ ( .CLK(CLK), .D(\__muladd_madd_140.madd._madd ), .Q(\__muladd_madd_140.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49092_ ( .CLK(CLK), .D(__delay_data_661), .Q(\__muladd_madd_140.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49093_ ( .CLK(CLK), .D(\__muladd_madd_140.madd._pipe_madd0 ), .Q(\__muladd_madd_140.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49096_ ( .CLK(CLK), .D(_cond_data_153), .Q(\__muladd_madd_155.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49097_ ( .CLK(CLK), .D(__delay_data_681), .Q(\__muladd_madd_155.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49098_ ( .CLK(CLK), .D(\__muladd_madd_155.madd._madd ), .Q(\__muladd_madd_155.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49099_ ( .CLK(CLK), .D(__delay_data_678), .Q(\__muladd_madd_155.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49100_ ( .CLK(CLK), .D(\__muladd_madd_155.madd._pipe_madd0 ), .Q(\__muladd_madd_155.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49103_ ( .CLK(CLK), .D(_cond_data_168), .Q(\__muladd_madd_170.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49104_ ( .CLK(CLK), .D(__delay_data_698), .Q(\__muladd_madd_170.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49105_ ( .CLK(CLK), .D(\__muladd_madd_170.madd._madd ), .Q(\__muladd_madd_170.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49106_ ( .CLK(CLK), .D(__delay_data_695), .Q(\__muladd_madd_170.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49107_ ( .CLK(CLK), .D(\__muladd_madd_170.madd._pipe_madd0 ), .Q(\__muladd_madd_170.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49110_ ( .CLK(CLK), .D(_cond_data_183), .Q(\__muladd_madd_185.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49111_ ( .CLK(CLK), .D(__delay_data_715), .Q(\__muladd_madd_185.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49112_ ( .CLK(CLK), .D(\__muladd_madd_185.madd._madd ), .Q(\__muladd_madd_185.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49113_ ( .CLK(CLK), .D(__delay_data_712), .Q(\__muladd_madd_185.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49114_ ( .CLK(CLK), .D(\__muladd_madd_185.madd._pipe_madd0 ), .Q(\__muladd_madd_185.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49117_ ( .CLK(CLK), .D(_cond_data_63), .Q(\__muladd_madd_65.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49118_ ( .CLK(CLK), .D(__delay_data_579), .Q(\__muladd_madd_65.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49119_ ( .CLK(CLK), .D(\__muladd_madd_65.madd._madd ), .Q(\__muladd_madd_65.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49120_ ( .CLK(CLK), .D(__delay_data_576), .Q(\__muladd_madd_65.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49121_ ( .CLK(CLK), .D(\__muladd_madd_65.madd._pipe_madd0 ), .Q(\__muladd_madd_65.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49124_ ( .CLK(CLK), .D(_cond_data_78), .Q(\__muladd_madd_80.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49125_ ( .CLK(CLK), .D(__delay_data_596), .Q(\__muladd_madd_80.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49126_ ( .CLK(CLK), .D(\__muladd_madd_80.madd._madd ), .Q(\__muladd_madd_80.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49127_ ( .CLK(CLK), .D(__delay_data_593), .Q(\__muladd_madd_80.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49128_ ( .CLK(CLK), .D(\__muladd_madd_80.madd._pipe_madd0 ), .Q(\__muladd_madd_80.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49131_ ( .CLK(CLK), .D(_cond_data_93), .Q(\__muladd_madd_95.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49132_ ( .CLK(CLK), .D(__delay_data_613), .Q(\__muladd_madd_95.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49133_ ( .CLK(CLK), .D(\__muladd_madd_95.madd._madd ), .Q(\__muladd_madd_95.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49134_ ( .CLK(CLK), .D(__delay_data_610), .Q(\__muladd_madd_95.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(16) ) _49135_ ( .CLK(CLK), .D(\__muladd_madd_95.madd._pipe_madd0 ), .Q(\__muladd_madd_95.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _49137_ ( .CLK(CLK), .D(__variable_wdata_37), .Q(\_times_mul_39.mult._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _49138_ ( .CLK(CLK), .D(__variable_wdata_36), .Q(\_times_mul_39.mult._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(40) ) _49139_ ( .CLK(CLK), .D(\_times_mul_39.mult._mul ), .Q(\_times_mul_39.mult._pipe_mul0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(40) ) _49140_ ( .CLK(CLK), .D(\_times_mul_39.mult._pipe_mul0 ), .Q(\_times_mul_39.mult._pipe_mul1 ) );
  ram_w32_l128_id0 inst_ram_w32_l128_id0 ( .CLK(CLK), .ram_w32_l128_id0_0_addr(ram_w32_l128_id0_0_addr), .ram_w32_l128_id0_0_rdata(ram_w32_l128_id0_0_rdata), .ram_w32_l128_id0_0_wdata(0), .ram_w32_l128_id0_0_wenable(1'h0), .ram_w32_l128_id0_1_addr(ram_w32_l128_id0_1_addr), .ram_w32_l128_id0_1_rdata(ram_w32_l128_id0_1_rdata), .ram_w32_l128_id0_1_wdata(ram_w32_l128_id0_1_wdata), .ram_w32_l128_id0_1_wenable(ram_w32_l128_id0_1_wenable) );
  ram_w8_l2048_id0_0 inst_ram_w8_l2048_id0_0 ( .CLK(CLK), .ram_w8_l2048_id0_0_0_addr(ram_w8_l2048_id0_0_0_addr), .ram_w8_l2048_id0_0_0_rdata(ram_w8_l2048_id0_0_0_rdata), .ram_w8_l2048_id0_0_0_wdata(ram_w8_l2048_id0_0_0_wdata), .ram_w8_l2048_id0_0_0_wenable(ram_w8_l2048_id0_0_0_wenable), .ram_w8_l2048_id0_0_1_addr(ram_w8_l2048_id0_0_1_addr), .ram_w8_l2048_id0_0_1_rdata(ram_w8_l2048_id0_0_1_rdata), .ram_w8_l2048_id0_0_1_wdata(ram_w8_l2048_id0_0_1_wdata), .ram_w8_l2048_id0_0_1_wenable(ram_w8_l2048_id0_0_1_wenable) );
  ram_w8_l2048_id0_1 inst_ram_w8_l2048_id0_1 ( .CLK(CLK), .ram_w8_l2048_id0_1_0_addr(ram_w8_l2048_id0_1_0_addr), .ram_w8_l2048_id0_1_0_rdata(ram_w8_l2048_id0_1_0_rdata), .ram_w8_l2048_id0_1_0_wdata(ram_w8_l2048_id0_1_0_wdata), .ram_w8_l2048_id0_1_0_wenable(ram_w8_l2048_id0_1_0_wenable), .ram_w8_l2048_id0_1_1_addr(ram_w8_l2048_id0_1_1_addr), .ram_w8_l2048_id0_1_1_rdata(ram_w8_l2048_id0_1_1_rdata), .ram_w8_l2048_id0_1_1_wdata(ram_w8_l2048_id0_1_1_wdata), .ram_w8_l2048_id0_1_1_wenable(ram_w8_l2048_id0_1_1_wenable) );
  ram_w8_l2048_id0_2 inst_ram_w8_l2048_id0_2 ( .CLK(CLK), .ram_w8_l2048_id0_2_0_addr(ram_w8_l2048_id0_2_0_addr), .ram_w8_l2048_id0_2_0_rdata(ram_w8_l2048_id0_2_0_rdata), .ram_w8_l2048_id0_2_0_wdata(ram_w8_l2048_id0_2_0_wdata), .ram_w8_l2048_id0_2_0_wenable(ram_w8_l2048_id0_2_0_wenable), .ram_w8_l2048_id0_2_1_addr(ram_w8_l2048_id0_2_1_addr), .ram_w8_l2048_id0_2_1_rdata(ram_w8_l2048_id0_2_1_rdata), .ram_w8_l2048_id0_2_1_wdata(ram_w8_l2048_id0_2_1_wdata), .ram_w8_l2048_id0_2_1_wenable(ram_w8_l2048_id0_2_1_wenable) );
  ram_w8_l2048_id0_3 inst_ram_w8_l2048_id0_3 ( .CLK(CLK), .ram_w8_l2048_id0_3_0_addr(ram_w8_l2048_id0_3_0_addr), .ram_w8_l2048_id0_3_0_rdata(ram_w8_l2048_id0_3_0_rdata), .ram_w8_l2048_id0_3_0_wdata(ram_w8_l2048_id0_3_0_wdata), .ram_w8_l2048_id0_3_0_wenable(ram_w8_l2048_id0_3_0_wenable), .ram_w8_l2048_id0_3_1_addr(ram_w8_l2048_id0_3_1_addr), .ram_w8_l2048_id0_3_1_rdata(ram_w8_l2048_id0_3_1_rdata), .ram_w8_l2048_id0_3_1_wdata(ram_w8_l2048_id0_3_1_wdata), .ram_w8_l2048_id0_3_1_wenable(ram_w8_l2048_id0_3_1_wenable) );
  ram_w8_l2048_id10_0 inst_ram_w8_l2048_id10_0 ( .CLK(CLK), .ram_w8_l2048_id10_0_0_addr(ram_w8_l2048_id10_0_0_addr), .ram_w8_l2048_id10_0_0_rdata(ram_w8_l2048_id10_0_0_rdata), .ram_w8_l2048_id10_0_0_wdata(8'h00), .ram_w8_l2048_id10_0_0_wenable(1'h0), .ram_w8_l2048_id10_0_1_addr(ram_w8_l2048_id10_0_1_addr), .ram_w8_l2048_id10_0_1_rdata(ram_w8_l2048_id10_0_1_rdata), .ram_w8_l2048_id10_0_1_wdata(ram_w8_l2048_id10_0_1_wdata), .ram_w8_l2048_id10_0_1_wenable(ram_w8_l2048_id10_0_1_wenable) );
  ram_w8_l2048_id10_1 inst_ram_w8_l2048_id10_1 ( .CLK(CLK), .ram_w8_l2048_id10_1_0_addr(ram_w8_l2048_id10_1_0_addr), .ram_w8_l2048_id10_1_0_rdata(ram_w8_l2048_id10_1_0_rdata), .ram_w8_l2048_id10_1_0_wdata(8'h00), .ram_w8_l2048_id10_1_0_wenable(1'h0), .ram_w8_l2048_id10_1_1_addr(ram_w8_l2048_id10_1_1_addr), .ram_w8_l2048_id10_1_1_rdata(ram_w8_l2048_id10_1_1_rdata), .ram_w8_l2048_id10_1_1_wdata(ram_w8_l2048_id10_1_1_wdata), .ram_w8_l2048_id10_1_1_wenable(ram_w8_l2048_id10_1_1_wenable) );
  ram_w8_l2048_id10_2 inst_ram_w8_l2048_id10_2 ( .CLK(CLK), .ram_w8_l2048_id10_2_0_addr(ram_w8_l2048_id10_2_0_addr), .ram_w8_l2048_id10_2_0_rdata(ram_w8_l2048_id10_2_0_rdata), .ram_w8_l2048_id10_2_0_wdata(8'h00), .ram_w8_l2048_id10_2_0_wenable(1'h0), .ram_w8_l2048_id10_2_1_addr(ram_w8_l2048_id10_2_1_addr), .ram_w8_l2048_id10_2_1_rdata(ram_w8_l2048_id10_2_1_rdata), .ram_w8_l2048_id10_2_1_wdata(ram_w8_l2048_id10_2_1_wdata), .ram_w8_l2048_id10_2_1_wenable(ram_w8_l2048_id10_2_1_wenable) );
  ram_w8_l2048_id10_3 inst_ram_w8_l2048_id10_3 ( .CLK(CLK), .ram_w8_l2048_id10_3_0_addr(ram_w8_l2048_id10_3_0_addr), .ram_w8_l2048_id10_3_0_rdata(ram_w8_l2048_id10_3_0_rdata), .ram_w8_l2048_id10_3_0_wdata(8'h00), .ram_w8_l2048_id10_3_0_wenable(1'h0), .ram_w8_l2048_id10_3_1_addr(ram_w8_l2048_id10_3_1_addr), .ram_w8_l2048_id10_3_1_rdata(ram_w8_l2048_id10_3_1_rdata), .ram_w8_l2048_id10_3_1_wdata(ram_w8_l2048_id10_3_1_wdata), .ram_w8_l2048_id10_3_1_wenable(ram_w8_l2048_id10_3_1_wenable) );
  ram_w8_l2048_id11_0 inst_ram_w8_l2048_id11_0 ( .CLK(CLK), .ram_w8_l2048_id11_0_0_addr(ram_w8_l2048_id11_0_0_addr), .ram_w8_l2048_id11_0_0_rdata(ram_w8_l2048_id11_0_0_rdata), .ram_w8_l2048_id11_0_0_wdata(8'h00), .ram_w8_l2048_id11_0_0_wenable(1'h0), .ram_w8_l2048_id11_0_1_addr(ram_w8_l2048_id11_0_1_addr), .ram_w8_l2048_id11_0_1_rdata(ram_w8_l2048_id11_0_1_rdata), .ram_w8_l2048_id11_0_1_wdata(ram_w8_l2048_id11_0_1_wdata), .ram_w8_l2048_id11_0_1_wenable(ram_w8_l2048_id11_0_1_wenable) );
  ram_w8_l2048_id11_1 inst_ram_w8_l2048_id11_1 ( .CLK(CLK), .ram_w8_l2048_id11_1_0_addr(ram_w8_l2048_id11_1_0_addr), .ram_w8_l2048_id11_1_0_rdata(ram_w8_l2048_id11_1_0_rdata), .ram_w8_l2048_id11_1_0_wdata(8'h00), .ram_w8_l2048_id11_1_0_wenable(1'h0), .ram_w8_l2048_id11_1_1_addr(ram_w8_l2048_id11_1_1_addr), .ram_w8_l2048_id11_1_1_rdata(ram_w8_l2048_id11_1_1_rdata), .ram_w8_l2048_id11_1_1_wdata(ram_w8_l2048_id11_1_1_wdata), .ram_w8_l2048_id11_1_1_wenable(ram_w8_l2048_id11_1_1_wenable) );
  ram_w8_l2048_id11_2 inst_ram_w8_l2048_id11_2 ( .CLK(CLK), .ram_w8_l2048_id11_2_0_addr(ram_w8_l2048_id11_2_0_addr), .ram_w8_l2048_id11_2_0_rdata(ram_w8_l2048_id11_2_0_rdata), .ram_w8_l2048_id11_2_0_wdata(8'h00), .ram_w8_l2048_id11_2_0_wenable(1'h0), .ram_w8_l2048_id11_2_1_addr(ram_w8_l2048_id11_2_1_addr), .ram_w8_l2048_id11_2_1_rdata(ram_w8_l2048_id11_2_1_rdata), .ram_w8_l2048_id11_2_1_wdata(ram_w8_l2048_id11_2_1_wdata), .ram_w8_l2048_id11_2_1_wenable(ram_w8_l2048_id11_2_1_wenable) );
  ram_w8_l2048_id11_3 inst_ram_w8_l2048_id11_3 ( .CLK(CLK), .ram_w8_l2048_id11_3_0_addr(ram_w8_l2048_id11_3_0_addr), .ram_w8_l2048_id11_3_0_rdata(ram_w8_l2048_id11_3_0_rdata), .ram_w8_l2048_id11_3_0_wdata(8'h00), .ram_w8_l2048_id11_3_0_wenable(1'h0), .ram_w8_l2048_id11_3_1_addr(ram_w8_l2048_id11_3_1_addr), .ram_w8_l2048_id11_3_1_rdata(ram_w8_l2048_id11_3_1_rdata), .ram_w8_l2048_id11_3_1_wdata(ram_w8_l2048_id11_3_1_wdata), .ram_w8_l2048_id11_3_1_wenable(ram_w8_l2048_id11_3_1_wenable) );
  ram_w8_l2048_id12_0 inst_ram_w8_l2048_id12_0 ( .CLK(CLK), .ram_w8_l2048_id12_0_0_addr(ram_w8_l2048_id12_0_0_addr), .ram_w8_l2048_id12_0_0_rdata(ram_w8_l2048_id12_0_0_rdata), .ram_w8_l2048_id12_0_0_wdata(8'h00), .ram_w8_l2048_id12_0_0_wenable(1'h0), .ram_w8_l2048_id12_0_1_addr(ram_w8_l2048_id12_0_1_addr), .ram_w8_l2048_id12_0_1_rdata(ram_w8_l2048_id12_0_1_rdata), .ram_w8_l2048_id12_0_1_wdata(ram_w8_l2048_id12_0_1_wdata), .ram_w8_l2048_id12_0_1_wenable(ram_w8_l2048_id12_0_1_wenable) );
  ram_w8_l2048_id12_1 inst_ram_w8_l2048_id12_1 ( .CLK(CLK), .ram_w8_l2048_id12_1_0_addr(ram_w8_l2048_id12_1_0_addr), .ram_w8_l2048_id12_1_0_rdata(ram_w8_l2048_id12_1_0_rdata), .ram_w8_l2048_id12_1_0_wdata(8'h00), .ram_w8_l2048_id12_1_0_wenable(1'h0), .ram_w8_l2048_id12_1_1_addr(ram_w8_l2048_id12_1_1_addr), .ram_w8_l2048_id12_1_1_rdata(ram_w8_l2048_id12_1_1_rdata), .ram_w8_l2048_id12_1_1_wdata(ram_w8_l2048_id12_1_1_wdata), .ram_w8_l2048_id12_1_1_wenable(ram_w8_l2048_id12_1_1_wenable) );
  ram_w8_l2048_id12_2 inst_ram_w8_l2048_id12_2 ( .CLK(CLK), .ram_w8_l2048_id12_2_0_addr(ram_w8_l2048_id12_2_0_addr), .ram_w8_l2048_id12_2_0_rdata(ram_w8_l2048_id12_2_0_rdata), .ram_w8_l2048_id12_2_0_wdata(8'h00), .ram_w8_l2048_id12_2_0_wenable(1'h0), .ram_w8_l2048_id12_2_1_addr(ram_w8_l2048_id12_2_1_addr), .ram_w8_l2048_id12_2_1_rdata(ram_w8_l2048_id12_2_1_rdata), .ram_w8_l2048_id12_2_1_wdata(ram_w8_l2048_id12_2_1_wdata), .ram_w8_l2048_id12_2_1_wenable(ram_w8_l2048_id12_2_1_wenable) );
  ram_w8_l2048_id12_3 inst_ram_w8_l2048_id12_3 ( .CLK(CLK), .ram_w8_l2048_id12_3_0_addr(ram_w8_l2048_id12_3_0_addr), .ram_w8_l2048_id12_3_0_rdata(ram_w8_l2048_id12_3_0_rdata), .ram_w8_l2048_id12_3_0_wdata(8'h00), .ram_w8_l2048_id12_3_0_wenable(1'h0), .ram_w8_l2048_id12_3_1_addr(ram_w8_l2048_id12_3_1_addr), .ram_w8_l2048_id12_3_1_rdata(ram_w8_l2048_id12_3_1_rdata), .ram_w8_l2048_id12_3_1_wdata(ram_w8_l2048_id12_3_1_wdata), .ram_w8_l2048_id12_3_1_wenable(ram_w8_l2048_id12_3_1_wenable) );
  ram_w8_l2048_id13_0 inst_ram_w8_l2048_id13_0 ( .CLK(CLK), .ram_w8_l2048_id13_0_0_addr(ram_w8_l2048_id13_0_0_addr), .ram_w8_l2048_id13_0_0_rdata(ram_w8_l2048_id13_0_0_rdata), .ram_w8_l2048_id13_0_0_wdata(8'h00), .ram_w8_l2048_id13_0_0_wenable(1'h0), .ram_w8_l2048_id13_0_1_addr(ram_w8_l2048_id13_0_1_addr), .ram_w8_l2048_id13_0_1_rdata(ram_w8_l2048_id13_0_1_rdata), .ram_w8_l2048_id13_0_1_wdata(ram_w8_l2048_id13_0_1_wdata), .ram_w8_l2048_id13_0_1_wenable(ram_w8_l2048_id13_0_1_wenable) );
  ram_w8_l2048_id13_1 inst_ram_w8_l2048_id13_1 ( .CLK(CLK), .ram_w8_l2048_id13_1_0_addr(ram_w8_l2048_id13_1_0_addr), .ram_w8_l2048_id13_1_0_rdata(ram_w8_l2048_id13_1_0_rdata), .ram_w8_l2048_id13_1_0_wdata(8'h00), .ram_w8_l2048_id13_1_0_wenable(1'h0), .ram_w8_l2048_id13_1_1_addr(ram_w8_l2048_id13_1_1_addr), .ram_w8_l2048_id13_1_1_rdata(ram_w8_l2048_id13_1_1_rdata), .ram_w8_l2048_id13_1_1_wdata(ram_w8_l2048_id13_1_1_wdata), .ram_w8_l2048_id13_1_1_wenable(ram_w8_l2048_id13_1_1_wenable) );
  ram_w8_l2048_id13_2 inst_ram_w8_l2048_id13_2 ( .CLK(CLK), .ram_w8_l2048_id13_2_0_addr(ram_w8_l2048_id13_2_0_addr), .ram_w8_l2048_id13_2_0_rdata(ram_w8_l2048_id13_2_0_rdata), .ram_w8_l2048_id13_2_0_wdata(8'h00), .ram_w8_l2048_id13_2_0_wenable(1'h0), .ram_w8_l2048_id13_2_1_addr(ram_w8_l2048_id13_2_1_addr), .ram_w8_l2048_id13_2_1_rdata(ram_w8_l2048_id13_2_1_rdata), .ram_w8_l2048_id13_2_1_wdata(ram_w8_l2048_id13_2_1_wdata), .ram_w8_l2048_id13_2_1_wenable(ram_w8_l2048_id13_2_1_wenable) );
  ram_w8_l2048_id13_3 inst_ram_w8_l2048_id13_3 ( .CLK(CLK), .ram_w8_l2048_id13_3_0_addr(ram_w8_l2048_id13_3_0_addr), .ram_w8_l2048_id13_3_0_rdata(ram_w8_l2048_id13_3_0_rdata), .ram_w8_l2048_id13_3_0_wdata(8'h00), .ram_w8_l2048_id13_3_0_wenable(1'h0), .ram_w8_l2048_id13_3_1_addr(ram_w8_l2048_id13_3_1_addr), .ram_w8_l2048_id13_3_1_rdata(ram_w8_l2048_id13_3_1_rdata), .ram_w8_l2048_id13_3_1_wdata(ram_w8_l2048_id13_3_1_wdata), .ram_w8_l2048_id13_3_1_wenable(ram_w8_l2048_id13_3_1_wenable) );
  ram_w8_l2048_id14_0 inst_ram_w8_l2048_id14_0 ( .CLK(CLK), .ram_w8_l2048_id14_0_0_addr(ram_w8_l2048_id14_0_0_addr), .ram_w8_l2048_id14_0_0_rdata(ram_w8_l2048_id14_0_0_rdata), .ram_w8_l2048_id14_0_0_wdata(8'h00), .ram_w8_l2048_id14_0_0_wenable(1'h0), .ram_w8_l2048_id14_0_1_addr(ram_w8_l2048_id14_0_1_addr), .ram_w8_l2048_id14_0_1_rdata(ram_w8_l2048_id14_0_1_rdata), .ram_w8_l2048_id14_0_1_wdata(ram_w8_l2048_id14_0_1_wdata), .ram_w8_l2048_id14_0_1_wenable(ram_w8_l2048_id14_0_1_wenable) );
  ram_w8_l2048_id14_1 inst_ram_w8_l2048_id14_1 ( .CLK(CLK), .ram_w8_l2048_id14_1_0_addr(ram_w8_l2048_id14_1_0_addr), .ram_w8_l2048_id14_1_0_rdata(ram_w8_l2048_id14_1_0_rdata), .ram_w8_l2048_id14_1_0_wdata(8'h00), .ram_w8_l2048_id14_1_0_wenable(1'h0), .ram_w8_l2048_id14_1_1_addr(ram_w8_l2048_id14_1_1_addr), .ram_w8_l2048_id14_1_1_rdata(ram_w8_l2048_id14_1_1_rdata), .ram_w8_l2048_id14_1_1_wdata(ram_w8_l2048_id14_1_1_wdata), .ram_w8_l2048_id14_1_1_wenable(ram_w8_l2048_id14_1_1_wenable) );
  ram_w8_l2048_id14_2 inst_ram_w8_l2048_id14_2 ( .CLK(CLK), .ram_w8_l2048_id14_2_0_addr(ram_w8_l2048_id14_2_0_addr), .ram_w8_l2048_id14_2_0_rdata(ram_w8_l2048_id14_2_0_rdata), .ram_w8_l2048_id14_2_0_wdata(8'h00), .ram_w8_l2048_id14_2_0_wenable(1'h0), .ram_w8_l2048_id14_2_1_addr(ram_w8_l2048_id14_2_1_addr), .ram_w8_l2048_id14_2_1_rdata(ram_w8_l2048_id14_2_1_rdata), .ram_w8_l2048_id14_2_1_wdata(ram_w8_l2048_id14_2_1_wdata), .ram_w8_l2048_id14_2_1_wenable(ram_w8_l2048_id14_2_1_wenable) );
  ram_w8_l2048_id14_3 inst_ram_w8_l2048_id14_3 ( .CLK(CLK), .ram_w8_l2048_id14_3_0_addr(ram_w8_l2048_id14_3_0_addr), .ram_w8_l2048_id14_3_0_rdata(ram_w8_l2048_id14_3_0_rdata), .ram_w8_l2048_id14_3_0_wdata(8'h00), .ram_w8_l2048_id14_3_0_wenable(1'h0), .ram_w8_l2048_id14_3_1_addr(ram_w8_l2048_id14_3_1_addr), .ram_w8_l2048_id14_3_1_rdata(ram_w8_l2048_id14_3_1_rdata), .ram_w8_l2048_id14_3_1_wdata(ram_w8_l2048_id14_3_1_wdata), .ram_w8_l2048_id14_3_1_wenable(ram_w8_l2048_id14_3_1_wenable) );
  ram_w8_l2048_id15_0 inst_ram_w8_l2048_id15_0 ( .CLK(CLK), .ram_w8_l2048_id15_0_0_addr(ram_w8_l2048_id15_0_0_addr), .ram_w8_l2048_id15_0_0_rdata(ram_w8_l2048_id15_0_0_rdata), .ram_w8_l2048_id15_0_0_wdata(8'h00), .ram_w8_l2048_id15_0_0_wenable(1'h0), .ram_w8_l2048_id15_0_1_addr(ram_w8_l2048_id15_0_1_addr), .ram_w8_l2048_id15_0_1_rdata(ram_w8_l2048_id15_0_1_rdata), .ram_w8_l2048_id15_0_1_wdata(ram_w8_l2048_id15_0_1_wdata), .ram_w8_l2048_id15_0_1_wenable(ram_w8_l2048_id15_0_1_wenable) );
  ram_w8_l2048_id15_1 inst_ram_w8_l2048_id15_1 ( .CLK(CLK), .ram_w8_l2048_id15_1_0_addr(ram_w8_l2048_id15_1_0_addr), .ram_w8_l2048_id15_1_0_rdata(ram_w8_l2048_id15_1_0_rdata), .ram_w8_l2048_id15_1_0_wdata(8'h00), .ram_w8_l2048_id15_1_0_wenable(1'h0), .ram_w8_l2048_id15_1_1_addr(ram_w8_l2048_id15_1_1_addr), .ram_w8_l2048_id15_1_1_rdata(ram_w8_l2048_id15_1_1_rdata), .ram_w8_l2048_id15_1_1_wdata(ram_w8_l2048_id15_1_1_wdata), .ram_w8_l2048_id15_1_1_wenable(ram_w8_l2048_id15_1_1_wenable) );
  ram_w8_l2048_id15_2 inst_ram_w8_l2048_id15_2 ( .CLK(CLK), .ram_w8_l2048_id15_2_0_addr(ram_w8_l2048_id15_2_0_addr), .ram_w8_l2048_id15_2_0_rdata(ram_w8_l2048_id15_2_0_rdata), .ram_w8_l2048_id15_2_0_wdata(8'h00), .ram_w8_l2048_id15_2_0_wenable(1'h0), .ram_w8_l2048_id15_2_1_addr(ram_w8_l2048_id15_2_1_addr), .ram_w8_l2048_id15_2_1_rdata(ram_w8_l2048_id15_2_1_rdata), .ram_w8_l2048_id15_2_1_wdata(ram_w8_l2048_id15_2_1_wdata), .ram_w8_l2048_id15_2_1_wenable(ram_w8_l2048_id15_2_1_wenable) );
  ram_w8_l2048_id15_3 inst_ram_w8_l2048_id15_3 ( .CLK(CLK), .ram_w8_l2048_id15_3_0_addr(ram_w8_l2048_id15_3_0_addr), .ram_w8_l2048_id15_3_0_rdata(ram_w8_l2048_id15_3_0_rdata), .ram_w8_l2048_id15_3_0_wdata(8'h00), .ram_w8_l2048_id15_3_0_wenable(1'h0), .ram_w8_l2048_id15_3_1_addr(ram_w8_l2048_id15_3_1_addr), .ram_w8_l2048_id15_3_1_rdata(ram_w8_l2048_id15_3_1_rdata), .ram_w8_l2048_id15_3_1_wdata(ram_w8_l2048_id15_3_1_wdata), .ram_w8_l2048_id15_3_1_wenable(ram_w8_l2048_id15_3_1_wenable) );
  ram_w8_l2048_id16_0 inst_ram_w8_l2048_id16_0 ( .CLK(CLK), .ram_w8_l2048_id16_0_0_addr(ram_w8_l2048_id16_0_0_addr), .ram_w8_l2048_id16_0_0_rdata(ram_w8_l2048_id16_0_0_rdata), .ram_w8_l2048_id16_0_0_wdata(8'h00), .ram_w8_l2048_id16_0_0_wenable(1'h0), .ram_w8_l2048_id16_0_1_addr(ram_w8_l2048_id16_0_1_addr), .ram_w8_l2048_id16_0_1_rdata(ram_w8_l2048_id16_0_1_rdata), .ram_w8_l2048_id16_0_1_wdata(ram_w8_l2048_id16_0_1_wdata), .ram_w8_l2048_id16_0_1_wenable(ram_w8_l2048_id16_0_1_wenable) );
  ram_w8_l2048_id16_1 inst_ram_w8_l2048_id16_1 ( .CLK(CLK), .ram_w8_l2048_id16_1_0_addr(ram_w8_l2048_id16_1_0_addr), .ram_w8_l2048_id16_1_0_rdata(ram_w8_l2048_id16_1_0_rdata), .ram_w8_l2048_id16_1_0_wdata(8'h00), .ram_w8_l2048_id16_1_0_wenable(1'h0), .ram_w8_l2048_id16_1_1_addr(ram_w8_l2048_id16_1_1_addr), .ram_w8_l2048_id16_1_1_rdata(ram_w8_l2048_id16_1_1_rdata), .ram_w8_l2048_id16_1_1_wdata(ram_w8_l2048_id16_1_1_wdata), .ram_w8_l2048_id16_1_1_wenable(ram_w8_l2048_id16_1_1_wenable) );
  ram_w8_l2048_id16_2 inst_ram_w8_l2048_id16_2 ( .CLK(CLK), .ram_w8_l2048_id16_2_0_addr(ram_w8_l2048_id16_2_0_addr), .ram_w8_l2048_id16_2_0_rdata(ram_w8_l2048_id16_2_0_rdata), .ram_w8_l2048_id16_2_0_wdata(8'h00), .ram_w8_l2048_id16_2_0_wenable(1'h0), .ram_w8_l2048_id16_2_1_addr(ram_w8_l2048_id16_2_1_addr), .ram_w8_l2048_id16_2_1_rdata(ram_w8_l2048_id16_2_1_rdata), .ram_w8_l2048_id16_2_1_wdata(ram_w8_l2048_id16_2_1_wdata), .ram_w8_l2048_id16_2_1_wenable(ram_w8_l2048_id16_2_1_wenable) );
  ram_w8_l2048_id16_3 inst_ram_w8_l2048_id16_3 ( .CLK(CLK), .ram_w8_l2048_id16_3_0_addr(ram_w8_l2048_id16_3_0_addr), .ram_w8_l2048_id16_3_0_rdata(ram_w8_l2048_id16_3_0_rdata), .ram_w8_l2048_id16_3_0_wdata(8'h00), .ram_w8_l2048_id16_3_0_wenable(1'h0), .ram_w8_l2048_id16_3_1_addr(ram_w8_l2048_id16_3_1_addr), .ram_w8_l2048_id16_3_1_rdata(ram_w8_l2048_id16_3_1_rdata), .ram_w8_l2048_id16_3_1_wdata(ram_w8_l2048_id16_3_1_wdata), .ram_w8_l2048_id16_3_1_wenable(ram_w8_l2048_id16_3_1_wenable) );
  ram_w8_l2048_id17_0 inst_ram_w8_l2048_id17_0 ( .CLK(CLK), .ram_w8_l2048_id17_0_0_addr(ram_w8_l2048_id17_0_0_addr), .ram_w8_l2048_id17_0_0_rdata(ram_w8_l2048_id17_0_0_rdata), .ram_w8_l2048_id17_0_0_wdata(8'h00), .ram_w8_l2048_id17_0_0_wenable(1'h0), .ram_w8_l2048_id17_0_1_addr(ram_w8_l2048_id17_0_1_addr), .ram_w8_l2048_id17_0_1_rdata(ram_w8_l2048_id17_0_1_rdata), .ram_w8_l2048_id17_0_1_wdata(ram_w8_l2048_id17_0_1_wdata), .ram_w8_l2048_id17_0_1_wenable(ram_w8_l2048_id17_0_1_wenable) );
  ram_w8_l2048_id17_1 inst_ram_w8_l2048_id17_1 ( .CLK(CLK), .ram_w8_l2048_id17_1_0_addr(ram_w8_l2048_id17_1_0_addr), .ram_w8_l2048_id17_1_0_rdata(ram_w8_l2048_id17_1_0_rdata), .ram_w8_l2048_id17_1_0_wdata(8'h00), .ram_w8_l2048_id17_1_0_wenable(1'h0), .ram_w8_l2048_id17_1_1_addr(ram_w8_l2048_id17_1_1_addr), .ram_w8_l2048_id17_1_1_rdata(ram_w8_l2048_id17_1_1_rdata), .ram_w8_l2048_id17_1_1_wdata(ram_w8_l2048_id17_1_1_wdata), .ram_w8_l2048_id17_1_1_wenable(ram_w8_l2048_id17_1_1_wenable) );
  ram_w8_l2048_id17_2 inst_ram_w8_l2048_id17_2 ( .CLK(CLK), .ram_w8_l2048_id17_2_0_addr(ram_w8_l2048_id17_2_0_addr), .ram_w8_l2048_id17_2_0_rdata(ram_w8_l2048_id17_2_0_rdata), .ram_w8_l2048_id17_2_0_wdata(8'h00), .ram_w8_l2048_id17_2_0_wenable(1'h0), .ram_w8_l2048_id17_2_1_addr(ram_w8_l2048_id17_2_1_addr), .ram_w8_l2048_id17_2_1_rdata(ram_w8_l2048_id17_2_1_rdata), .ram_w8_l2048_id17_2_1_wdata(ram_w8_l2048_id17_2_1_wdata), .ram_w8_l2048_id17_2_1_wenable(ram_w8_l2048_id17_2_1_wenable) );
  ram_w8_l2048_id17_3 inst_ram_w8_l2048_id17_3 ( .CLK(CLK), .ram_w8_l2048_id17_3_0_addr(ram_w8_l2048_id17_3_0_addr), .ram_w8_l2048_id17_3_0_rdata(ram_w8_l2048_id17_3_0_rdata), .ram_w8_l2048_id17_3_0_wdata(8'h00), .ram_w8_l2048_id17_3_0_wenable(1'h0), .ram_w8_l2048_id17_3_1_addr(ram_w8_l2048_id17_3_1_addr), .ram_w8_l2048_id17_3_1_rdata(ram_w8_l2048_id17_3_1_rdata), .ram_w8_l2048_id17_3_1_wdata(ram_w8_l2048_id17_3_1_wdata), .ram_w8_l2048_id17_3_1_wenable(ram_w8_l2048_id17_3_1_wenable) );
  ram_w8_l2048_id18_0 inst_ram_w8_l2048_id18_0 ( .CLK(CLK), .ram_w8_l2048_id18_0_0_addr(ram_w8_l2048_id18_0_0_addr), .ram_w8_l2048_id18_0_0_rdata(ram_w8_l2048_id18_0_0_rdata), .ram_w8_l2048_id18_0_0_wdata(8'h00), .ram_w8_l2048_id18_0_0_wenable(1'h0), .ram_w8_l2048_id18_0_1_addr(ram_w8_l2048_id18_0_1_addr), .ram_w8_l2048_id18_0_1_rdata(ram_w8_l2048_id18_0_1_rdata), .ram_w8_l2048_id18_0_1_wdata(ram_w8_l2048_id18_0_1_wdata), .ram_w8_l2048_id18_0_1_wenable(ram_w8_l2048_id18_0_1_wenable) );
  ram_w8_l2048_id18_1 inst_ram_w8_l2048_id18_1 ( .CLK(CLK), .ram_w8_l2048_id18_1_0_addr(ram_w8_l2048_id18_1_0_addr), .ram_w8_l2048_id18_1_0_rdata(ram_w8_l2048_id18_1_0_rdata), .ram_w8_l2048_id18_1_0_wdata(8'h00), .ram_w8_l2048_id18_1_0_wenable(1'h0), .ram_w8_l2048_id18_1_1_addr(ram_w8_l2048_id18_1_1_addr), .ram_w8_l2048_id18_1_1_rdata(ram_w8_l2048_id18_1_1_rdata), .ram_w8_l2048_id18_1_1_wdata(ram_w8_l2048_id18_1_1_wdata), .ram_w8_l2048_id18_1_1_wenable(ram_w8_l2048_id18_1_1_wenable) );
  ram_w8_l2048_id18_2 inst_ram_w8_l2048_id18_2 ( .CLK(CLK), .ram_w8_l2048_id18_2_0_addr(ram_w8_l2048_id18_2_0_addr), .ram_w8_l2048_id18_2_0_rdata(ram_w8_l2048_id18_2_0_rdata), .ram_w8_l2048_id18_2_0_wdata(8'h00), .ram_w8_l2048_id18_2_0_wenable(1'h0), .ram_w8_l2048_id18_2_1_addr(ram_w8_l2048_id18_2_1_addr), .ram_w8_l2048_id18_2_1_rdata(ram_w8_l2048_id18_2_1_rdata), .ram_w8_l2048_id18_2_1_wdata(ram_w8_l2048_id18_2_1_wdata), .ram_w8_l2048_id18_2_1_wenable(ram_w8_l2048_id18_2_1_wenable) );
  ram_w8_l2048_id18_3 inst_ram_w8_l2048_id18_3 ( .CLK(CLK), .ram_w8_l2048_id18_3_0_addr(ram_w8_l2048_id18_3_0_addr), .ram_w8_l2048_id18_3_0_rdata(ram_w8_l2048_id18_3_0_rdata), .ram_w8_l2048_id18_3_0_wdata(8'h00), .ram_w8_l2048_id18_3_0_wenable(1'h0), .ram_w8_l2048_id18_3_1_addr(ram_w8_l2048_id18_3_1_addr), .ram_w8_l2048_id18_3_1_rdata(ram_w8_l2048_id18_3_1_rdata), .ram_w8_l2048_id18_3_1_wdata(ram_w8_l2048_id18_3_1_wdata), .ram_w8_l2048_id18_3_1_wenable(ram_w8_l2048_id18_3_1_wenable) );
  ram_w8_l2048_id19_0 inst_ram_w8_l2048_id19_0 ( .CLK(CLK), .ram_w8_l2048_id19_0_0_addr(ram_w8_l2048_id19_0_0_addr), .ram_w8_l2048_id19_0_0_rdata(ram_w8_l2048_id19_0_0_rdata), .ram_w8_l2048_id19_0_0_wdata(ram_w8_l2048_id19_0_0_wdata), .ram_w8_l2048_id19_0_0_wenable(ram_w8_l2048_id19_0_0_wenable), .ram_w8_l2048_id19_0_1_addr(ram_w8_l2048_id19_0_1_addr), .ram_w8_l2048_id19_0_1_rdata(ram_w8_l2048_id19_0_1_rdata), .ram_w8_l2048_id19_0_1_wdata(8'h00), .ram_w8_l2048_id19_0_1_wenable(1'h0) );
  ram_w8_l2048_id19_1 inst_ram_w8_l2048_id19_1 ( .CLK(CLK), .ram_w8_l2048_id19_1_0_addr(ram_w8_l2048_id19_1_0_addr), .ram_w8_l2048_id19_1_0_rdata(ram_w8_l2048_id19_1_0_rdata), .ram_w8_l2048_id19_1_0_wdata(ram_w8_l2048_id19_1_0_wdata), .ram_w8_l2048_id19_1_0_wenable(ram_w8_l2048_id19_1_0_wenable), .ram_w8_l2048_id19_1_1_addr(ram_w8_l2048_id19_1_1_addr), .ram_w8_l2048_id19_1_1_rdata(ram_w8_l2048_id19_1_1_rdata), .ram_w8_l2048_id19_1_1_wdata(8'h00), .ram_w8_l2048_id19_1_1_wenable(1'h0) );
  ram_w8_l2048_id19_2 inst_ram_w8_l2048_id19_2 ( .CLK(CLK), .ram_w8_l2048_id19_2_0_addr(ram_w8_l2048_id19_2_0_addr), .ram_w8_l2048_id19_2_0_rdata(ram_w8_l2048_id19_2_0_rdata), .ram_w8_l2048_id19_2_0_wdata(ram_w8_l2048_id19_2_0_wdata), .ram_w8_l2048_id19_2_0_wenable(ram_w8_l2048_id19_2_0_wenable), .ram_w8_l2048_id19_2_1_addr(ram_w8_l2048_id19_2_1_addr), .ram_w8_l2048_id19_2_1_rdata(ram_w8_l2048_id19_2_1_rdata), .ram_w8_l2048_id19_2_1_wdata(8'h00), .ram_w8_l2048_id19_2_1_wenable(1'h0) );
  ram_w8_l2048_id19_3 inst_ram_w8_l2048_id19_3 ( .CLK(CLK), .ram_w8_l2048_id19_3_0_addr(ram_w8_l2048_id19_3_0_addr), .ram_w8_l2048_id19_3_0_rdata(ram_w8_l2048_id19_3_0_rdata), .ram_w8_l2048_id19_3_0_wdata(ram_w8_l2048_id19_3_0_wdata), .ram_w8_l2048_id19_3_0_wenable(ram_w8_l2048_id19_3_0_wenable), .ram_w8_l2048_id19_3_1_addr(ram_w8_l2048_id19_3_1_addr), .ram_w8_l2048_id19_3_1_rdata(ram_w8_l2048_id19_3_1_rdata), .ram_w8_l2048_id19_3_1_wdata(8'h00), .ram_w8_l2048_id19_3_1_wenable(1'h0) );
  ram_w8_l2048_id1_0 inst_ram_w8_l2048_id1_0 ( .CLK(CLK), .ram_w8_l2048_id1_0_0_addr(ram_w8_l2048_id1_0_0_addr), .ram_w8_l2048_id1_0_0_rdata(ram_w8_l2048_id1_0_0_rdata), .ram_w8_l2048_id1_0_0_wdata(ram_w8_l2048_id1_0_0_wdata), .ram_w8_l2048_id1_0_0_wenable(ram_w8_l2048_id1_0_0_wenable), .ram_w8_l2048_id1_0_1_addr(ram_w8_l2048_id1_0_1_addr), .ram_w8_l2048_id1_0_1_rdata(ram_w8_l2048_id1_0_1_rdata), .ram_w8_l2048_id1_0_1_wdata(ram_w8_l2048_id1_0_1_wdata), .ram_w8_l2048_id1_0_1_wenable(ram_w8_l2048_id1_0_1_wenable) );
  ram_w8_l2048_id1_1 inst_ram_w8_l2048_id1_1 ( .CLK(CLK), .ram_w8_l2048_id1_1_0_addr(ram_w8_l2048_id1_1_0_addr), .ram_w8_l2048_id1_1_0_rdata(ram_w8_l2048_id1_1_0_rdata), .ram_w8_l2048_id1_1_0_wdata(ram_w8_l2048_id1_1_0_wdata), .ram_w8_l2048_id1_1_0_wenable(ram_w8_l2048_id1_1_0_wenable), .ram_w8_l2048_id1_1_1_addr(ram_w8_l2048_id1_1_1_addr), .ram_w8_l2048_id1_1_1_rdata(ram_w8_l2048_id1_1_1_rdata), .ram_w8_l2048_id1_1_1_wdata(ram_w8_l2048_id1_1_1_wdata), .ram_w8_l2048_id1_1_1_wenable(ram_w8_l2048_id1_1_1_wenable) );
  ram_w8_l2048_id1_2 inst_ram_w8_l2048_id1_2 ( .CLK(CLK), .ram_w8_l2048_id1_2_0_addr(ram_w8_l2048_id1_2_0_addr), .ram_w8_l2048_id1_2_0_rdata(ram_w8_l2048_id1_2_0_rdata), .ram_w8_l2048_id1_2_0_wdata(ram_w8_l2048_id1_2_0_wdata), .ram_w8_l2048_id1_2_0_wenable(ram_w8_l2048_id1_2_0_wenable), .ram_w8_l2048_id1_2_1_addr(ram_w8_l2048_id1_2_1_addr), .ram_w8_l2048_id1_2_1_rdata(ram_w8_l2048_id1_2_1_rdata), .ram_w8_l2048_id1_2_1_wdata(ram_w8_l2048_id1_2_1_wdata), .ram_w8_l2048_id1_2_1_wenable(ram_w8_l2048_id1_2_1_wenable) );
  ram_w8_l2048_id1_3 inst_ram_w8_l2048_id1_3 ( .CLK(CLK), .ram_w8_l2048_id1_3_0_addr(ram_w8_l2048_id1_3_0_addr), .ram_w8_l2048_id1_3_0_rdata(ram_w8_l2048_id1_3_0_rdata), .ram_w8_l2048_id1_3_0_wdata(ram_w8_l2048_id1_3_0_wdata), .ram_w8_l2048_id1_3_0_wenable(ram_w8_l2048_id1_3_0_wenable), .ram_w8_l2048_id1_3_1_addr(ram_w8_l2048_id1_3_1_addr), .ram_w8_l2048_id1_3_1_rdata(ram_w8_l2048_id1_3_1_rdata), .ram_w8_l2048_id1_3_1_wdata(ram_w8_l2048_id1_3_1_wdata), .ram_w8_l2048_id1_3_1_wenable(ram_w8_l2048_id1_3_1_wenable) );
  ram_w8_l2048_id2_0 inst_ram_w8_l2048_id2_0 ( .CLK(CLK), .ram_w8_l2048_id2_0_0_addr(ram_w8_l2048_id2_0_0_addr), .ram_w8_l2048_id2_0_0_rdata(ram_w8_l2048_id2_0_0_rdata), .ram_w8_l2048_id2_0_0_wdata(8'h00), .ram_w8_l2048_id2_0_0_wenable(1'h0), .ram_w8_l2048_id2_0_1_addr(ram_w8_l2048_id2_0_1_addr), .ram_w8_l2048_id2_0_1_rdata(ram_w8_l2048_id2_0_1_rdata), .ram_w8_l2048_id2_0_1_wdata(ram_w8_l2048_id2_0_1_wdata), .ram_w8_l2048_id2_0_1_wenable(ram_w8_l2048_id2_0_1_wenable) );
  ram_w8_l2048_id2_1 inst_ram_w8_l2048_id2_1 ( .CLK(CLK), .ram_w8_l2048_id2_1_0_addr(ram_w8_l2048_id2_1_0_addr), .ram_w8_l2048_id2_1_0_rdata(ram_w8_l2048_id2_1_0_rdata), .ram_w8_l2048_id2_1_0_wdata(8'h00), .ram_w8_l2048_id2_1_0_wenable(1'h0), .ram_w8_l2048_id2_1_1_addr(ram_w8_l2048_id2_1_1_addr), .ram_w8_l2048_id2_1_1_rdata(ram_w8_l2048_id2_1_1_rdata), .ram_w8_l2048_id2_1_1_wdata(ram_w8_l2048_id2_1_1_wdata), .ram_w8_l2048_id2_1_1_wenable(ram_w8_l2048_id2_1_1_wenable) );
  ram_w8_l2048_id2_2 inst_ram_w8_l2048_id2_2 ( .CLK(CLK), .ram_w8_l2048_id2_2_0_addr(ram_w8_l2048_id2_2_0_addr), .ram_w8_l2048_id2_2_0_rdata(ram_w8_l2048_id2_2_0_rdata), .ram_w8_l2048_id2_2_0_wdata(8'h00), .ram_w8_l2048_id2_2_0_wenable(1'h0), .ram_w8_l2048_id2_2_1_addr(ram_w8_l2048_id2_2_1_addr), .ram_w8_l2048_id2_2_1_rdata(ram_w8_l2048_id2_2_1_rdata), .ram_w8_l2048_id2_2_1_wdata(ram_w8_l2048_id2_2_1_wdata), .ram_w8_l2048_id2_2_1_wenable(ram_w8_l2048_id2_2_1_wenable) );
  ram_w8_l2048_id2_3 inst_ram_w8_l2048_id2_3 ( .CLK(CLK), .ram_w8_l2048_id2_3_0_addr(ram_w8_l2048_id2_3_0_addr), .ram_w8_l2048_id2_3_0_rdata(ram_w8_l2048_id2_3_0_rdata), .ram_w8_l2048_id2_3_0_wdata(8'h00), .ram_w8_l2048_id2_3_0_wenable(1'h0), .ram_w8_l2048_id2_3_1_addr(ram_w8_l2048_id2_3_1_addr), .ram_w8_l2048_id2_3_1_rdata(ram_w8_l2048_id2_3_1_rdata), .ram_w8_l2048_id2_3_1_wdata(ram_w8_l2048_id2_3_1_wdata), .ram_w8_l2048_id2_3_1_wenable(ram_w8_l2048_id2_3_1_wenable) );
  ram_w8_l2048_id3_0 inst_ram_w8_l2048_id3_0 ( .CLK(CLK), .ram_w8_l2048_id3_0_0_addr(ram_w8_l2048_id3_0_0_addr), .ram_w8_l2048_id3_0_0_rdata(ram_w8_l2048_id3_0_0_rdata), .ram_w8_l2048_id3_0_0_wdata(8'h00), .ram_w8_l2048_id3_0_0_wenable(1'h0), .ram_w8_l2048_id3_0_1_addr(ram_w8_l2048_id3_0_1_addr), .ram_w8_l2048_id3_0_1_rdata(ram_w8_l2048_id3_0_1_rdata), .ram_w8_l2048_id3_0_1_wdata(ram_w8_l2048_id3_0_1_wdata), .ram_w8_l2048_id3_0_1_wenable(ram_w8_l2048_id3_0_1_wenable) );
  ram_w8_l2048_id3_1 inst_ram_w8_l2048_id3_1 ( .CLK(CLK), .ram_w8_l2048_id3_1_0_addr(ram_w8_l2048_id3_1_0_addr), .ram_w8_l2048_id3_1_0_rdata(ram_w8_l2048_id3_1_0_rdata), .ram_w8_l2048_id3_1_0_wdata(8'h00), .ram_w8_l2048_id3_1_0_wenable(1'h0), .ram_w8_l2048_id3_1_1_addr(ram_w8_l2048_id3_1_1_addr), .ram_w8_l2048_id3_1_1_rdata(ram_w8_l2048_id3_1_1_rdata), .ram_w8_l2048_id3_1_1_wdata(ram_w8_l2048_id3_1_1_wdata), .ram_w8_l2048_id3_1_1_wenable(ram_w8_l2048_id3_1_1_wenable) );
  ram_w8_l2048_id3_2 inst_ram_w8_l2048_id3_2 ( .CLK(CLK), .ram_w8_l2048_id3_2_0_addr(ram_w8_l2048_id3_2_0_addr), .ram_w8_l2048_id3_2_0_rdata(ram_w8_l2048_id3_2_0_rdata), .ram_w8_l2048_id3_2_0_wdata(8'h00), .ram_w8_l2048_id3_2_0_wenable(1'h0), .ram_w8_l2048_id3_2_1_addr(ram_w8_l2048_id3_2_1_addr), .ram_w8_l2048_id3_2_1_rdata(ram_w8_l2048_id3_2_1_rdata), .ram_w8_l2048_id3_2_1_wdata(ram_w8_l2048_id3_2_1_wdata), .ram_w8_l2048_id3_2_1_wenable(ram_w8_l2048_id3_2_1_wenable) );
  ram_w8_l2048_id3_3 inst_ram_w8_l2048_id3_3 ( .CLK(CLK), .ram_w8_l2048_id3_3_0_addr(ram_w8_l2048_id3_3_0_addr), .ram_w8_l2048_id3_3_0_rdata(ram_w8_l2048_id3_3_0_rdata), .ram_w8_l2048_id3_3_0_wdata(8'h00), .ram_w8_l2048_id3_3_0_wenable(1'h0), .ram_w8_l2048_id3_3_1_addr(ram_w8_l2048_id3_3_1_addr), .ram_w8_l2048_id3_3_1_rdata(ram_w8_l2048_id3_3_1_rdata), .ram_w8_l2048_id3_3_1_wdata(ram_w8_l2048_id3_3_1_wdata), .ram_w8_l2048_id3_3_1_wenable(ram_w8_l2048_id3_3_1_wenable) );
  ram_w8_l2048_id4_0 inst_ram_w8_l2048_id4_0 ( .CLK(CLK), .ram_w8_l2048_id4_0_0_addr(ram_w8_l2048_id4_0_0_addr), .ram_w8_l2048_id4_0_0_rdata(ram_w8_l2048_id4_0_0_rdata), .ram_w8_l2048_id4_0_0_wdata(8'h00), .ram_w8_l2048_id4_0_0_wenable(1'h0), .ram_w8_l2048_id4_0_1_addr(ram_w8_l2048_id4_0_1_addr), .ram_w8_l2048_id4_0_1_rdata(ram_w8_l2048_id4_0_1_rdata), .ram_w8_l2048_id4_0_1_wdata(ram_w8_l2048_id4_0_1_wdata), .ram_w8_l2048_id4_0_1_wenable(ram_w8_l2048_id4_0_1_wenable) );
  ram_w8_l2048_id4_1 inst_ram_w8_l2048_id4_1 ( .CLK(CLK), .ram_w8_l2048_id4_1_0_addr(ram_w8_l2048_id4_1_0_addr), .ram_w8_l2048_id4_1_0_rdata(ram_w8_l2048_id4_1_0_rdata), .ram_w8_l2048_id4_1_0_wdata(8'h00), .ram_w8_l2048_id4_1_0_wenable(1'h0), .ram_w8_l2048_id4_1_1_addr(ram_w8_l2048_id4_1_1_addr), .ram_w8_l2048_id4_1_1_rdata(ram_w8_l2048_id4_1_1_rdata), .ram_w8_l2048_id4_1_1_wdata(ram_w8_l2048_id4_1_1_wdata), .ram_w8_l2048_id4_1_1_wenable(ram_w8_l2048_id4_1_1_wenable) );
  ram_w8_l2048_id4_2 inst_ram_w8_l2048_id4_2 ( .CLK(CLK), .ram_w8_l2048_id4_2_0_addr(ram_w8_l2048_id4_2_0_addr), .ram_w8_l2048_id4_2_0_rdata(ram_w8_l2048_id4_2_0_rdata), .ram_w8_l2048_id4_2_0_wdata(8'h00), .ram_w8_l2048_id4_2_0_wenable(1'h0), .ram_w8_l2048_id4_2_1_addr(ram_w8_l2048_id4_2_1_addr), .ram_w8_l2048_id4_2_1_rdata(ram_w8_l2048_id4_2_1_rdata), .ram_w8_l2048_id4_2_1_wdata(ram_w8_l2048_id4_2_1_wdata), .ram_w8_l2048_id4_2_1_wenable(ram_w8_l2048_id4_2_1_wenable) );
  ram_w8_l2048_id4_3 inst_ram_w8_l2048_id4_3 ( .CLK(CLK), .ram_w8_l2048_id4_3_0_addr(ram_w8_l2048_id4_3_0_addr), .ram_w8_l2048_id4_3_0_rdata(ram_w8_l2048_id4_3_0_rdata), .ram_w8_l2048_id4_3_0_wdata(8'h00), .ram_w8_l2048_id4_3_0_wenable(1'h0), .ram_w8_l2048_id4_3_1_addr(ram_w8_l2048_id4_3_1_addr), .ram_w8_l2048_id4_3_1_rdata(ram_w8_l2048_id4_3_1_rdata), .ram_w8_l2048_id4_3_1_wdata(ram_w8_l2048_id4_3_1_wdata), .ram_w8_l2048_id4_3_1_wenable(ram_w8_l2048_id4_3_1_wenable) );
  ram_w8_l2048_id5_0 inst_ram_w8_l2048_id5_0 ( .CLK(CLK), .ram_w8_l2048_id5_0_0_addr(ram_w8_l2048_id5_0_0_addr), .ram_w8_l2048_id5_0_0_rdata(ram_w8_l2048_id5_0_0_rdata), .ram_w8_l2048_id5_0_0_wdata(8'h00), .ram_w8_l2048_id5_0_0_wenable(1'h0), .ram_w8_l2048_id5_0_1_addr(ram_w8_l2048_id5_0_1_addr), .ram_w8_l2048_id5_0_1_rdata(ram_w8_l2048_id5_0_1_rdata), .ram_w8_l2048_id5_0_1_wdata(ram_w8_l2048_id5_0_1_wdata), .ram_w8_l2048_id5_0_1_wenable(ram_w8_l2048_id5_0_1_wenable) );
  ram_w8_l2048_id5_1 inst_ram_w8_l2048_id5_1 ( .CLK(CLK), .ram_w8_l2048_id5_1_0_addr(ram_w8_l2048_id5_1_0_addr), .ram_w8_l2048_id5_1_0_rdata(ram_w8_l2048_id5_1_0_rdata), .ram_w8_l2048_id5_1_0_wdata(8'h00), .ram_w8_l2048_id5_1_0_wenable(1'h0), .ram_w8_l2048_id5_1_1_addr(ram_w8_l2048_id5_1_1_addr), .ram_w8_l2048_id5_1_1_rdata(ram_w8_l2048_id5_1_1_rdata), .ram_w8_l2048_id5_1_1_wdata(ram_w8_l2048_id5_1_1_wdata), .ram_w8_l2048_id5_1_1_wenable(ram_w8_l2048_id5_1_1_wenable) );
  ram_w8_l2048_id5_2 inst_ram_w8_l2048_id5_2 ( .CLK(CLK), .ram_w8_l2048_id5_2_0_addr(ram_w8_l2048_id5_2_0_addr), .ram_w8_l2048_id5_2_0_rdata(ram_w8_l2048_id5_2_0_rdata), .ram_w8_l2048_id5_2_0_wdata(8'h00), .ram_w8_l2048_id5_2_0_wenable(1'h0), .ram_w8_l2048_id5_2_1_addr(ram_w8_l2048_id5_2_1_addr), .ram_w8_l2048_id5_2_1_rdata(ram_w8_l2048_id5_2_1_rdata), .ram_w8_l2048_id5_2_1_wdata(ram_w8_l2048_id5_2_1_wdata), .ram_w8_l2048_id5_2_1_wenable(ram_w8_l2048_id5_2_1_wenable) );
  ram_w8_l2048_id5_3 inst_ram_w8_l2048_id5_3 ( .CLK(CLK), .ram_w8_l2048_id5_3_0_addr(ram_w8_l2048_id5_3_0_addr), .ram_w8_l2048_id5_3_0_rdata(ram_w8_l2048_id5_3_0_rdata), .ram_w8_l2048_id5_3_0_wdata(8'h00), .ram_w8_l2048_id5_3_0_wenable(1'h0), .ram_w8_l2048_id5_3_1_addr(ram_w8_l2048_id5_3_1_addr), .ram_w8_l2048_id5_3_1_rdata(ram_w8_l2048_id5_3_1_rdata), .ram_w8_l2048_id5_3_1_wdata(ram_w8_l2048_id5_3_1_wdata), .ram_w8_l2048_id5_3_1_wenable(ram_w8_l2048_id5_3_1_wenable) );
  ram_w8_l2048_id6_0 inst_ram_w8_l2048_id6_0 ( .CLK(CLK), .ram_w8_l2048_id6_0_0_addr(ram_w8_l2048_id6_0_0_addr), .ram_w8_l2048_id6_0_0_rdata(ram_w8_l2048_id6_0_0_rdata), .ram_w8_l2048_id6_0_0_wdata(8'h00), .ram_w8_l2048_id6_0_0_wenable(1'h0), .ram_w8_l2048_id6_0_1_addr(ram_w8_l2048_id6_0_1_addr), .ram_w8_l2048_id6_0_1_rdata(ram_w8_l2048_id6_0_1_rdata), .ram_w8_l2048_id6_0_1_wdata(ram_w8_l2048_id6_0_1_wdata), .ram_w8_l2048_id6_0_1_wenable(ram_w8_l2048_id6_0_1_wenable) );
  ram_w8_l2048_id6_1 inst_ram_w8_l2048_id6_1 ( .CLK(CLK), .ram_w8_l2048_id6_1_0_addr(ram_w8_l2048_id6_1_0_addr), .ram_w8_l2048_id6_1_0_rdata(ram_w8_l2048_id6_1_0_rdata), .ram_w8_l2048_id6_1_0_wdata(8'h00), .ram_w8_l2048_id6_1_0_wenable(1'h0), .ram_w8_l2048_id6_1_1_addr(ram_w8_l2048_id6_1_1_addr), .ram_w8_l2048_id6_1_1_rdata(ram_w8_l2048_id6_1_1_rdata), .ram_w8_l2048_id6_1_1_wdata(ram_w8_l2048_id6_1_1_wdata), .ram_w8_l2048_id6_1_1_wenable(ram_w8_l2048_id6_1_1_wenable) );
  ram_w8_l2048_id6_2 inst_ram_w8_l2048_id6_2 ( .CLK(CLK), .ram_w8_l2048_id6_2_0_addr(ram_w8_l2048_id6_2_0_addr), .ram_w8_l2048_id6_2_0_rdata(ram_w8_l2048_id6_2_0_rdata), .ram_w8_l2048_id6_2_0_wdata(8'h00), .ram_w8_l2048_id6_2_0_wenable(1'h0), .ram_w8_l2048_id6_2_1_addr(ram_w8_l2048_id6_2_1_addr), .ram_w8_l2048_id6_2_1_rdata(ram_w8_l2048_id6_2_1_rdata), .ram_w8_l2048_id6_2_1_wdata(ram_w8_l2048_id6_2_1_wdata), .ram_w8_l2048_id6_2_1_wenable(ram_w8_l2048_id6_2_1_wenable) );
  ram_w8_l2048_id6_3 inst_ram_w8_l2048_id6_3 ( .CLK(CLK), .ram_w8_l2048_id6_3_0_addr(ram_w8_l2048_id6_3_0_addr), .ram_w8_l2048_id6_3_0_rdata(ram_w8_l2048_id6_3_0_rdata), .ram_w8_l2048_id6_3_0_wdata(8'h00), .ram_w8_l2048_id6_3_0_wenable(1'h0), .ram_w8_l2048_id6_3_1_addr(ram_w8_l2048_id6_3_1_addr), .ram_w8_l2048_id6_3_1_rdata(ram_w8_l2048_id6_3_1_rdata), .ram_w8_l2048_id6_3_1_wdata(ram_w8_l2048_id6_3_1_wdata), .ram_w8_l2048_id6_3_1_wenable(ram_w8_l2048_id6_3_1_wenable) );
  ram_w8_l2048_id7_0 inst_ram_w8_l2048_id7_0 ( .CLK(CLK), .ram_w8_l2048_id7_0_0_addr(ram_w8_l2048_id7_0_0_addr), .ram_w8_l2048_id7_0_0_rdata(ram_w8_l2048_id7_0_0_rdata), .ram_w8_l2048_id7_0_0_wdata(8'h00), .ram_w8_l2048_id7_0_0_wenable(1'h0), .ram_w8_l2048_id7_0_1_addr(ram_w8_l2048_id7_0_1_addr), .ram_w8_l2048_id7_0_1_rdata(ram_w8_l2048_id7_0_1_rdata), .ram_w8_l2048_id7_0_1_wdata(ram_w8_l2048_id7_0_1_wdata), .ram_w8_l2048_id7_0_1_wenable(ram_w8_l2048_id7_0_1_wenable) );
  ram_w8_l2048_id7_1 inst_ram_w8_l2048_id7_1 ( .CLK(CLK), .ram_w8_l2048_id7_1_0_addr(ram_w8_l2048_id7_1_0_addr), .ram_w8_l2048_id7_1_0_rdata(ram_w8_l2048_id7_1_0_rdata), .ram_w8_l2048_id7_1_0_wdata(8'h00), .ram_w8_l2048_id7_1_0_wenable(1'h0), .ram_w8_l2048_id7_1_1_addr(ram_w8_l2048_id7_1_1_addr), .ram_w8_l2048_id7_1_1_rdata(ram_w8_l2048_id7_1_1_rdata), .ram_w8_l2048_id7_1_1_wdata(ram_w8_l2048_id7_1_1_wdata), .ram_w8_l2048_id7_1_1_wenable(ram_w8_l2048_id7_1_1_wenable) );
  ram_w8_l2048_id7_2 inst_ram_w8_l2048_id7_2 ( .CLK(CLK), .ram_w8_l2048_id7_2_0_addr(ram_w8_l2048_id7_2_0_addr), .ram_w8_l2048_id7_2_0_rdata(ram_w8_l2048_id7_2_0_rdata), .ram_w8_l2048_id7_2_0_wdata(8'h00), .ram_w8_l2048_id7_2_0_wenable(1'h0), .ram_w8_l2048_id7_2_1_addr(ram_w8_l2048_id7_2_1_addr), .ram_w8_l2048_id7_2_1_rdata(ram_w8_l2048_id7_2_1_rdata), .ram_w8_l2048_id7_2_1_wdata(ram_w8_l2048_id7_2_1_wdata), .ram_w8_l2048_id7_2_1_wenable(ram_w8_l2048_id7_2_1_wenable) );
  ram_w8_l2048_id7_3 inst_ram_w8_l2048_id7_3 ( .CLK(CLK), .ram_w8_l2048_id7_3_0_addr(ram_w8_l2048_id7_3_0_addr), .ram_w8_l2048_id7_3_0_rdata(ram_w8_l2048_id7_3_0_rdata), .ram_w8_l2048_id7_3_0_wdata(8'h00), .ram_w8_l2048_id7_3_0_wenable(1'h0), .ram_w8_l2048_id7_3_1_addr(ram_w8_l2048_id7_3_1_addr), .ram_w8_l2048_id7_3_1_rdata(ram_w8_l2048_id7_3_1_rdata), .ram_w8_l2048_id7_3_1_wdata(ram_w8_l2048_id7_3_1_wdata), .ram_w8_l2048_id7_3_1_wenable(ram_w8_l2048_id7_3_1_wenable) );
  ram_w8_l2048_id8_0 inst_ram_w8_l2048_id8_0 ( .CLK(CLK), .ram_w8_l2048_id8_0_0_addr(ram_w8_l2048_id8_0_0_addr), .ram_w8_l2048_id8_0_0_rdata(ram_w8_l2048_id8_0_0_rdata), .ram_w8_l2048_id8_0_0_wdata(8'h00), .ram_w8_l2048_id8_0_0_wenable(1'h0), .ram_w8_l2048_id8_0_1_addr(ram_w8_l2048_id8_0_1_addr), .ram_w8_l2048_id8_0_1_rdata(ram_w8_l2048_id8_0_1_rdata), .ram_w8_l2048_id8_0_1_wdata(ram_w8_l2048_id8_0_1_wdata), .ram_w8_l2048_id8_0_1_wenable(ram_w8_l2048_id8_0_1_wenable) );
  ram_w8_l2048_id8_1 inst_ram_w8_l2048_id8_1 ( .CLK(CLK), .ram_w8_l2048_id8_1_0_addr(ram_w8_l2048_id8_1_0_addr), .ram_w8_l2048_id8_1_0_rdata(ram_w8_l2048_id8_1_0_rdata), .ram_w8_l2048_id8_1_0_wdata(8'h00), .ram_w8_l2048_id8_1_0_wenable(1'h0), .ram_w8_l2048_id8_1_1_addr(ram_w8_l2048_id8_1_1_addr), .ram_w8_l2048_id8_1_1_rdata(ram_w8_l2048_id8_1_1_rdata), .ram_w8_l2048_id8_1_1_wdata(ram_w8_l2048_id8_1_1_wdata), .ram_w8_l2048_id8_1_1_wenable(ram_w8_l2048_id8_1_1_wenable) );
  ram_w8_l2048_id8_2 inst_ram_w8_l2048_id8_2 ( .CLK(CLK), .ram_w8_l2048_id8_2_0_addr(ram_w8_l2048_id8_2_0_addr), .ram_w8_l2048_id8_2_0_rdata(ram_w8_l2048_id8_2_0_rdata), .ram_w8_l2048_id8_2_0_wdata(8'h00), .ram_w8_l2048_id8_2_0_wenable(1'h0), .ram_w8_l2048_id8_2_1_addr(ram_w8_l2048_id8_2_1_addr), .ram_w8_l2048_id8_2_1_rdata(ram_w8_l2048_id8_2_1_rdata), .ram_w8_l2048_id8_2_1_wdata(ram_w8_l2048_id8_2_1_wdata), .ram_w8_l2048_id8_2_1_wenable(ram_w8_l2048_id8_2_1_wenable) );
  ram_w8_l2048_id8_3 inst_ram_w8_l2048_id8_3 ( .CLK(CLK), .ram_w8_l2048_id8_3_0_addr(ram_w8_l2048_id8_3_0_addr), .ram_w8_l2048_id8_3_0_rdata(ram_w8_l2048_id8_3_0_rdata), .ram_w8_l2048_id8_3_0_wdata(8'h00), .ram_w8_l2048_id8_3_0_wenable(1'h0), .ram_w8_l2048_id8_3_1_addr(ram_w8_l2048_id8_3_1_addr), .ram_w8_l2048_id8_3_1_rdata(ram_w8_l2048_id8_3_1_rdata), .ram_w8_l2048_id8_3_1_wdata(ram_w8_l2048_id8_3_1_wdata), .ram_w8_l2048_id8_3_1_wenable(ram_w8_l2048_id8_3_1_wenable) );
  ram_w8_l2048_id9_0 inst_ram_w8_l2048_id9_0 ( .CLK(CLK), .ram_w8_l2048_id9_0_0_addr(ram_w8_l2048_id9_0_0_addr), .ram_w8_l2048_id9_0_0_rdata(ram_w8_l2048_id9_0_0_rdata), .ram_w8_l2048_id9_0_0_wdata(8'h00), .ram_w8_l2048_id9_0_0_wenable(1'h0), .ram_w8_l2048_id9_0_1_addr(ram_w8_l2048_id9_0_1_addr), .ram_w8_l2048_id9_0_1_rdata(ram_w8_l2048_id9_0_1_rdata), .ram_w8_l2048_id9_0_1_wdata(ram_w8_l2048_id9_0_1_wdata), .ram_w8_l2048_id9_0_1_wenable(ram_w8_l2048_id9_0_1_wenable) );
  ram_w8_l2048_id9_1 inst_ram_w8_l2048_id9_1 ( .CLK(CLK), .ram_w8_l2048_id9_1_0_addr(ram_w8_l2048_id9_1_0_addr), .ram_w8_l2048_id9_1_0_rdata(ram_w8_l2048_id9_1_0_rdata), .ram_w8_l2048_id9_1_0_wdata(8'h00), .ram_w8_l2048_id9_1_0_wenable(1'h0), .ram_w8_l2048_id9_1_1_addr(ram_w8_l2048_id9_1_1_addr), .ram_w8_l2048_id9_1_1_rdata(ram_w8_l2048_id9_1_1_rdata), .ram_w8_l2048_id9_1_1_wdata(ram_w8_l2048_id9_1_1_wdata), .ram_w8_l2048_id9_1_1_wenable(ram_w8_l2048_id9_1_1_wenable) );
  ram_w8_l2048_id9_2 inst_ram_w8_l2048_id9_2 ( .CLK(CLK), .ram_w8_l2048_id9_2_0_addr(ram_w8_l2048_id9_2_0_addr), .ram_w8_l2048_id9_2_0_rdata(ram_w8_l2048_id9_2_0_rdata), .ram_w8_l2048_id9_2_0_wdata(8'h00), .ram_w8_l2048_id9_2_0_wenable(1'h0), .ram_w8_l2048_id9_2_1_addr(ram_w8_l2048_id9_2_1_addr), .ram_w8_l2048_id9_2_1_rdata(ram_w8_l2048_id9_2_1_rdata), .ram_w8_l2048_id9_2_1_wdata(ram_w8_l2048_id9_2_1_wdata), .ram_w8_l2048_id9_2_1_wenable(ram_w8_l2048_id9_2_1_wenable) );
  ram_w8_l2048_id9_3 inst_ram_w8_l2048_id9_3 ( .CLK(CLK), .ram_w8_l2048_id9_3_0_addr(ram_w8_l2048_id9_3_0_addr), .ram_w8_l2048_id9_3_0_rdata(ram_w8_l2048_id9_3_0_rdata), .ram_w8_l2048_id9_3_0_wdata(8'h00), .ram_w8_l2048_id9_3_0_wenable(1'h0), .ram_w8_l2048_id9_3_1_addr(ram_w8_l2048_id9_3_1_addr), .ram_w8_l2048_id9_3_1_rdata(ram_w8_l2048_id9_3_1_rdata), .ram_w8_l2048_id9_3_1_wdata(ram_w8_l2048_id9_3_1_wdata), .ram_w8_l2048_id9_3_1_wenable(ram_w8_l2048_id9_3_1_wenable) );
  ram_w8_l4096_id0_0 inst_ram_w8_l4096_id0_0 ( .CLK(CLK), .ram_w8_l4096_id0_0_0_addr(ram_w8_l4096_id0_0_0_addr), .ram_w8_l4096_id0_0_0_rdata(ram_w8_l4096_id0_0_0_rdata), .ram_w8_l4096_id0_0_0_wdata(8'h00), .ram_w8_l4096_id0_0_0_wenable(1'h0), .ram_w8_l4096_id0_0_1_addr(ram_w8_l4096_id0_0_1_addr), .ram_w8_l4096_id0_0_1_rdata(ram_w8_l4096_id0_0_1_rdata), .ram_w8_l4096_id0_0_1_wdata(ram_w8_l4096_id0_0_1_wdata), .ram_w8_l4096_id0_0_1_wenable(ram_w8_l4096_id0_0_1_wenable) );
  ram_w8_l4096_id0_1 inst_ram_w8_l4096_id0_1 ( .CLK(CLK), .ram_w8_l4096_id0_1_0_addr(ram_w8_l4096_id0_1_0_addr), .ram_w8_l4096_id0_1_0_rdata(ram_w8_l4096_id0_1_0_rdata), .ram_w8_l4096_id0_1_0_wdata(8'h00), .ram_w8_l4096_id0_1_0_wenable(1'h0), .ram_w8_l4096_id0_1_1_addr(ram_w8_l4096_id0_1_1_addr), .ram_w8_l4096_id0_1_1_rdata(ram_w8_l4096_id0_1_1_rdata), .ram_w8_l4096_id0_1_1_wdata(ram_w8_l4096_id0_1_1_wdata), .ram_w8_l4096_id0_1_1_wenable(ram_w8_l4096_id0_1_1_wenable) );
  ram_w8_l4096_id0_2 inst_ram_w8_l4096_id0_2 ( .CLK(CLK), .ram_w8_l4096_id0_2_0_addr(ram_w8_l4096_id0_2_0_addr), .ram_w8_l4096_id0_2_0_rdata(ram_w8_l4096_id0_2_0_rdata), .ram_w8_l4096_id0_2_0_wdata(8'h00), .ram_w8_l4096_id0_2_0_wenable(1'h0), .ram_w8_l4096_id0_2_1_addr(ram_w8_l4096_id0_2_1_addr), .ram_w8_l4096_id0_2_1_rdata(ram_w8_l4096_id0_2_1_rdata), .ram_w8_l4096_id0_2_1_wdata(ram_w8_l4096_id0_2_1_wdata), .ram_w8_l4096_id0_2_1_wenable(ram_w8_l4096_id0_2_1_wenable) );
  ram_w8_l4096_id0_3 inst_ram_w8_l4096_id0_3 ( .CLK(CLK), .ram_w8_l4096_id0_3_0_addr(ram_w8_l4096_id0_3_0_addr), .ram_w8_l4096_id0_3_0_rdata(ram_w8_l4096_id0_3_0_rdata), .ram_w8_l4096_id0_3_0_wdata(8'h00), .ram_w8_l4096_id0_3_0_wenable(1'h0), .ram_w8_l4096_id0_3_1_addr(ram_w8_l4096_id0_3_1_addr), .ram_w8_l4096_id0_3_1_rdata(ram_w8_l4096_id0_3_1_rdata), .ram_w8_l4096_id0_3_1_wdata(ram_w8_l4096_id0_3_1_wdata), .ram_w8_l4096_id0_3_1_wenable(ram_w8_l4096_id0_3_1_wenable) );
endmodule
