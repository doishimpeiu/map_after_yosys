

module nngenmod
(
  input CLK,
  input RESETN,
  output reg [32-1:0] maxi_awaddr,
  output reg [8-1:0] maxi_awlen,
  output [3-1:0] maxi_awsize,
  output [2-1:0] maxi_awburst,
  output [1-1:0] maxi_awlock,
  output [4-1:0] maxi_awcache,
  output [3-1:0] maxi_awprot,
  output [4-1:0] maxi_awqos,
  output [2-1:0] maxi_awuser,
  output reg maxi_awvalid,
  input maxi_awready,
  output reg [32-1:0] maxi_wdata,
  output reg [4-1:0] maxi_wstrb,
  output reg maxi_wlast,
  output reg maxi_wvalid,
  input maxi_wready,
  input [2-1:0] maxi_bresp,
  input maxi_bvalid,
  output maxi_bready,
  output reg [32-1:0] maxi_araddr,
  output reg [8-1:0] maxi_arlen,
  output [3-1:0] maxi_arsize,
  output [2-1:0] maxi_arburst,
  output [1-1:0] maxi_arlock,
  output [4-1:0] maxi_arcache,
  output [3-1:0] maxi_arprot,
  output [4-1:0] maxi_arqos,
  output [2-1:0] maxi_aruser,
  output reg maxi_arvalid,
  input maxi_arready,
  input [32-1:0] maxi_rdata,
  input [2-1:0] maxi_rresp,
  input maxi_rlast,
  input maxi_rvalid,
  output maxi_rready,
  input [6-1:0] saxi_awaddr,
  input [4-1:0] saxi_awcache,
  input [3-1:0] saxi_awprot,
  input saxi_awvalid,
  output saxi_awready,
  input [32-1:0] saxi_wdata,
  input [4-1:0] saxi_wstrb,
  input saxi_wvalid,
  output saxi_wready,
  output [2-1:0] saxi_bresp,
  output reg saxi_bvalid,
  input saxi_bready,
  input [6-1:0] saxi_araddr,
  input [4-1:0] saxi_arcache,
  input [3-1:0] saxi_arprot,
  input saxi_arvalid,
  output saxi_arready,
  output reg [32-1:0] saxi_rdata,
  output [2-1:0] saxi_rresp,
  output reg saxi_rvalid,
  input saxi_rready
);

  wire RESETN_inv;
  assign RESETN_inv = !RESETN;
  wire RESETN_inv_buf;
  reg _RESETN_inv_1;
  reg _RESETN_inv_2;
  assign RESETN_inv_buf = _RESETN_inv_2;
  assign maxi_awsize = 2;
  assign maxi_awburst = 1;
  assign maxi_awlock = 0;
  assign maxi_awcache = 3;
  assign maxi_awprot = 0;
  assign maxi_awqos = 0;
  assign maxi_awuser = 0;
  assign maxi_bready = 1;
  assign maxi_arsize = 2;
  assign maxi_arburst = 1;
  assign maxi_arlock = 0;
  assign maxi_arcache = 3;
  assign maxi_arprot = 0;
  assign maxi_arqos = 0;
  assign maxi_aruser = 0;
  reg _maxi_read_start;
  reg [8-1:0] _maxi_read_op_sel;
  reg [32-1:0] _maxi_read_local_addr;
  reg [32-1:0] _maxi_read_global_addr;
  reg [33-1:0] _maxi_read_size;
  reg [32-1:0] _maxi_read_local_stride;
  reg _maxi_read_idle;
  reg _maxi_write_start;
  reg [8-1:0] _maxi_write_op_sel;
  reg [32-1:0] _maxi_write_local_addr;
  reg [32-1:0] _maxi_write_global_addr;
  reg [33-1:0] _maxi_write_size;
  reg [32-1:0] _maxi_write_local_stride;
  reg _maxi_write_idle;
  reg [32-1:0] _maxi_global_base_addr;
  wire _maxi_write_data_done;
  assign saxi_bresp = 0;
  assign saxi_rresp = 0;
  reg signed [32-1:0] _saxi_register_0;
  reg signed [32-1:0] _saxi_register_1;
  reg signed [32-1:0] _saxi_register_2;
  reg signed [32-1:0] _saxi_register_3;
  reg signed [32-1:0] _saxi_register_4;
  reg signed [32-1:0] _saxi_register_5;
  reg signed [32-1:0] _saxi_register_6;
  reg signed [32-1:0] _saxi_register_7;
  reg signed [32-1:0] _saxi_register_8;
  reg signed [32-1:0] _saxi_register_9;
  reg signed [32-1:0] _saxi_register_10;
  reg signed [32-1:0] _saxi_register_11;
  reg signed [32-1:0] _saxi_register_12;
  reg signed [32-1:0] _saxi_register_13;
  reg _saxi_flag_0;
  reg _saxi_flag_1;
  reg _saxi_flag_2;
  reg _saxi_flag_3;
  reg _saxi_flag_4;
  reg _saxi_flag_5;
  reg _saxi_flag_6;
  reg _saxi_flag_7;
  reg _saxi_flag_8;
  reg _saxi_flag_9;
  reg _saxi_flag_10;
  reg _saxi_flag_11;
  reg _saxi_flag_12;
  reg _saxi_flag_13;
  reg signed [32-1:0] _saxi_resetval_0;
  reg signed [32-1:0] _saxi_resetval_1;
  reg signed [32-1:0] _saxi_resetval_2;
  reg signed [32-1:0] _saxi_resetval_3;
  reg signed [32-1:0] _saxi_resetval_4;
  reg signed [32-1:0] _saxi_resetval_5;
  reg signed [32-1:0] _saxi_resetval_6;
  reg signed [32-1:0] _saxi_resetval_7;
  reg signed [32-1:0] _saxi_resetval_8;
  reg signed [32-1:0] _saxi_resetval_9;
  reg signed [32-1:0] _saxi_resetval_10;
  reg signed [32-1:0] _saxi_resetval_11;
  reg signed [32-1:0] _saxi_resetval_12;
  reg signed [32-1:0] _saxi_resetval_13;
  localparam _saxi_maskwidth = 4;
  localparam _saxi_mask = { _saxi_maskwidth{ 1'd1 } };
  localparam _saxi_shift = 2;
  reg [32-1:0] _saxi_register_fsm;
  localparam _saxi_register_fsm_init = 0;
  reg [6-1:0] _tmp_0;
  reg _tmp_1;
  reg _tmp_2;
  reg _tmp_3;
  reg _tmp_4;
  assign saxi_awready = (_saxi_register_fsm == 0) && !_tmp_1 && !_tmp_2 && !saxi_bvalid && _tmp_3;
  assign saxi_arready = (_saxi_register_fsm == 0) && !_tmp_2 && !_tmp_1 && _tmp_4;
  reg [_saxi_maskwidth-1:0] _tmp_5;
  wire signed [32-1:0] _tmp_6;
  assign _tmp_6 = (_tmp_5 == 0)? _saxi_register_0 : 
                  (_tmp_5 == 1)? _saxi_register_1 : 
                  (_tmp_5 == 2)? _saxi_register_2 : 
                  (_tmp_5 == 3)? _saxi_register_3 : 
                  (_tmp_5 == 4)? _saxi_register_4 : 
                  (_tmp_5 == 5)? _saxi_register_5 : 
                  (_tmp_5 == 6)? _saxi_register_6 : 
                  (_tmp_5 == 7)? _saxi_register_7 : 
                  (_tmp_5 == 8)? _saxi_register_8 : 
                  (_tmp_5 == 9)? _saxi_register_9 : 
                  (_tmp_5 == 10)? _saxi_register_10 : 
                  (_tmp_5 == 11)? _saxi_register_11 : 
                  (_tmp_5 == 12)? _saxi_register_12 : 
                  (_tmp_5 == 13)? _saxi_register_13 : 'hx;
  wire _tmp_7;
  assign _tmp_7 = (_tmp_5 == 0)? _saxi_flag_0 : 
                  (_tmp_5 == 1)? _saxi_flag_1 : 
                  (_tmp_5 == 2)? _saxi_flag_2 : 
                  (_tmp_5 == 3)? _saxi_flag_3 : 
                  (_tmp_5 == 4)? _saxi_flag_4 : 
                  (_tmp_5 == 5)? _saxi_flag_5 : 
                  (_tmp_5 == 6)? _saxi_flag_6 : 
                  (_tmp_5 == 7)? _saxi_flag_7 : 
                  (_tmp_5 == 8)? _saxi_flag_8 : 
                  (_tmp_5 == 9)? _saxi_flag_9 : 
                  (_tmp_5 == 10)? _saxi_flag_10 : 
                  (_tmp_5 == 11)? _saxi_flag_11 : 
                  (_tmp_5 == 12)? _saxi_flag_12 : 
                  (_tmp_5 == 13)? _saxi_flag_13 : 'hx;
  wire signed [32-1:0] _tmp_8;
  assign _tmp_8 = (_tmp_5 == 0)? _saxi_resetval_0 : 
                  (_tmp_5 == 1)? _saxi_resetval_1 : 
                  (_tmp_5 == 2)? _saxi_resetval_2 : 
                  (_tmp_5 == 3)? _saxi_resetval_3 : 
                  (_tmp_5 == 4)? _saxi_resetval_4 : 
                  (_tmp_5 == 5)? _saxi_resetval_5 : 
                  (_tmp_5 == 6)? _saxi_resetval_6 : 
                  (_tmp_5 == 7)? _saxi_resetval_7 : 
                  (_tmp_5 == 8)? _saxi_resetval_8 : 
                  (_tmp_5 == 9)? _saxi_resetval_9 : 
                  (_tmp_5 == 10)? _saxi_resetval_10 : 
                  (_tmp_5 == 11)? _saxi_resetval_11 : 
                  (_tmp_5 == 12)? _saxi_resetval_12 : 
                  (_tmp_5 == 13)? _saxi_resetval_13 : 'hx;
  reg _saxi_cond_0_1;
  assign saxi_wready = _saxi_register_fsm == 2;
  wire maxi_idle;
  assign maxi_idle = _maxi_write_idle & _maxi_read_idle;
  wire sw_rst_logic;
  assign sw_rst_logic = maxi_idle & _saxi_register_6;
  wire rst_logic;
  assign rst_logic = RESETN_inv_buf | sw_rst_logic;
  reg RST;
  reg _rst_logic_1;
  reg _rst_logic_2;
  reg [10-1:0] ram_w4_l8192_id0_0_0_addr;
  wire [4-1:0] ram_w4_l8192_id0_0_0_rdata;
  reg [4-1:0] ram_w4_l8192_id0_0_0_wdata;
  reg ram_w4_l8192_id0_0_0_wenable;
  reg [10-1:0] ram_w4_l8192_id0_0_1_addr;
  wire [4-1:0] ram_w4_l8192_id0_0_1_rdata;
  reg [4-1:0] ram_w4_l8192_id0_0_1_wdata;
  reg ram_w4_l8192_id0_0_1_wenable;

  ram_w4_l8192_id0_0
  inst_ram_w4_l8192_id0_0
  (
    .CLK(CLK),
    .ram_w4_l8192_id0_0_0_addr(ram_w4_l8192_id0_0_0_addr),
    .ram_w4_l8192_id0_0_0_rdata(ram_w4_l8192_id0_0_0_rdata),
    .ram_w4_l8192_id0_0_0_wdata(ram_w4_l8192_id0_0_0_wdata),
    .ram_w4_l8192_id0_0_0_wenable(ram_w4_l8192_id0_0_0_wenable),
    .ram_w4_l8192_id0_0_1_addr(ram_w4_l8192_id0_0_1_addr),
    .ram_w4_l8192_id0_0_1_rdata(ram_w4_l8192_id0_0_1_rdata),
    .ram_w4_l8192_id0_0_1_wdata(ram_w4_l8192_id0_0_1_wdata),
    .ram_w4_l8192_id0_0_1_wenable(ram_w4_l8192_id0_0_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id0_1_0_addr;
  wire [4-1:0] ram_w4_l8192_id0_1_0_rdata;
  reg [4-1:0] ram_w4_l8192_id0_1_0_wdata;
  reg ram_w4_l8192_id0_1_0_wenable;
  reg [10-1:0] ram_w4_l8192_id0_1_1_addr;
  wire [4-1:0] ram_w4_l8192_id0_1_1_rdata;
  reg [4-1:0] ram_w4_l8192_id0_1_1_wdata;
  reg ram_w4_l8192_id0_1_1_wenable;

  ram_w4_l8192_id0_1
  inst_ram_w4_l8192_id0_1
  (
    .CLK(CLK),
    .ram_w4_l8192_id0_1_0_addr(ram_w4_l8192_id0_1_0_addr),
    .ram_w4_l8192_id0_1_0_rdata(ram_w4_l8192_id0_1_0_rdata),
    .ram_w4_l8192_id0_1_0_wdata(ram_w4_l8192_id0_1_0_wdata),
    .ram_w4_l8192_id0_1_0_wenable(ram_w4_l8192_id0_1_0_wenable),
    .ram_w4_l8192_id0_1_1_addr(ram_w4_l8192_id0_1_1_addr),
    .ram_w4_l8192_id0_1_1_rdata(ram_w4_l8192_id0_1_1_rdata),
    .ram_w4_l8192_id0_1_1_wdata(ram_w4_l8192_id0_1_1_wdata),
    .ram_w4_l8192_id0_1_1_wenable(ram_w4_l8192_id0_1_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id0_2_0_addr;
  wire [4-1:0] ram_w4_l8192_id0_2_0_rdata;
  reg [4-1:0] ram_w4_l8192_id0_2_0_wdata;
  reg ram_w4_l8192_id0_2_0_wenable;
  reg [10-1:0] ram_w4_l8192_id0_2_1_addr;
  wire [4-1:0] ram_w4_l8192_id0_2_1_rdata;
  reg [4-1:0] ram_w4_l8192_id0_2_1_wdata;
  reg ram_w4_l8192_id0_2_1_wenable;

  ram_w4_l8192_id0_2
  inst_ram_w4_l8192_id0_2
  (
    .CLK(CLK),
    .ram_w4_l8192_id0_2_0_addr(ram_w4_l8192_id0_2_0_addr),
    .ram_w4_l8192_id0_2_0_rdata(ram_w4_l8192_id0_2_0_rdata),
    .ram_w4_l8192_id0_2_0_wdata(ram_w4_l8192_id0_2_0_wdata),
    .ram_w4_l8192_id0_2_0_wenable(ram_w4_l8192_id0_2_0_wenable),
    .ram_w4_l8192_id0_2_1_addr(ram_w4_l8192_id0_2_1_addr),
    .ram_w4_l8192_id0_2_1_rdata(ram_w4_l8192_id0_2_1_rdata),
    .ram_w4_l8192_id0_2_1_wdata(ram_w4_l8192_id0_2_1_wdata),
    .ram_w4_l8192_id0_2_1_wenable(ram_w4_l8192_id0_2_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id0_3_0_addr;
  wire [4-1:0] ram_w4_l8192_id0_3_0_rdata;
  reg [4-1:0] ram_w4_l8192_id0_3_0_wdata;
  reg ram_w4_l8192_id0_3_0_wenable;
  reg [10-1:0] ram_w4_l8192_id0_3_1_addr;
  wire [4-1:0] ram_w4_l8192_id0_3_1_rdata;
  reg [4-1:0] ram_w4_l8192_id0_3_1_wdata;
  reg ram_w4_l8192_id0_3_1_wenable;

  ram_w4_l8192_id0_3
  inst_ram_w4_l8192_id0_3
  (
    .CLK(CLK),
    .ram_w4_l8192_id0_3_0_addr(ram_w4_l8192_id0_3_0_addr),
    .ram_w4_l8192_id0_3_0_rdata(ram_w4_l8192_id0_3_0_rdata),
    .ram_w4_l8192_id0_3_0_wdata(ram_w4_l8192_id0_3_0_wdata),
    .ram_w4_l8192_id0_3_0_wenable(ram_w4_l8192_id0_3_0_wenable),
    .ram_w4_l8192_id0_3_1_addr(ram_w4_l8192_id0_3_1_addr),
    .ram_w4_l8192_id0_3_1_rdata(ram_w4_l8192_id0_3_1_rdata),
    .ram_w4_l8192_id0_3_1_wdata(ram_w4_l8192_id0_3_1_wdata),
    .ram_w4_l8192_id0_3_1_wenable(ram_w4_l8192_id0_3_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id0_4_0_addr;
  wire [4-1:0] ram_w4_l8192_id0_4_0_rdata;
  reg [4-1:0] ram_w4_l8192_id0_4_0_wdata;
  reg ram_w4_l8192_id0_4_0_wenable;
  reg [10-1:0] ram_w4_l8192_id0_4_1_addr;
  wire [4-1:0] ram_w4_l8192_id0_4_1_rdata;
  reg [4-1:0] ram_w4_l8192_id0_4_1_wdata;
  reg ram_w4_l8192_id0_4_1_wenable;

  ram_w4_l8192_id0_4
  inst_ram_w4_l8192_id0_4
  (
    .CLK(CLK),
    .ram_w4_l8192_id0_4_0_addr(ram_w4_l8192_id0_4_0_addr),
    .ram_w4_l8192_id0_4_0_rdata(ram_w4_l8192_id0_4_0_rdata),
    .ram_w4_l8192_id0_4_0_wdata(ram_w4_l8192_id0_4_0_wdata),
    .ram_w4_l8192_id0_4_0_wenable(ram_w4_l8192_id0_4_0_wenable),
    .ram_w4_l8192_id0_4_1_addr(ram_w4_l8192_id0_4_1_addr),
    .ram_w4_l8192_id0_4_1_rdata(ram_w4_l8192_id0_4_1_rdata),
    .ram_w4_l8192_id0_4_1_wdata(ram_w4_l8192_id0_4_1_wdata),
    .ram_w4_l8192_id0_4_1_wenable(ram_w4_l8192_id0_4_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id0_5_0_addr;
  wire [4-1:0] ram_w4_l8192_id0_5_0_rdata;
  reg [4-1:0] ram_w4_l8192_id0_5_0_wdata;
  reg ram_w4_l8192_id0_5_0_wenable;
  reg [10-1:0] ram_w4_l8192_id0_5_1_addr;
  wire [4-1:0] ram_w4_l8192_id0_5_1_rdata;
  reg [4-1:0] ram_w4_l8192_id0_5_1_wdata;
  reg ram_w4_l8192_id0_5_1_wenable;

  ram_w4_l8192_id0_5
  inst_ram_w4_l8192_id0_5
  (
    .CLK(CLK),
    .ram_w4_l8192_id0_5_0_addr(ram_w4_l8192_id0_5_0_addr),
    .ram_w4_l8192_id0_5_0_rdata(ram_w4_l8192_id0_5_0_rdata),
    .ram_w4_l8192_id0_5_0_wdata(ram_w4_l8192_id0_5_0_wdata),
    .ram_w4_l8192_id0_5_0_wenable(ram_w4_l8192_id0_5_0_wenable),
    .ram_w4_l8192_id0_5_1_addr(ram_w4_l8192_id0_5_1_addr),
    .ram_w4_l8192_id0_5_1_rdata(ram_w4_l8192_id0_5_1_rdata),
    .ram_w4_l8192_id0_5_1_wdata(ram_w4_l8192_id0_5_1_wdata),
    .ram_w4_l8192_id0_5_1_wenable(ram_w4_l8192_id0_5_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id0_6_0_addr;
  wire [4-1:0] ram_w4_l8192_id0_6_0_rdata;
  reg [4-1:0] ram_w4_l8192_id0_6_0_wdata;
  reg ram_w4_l8192_id0_6_0_wenable;
  reg [10-1:0] ram_w4_l8192_id0_6_1_addr;
  wire [4-1:0] ram_w4_l8192_id0_6_1_rdata;
  reg [4-1:0] ram_w4_l8192_id0_6_1_wdata;
  reg ram_w4_l8192_id0_6_1_wenable;

  ram_w4_l8192_id0_6
  inst_ram_w4_l8192_id0_6
  (
    .CLK(CLK),
    .ram_w4_l8192_id0_6_0_addr(ram_w4_l8192_id0_6_0_addr),
    .ram_w4_l8192_id0_6_0_rdata(ram_w4_l8192_id0_6_0_rdata),
    .ram_w4_l8192_id0_6_0_wdata(ram_w4_l8192_id0_6_0_wdata),
    .ram_w4_l8192_id0_6_0_wenable(ram_w4_l8192_id0_6_0_wenable),
    .ram_w4_l8192_id0_6_1_addr(ram_w4_l8192_id0_6_1_addr),
    .ram_w4_l8192_id0_6_1_rdata(ram_w4_l8192_id0_6_1_rdata),
    .ram_w4_l8192_id0_6_1_wdata(ram_w4_l8192_id0_6_1_wdata),
    .ram_w4_l8192_id0_6_1_wenable(ram_w4_l8192_id0_6_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id0_7_0_addr;
  wire [4-1:0] ram_w4_l8192_id0_7_0_rdata;
  reg [4-1:0] ram_w4_l8192_id0_7_0_wdata;
  reg ram_w4_l8192_id0_7_0_wenable;
  reg [10-1:0] ram_w4_l8192_id0_7_1_addr;
  wire [4-1:0] ram_w4_l8192_id0_7_1_rdata;
  reg [4-1:0] ram_w4_l8192_id0_7_1_wdata;
  reg ram_w4_l8192_id0_7_1_wenable;

  ram_w4_l8192_id0_7
  inst_ram_w4_l8192_id0_7
  (
    .CLK(CLK),
    .ram_w4_l8192_id0_7_0_addr(ram_w4_l8192_id0_7_0_addr),
    .ram_w4_l8192_id0_7_0_rdata(ram_w4_l8192_id0_7_0_rdata),
    .ram_w4_l8192_id0_7_0_wdata(ram_w4_l8192_id0_7_0_wdata),
    .ram_w4_l8192_id0_7_0_wenable(ram_w4_l8192_id0_7_0_wenable),
    .ram_w4_l8192_id0_7_1_addr(ram_w4_l8192_id0_7_1_addr),
    .ram_w4_l8192_id0_7_1_rdata(ram_w4_l8192_id0_7_1_rdata),
    .ram_w4_l8192_id0_7_1_wdata(ram_w4_l8192_id0_7_1_wdata),
    .ram_w4_l8192_id0_7_1_wenable(ram_w4_l8192_id0_7_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id1_0_0_addr;
  wire [4-1:0] ram_w4_l8192_id1_0_0_rdata;
  reg [4-1:0] ram_w4_l8192_id1_0_0_wdata;
  reg ram_w4_l8192_id1_0_0_wenable;
  reg [10-1:0] ram_w4_l8192_id1_0_1_addr;
  wire [4-1:0] ram_w4_l8192_id1_0_1_rdata;
  reg [4-1:0] ram_w4_l8192_id1_0_1_wdata;
  reg ram_w4_l8192_id1_0_1_wenable;

  ram_w4_l8192_id1_0
  inst_ram_w4_l8192_id1_0
  (
    .CLK(CLK),
    .ram_w4_l8192_id1_0_0_addr(ram_w4_l8192_id1_0_0_addr),
    .ram_w4_l8192_id1_0_0_rdata(ram_w4_l8192_id1_0_0_rdata),
    .ram_w4_l8192_id1_0_0_wdata(ram_w4_l8192_id1_0_0_wdata),
    .ram_w4_l8192_id1_0_0_wenable(ram_w4_l8192_id1_0_0_wenable),
    .ram_w4_l8192_id1_0_1_addr(ram_w4_l8192_id1_0_1_addr),
    .ram_w4_l8192_id1_0_1_rdata(ram_w4_l8192_id1_0_1_rdata),
    .ram_w4_l8192_id1_0_1_wdata(ram_w4_l8192_id1_0_1_wdata),
    .ram_w4_l8192_id1_0_1_wenable(ram_w4_l8192_id1_0_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id1_1_0_addr;
  wire [4-1:0] ram_w4_l8192_id1_1_0_rdata;
  reg [4-1:0] ram_w4_l8192_id1_1_0_wdata;
  reg ram_w4_l8192_id1_1_0_wenable;
  reg [10-1:0] ram_w4_l8192_id1_1_1_addr;
  wire [4-1:0] ram_w4_l8192_id1_1_1_rdata;
  reg [4-1:0] ram_w4_l8192_id1_1_1_wdata;
  reg ram_w4_l8192_id1_1_1_wenable;

  ram_w4_l8192_id1_1
  inst_ram_w4_l8192_id1_1
  (
    .CLK(CLK),
    .ram_w4_l8192_id1_1_0_addr(ram_w4_l8192_id1_1_0_addr),
    .ram_w4_l8192_id1_1_0_rdata(ram_w4_l8192_id1_1_0_rdata),
    .ram_w4_l8192_id1_1_0_wdata(ram_w4_l8192_id1_1_0_wdata),
    .ram_w4_l8192_id1_1_0_wenable(ram_w4_l8192_id1_1_0_wenable),
    .ram_w4_l8192_id1_1_1_addr(ram_w4_l8192_id1_1_1_addr),
    .ram_w4_l8192_id1_1_1_rdata(ram_w4_l8192_id1_1_1_rdata),
    .ram_w4_l8192_id1_1_1_wdata(ram_w4_l8192_id1_1_1_wdata),
    .ram_w4_l8192_id1_1_1_wenable(ram_w4_l8192_id1_1_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id1_2_0_addr;
  wire [4-1:0] ram_w4_l8192_id1_2_0_rdata;
  reg [4-1:0] ram_w4_l8192_id1_2_0_wdata;
  reg ram_w4_l8192_id1_2_0_wenable;
  reg [10-1:0] ram_w4_l8192_id1_2_1_addr;
  wire [4-1:0] ram_w4_l8192_id1_2_1_rdata;
  reg [4-1:0] ram_w4_l8192_id1_2_1_wdata;
  reg ram_w4_l8192_id1_2_1_wenable;

  ram_w4_l8192_id1_2
  inst_ram_w4_l8192_id1_2
  (
    .CLK(CLK),
    .ram_w4_l8192_id1_2_0_addr(ram_w4_l8192_id1_2_0_addr),
    .ram_w4_l8192_id1_2_0_rdata(ram_w4_l8192_id1_2_0_rdata),
    .ram_w4_l8192_id1_2_0_wdata(ram_w4_l8192_id1_2_0_wdata),
    .ram_w4_l8192_id1_2_0_wenable(ram_w4_l8192_id1_2_0_wenable),
    .ram_w4_l8192_id1_2_1_addr(ram_w4_l8192_id1_2_1_addr),
    .ram_w4_l8192_id1_2_1_rdata(ram_w4_l8192_id1_2_1_rdata),
    .ram_w4_l8192_id1_2_1_wdata(ram_w4_l8192_id1_2_1_wdata),
    .ram_w4_l8192_id1_2_1_wenable(ram_w4_l8192_id1_2_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id1_3_0_addr;
  wire [4-1:0] ram_w4_l8192_id1_3_0_rdata;
  reg [4-1:0] ram_w4_l8192_id1_3_0_wdata;
  reg ram_w4_l8192_id1_3_0_wenable;
  reg [10-1:0] ram_w4_l8192_id1_3_1_addr;
  wire [4-1:0] ram_w4_l8192_id1_3_1_rdata;
  reg [4-1:0] ram_w4_l8192_id1_3_1_wdata;
  reg ram_w4_l8192_id1_3_1_wenable;

  ram_w4_l8192_id1_3
  inst_ram_w4_l8192_id1_3
  (
    .CLK(CLK),
    .ram_w4_l8192_id1_3_0_addr(ram_w4_l8192_id1_3_0_addr),
    .ram_w4_l8192_id1_3_0_rdata(ram_w4_l8192_id1_3_0_rdata),
    .ram_w4_l8192_id1_3_0_wdata(ram_w4_l8192_id1_3_0_wdata),
    .ram_w4_l8192_id1_3_0_wenable(ram_w4_l8192_id1_3_0_wenable),
    .ram_w4_l8192_id1_3_1_addr(ram_w4_l8192_id1_3_1_addr),
    .ram_w4_l8192_id1_3_1_rdata(ram_w4_l8192_id1_3_1_rdata),
    .ram_w4_l8192_id1_3_1_wdata(ram_w4_l8192_id1_3_1_wdata),
    .ram_w4_l8192_id1_3_1_wenable(ram_w4_l8192_id1_3_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id1_4_0_addr;
  wire [4-1:0] ram_w4_l8192_id1_4_0_rdata;
  reg [4-1:0] ram_w4_l8192_id1_4_0_wdata;
  reg ram_w4_l8192_id1_4_0_wenable;
  reg [10-1:0] ram_w4_l8192_id1_4_1_addr;
  wire [4-1:0] ram_w4_l8192_id1_4_1_rdata;
  reg [4-1:0] ram_w4_l8192_id1_4_1_wdata;
  reg ram_w4_l8192_id1_4_1_wenable;

  ram_w4_l8192_id1_4
  inst_ram_w4_l8192_id1_4
  (
    .CLK(CLK),
    .ram_w4_l8192_id1_4_0_addr(ram_w4_l8192_id1_4_0_addr),
    .ram_w4_l8192_id1_4_0_rdata(ram_w4_l8192_id1_4_0_rdata),
    .ram_w4_l8192_id1_4_0_wdata(ram_w4_l8192_id1_4_0_wdata),
    .ram_w4_l8192_id1_4_0_wenable(ram_w4_l8192_id1_4_0_wenable),
    .ram_w4_l8192_id1_4_1_addr(ram_w4_l8192_id1_4_1_addr),
    .ram_w4_l8192_id1_4_1_rdata(ram_w4_l8192_id1_4_1_rdata),
    .ram_w4_l8192_id1_4_1_wdata(ram_w4_l8192_id1_4_1_wdata),
    .ram_w4_l8192_id1_4_1_wenable(ram_w4_l8192_id1_4_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id1_5_0_addr;
  wire [4-1:0] ram_w4_l8192_id1_5_0_rdata;
  reg [4-1:0] ram_w4_l8192_id1_5_0_wdata;
  reg ram_w4_l8192_id1_5_0_wenable;
  reg [10-1:0] ram_w4_l8192_id1_5_1_addr;
  wire [4-1:0] ram_w4_l8192_id1_5_1_rdata;
  reg [4-1:0] ram_w4_l8192_id1_5_1_wdata;
  reg ram_w4_l8192_id1_5_1_wenable;

  ram_w4_l8192_id1_5
  inst_ram_w4_l8192_id1_5
  (
    .CLK(CLK),
    .ram_w4_l8192_id1_5_0_addr(ram_w4_l8192_id1_5_0_addr),
    .ram_w4_l8192_id1_5_0_rdata(ram_w4_l8192_id1_5_0_rdata),
    .ram_w4_l8192_id1_5_0_wdata(ram_w4_l8192_id1_5_0_wdata),
    .ram_w4_l8192_id1_5_0_wenable(ram_w4_l8192_id1_5_0_wenable),
    .ram_w4_l8192_id1_5_1_addr(ram_w4_l8192_id1_5_1_addr),
    .ram_w4_l8192_id1_5_1_rdata(ram_w4_l8192_id1_5_1_rdata),
    .ram_w4_l8192_id1_5_1_wdata(ram_w4_l8192_id1_5_1_wdata),
    .ram_w4_l8192_id1_5_1_wenable(ram_w4_l8192_id1_5_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id1_6_0_addr;
  wire [4-1:0] ram_w4_l8192_id1_6_0_rdata;
  reg [4-1:0] ram_w4_l8192_id1_6_0_wdata;
  reg ram_w4_l8192_id1_6_0_wenable;
  reg [10-1:0] ram_w4_l8192_id1_6_1_addr;
  wire [4-1:0] ram_w4_l8192_id1_6_1_rdata;
  reg [4-1:0] ram_w4_l8192_id1_6_1_wdata;
  reg ram_w4_l8192_id1_6_1_wenable;

  ram_w4_l8192_id1_6
  inst_ram_w4_l8192_id1_6
  (
    .CLK(CLK),
    .ram_w4_l8192_id1_6_0_addr(ram_w4_l8192_id1_6_0_addr),
    .ram_w4_l8192_id1_6_0_rdata(ram_w4_l8192_id1_6_0_rdata),
    .ram_w4_l8192_id1_6_0_wdata(ram_w4_l8192_id1_6_0_wdata),
    .ram_w4_l8192_id1_6_0_wenable(ram_w4_l8192_id1_6_0_wenable),
    .ram_w4_l8192_id1_6_1_addr(ram_w4_l8192_id1_6_1_addr),
    .ram_w4_l8192_id1_6_1_rdata(ram_w4_l8192_id1_6_1_rdata),
    .ram_w4_l8192_id1_6_1_wdata(ram_w4_l8192_id1_6_1_wdata),
    .ram_w4_l8192_id1_6_1_wenable(ram_w4_l8192_id1_6_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id1_7_0_addr;
  wire [4-1:0] ram_w4_l8192_id1_7_0_rdata;
  reg [4-1:0] ram_w4_l8192_id1_7_0_wdata;
  reg ram_w4_l8192_id1_7_0_wenable;
  reg [10-1:0] ram_w4_l8192_id1_7_1_addr;
  wire [4-1:0] ram_w4_l8192_id1_7_1_rdata;
  reg [4-1:0] ram_w4_l8192_id1_7_1_wdata;
  reg ram_w4_l8192_id1_7_1_wenable;

  ram_w4_l8192_id1_7
  inst_ram_w4_l8192_id1_7
  (
    .CLK(CLK),
    .ram_w4_l8192_id1_7_0_addr(ram_w4_l8192_id1_7_0_addr),
    .ram_w4_l8192_id1_7_0_rdata(ram_w4_l8192_id1_7_0_rdata),
    .ram_w4_l8192_id1_7_0_wdata(ram_w4_l8192_id1_7_0_wdata),
    .ram_w4_l8192_id1_7_0_wenable(ram_w4_l8192_id1_7_0_wenable),
    .ram_w4_l8192_id1_7_1_addr(ram_w4_l8192_id1_7_1_addr),
    .ram_w4_l8192_id1_7_1_rdata(ram_w4_l8192_id1_7_1_rdata),
    .ram_w4_l8192_id1_7_1_wdata(ram_w4_l8192_id1_7_1_wdata),
    .ram_w4_l8192_id1_7_1_wenable(ram_w4_l8192_id1_7_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id2_0_0_addr;
  wire [4-1:0] ram_w4_l8192_id2_0_0_rdata;
  reg [4-1:0] ram_w4_l8192_id2_0_0_wdata;
  reg ram_w4_l8192_id2_0_0_wenable;
  reg [10-1:0] ram_w4_l8192_id2_0_1_addr;
  wire [4-1:0] ram_w4_l8192_id2_0_1_rdata;
  reg [4-1:0] ram_w4_l8192_id2_0_1_wdata;
  reg ram_w4_l8192_id2_0_1_wenable;

  ram_w4_l8192_id2_0
  inst_ram_w4_l8192_id2_0
  (
    .CLK(CLK),
    .ram_w4_l8192_id2_0_0_addr(ram_w4_l8192_id2_0_0_addr),
    .ram_w4_l8192_id2_0_0_rdata(ram_w4_l8192_id2_0_0_rdata),
    .ram_w4_l8192_id2_0_0_wdata(ram_w4_l8192_id2_0_0_wdata),
    .ram_w4_l8192_id2_0_0_wenable(ram_w4_l8192_id2_0_0_wenable),
    .ram_w4_l8192_id2_0_1_addr(ram_w4_l8192_id2_0_1_addr),
    .ram_w4_l8192_id2_0_1_rdata(ram_w4_l8192_id2_0_1_rdata),
    .ram_w4_l8192_id2_0_1_wdata(ram_w4_l8192_id2_0_1_wdata),
    .ram_w4_l8192_id2_0_1_wenable(ram_w4_l8192_id2_0_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id2_1_0_addr;
  wire [4-1:0] ram_w4_l8192_id2_1_0_rdata;
  reg [4-1:0] ram_w4_l8192_id2_1_0_wdata;
  reg ram_w4_l8192_id2_1_0_wenable;
  reg [10-1:0] ram_w4_l8192_id2_1_1_addr;
  wire [4-1:0] ram_w4_l8192_id2_1_1_rdata;
  reg [4-1:0] ram_w4_l8192_id2_1_1_wdata;
  reg ram_w4_l8192_id2_1_1_wenable;

  ram_w4_l8192_id2_1
  inst_ram_w4_l8192_id2_1
  (
    .CLK(CLK),
    .ram_w4_l8192_id2_1_0_addr(ram_w4_l8192_id2_1_0_addr),
    .ram_w4_l8192_id2_1_0_rdata(ram_w4_l8192_id2_1_0_rdata),
    .ram_w4_l8192_id2_1_0_wdata(ram_w4_l8192_id2_1_0_wdata),
    .ram_w4_l8192_id2_1_0_wenable(ram_w4_l8192_id2_1_0_wenable),
    .ram_w4_l8192_id2_1_1_addr(ram_w4_l8192_id2_1_1_addr),
    .ram_w4_l8192_id2_1_1_rdata(ram_w4_l8192_id2_1_1_rdata),
    .ram_w4_l8192_id2_1_1_wdata(ram_w4_l8192_id2_1_1_wdata),
    .ram_w4_l8192_id2_1_1_wenable(ram_w4_l8192_id2_1_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id2_2_0_addr;
  wire [4-1:0] ram_w4_l8192_id2_2_0_rdata;
  reg [4-1:0] ram_w4_l8192_id2_2_0_wdata;
  reg ram_w4_l8192_id2_2_0_wenable;
  reg [10-1:0] ram_w4_l8192_id2_2_1_addr;
  wire [4-1:0] ram_w4_l8192_id2_2_1_rdata;
  reg [4-1:0] ram_w4_l8192_id2_2_1_wdata;
  reg ram_w4_l8192_id2_2_1_wenable;

  ram_w4_l8192_id2_2
  inst_ram_w4_l8192_id2_2
  (
    .CLK(CLK),
    .ram_w4_l8192_id2_2_0_addr(ram_w4_l8192_id2_2_0_addr),
    .ram_w4_l8192_id2_2_0_rdata(ram_w4_l8192_id2_2_0_rdata),
    .ram_w4_l8192_id2_2_0_wdata(ram_w4_l8192_id2_2_0_wdata),
    .ram_w4_l8192_id2_2_0_wenable(ram_w4_l8192_id2_2_0_wenable),
    .ram_w4_l8192_id2_2_1_addr(ram_w4_l8192_id2_2_1_addr),
    .ram_w4_l8192_id2_2_1_rdata(ram_w4_l8192_id2_2_1_rdata),
    .ram_w4_l8192_id2_2_1_wdata(ram_w4_l8192_id2_2_1_wdata),
    .ram_w4_l8192_id2_2_1_wenable(ram_w4_l8192_id2_2_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id2_3_0_addr;
  wire [4-1:0] ram_w4_l8192_id2_3_0_rdata;
  reg [4-1:0] ram_w4_l8192_id2_3_0_wdata;
  reg ram_w4_l8192_id2_3_0_wenable;
  reg [10-1:0] ram_w4_l8192_id2_3_1_addr;
  wire [4-1:0] ram_w4_l8192_id2_3_1_rdata;
  reg [4-1:0] ram_w4_l8192_id2_3_1_wdata;
  reg ram_w4_l8192_id2_3_1_wenable;

  ram_w4_l8192_id2_3
  inst_ram_w4_l8192_id2_3
  (
    .CLK(CLK),
    .ram_w4_l8192_id2_3_0_addr(ram_w4_l8192_id2_3_0_addr),
    .ram_w4_l8192_id2_3_0_rdata(ram_w4_l8192_id2_3_0_rdata),
    .ram_w4_l8192_id2_3_0_wdata(ram_w4_l8192_id2_3_0_wdata),
    .ram_w4_l8192_id2_3_0_wenable(ram_w4_l8192_id2_3_0_wenable),
    .ram_w4_l8192_id2_3_1_addr(ram_w4_l8192_id2_3_1_addr),
    .ram_w4_l8192_id2_3_1_rdata(ram_w4_l8192_id2_3_1_rdata),
    .ram_w4_l8192_id2_3_1_wdata(ram_w4_l8192_id2_3_1_wdata),
    .ram_w4_l8192_id2_3_1_wenable(ram_w4_l8192_id2_3_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id2_4_0_addr;
  wire [4-1:0] ram_w4_l8192_id2_4_0_rdata;
  reg [4-1:0] ram_w4_l8192_id2_4_0_wdata;
  reg ram_w4_l8192_id2_4_0_wenable;
  reg [10-1:0] ram_w4_l8192_id2_4_1_addr;
  wire [4-1:0] ram_w4_l8192_id2_4_1_rdata;
  reg [4-1:0] ram_w4_l8192_id2_4_1_wdata;
  reg ram_w4_l8192_id2_4_1_wenable;

  ram_w4_l8192_id2_4
  inst_ram_w4_l8192_id2_4
  (
    .CLK(CLK),
    .ram_w4_l8192_id2_4_0_addr(ram_w4_l8192_id2_4_0_addr),
    .ram_w4_l8192_id2_4_0_rdata(ram_w4_l8192_id2_4_0_rdata),
    .ram_w4_l8192_id2_4_0_wdata(ram_w4_l8192_id2_4_0_wdata),
    .ram_w4_l8192_id2_4_0_wenable(ram_w4_l8192_id2_4_0_wenable),
    .ram_w4_l8192_id2_4_1_addr(ram_w4_l8192_id2_4_1_addr),
    .ram_w4_l8192_id2_4_1_rdata(ram_w4_l8192_id2_4_1_rdata),
    .ram_w4_l8192_id2_4_1_wdata(ram_w4_l8192_id2_4_1_wdata),
    .ram_w4_l8192_id2_4_1_wenable(ram_w4_l8192_id2_4_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id2_5_0_addr;
  wire [4-1:0] ram_w4_l8192_id2_5_0_rdata;
  reg [4-1:0] ram_w4_l8192_id2_5_0_wdata;
  reg ram_w4_l8192_id2_5_0_wenable;
  reg [10-1:0] ram_w4_l8192_id2_5_1_addr;
  wire [4-1:0] ram_w4_l8192_id2_5_1_rdata;
  reg [4-1:0] ram_w4_l8192_id2_5_1_wdata;
  reg ram_w4_l8192_id2_5_1_wenable;

  ram_w4_l8192_id2_5
  inst_ram_w4_l8192_id2_5
  (
    .CLK(CLK),
    .ram_w4_l8192_id2_5_0_addr(ram_w4_l8192_id2_5_0_addr),
    .ram_w4_l8192_id2_5_0_rdata(ram_w4_l8192_id2_5_0_rdata),
    .ram_w4_l8192_id2_5_0_wdata(ram_w4_l8192_id2_5_0_wdata),
    .ram_w4_l8192_id2_5_0_wenable(ram_w4_l8192_id2_5_0_wenable),
    .ram_w4_l8192_id2_5_1_addr(ram_w4_l8192_id2_5_1_addr),
    .ram_w4_l8192_id2_5_1_rdata(ram_w4_l8192_id2_5_1_rdata),
    .ram_w4_l8192_id2_5_1_wdata(ram_w4_l8192_id2_5_1_wdata),
    .ram_w4_l8192_id2_5_1_wenable(ram_w4_l8192_id2_5_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id2_6_0_addr;
  wire [4-1:0] ram_w4_l8192_id2_6_0_rdata;
  reg [4-1:0] ram_w4_l8192_id2_6_0_wdata;
  reg ram_w4_l8192_id2_6_0_wenable;
  reg [10-1:0] ram_w4_l8192_id2_6_1_addr;
  wire [4-1:0] ram_w4_l8192_id2_6_1_rdata;
  reg [4-1:0] ram_w4_l8192_id2_6_1_wdata;
  reg ram_w4_l8192_id2_6_1_wenable;

  ram_w4_l8192_id2_6
  inst_ram_w4_l8192_id2_6
  (
    .CLK(CLK),
    .ram_w4_l8192_id2_6_0_addr(ram_w4_l8192_id2_6_0_addr),
    .ram_w4_l8192_id2_6_0_rdata(ram_w4_l8192_id2_6_0_rdata),
    .ram_w4_l8192_id2_6_0_wdata(ram_w4_l8192_id2_6_0_wdata),
    .ram_w4_l8192_id2_6_0_wenable(ram_w4_l8192_id2_6_0_wenable),
    .ram_w4_l8192_id2_6_1_addr(ram_w4_l8192_id2_6_1_addr),
    .ram_w4_l8192_id2_6_1_rdata(ram_w4_l8192_id2_6_1_rdata),
    .ram_w4_l8192_id2_6_1_wdata(ram_w4_l8192_id2_6_1_wdata),
    .ram_w4_l8192_id2_6_1_wenable(ram_w4_l8192_id2_6_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id2_7_0_addr;
  wire [4-1:0] ram_w4_l8192_id2_7_0_rdata;
  reg [4-1:0] ram_w4_l8192_id2_7_0_wdata;
  reg ram_w4_l8192_id2_7_0_wenable;
  reg [10-1:0] ram_w4_l8192_id2_7_1_addr;
  wire [4-1:0] ram_w4_l8192_id2_7_1_rdata;
  reg [4-1:0] ram_w4_l8192_id2_7_1_wdata;
  reg ram_w4_l8192_id2_7_1_wenable;

  ram_w4_l8192_id2_7
  inst_ram_w4_l8192_id2_7
  (
    .CLK(CLK),
    .ram_w4_l8192_id2_7_0_addr(ram_w4_l8192_id2_7_0_addr),
    .ram_w4_l8192_id2_7_0_rdata(ram_w4_l8192_id2_7_0_rdata),
    .ram_w4_l8192_id2_7_0_wdata(ram_w4_l8192_id2_7_0_wdata),
    .ram_w4_l8192_id2_7_0_wenable(ram_w4_l8192_id2_7_0_wenable),
    .ram_w4_l8192_id2_7_1_addr(ram_w4_l8192_id2_7_1_addr),
    .ram_w4_l8192_id2_7_1_rdata(ram_w4_l8192_id2_7_1_rdata),
    .ram_w4_l8192_id2_7_1_wdata(ram_w4_l8192_id2_7_1_wdata),
    .ram_w4_l8192_id2_7_1_wenable(ram_w4_l8192_id2_7_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id3_0_0_addr;
  wire [4-1:0] ram_w4_l8192_id3_0_0_rdata;
  reg [4-1:0] ram_w4_l8192_id3_0_0_wdata;
  reg ram_w4_l8192_id3_0_0_wenable;
  reg [10-1:0] ram_w4_l8192_id3_0_1_addr;
  wire [4-1:0] ram_w4_l8192_id3_0_1_rdata;
  reg [4-1:0] ram_w4_l8192_id3_0_1_wdata;
  reg ram_w4_l8192_id3_0_1_wenable;

  ram_w4_l8192_id3_0
  inst_ram_w4_l8192_id3_0
  (
    .CLK(CLK),
    .ram_w4_l8192_id3_0_0_addr(ram_w4_l8192_id3_0_0_addr),
    .ram_w4_l8192_id3_0_0_rdata(ram_w4_l8192_id3_0_0_rdata),
    .ram_w4_l8192_id3_0_0_wdata(ram_w4_l8192_id3_0_0_wdata),
    .ram_w4_l8192_id3_0_0_wenable(ram_w4_l8192_id3_0_0_wenable),
    .ram_w4_l8192_id3_0_1_addr(ram_w4_l8192_id3_0_1_addr),
    .ram_w4_l8192_id3_0_1_rdata(ram_w4_l8192_id3_0_1_rdata),
    .ram_w4_l8192_id3_0_1_wdata(ram_w4_l8192_id3_0_1_wdata),
    .ram_w4_l8192_id3_0_1_wenable(ram_w4_l8192_id3_0_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id3_1_0_addr;
  wire [4-1:0] ram_w4_l8192_id3_1_0_rdata;
  reg [4-1:0] ram_w4_l8192_id3_1_0_wdata;
  reg ram_w4_l8192_id3_1_0_wenable;
  reg [10-1:0] ram_w4_l8192_id3_1_1_addr;
  wire [4-1:0] ram_w4_l8192_id3_1_1_rdata;
  reg [4-1:0] ram_w4_l8192_id3_1_1_wdata;
  reg ram_w4_l8192_id3_1_1_wenable;

  ram_w4_l8192_id3_1
  inst_ram_w4_l8192_id3_1
  (
    .CLK(CLK),
    .ram_w4_l8192_id3_1_0_addr(ram_w4_l8192_id3_1_0_addr),
    .ram_w4_l8192_id3_1_0_rdata(ram_w4_l8192_id3_1_0_rdata),
    .ram_w4_l8192_id3_1_0_wdata(ram_w4_l8192_id3_1_0_wdata),
    .ram_w4_l8192_id3_1_0_wenable(ram_w4_l8192_id3_1_0_wenable),
    .ram_w4_l8192_id3_1_1_addr(ram_w4_l8192_id3_1_1_addr),
    .ram_w4_l8192_id3_1_1_rdata(ram_w4_l8192_id3_1_1_rdata),
    .ram_w4_l8192_id3_1_1_wdata(ram_w4_l8192_id3_1_1_wdata),
    .ram_w4_l8192_id3_1_1_wenable(ram_w4_l8192_id3_1_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id3_2_0_addr;
  wire [4-1:0] ram_w4_l8192_id3_2_0_rdata;
  reg [4-1:0] ram_w4_l8192_id3_2_0_wdata;
  reg ram_w4_l8192_id3_2_0_wenable;
  reg [10-1:0] ram_w4_l8192_id3_2_1_addr;
  wire [4-1:0] ram_w4_l8192_id3_2_1_rdata;
  reg [4-1:0] ram_w4_l8192_id3_2_1_wdata;
  reg ram_w4_l8192_id3_2_1_wenable;

  ram_w4_l8192_id3_2
  inst_ram_w4_l8192_id3_2
  (
    .CLK(CLK),
    .ram_w4_l8192_id3_2_0_addr(ram_w4_l8192_id3_2_0_addr),
    .ram_w4_l8192_id3_2_0_rdata(ram_w4_l8192_id3_2_0_rdata),
    .ram_w4_l8192_id3_2_0_wdata(ram_w4_l8192_id3_2_0_wdata),
    .ram_w4_l8192_id3_2_0_wenable(ram_w4_l8192_id3_2_0_wenable),
    .ram_w4_l8192_id3_2_1_addr(ram_w4_l8192_id3_2_1_addr),
    .ram_w4_l8192_id3_2_1_rdata(ram_w4_l8192_id3_2_1_rdata),
    .ram_w4_l8192_id3_2_1_wdata(ram_w4_l8192_id3_2_1_wdata),
    .ram_w4_l8192_id3_2_1_wenable(ram_w4_l8192_id3_2_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id3_3_0_addr;
  wire [4-1:0] ram_w4_l8192_id3_3_0_rdata;
  reg [4-1:0] ram_w4_l8192_id3_3_0_wdata;
  reg ram_w4_l8192_id3_3_0_wenable;
  reg [10-1:0] ram_w4_l8192_id3_3_1_addr;
  wire [4-1:0] ram_w4_l8192_id3_3_1_rdata;
  reg [4-1:0] ram_w4_l8192_id3_3_1_wdata;
  reg ram_w4_l8192_id3_3_1_wenable;

  ram_w4_l8192_id3_3
  inst_ram_w4_l8192_id3_3
  (
    .CLK(CLK),
    .ram_w4_l8192_id3_3_0_addr(ram_w4_l8192_id3_3_0_addr),
    .ram_w4_l8192_id3_3_0_rdata(ram_w4_l8192_id3_3_0_rdata),
    .ram_w4_l8192_id3_3_0_wdata(ram_w4_l8192_id3_3_0_wdata),
    .ram_w4_l8192_id3_3_0_wenable(ram_w4_l8192_id3_3_0_wenable),
    .ram_w4_l8192_id3_3_1_addr(ram_w4_l8192_id3_3_1_addr),
    .ram_w4_l8192_id3_3_1_rdata(ram_w4_l8192_id3_3_1_rdata),
    .ram_w4_l8192_id3_3_1_wdata(ram_w4_l8192_id3_3_1_wdata),
    .ram_w4_l8192_id3_3_1_wenable(ram_w4_l8192_id3_3_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id3_4_0_addr;
  wire [4-1:0] ram_w4_l8192_id3_4_0_rdata;
  reg [4-1:0] ram_w4_l8192_id3_4_0_wdata;
  reg ram_w4_l8192_id3_4_0_wenable;
  reg [10-1:0] ram_w4_l8192_id3_4_1_addr;
  wire [4-1:0] ram_w4_l8192_id3_4_1_rdata;
  reg [4-1:0] ram_w4_l8192_id3_4_1_wdata;
  reg ram_w4_l8192_id3_4_1_wenable;

  ram_w4_l8192_id3_4
  inst_ram_w4_l8192_id3_4
  (
    .CLK(CLK),
    .ram_w4_l8192_id3_4_0_addr(ram_w4_l8192_id3_4_0_addr),
    .ram_w4_l8192_id3_4_0_rdata(ram_w4_l8192_id3_4_0_rdata),
    .ram_w4_l8192_id3_4_0_wdata(ram_w4_l8192_id3_4_0_wdata),
    .ram_w4_l8192_id3_4_0_wenable(ram_w4_l8192_id3_4_0_wenable),
    .ram_w4_l8192_id3_4_1_addr(ram_w4_l8192_id3_4_1_addr),
    .ram_w4_l8192_id3_4_1_rdata(ram_w4_l8192_id3_4_1_rdata),
    .ram_w4_l8192_id3_4_1_wdata(ram_w4_l8192_id3_4_1_wdata),
    .ram_w4_l8192_id3_4_1_wenable(ram_w4_l8192_id3_4_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id3_5_0_addr;
  wire [4-1:0] ram_w4_l8192_id3_5_0_rdata;
  reg [4-1:0] ram_w4_l8192_id3_5_0_wdata;
  reg ram_w4_l8192_id3_5_0_wenable;
  reg [10-1:0] ram_w4_l8192_id3_5_1_addr;
  wire [4-1:0] ram_w4_l8192_id3_5_1_rdata;
  reg [4-1:0] ram_w4_l8192_id3_5_1_wdata;
  reg ram_w4_l8192_id3_5_1_wenable;

  ram_w4_l8192_id3_5
  inst_ram_w4_l8192_id3_5
  (
    .CLK(CLK),
    .ram_w4_l8192_id3_5_0_addr(ram_w4_l8192_id3_5_0_addr),
    .ram_w4_l8192_id3_5_0_rdata(ram_w4_l8192_id3_5_0_rdata),
    .ram_w4_l8192_id3_5_0_wdata(ram_w4_l8192_id3_5_0_wdata),
    .ram_w4_l8192_id3_5_0_wenable(ram_w4_l8192_id3_5_0_wenable),
    .ram_w4_l8192_id3_5_1_addr(ram_w4_l8192_id3_5_1_addr),
    .ram_w4_l8192_id3_5_1_rdata(ram_w4_l8192_id3_5_1_rdata),
    .ram_w4_l8192_id3_5_1_wdata(ram_w4_l8192_id3_5_1_wdata),
    .ram_w4_l8192_id3_5_1_wenable(ram_w4_l8192_id3_5_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id3_6_0_addr;
  wire [4-1:0] ram_w4_l8192_id3_6_0_rdata;
  reg [4-1:0] ram_w4_l8192_id3_6_0_wdata;
  reg ram_w4_l8192_id3_6_0_wenable;
  reg [10-1:0] ram_w4_l8192_id3_6_1_addr;
  wire [4-1:0] ram_w4_l8192_id3_6_1_rdata;
  reg [4-1:0] ram_w4_l8192_id3_6_1_wdata;
  reg ram_w4_l8192_id3_6_1_wenable;

  ram_w4_l8192_id3_6
  inst_ram_w4_l8192_id3_6
  (
    .CLK(CLK),
    .ram_w4_l8192_id3_6_0_addr(ram_w4_l8192_id3_6_0_addr),
    .ram_w4_l8192_id3_6_0_rdata(ram_w4_l8192_id3_6_0_rdata),
    .ram_w4_l8192_id3_6_0_wdata(ram_w4_l8192_id3_6_0_wdata),
    .ram_w4_l8192_id3_6_0_wenable(ram_w4_l8192_id3_6_0_wenable),
    .ram_w4_l8192_id3_6_1_addr(ram_w4_l8192_id3_6_1_addr),
    .ram_w4_l8192_id3_6_1_rdata(ram_w4_l8192_id3_6_1_rdata),
    .ram_w4_l8192_id3_6_1_wdata(ram_w4_l8192_id3_6_1_wdata),
    .ram_w4_l8192_id3_6_1_wenable(ram_w4_l8192_id3_6_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id3_7_0_addr;
  wire [4-1:0] ram_w4_l8192_id3_7_0_rdata;
  reg [4-1:0] ram_w4_l8192_id3_7_0_wdata;
  reg ram_w4_l8192_id3_7_0_wenable;
  reg [10-1:0] ram_w4_l8192_id3_7_1_addr;
  wire [4-1:0] ram_w4_l8192_id3_7_1_rdata;
  reg [4-1:0] ram_w4_l8192_id3_7_1_wdata;
  reg ram_w4_l8192_id3_7_1_wenable;

  ram_w4_l8192_id3_7
  inst_ram_w4_l8192_id3_7
  (
    .CLK(CLK),
    .ram_w4_l8192_id3_7_0_addr(ram_w4_l8192_id3_7_0_addr),
    .ram_w4_l8192_id3_7_0_rdata(ram_w4_l8192_id3_7_0_rdata),
    .ram_w4_l8192_id3_7_0_wdata(ram_w4_l8192_id3_7_0_wdata),
    .ram_w4_l8192_id3_7_0_wenable(ram_w4_l8192_id3_7_0_wenable),
    .ram_w4_l8192_id3_7_1_addr(ram_w4_l8192_id3_7_1_addr),
    .ram_w4_l8192_id3_7_1_rdata(ram_w4_l8192_id3_7_1_rdata),
    .ram_w4_l8192_id3_7_1_wdata(ram_w4_l8192_id3_7_1_wdata),
    .ram_w4_l8192_id3_7_1_wenable(ram_w4_l8192_id3_7_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id4_0_0_addr;
  wire [4-1:0] ram_w4_l8192_id4_0_0_rdata;
  reg [4-1:0] ram_w4_l8192_id4_0_0_wdata;
  reg ram_w4_l8192_id4_0_0_wenable;
  reg [10-1:0] ram_w4_l8192_id4_0_1_addr;
  wire [4-1:0] ram_w4_l8192_id4_0_1_rdata;
  reg [4-1:0] ram_w4_l8192_id4_0_1_wdata;
  reg ram_w4_l8192_id4_0_1_wenable;

  ram_w4_l8192_id4_0
  inst_ram_w4_l8192_id4_0
  (
    .CLK(CLK),
    .ram_w4_l8192_id4_0_0_addr(ram_w4_l8192_id4_0_0_addr),
    .ram_w4_l8192_id4_0_0_rdata(ram_w4_l8192_id4_0_0_rdata),
    .ram_w4_l8192_id4_0_0_wdata(ram_w4_l8192_id4_0_0_wdata),
    .ram_w4_l8192_id4_0_0_wenable(ram_w4_l8192_id4_0_0_wenable),
    .ram_w4_l8192_id4_0_1_addr(ram_w4_l8192_id4_0_1_addr),
    .ram_w4_l8192_id4_0_1_rdata(ram_w4_l8192_id4_0_1_rdata),
    .ram_w4_l8192_id4_0_1_wdata(ram_w4_l8192_id4_0_1_wdata),
    .ram_w4_l8192_id4_0_1_wenable(ram_w4_l8192_id4_0_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id4_1_0_addr;
  wire [4-1:0] ram_w4_l8192_id4_1_0_rdata;
  reg [4-1:0] ram_w4_l8192_id4_1_0_wdata;
  reg ram_w4_l8192_id4_1_0_wenable;
  reg [10-1:0] ram_w4_l8192_id4_1_1_addr;
  wire [4-1:0] ram_w4_l8192_id4_1_1_rdata;
  reg [4-1:0] ram_w4_l8192_id4_1_1_wdata;
  reg ram_w4_l8192_id4_1_1_wenable;

  ram_w4_l8192_id4_1
  inst_ram_w4_l8192_id4_1
  (
    .CLK(CLK),
    .ram_w4_l8192_id4_1_0_addr(ram_w4_l8192_id4_1_0_addr),
    .ram_w4_l8192_id4_1_0_rdata(ram_w4_l8192_id4_1_0_rdata),
    .ram_w4_l8192_id4_1_0_wdata(ram_w4_l8192_id4_1_0_wdata),
    .ram_w4_l8192_id4_1_0_wenable(ram_w4_l8192_id4_1_0_wenable),
    .ram_w4_l8192_id4_1_1_addr(ram_w4_l8192_id4_1_1_addr),
    .ram_w4_l8192_id4_1_1_rdata(ram_w4_l8192_id4_1_1_rdata),
    .ram_w4_l8192_id4_1_1_wdata(ram_w4_l8192_id4_1_1_wdata),
    .ram_w4_l8192_id4_1_1_wenable(ram_w4_l8192_id4_1_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id4_2_0_addr;
  wire [4-1:0] ram_w4_l8192_id4_2_0_rdata;
  reg [4-1:0] ram_w4_l8192_id4_2_0_wdata;
  reg ram_w4_l8192_id4_2_0_wenable;
  reg [10-1:0] ram_w4_l8192_id4_2_1_addr;
  wire [4-1:0] ram_w4_l8192_id4_2_1_rdata;
  reg [4-1:0] ram_w4_l8192_id4_2_1_wdata;
  reg ram_w4_l8192_id4_2_1_wenable;

  ram_w4_l8192_id4_2
  inst_ram_w4_l8192_id4_2
  (
    .CLK(CLK),
    .ram_w4_l8192_id4_2_0_addr(ram_w4_l8192_id4_2_0_addr),
    .ram_w4_l8192_id4_2_0_rdata(ram_w4_l8192_id4_2_0_rdata),
    .ram_w4_l8192_id4_2_0_wdata(ram_w4_l8192_id4_2_0_wdata),
    .ram_w4_l8192_id4_2_0_wenable(ram_w4_l8192_id4_2_0_wenable),
    .ram_w4_l8192_id4_2_1_addr(ram_w4_l8192_id4_2_1_addr),
    .ram_w4_l8192_id4_2_1_rdata(ram_w4_l8192_id4_2_1_rdata),
    .ram_w4_l8192_id4_2_1_wdata(ram_w4_l8192_id4_2_1_wdata),
    .ram_w4_l8192_id4_2_1_wenable(ram_w4_l8192_id4_2_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id4_3_0_addr;
  wire [4-1:0] ram_w4_l8192_id4_3_0_rdata;
  reg [4-1:0] ram_w4_l8192_id4_3_0_wdata;
  reg ram_w4_l8192_id4_3_0_wenable;
  reg [10-1:0] ram_w4_l8192_id4_3_1_addr;
  wire [4-1:0] ram_w4_l8192_id4_3_1_rdata;
  reg [4-1:0] ram_w4_l8192_id4_3_1_wdata;
  reg ram_w4_l8192_id4_3_1_wenable;

  ram_w4_l8192_id4_3
  inst_ram_w4_l8192_id4_3
  (
    .CLK(CLK),
    .ram_w4_l8192_id4_3_0_addr(ram_w4_l8192_id4_3_0_addr),
    .ram_w4_l8192_id4_3_0_rdata(ram_w4_l8192_id4_3_0_rdata),
    .ram_w4_l8192_id4_3_0_wdata(ram_w4_l8192_id4_3_0_wdata),
    .ram_w4_l8192_id4_3_0_wenable(ram_w4_l8192_id4_3_0_wenable),
    .ram_w4_l8192_id4_3_1_addr(ram_w4_l8192_id4_3_1_addr),
    .ram_w4_l8192_id4_3_1_rdata(ram_w4_l8192_id4_3_1_rdata),
    .ram_w4_l8192_id4_3_1_wdata(ram_w4_l8192_id4_3_1_wdata),
    .ram_w4_l8192_id4_3_1_wenable(ram_w4_l8192_id4_3_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id4_4_0_addr;
  wire [4-1:0] ram_w4_l8192_id4_4_0_rdata;
  reg [4-1:0] ram_w4_l8192_id4_4_0_wdata;
  reg ram_w4_l8192_id4_4_0_wenable;
  reg [10-1:0] ram_w4_l8192_id4_4_1_addr;
  wire [4-1:0] ram_w4_l8192_id4_4_1_rdata;
  reg [4-1:0] ram_w4_l8192_id4_4_1_wdata;
  reg ram_w4_l8192_id4_4_1_wenable;

  ram_w4_l8192_id4_4
  inst_ram_w4_l8192_id4_4
  (
    .CLK(CLK),
    .ram_w4_l8192_id4_4_0_addr(ram_w4_l8192_id4_4_0_addr),
    .ram_w4_l8192_id4_4_0_rdata(ram_w4_l8192_id4_4_0_rdata),
    .ram_w4_l8192_id4_4_0_wdata(ram_w4_l8192_id4_4_0_wdata),
    .ram_w4_l8192_id4_4_0_wenable(ram_w4_l8192_id4_4_0_wenable),
    .ram_w4_l8192_id4_4_1_addr(ram_w4_l8192_id4_4_1_addr),
    .ram_w4_l8192_id4_4_1_rdata(ram_w4_l8192_id4_4_1_rdata),
    .ram_w4_l8192_id4_4_1_wdata(ram_w4_l8192_id4_4_1_wdata),
    .ram_w4_l8192_id4_4_1_wenable(ram_w4_l8192_id4_4_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id4_5_0_addr;
  wire [4-1:0] ram_w4_l8192_id4_5_0_rdata;
  reg [4-1:0] ram_w4_l8192_id4_5_0_wdata;
  reg ram_w4_l8192_id4_5_0_wenable;
  reg [10-1:0] ram_w4_l8192_id4_5_1_addr;
  wire [4-1:0] ram_w4_l8192_id4_5_1_rdata;
  reg [4-1:0] ram_w4_l8192_id4_5_1_wdata;
  reg ram_w4_l8192_id4_5_1_wenable;

  ram_w4_l8192_id4_5
  inst_ram_w4_l8192_id4_5
  (
    .CLK(CLK),
    .ram_w4_l8192_id4_5_0_addr(ram_w4_l8192_id4_5_0_addr),
    .ram_w4_l8192_id4_5_0_rdata(ram_w4_l8192_id4_5_0_rdata),
    .ram_w4_l8192_id4_5_0_wdata(ram_w4_l8192_id4_5_0_wdata),
    .ram_w4_l8192_id4_5_0_wenable(ram_w4_l8192_id4_5_0_wenable),
    .ram_w4_l8192_id4_5_1_addr(ram_w4_l8192_id4_5_1_addr),
    .ram_w4_l8192_id4_5_1_rdata(ram_w4_l8192_id4_5_1_rdata),
    .ram_w4_l8192_id4_5_1_wdata(ram_w4_l8192_id4_5_1_wdata),
    .ram_w4_l8192_id4_5_1_wenable(ram_w4_l8192_id4_5_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id4_6_0_addr;
  wire [4-1:0] ram_w4_l8192_id4_6_0_rdata;
  reg [4-1:0] ram_w4_l8192_id4_6_0_wdata;
  reg ram_w4_l8192_id4_6_0_wenable;
  reg [10-1:0] ram_w4_l8192_id4_6_1_addr;
  wire [4-1:0] ram_w4_l8192_id4_6_1_rdata;
  reg [4-1:0] ram_w4_l8192_id4_6_1_wdata;
  reg ram_w4_l8192_id4_6_1_wenable;

  ram_w4_l8192_id4_6
  inst_ram_w4_l8192_id4_6
  (
    .CLK(CLK),
    .ram_w4_l8192_id4_6_0_addr(ram_w4_l8192_id4_6_0_addr),
    .ram_w4_l8192_id4_6_0_rdata(ram_w4_l8192_id4_6_0_rdata),
    .ram_w4_l8192_id4_6_0_wdata(ram_w4_l8192_id4_6_0_wdata),
    .ram_w4_l8192_id4_6_0_wenable(ram_w4_l8192_id4_6_0_wenable),
    .ram_w4_l8192_id4_6_1_addr(ram_w4_l8192_id4_6_1_addr),
    .ram_w4_l8192_id4_6_1_rdata(ram_w4_l8192_id4_6_1_rdata),
    .ram_w4_l8192_id4_6_1_wdata(ram_w4_l8192_id4_6_1_wdata),
    .ram_w4_l8192_id4_6_1_wenable(ram_w4_l8192_id4_6_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id4_7_0_addr;
  wire [4-1:0] ram_w4_l8192_id4_7_0_rdata;
  reg [4-1:0] ram_w4_l8192_id4_7_0_wdata;
  reg ram_w4_l8192_id4_7_0_wenable;
  reg [10-1:0] ram_w4_l8192_id4_7_1_addr;
  wire [4-1:0] ram_w4_l8192_id4_7_1_rdata;
  reg [4-1:0] ram_w4_l8192_id4_7_1_wdata;
  reg ram_w4_l8192_id4_7_1_wenable;

  ram_w4_l8192_id4_7
  inst_ram_w4_l8192_id4_7
  (
    .CLK(CLK),
    .ram_w4_l8192_id4_7_0_addr(ram_w4_l8192_id4_7_0_addr),
    .ram_w4_l8192_id4_7_0_rdata(ram_w4_l8192_id4_7_0_rdata),
    .ram_w4_l8192_id4_7_0_wdata(ram_w4_l8192_id4_7_0_wdata),
    .ram_w4_l8192_id4_7_0_wenable(ram_w4_l8192_id4_7_0_wenable),
    .ram_w4_l8192_id4_7_1_addr(ram_w4_l8192_id4_7_1_addr),
    .ram_w4_l8192_id4_7_1_rdata(ram_w4_l8192_id4_7_1_rdata),
    .ram_w4_l8192_id4_7_1_wdata(ram_w4_l8192_id4_7_1_wdata),
    .ram_w4_l8192_id4_7_1_wenable(ram_w4_l8192_id4_7_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id5_0_0_addr;
  wire [4-1:0] ram_w4_l8192_id5_0_0_rdata;
  reg [4-1:0] ram_w4_l8192_id5_0_0_wdata;
  reg ram_w4_l8192_id5_0_0_wenable;
  reg [10-1:0] ram_w4_l8192_id5_0_1_addr;
  wire [4-1:0] ram_w4_l8192_id5_0_1_rdata;
  reg [4-1:0] ram_w4_l8192_id5_0_1_wdata;
  reg ram_w4_l8192_id5_0_1_wenable;

  ram_w4_l8192_id5_0
  inst_ram_w4_l8192_id5_0
  (
    .CLK(CLK),
    .ram_w4_l8192_id5_0_0_addr(ram_w4_l8192_id5_0_0_addr),
    .ram_w4_l8192_id5_0_0_rdata(ram_w4_l8192_id5_0_0_rdata),
    .ram_w4_l8192_id5_0_0_wdata(ram_w4_l8192_id5_0_0_wdata),
    .ram_w4_l8192_id5_0_0_wenable(ram_w4_l8192_id5_0_0_wenable),
    .ram_w4_l8192_id5_0_1_addr(ram_w4_l8192_id5_0_1_addr),
    .ram_w4_l8192_id5_0_1_rdata(ram_w4_l8192_id5_0_1_rdata),
    .ram_w4_l8192_id5_0_1_wdata(ram_w4_l8192_id5_0_1_wdata),
    .ram_w4_l8192_id5_0_1_wenable(ram_w4_l8192_id5_0_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id5_1_0_addr;
  wire [4-1:0] ram_w4_l8192_id5_1_0_rdata;
  reg [4-1:0] ram_w4_l8192_id5_1_0_wdata;
  reg ram_w4_l8192_id5_1_0_wenable;
  reg [10-1:0] ram_w4_l8192_id5_1_1_addr;
  wire [4-1:0] ram_w4_l8192_id5_1_1_rdata;
  reg [4-1:0] ram_w4_l8192_id5_1_1_wdata;
  reg ram_w4_l8192_id5_1_1_wenable;

  ram_w4_l8192_id5_1
  inst_ram_w4_l8192_id5_1
  (
    .CLK(CLK),
    .ram_w4_l8192_id5_1_0_addr(ram_w4_l8192_id5_1_0_addr),
    .ram_w4_l8192_id5_1_0_rdata(ram_w4_l8192_id5_1_0_rdata),
    .ram_w4_l8192_id5_1_0_wdata(ram_w4_l8192_id5_1_0_wdata),
    .ram_w4_l8192_id5_1_0_wenable(ram_w4_l8192_id5_1_0_wenable),
    .ram_w4_l8192_id5_1_1_addr(ram_w4_l8192_id5_1_1_addr),
    .ram_w4_l8192_id5_1_1_rdata(ram_w4_l8192_id5_1_1_rdata),
    .ram_w4_l8192_id5_1_1_wdata(ram_w4_l8192_id5_1_1_wdata),
    .ram_w4_l8192_id5_1_1_wenable(ram_w4_l8192_id5_1_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id5_2_0_addr;
  wire [4-1:0] ram_w4_l8192_id5_2_0_rdata;
  reg [4-1:0] ram_w4_l8192_id5_2_0_wdata;
  reg ram_w4_l8192_id5_2_0_wenable;
  reg [10-1:0] ram_w4_l8192_id5_2_1_addr;
  wire [4-1:0] ram_w4_l8192_id5_2_1_rdata;
  reg [4-1:0] ram_w4_l8192_id5_2_1_wdata;
  reg ram_w4_l8192_id5_2_1_wenable;

  ram_w4_l8192_id5_2
  inst_ram_w4_l8192_id5_2
  (
    .CLK(CLK),
    .ram_w4_l8192_id5_2_0_addr(ram_w4_l8192_id5_2_0_addr),
    .ram_w4_l8192_id5_2_0_rdata(ram_w4_l8192_id5_2_0_rdata),
    .ram_w4_l8192_id5_2_0_wdata(ram_w4_l8192_id5_2_0_wdata),
    .ram_w4_l8192_id5_2_0_wenable(ram_w4_l8192_id5_2_0_wenable),
    .ram_w4_l8192_id5_2_1_addr(ram_w4_l8192_id5_2_1_addr),
    .ram_w4_l8192_id5_2_1_rdata(ram_w4_l8192_id5_2_1_rdata),
    .ram_w4_l8192_id5_2_1_wdata(ram_w4_l8192_id5_2_1_wdata),
    .ram_w4_l8192_id5_2_1_wenable(ram_w4_l8192_id5_2_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id5_3_0_addr;
  wire [4-1:0] ram_w4_l8192_id5_3_0_rdata;
  reg [4-1:0] ram_w4_l8192_id5_3_0_wdata;
  reg ram_w4_l8192_id5_3_0_wenable;
  reg [10-1:0] ram_w4_l8192_id5_3_1_addr;
  wire [4-1:0] ram_w4_l8192_id5_3_1_rdata;
  reg [4-1:0] ram_w4_l8192_id5_3_1_wdata;
  reg ram_w4_l8192_id5_3_1_wenable;

  ram_w4_l8192_id5_3
  inst_ram_w4_l8192_id5_3
  (
    .CLK(CLK),
    .ram_w4_l8192_id5_3_0_addr(ram_w4_l8192_id5_3_0_addr),
    .ram_w4_l8192_id5_3_0_rdata(ram_w4_l8192_id5_3_0_rdata),
    .ram_w4_l8192_id5_3_0_wdata(ram_w4_l8192_id5_3_0_wdata),
    .ram_w4_l8192_id5_3_0_wenable(ram_w4_l8192_id5_3_0_wenable),
    .ram_w4_l8192_id5_3_1_addr(ram_w4_l8192_id5_3_1_addr),
    .ram_w4_l8192_id5_3_1_rdata(ram_w4_l8192_id5_3_1_rdata),
    .ram_w4_l8192_id5_3_1_wdata(ram_w4_l8192_id5_3_1_wdata),
    .ram_w4_l8192_id5_3_1_wenable(ram_w4_l8192_id5_3_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id5_4_0_addr;
  wire [4-1:0] ram_w4_l8192_id5_4_0_rdata;
  reg [4-1:0] ram_w4_l8192_id5_4_0_wdata;
  reg ram_w4_l8192_id5_4_0_wenable;
  reg [10-1:0] ram_w4_l8192_id5_4_1_addr;
  wire [4-1:0] ram_w4_l8192_id5_4_1_rdata;
  reg [4-1:0] ram_w4_l8192_id5_4_1_wdata;
  reg ram_w4_l8192_id5_4_1_wenable;

  ram_w4_l8192_id5_4
  inst_ram_w4_l8192_id5_4
  (
    .CLK(CLK),
    .ram_w4_l8192_id5_4_0_addr(ram_w4_l8192_id5_4_0_addr),
    .ram_w4_l8192_id5_4_0_rdata(ram_w4_l8192_id5_4_0_rdata),
    .ram_w4_l8192_id5_4_0_wdata(ram_w4_l8192_id5_4_0_wdata),
    .ram_w4_l8192_id5_4_0_wenable(ram_w4_l8192_id5_4_0_wenable),
    .ram_w4_l8192_id5_4_1_addr(ram_w4_l8192_id5_4_1_addr),
    .ram_w4_l8192_id5_4_1_rdata(ram_w4_l8192_id5_4_1_rdata),
    .ram_w4_l8192_id5_4_1_wdata(ram_w4_l8192_id5_4_1_wdata),
    .ram_w4_l8192_id5_4_1_wenable(ram_w4_l8192_id5_4_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id5_5_0_addr;
  wire [4-1:0] ram_w4_l8192_id5_5_0_rdata;
  reg [4-1:0] ram_w4_l8192_id5_5_0_wdata;
  reg ram_w4_l8192_id5_5_0_wenable;
  reg [10-1:0] ram_w4_l8192_id5_5_1_addr;
  wire [4-1:0] ram_w4_l8192_id5_5_1_rdata;
  reg [4-1:0] ram_w4_l8192_id5_5_1_wdata;
  reg ram_w4_l8192_id5_5_1_wenable;

  ram_w4_l8192_id5_5
  inst_ram_w4_l8192_id5_5
  (
    .CLK(CLK),
    .ram_w4_l8192_id5_5_0_addr(ram_w4_l8192_id5_5_0_addr),
    .ram_w4_l8192_id5_5_0_rdata(ram_w4_l8192_id5_5_0_rdata),
    .ram_w4_l8192_id5_5_0_wdata(ram_w4_l8192_id5_5_0_wdata),
    .ram_w4_l8192_id5_5_0_wenable(ram_w4_l8192_id5_5_0_wenable),
    .ram_w4_l8192_id5_5_1_addr(ram_w4_l8192_id5_5_1_addr),
    .ram_w4_l8192_id5_5_1_rdata(ram_w4_l8192_id5_5_1_rdata),
    .ram_w4_l8192_id5_5_1_wdata(ram_w4_l8192_id5_5_1_wdata),
    .ram_w4_l8192_id5_5_1_wenable(ram_w4_l8192_id5_5_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id5_6_0_addr;
  wire [4-1:0] ram_w4_l8192_id5_6_0_rdata;
  reg [4-1:0] ram_w4_l8192_id5_6_0_wdata;
  reg ram_w4_l8192_id5_6_0_wenable;
  reg [10-1:0] ram_w4_l8192_id5_6_1_addr;
  wire [4-1:0] ram_w4_l8192_id5_6_1_rdata;
  reg [4-1:0] ram_w4_l8192_id5_6_1_wdata;
  reg ram_w4_l8192_id5_6_1_wenable;

  ram_w4_l8192_id5_6
  inst_ram_w4_l8192_id5_6
  (
    .CLK(CLK),
    .ram_w4_l8192_id5_6_0_addr(ram_w4_l8192_id5_6_0_addr),
    .ram_w4_l8192_id5_6_0_rdata(ram_w4_l8192_id5_6_0_rdata),
    .ram_w4_l8192_id5_6_0_wdata(ram_w4_l8192_id5_6_0_wdata),
    .ram_w4_l8192_id5_6_0_wenable(ram_w4_l8192_id5_6_0_wenable),
    .ram_w4_l8192_id5_6_1_addr(ram_w4_l8192_id5_6_1_addr),
    .ram_w4_l8192_id5_6_1_rdata(ram_w4_l8192_id5_6_1_rdata),
    .ram_w4_l8192_id5_6_1_wdata(ram_w4_l8192_id5_6_1_wdata),
    .ram_w4_l8192_id5_6_1_wenable(ram_w4_l8192_id5_6_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id5_7_0_addr;
  wire [4-1:0] ram_w4_l8192_id5_7_0_rdata;
  reg [4-1:0] ram_w4_l8192_id5_7_0_wdata;
  reg ram_w4_l8192_id5_7_0_wenable;
  reg [10-1:0] ram_w4_l8192_id5_7_1_addr;
  wire [4-1:0] ram_w4_l8192_id5_7_1_rdata;
  reg [4-1:0] ram_w4_l8192_id5_7_1_wdata;
  reg ram_w4_l8192_id5_7_1_wenable;

  ram_w4_l8192_id5_7
  inst_ram_w4_l8192_id5_7
  (
    .CLK(CLK),
    .ram_w4_l8192_id5_7_0_addr(ram_w4_l8192_id5_7_0_addr),
    .ram_w4_l8192_id5_7_0_rdata(ram_w4_l8192_id5_7_0_rdata),
    .ram_w4_l8192_id5_7_0_wdata(ram_w4_l8192_id5_7_0_wdata),
    .ram_w4_l8192_id5_7_0_wenable(ram_w4_l8192_id5_7_0_wenable),
    .ram_w4_l8192_id5_7_1_addr(ram_w4_l8192_id5_7_1_addr),
    .ram_w4_l8192_id5_7_1_rdata(ram_w4_l8192_id5_7_1_rdata),
    .ram_w4_l8192_id5_7_1_wdata(ram_w4_l8192_id5_7_1_wdata),
    .ram_w4_l8192_id5_7_1_wenable(ram_w4_l8192_id5_7_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id6_0_0_addr;
  wire [4-1:0] ram_w4_l8192_id6_0_0_rdata;
  reg [4-1:0] ram_w4_l8192_id6_0_0_wdata;
  reg ram_w4_l8192_id6_0_0_wenable;
  reg [10-1:0] ram_w4_l8192_id6_0_1_addr;
  wire [4-1:0] ram_w4_l8192_id6_0_1_rdata;
  reg [4-1:0] ram_w4_l8192_id6_0_1_wdata;
  reg ram_w4_l8192_id6_0_1_wenable;

  ram_w4_l8192_id6_0
  inst_ram_w4_l8192_id6_0
  (
    .CLK(CLK),
    .ram_w4_l8192_id6_0_0_addr(ram_w4_l8192_id6_0_0_addr),
    .ram_w4_l8192_id6_0_0_rdata(ram_w4_l8192_id6_0_0_rdata),
    .ram_w4_l8192_id6_0_0_wdata(ram_w4_l8192_id6_0_0_wdata),
    .ram_w4_l8192_id6_0_0_wenable(ram_w4_l8192_id6_0_0_wenable),
    .ram_w4_l8192_id6_0_1_addr(ram_w4_l8192_id6_0_1_addr),
    .ram_w4_l8192_id6_0_1_rdata(ram_w4_l8192_id6_0_1_rdata),
    .ram_w4_l8192_id6_0_1_wdata(ram_w4_l8192_id6_0_1_wdata),
    .ram_w4_l8192_id6_0_1_wenable(ram_w4_l8192_id6_0_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id6_1_0_addr;
  wire [4-1:0] ram_w4_l8192_id6_1_0_rdata;
  reg [4-1:0] ram_w4_l8192_id6_1_0_wdata;
  reg ram_w4_l8192_id6_1_0_wenable;
  reg [10-1:0] ram_w4_l8192_id6_1_1_addr;
  wire [4-1:0] ram_w4_l8192_id6_1_1_rdata;
  reg [4-1:0] ram_w4_l8192_id6_1_1_wdata;
  reg ram_w4_l8192_id6_1_1_wenable;

  ram_w4_l8192_id6_1
  inst_ram_w4_l8192_id6_1
  (
    .CLK(CLK),
    .ram_w4_l8192_id6_1_0_addr(ram_w4_l8192_id6_1_0_addr),
    .ram_w4_l8192_id6_1_0_rdata(ram_w4_l8192_id6_1_0_rdata),
    .ram_w4_l8192_id6_1_0_wdata(ram_w4_l8192_id6_1_0_wdata),
    .ram_w4_l8192_id6_1_0_wenable(ram_w4_l8192_id6_1_0_wenable),
    .ram_w4_l8192_id6_1_1_addr(ram_w4_l8192_id6_1_1_addr),
    .ram_w4_l8192_id6_1_1_rdata(ram_w4_l8192_id6_1_1_rdata),
    .ram_w4_l8192_id6_1_1_wdata(ram_w4_l8192_id6_1_1_wdata),
    .ram_w4_l8192_id6_1_1_wenable(ram_w4_l8192_id6_1_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id6_2_0_addr;
  wire [4-1:0] ram_w4_l8192_id6_2_0_rdata;
  reg [4-1:0] ram_w4_l8192_id6_2_0_wdata;
  reg ram_w4_l8192_id6_2_0_wenable;
  reg [10-1:0] ram_w4_l8192_id6_2_1_addr;
  wire [4-1:0] ram_w4_l8192_id6_2_1_rdata;
  reg [4-1:0] ram_w4_l8192_id6_2_1_wdata;
  reg ram_w4_l8192_id6_2_1_wenable;

  ram_w4_l8192_id6_2
  inst_ram_w4_l8192_id6_2
  (
    .CLK(CLK),
    .ram_w4_l8192_id6_2_0_addr(ram_w4_l8192_id6_2_0_addr),
    .ram_w4_l8192_id6_2_0_rdata(ram_w4_l8192_id6_2_0_rdata),
    .ram_w4_l8192_id6_2_0_wdata(ram_w4_l8192_id6_2_0_wdata),
    .ram_w4_l8192_id6_2_0_wenable(ram_w4_l8192_id6_2_0_wenable),
    .ram_w4_l8192_id6_2_1_addr(ram_w4_l8192_id6_2_1_addr),
    .ram_w4_l8192_id6_2_1_rdata(ram_w4_l8192_id6_2_1_rdata),
    .ram_w4_l8192_id6_2_1_wdata(ram_w4_l8192_id6_2_1_wdata),
    .ram_w4_l8192_id6_2_1_wenable(ram_w4_l8192_id6_2_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id6_3_0_addr;
  wire [4-1:0] ram_w4_l8192_id6_3_0_rdata;
  reg [4-1:0] ram_w4_l8192_id6_3_0_wdata;
  reg ram_w4_l8192_id6_3_0_wenable;
  reg [10-1:0] ram_w4_l8192_id6_3_1_addr;
  wire [4-1:0] ram_w4_l8192_id6_3_1_rdata;
  reg [4-1:0] ram_w4_l8192_id6_3_1_wdata;
  reg ram_w4_l8192_id6_3_1_wenable;

  ram_w4_l8192_id6_3
  inst_ram_w4_l8192_id6_3
  (
    .CLK(CLK),
    .ram_w4_l8192_id6_3_0_addr(ram_w4_l8192_id6_3_0_addr),
    .ram_w4_l8192_id6_3_0_rdata(ram_w4_l8192_id6_3_0_rdata),
    .ram_w4_l8192_id6_3_0_wdata(ram_w4_l8192_id6_3_0_wdata),
    .ram_w4_l8192_id6_3_0_wenable(ram_w4_l8192_id6_3_0_wenable),
    .ram_w4_l8192_id6_3_1_addr(ram_w4_l8192_id6_3_1_addr),
    .ram_w4_l8192_id6_3_1_rdata(ram_w4_l8192_id6_3_1_rdata),
    .ram_w4_l8192_id6_3_1_wdata(ram_w4_l8192_id6_3_1_wdata),
    .ram_w4_l8192_id6_3_1_wenable(ram_w4_l8192_id6_3_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id6_4_0_addr;
  wire [4-1:0] ram_w4_l8192_id6_4_0_rdata;
  reg [4-1:0] ram_w4_l8192_id6_4_0_wdata;
  reg ram_w4_l8192_id6_4_0_wenable;
  reg [10-1:0] ram_w4_l8192_id6_4_1_addr;
  wire [4-1:0] ram_w4_l8192_id6_4_1_rdata;
  reg [4-1:0] ram_w4_l8192_id6_4_1_wdata;
  reg ram_w4_l8192_id6_4_1_wenable;

  ram_w4_l8192_id6_4
  inst_ram_w4_l8192_id6_4
  (
    .CLK(CLK),
    .ram_w4_l8192_id6_4_0_addr(ram_w4_l8192_id6_4_0_addr),
    .ram_w4_l8192_id6_4_0_rdata(ram_w4_l8192_id6_4_0_rdata),
    .ram_w4_l8192_id6_4_0_wdata(ram_w4_l8192_id6_4_0_wdata),
    .ram_w4_l8192_id6_4_0_wenable(ram_w4_l8192_id6_4_0_wenable),
    .ram_w4_l8192_id6_4_1_addr(ram_w4_l8192_id6_4_1_addr),
    .ram_w4_l8192_id6_4_1_rdata(ram_w4_l8192_id6_4_1_rdata),
    .ram_w4_l8192_id6_4_1_wdata(ram_w4_l8192_id6_4_1_wdata),
    .ram_w4_l8192_id6_4_1_wenable(ram_w4_l8192_id6_4_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id6_5_0_addr;
  wire [4-1:0] ram_w4_l8192_id6_5_0_rdata;
  reg [4-1:0] ram_w4_l8192_id6_5_0_wdata;
  reg ram_w4_l8192_id6_5_0_wenable;
  reg [10-1:0] ram_w4_l8192_id6_5_1_addr;
  wire [4-1:0] ram_w4_l8192_id6_5_1_rdata;
  reg [4-1:0] ram_w4_l8192_id6_5_1_wdata;
  reg ram_w4_l8192_id6_5_1_wenable;

  ram_w4_l8192_id6_5
  inst_ram_w4_l8192_id6_5
  (
    .CLK(CLK),
    .ram_w4_l8192_id6_5_0_addr(ram_w4_l8192_id6_5_0_addr),
    .ram_w4_l8192_id6_5_0_rdata(ram_w4_l8192_id6_5_0_rdata),
    .ram_w4_l8192_id6_5_0_wdata(ram_w4_l8192_id6_5_0_wdata),
    .ram_w4_l8192_id6_5_0_wenable(ram_w4_l8192_id6_5_0_wenable),
    .ram_w4_l8192_id6_5_1_addr(ram_w4_l8192_id6_5_1_addr),
    .ram_w4_l8192_id6_5_1_rdata(ram_w4_l8192_id6_5_1_rdata),
    .ram_w4_l8192_id6_5_1_wdata(ram_w4_l8192_id6_5_1_wdata),
    .ram_w4_l8192_id6_5_1_wenable(ram_w4_l8192_id6_5_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id6_6_0_addr;
  wire [4-1:0] ram_w4_l8192_id6_6_0_rdata;
  reg [4-1:0] ram_w4_l8192_id6_6_0_wdata;
  reg ram_w4_l8192_id6_6_0_wenable;
  reg [10-1:0] ram_w4_l8192_id6_6_1_addr;
  wire [4-1:0] ram_w4_l8192_id6_6_1_rdata;
  reg [4-1:0] ram_w4_l8192_id6_6_1_wdata;
  reg ram_w4_l8192_id6_6_1_wenable;

  ram_w4_l8192_id6_6
  inst_ram_w4_l8192_id6_6
  (
    .CLK(CLK),
    .ram_w4_l8192_id6_6_0_addr(ram_w4_l8192_id6_6_0_addr),
    .ram_w4_l8192_id6_6_0_rdata(ram_w4_l8192_id6_6_0_rdata),
    .ram_w4_l8192_id6_6_0_wdata(ram_w4_l8192_id6_6_0_wdata),
    .ram_w4_l8192_id6_6_0_wenable(ram_w4_l8192_id6_6_0_wenable),
    .ram_w4_l8192_id6_6_1_addr(ram_w4_l8192_id6_6_1_addr),
    .ram_w4_l8192_id6_6_1_rdata(ram_w4_l8192_id6_6_1_rdata),
    .ram_w4_l8192_id6_6_1_wdata(ram_w4_l8192_id6_6_1_wdata),
    .ram_w4_l8192_id6_6_1_wenable(ram_w4_l8192_id6_6_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id6_7_0_addr;
  wire [4-1:0] ram_w4_l8192_id6_7_0_rdata;
  reg [4-1:0] ram_w4_l8192_id6_7_0_wdata;
  reg ram_w4_l8192_id6_7_0_wenable;
  reg [10-1:0] ram_w4_l8192_id6_7_1_addr;
  wire [4-1:0] ram_w4_l8192_id6_7_1_rdata;
  reg [4-1:0] ram_w4_l8192_id6_7_1_wdata;
  reg ram_w4_l8192_id6_7_1_wenable;

  ram_w4_l8192_id6_7
  inst_ram_w4_l8192_id6_7
  (
    .CLK(CLK),
    .ram_w4_l8192_id6_7_0_addr(ram_w4_l8192_id6_7_0_addr),
    .ram_w4_l8192_id6_7_0_rdata(ram_w4_l8192_id6_7_0_rdata),
    .ram_w4_l8192_id6_7_0_wdata(ram_w4_l8192_id6_7_0_wdata),
    .ram_w4_l8192_id6_7_0_wenable(ram_w4_l8192_id6_7_0_wenable),
    .ram_w4_l8192_id6_7_1_addr(ram_w4_l8192_id6_7_1_addr),
    .ram_w4_l8192_id6_7_1_rdata(ram_w4_l8192_id6_7_1_rdata),
    .ram_w4_l8192_id6_7_1_wdata(ram_w4_l8192_id6_7_1_wdata),
    .ram_w4_l8192_id6_7_1_wenable(ram_w4_l8192_id6_7_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id7_0_0_addr;
  wire [4-1:0] ram_w4_l8192_id7_0_0_rdata;
  reg [4-1:0] ram_w4_l8192_id7_0_0_wdata;
  reg ram_w4_l8192_id7_0_0_wenable;
  reg [10-1:0] ram_w4_l8192_id7_0_1_addr;
  wire [4-1:0] ram_w4_l8192_id7_0_1_rdata;
  reg [4-1:0] ram_w4_l8192_id7_0_1_wdata;
  reg ram_w4_l8192_id7_0_1_wenable;

  ram_w4_l8192_id7_0
  inst_ram_w4_l8192_id7_0
  (
    .CLK(CLK),
    .ram_w4_l8192_id7_0_0_addr(ram_w4_l8192_id7_0_0_addr),
    .ram_w4_l8192_id7_0_0_rdata(ram_w4_l8192_id7_0_0_rdata),
    .ram_w4_l8192_id7_0_0_wdata(ram_w4_l8192_id7_0_0_wdata),
    .ram_w4_l8192_id7_0_0_wenable(ram_w4_l8192_id7_0_0_wenable),
    .ram_w4_l8192_id7_0_1_addr(ram_w4_l8192_id7_0_1_addr),
    .ram_w4_l8192_id7_0_1_rdata(ram_w4_l8192_id7_0_1_rdata),
    .ram_w4_l8192_id7_0_1_wdata(ram_w4_l8192_id7_0_1_wdata),
    .ram_w4_l8192_id7_0_1_wenable(ram_w4_l8192_id7_0_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id7_1_0_addr;
  wire [4-1:0] ram_w4_l8192_id7_1_0_rdata;
  reg [4-1:0] ram_w4_l8192_id7_1_0_wdata;
  reg ram_w4_l8192_id7_1_0_wenable;
  reg [10-1:0] ram_w4_l8192_id7_1_1_addr;
  wire [4-1:0] ram_w4_l8192_id7_1_1_rdata;
  reg [4-1:0] ram_w4_l8192_id7_1_1_wdata;
  reg ram_w4_l8192_id7_1_1_wenable;

  ram_w4_l8192_id7_1
  inst_ram_w4_l8192_id7_1
  (
    .CLK(CLK),
    .ram_w4_l8192_id7_1_0_addr(ram_w4_l8192_id7_1_0_addr),
    .ram_w4_l8192_id7_1_0_rdata(ram_w4_l8192_id7_1_0_rdata),
    .ram_w4_l8192_id7_1_0_wdata(ram_w4_l8192_id7_1_0_wdata),
    .ram_w4_l8192_id7_1_0_wenable(ram_w4_l8192_id7_1_0_wenable),
    .ram_w4_l8192_id7_1_1_addr(ram_w4_l8192_id7_1_1_addr),
    .ram_w4_l8192_id7_1_1_rdata(ram_w4_l8192_id7_1_1_rdata),
    .ram_w4_l8192_id7_1_1_wdata(ram_w4_l8192_id7_1_1_wdata),
    .ram_w4_l8192_id7_1_1_wenable(ram_w4_l8192_id7_1_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id7_2_0_addr;
  wire [4-1:0] ram_w4_l8192_id7_2_0_rdata;
  reg [4-1:0] ram_w4_l8192_id7_2_0_wdata;
  reg ram_w4_l8192_id7_2_0_wenable;
  reg [10-1:0] ram_w4_l8192_id7_2_1_addr;
  wire [4-1:0] ram_w4_l8192_id7_2_1_rdata;
  reg [4-1:0] ram_w4_l8192_id7_2_1_wdata;
  reg ram_w4_l8192_id7_2_1_wenable;

  ram_w4_l8192_id7_2
  inst_ram_w4_l8192_id7_2
  (
    .CLK(CLK),
    .ram_w4_l8192_id7_2_0_addr(ram_w4_l8192_id7_2_0_addr),
    .ram_w4_l8192_id7_2_0_rdata(ram_w4_l8192_id7_2_0_rdata),
    .ram_w4_l8192_id7_2_0_wdata(ram_w4_l8192_id7_2_0_wdata),
    .ram_w4_l8192_id7_2_0_wenable(ram_w4_l8192_id7_2_0_wenable),
    .ram_w4_l8192_id7_2_1_addr(ram_w4_l8192_id7_2_1_addr),
    .ram_w4_l8192_id7_2_1_rdata(ram_w4_l8192_id7_2_1_rdata),
    .ram_w4_l8192_id7_2_1_wdata(ram_w4_l8192_id7_2_1_wdata),
    .ram_w4_l8192_id7_2_1_wenable(ram_w4_l8192_id7_2_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id7_3_0_addr;
  wire [4-1:0] ram_w4_l8192_id7_3_0_rdata;
  reg [4-1:0] ram_w4_l8192_id7_3_0_wdata;
  reg ram_w4_l8192_id7_3_0_wenable;
  reg [10-1:0] ram_w4_l8192_id7_3_1_addr;
  wire [4-1:0] ram_w4_l8192_id7_3_1_rdata;
  reg [4-1:0] ram_w4_l8192_id7_3_1_wdata;
  reg ram_w4_l8192_id7_3_1_wenable;

  ram_w4_l8192_id7_3
  inst_ram_w4_l8192_id7_3
  (
    .CLK(CLK),
    .ram_w4_l8192_id7_3_0_addr(ram_w4_l8192_id7_3_0_addr),
    .ram_w4_l8192_id7_3_0_rdata(ram_w4_l8192_id7_3_0_rdata),
    .ram_w4_l8192_id7_3_0_wdata(ram_w4_l8192_id7_3_0_wdata),
    .ram_w4_l8192_id7_3_0_wenable(ram_w4_l8192_id7_3_0_wenable),
    .ram_w4_l8192_id7_3_1_addr(ram_w4_l8192_id7_3_1_addr),
    .ram_w4_l8192_id7_3_1_rdata(ram_w4_l8192_id7_3_1_rdata),
    .ram_w4_l8192_id7_3_1_wdata(ram_w4_l8192_id7_3_1_wdata),
    .ram_w4_l8192_id7_3_1_wenable(ram_w4_l8192_id7_3_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id7_4_0_addr;
  wire [4-1:0] ram_w4_l8192_id7_4_0_rdata;
  reg [4-1:0] ram_w4_l8192_id7_4_0_wdata;
  reg ram_w4_l8192_id7_4_0_wenable;
  reg [10-1:0] ram_w4_l8192_id7_4_1_addr;
  wire [4-1:0] ram_w4_l8192_id7_4_1_rdata;
  reg [4-1:0] ram_w4_l8192_id7_4_1_wdata;
  reg ram_w4_l8192_id7_4_1_wenable;

  ram_w4_l8192_id7_4
  inst_ram_w4_l8192_id7_4
  (
    .CLK(CLK),
    .ram_w4_l8192_id7_4_0_addr(ram_w4_l8192_id7_4_0_addr),
    .ram_w4_l8192_id7_4_0_rdata(ram_w4_l8192_id7_4_0_rdata),
    .ram_w4_l8192_id7_4_0_wdata(ram_w4_l8192_id7_4_0_wdata),
    .ram_w4_l8192_id7_4_0_wenable(ram_w4_l8192_id7_4_0_wenable),
    .ram_w4_l8192_id7_4_1_addr(ram_w4_l8192_id7_4_1_addr),
    .ram_w4_l8192_id7_4_1_rdata(ram_w4_l8192_id7_4_1_rdata),
    .ram_w4_l8192_id7_4_1_wdata(ram_w4_l8192_id7_4_1_wdata),
    .ram_w4_l8192_id7_4_1_wenable(ram_w4_l8192_id7_4_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id7_5_0_addr;
  wire [4-1:0] ram_w4_l8192_id7_5_0_rdata;
  reg [4-1:0] ram_w4_l8192_id7_5_0_wdata;
  reg ram_w4_l8192_id7_5_0_wenable;
  reg [10-1:0] ram_w4_l8192_id7_5_1_addr;
  wire [4-1:0] ram_w4_l8192_id7_5_1_rdata;
  reg [4-1:0] ram_w4_l8192_id7_5_1_wdata;
  reg ram_w4_l8192_id7_5_1_wenable;

  ram_w4_l8192_id7_5
  inst_ram_w4_l8192_id7_5
  (
    .CLK(CLK),
    .ram_w4_l8192_id7_5_0_addr(ram_w4_l8192_id7_5_0_addr),
    .ram_w4_l8192_id7_5_0_rdata(ram_w4_l8192_id7_5_0_rdata),
    .ram_w4_l8192_id7_5_0_wdata(ram_w4_l8192_id7_5_0_wdata),
    .ram_w4_l8192_id7_5_0_wenable(ram_w4_l8192_id7_5_0_wenable),
    .ram_w4_l8192_id7_5_1_addr(ram_w4_l8192_id7_5_1_addr),
    .ram_w4_l8192_id7_5_1_rdata(ram_w4_l8192_id7_5_1_rdata),
    .ram_w4_l8192_id7_5_1_wdata(ram_w4_l8192_id7_5_1_wdata),
    .ram_w4_l8192_id7_5_1_wenable(ram_w4_l8192_id7_5_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id7_6_0_addr;
  wire [4-1:0] ram_w4_l8192_id7_6_0_rdata;
  reg [4-1:0] ram_w4_l8192_id7_6_0_wdata;
  reg ram_w4_l8192_id7_6_0_wenable;
  reg [10-1:0] ram_w4_l8192_id7_6_1_addr;
  wire [4-1:0] ram_w4_l8192_id7_6_1_rdata;
  reg [4-1:0] ram_w4_l8192_id7_6_1_wdata;
  reg ram_w4_l8192_id7_6_1_wenable;

  ram_w4_l8192_id7_6
  inst_ram_w4_l8192_id7_6
  (
    .CLK(CLK),
    .ram_w4_l8192_id7_6_0_addr(ram_w4_l8192_id7_6_0_addr),
    .ram_w4_l8192_id7_6_0_rdata(ram_w4_l8192_id7_6_0_rdata),
    .ram_w4_l8192_id7_6_0_wdata(ram_w4_l8192_id7_6_0_wdata),
    .ram_w4_l8192_id7_6_0_wenable(ram_w4_l8192_id7_6_0_wenable),
    .ram_w4_l8192_id7_6_1_addr(ram_w4_l8192_id7_6_1_addr),
    .ram_w4_l8192_id7_6_1_rdata(ram_w4_l8192_id7_6_1_rdata),
    .ram_w4_l8192_id7_6_1_wdata(ram_w4_l8192_id7_6_1_wdata),
    .ram_w4_l8192_id7_6_1_wenable(ram_w4_l8192_id7_6_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id7_7_0_addr;
  wire [4-1:0] ram_w4_l8192_id7_7_0_rdata;
  reg [4-1:0] ram_w4_l8192_id7_7_0_wdata;
  reg ram_w4_l8192_id7_7_0_wenable;
  reg [10-1:0] ram_w4_l8192_id7_7_1_addr;
  wire [4-1:0] ram_w4_l8192_id7_7_1_rdata;
  reg [4-1:0] ram_w4_l8192_id7_7_1_wdata;
  reg ram_w4_l8192_id7_7_1_wenable;

  ram_w4_l8192_id7_7
  inst_ram_w4_l8192_id7_7
  (
    .CLK(CLK),
    .ram_w4_l8192_id7_7_0_addr(ram_w4_l8192_id7_7_0_addr),
    .ram_w4_l8192_id7_7_0_rdata(ram_w4_l8192_id7_7_0_rdata),
    .ram_w4_l8192_id7_7_0_wdata(ram_w4_l8192_id7_7_0_wdata),
    .ram_w4_l8192_id7_7_0_wenable(ram_w4_l8192_id7_7_0_wenable),
    .ram_w4_l8192_id7_7_1_addr(ram_w4_l8192_id7_7_1_addr),
    .ram_w4_l8192_id7_7_1_rdata(ram_w4_l8192_id7_7_1_rdata),
    .ram_w4_l8192_id7_7_1_wdata(ram_w4_l8192_id7_7_1_wdata),
    .ram_w4_l8192_id7_7_1_wenable(ram_w4_l8192_id7_7_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id8_0_0_addr;
  wire [4-1:0] ram_w4_l8192_id8_0_0_rdata;
  reg [4-1:0] ram_w4_l8192_id8_0_0_wdata;
  reg ram_w4_l8192_id8_0_0_wenable;
  reg [10-1:0] ram_w4_l8192_id8_0_1_addr;
  wire [4-1:0] ram_w4_l8192_id8_0_1_rdata;
  reg [4-1:0] ram_w4_l8192_id8_0_1_wdata;
  reg ram_w4_l8192_id8_0_1_wenable;

  ram_w4_l8192_id8_0
  inst_ram_w4_l8192_id8_0
  (
    .CLK(CLK),
    .ram_w4_l8192_id8_0_0_addr(ram_w4_l8192_id8_0_0_addr),
    .ram_w4_l8192_id8_0_0_rdata(ram_w4_l8192_id8_0_0_rdata),
    .ram_w4_l8192_id8_0_0_wdata(ram_w4_l8192_id8_0_0_wdata),
    .ram_w4_l8192_id8_0_0_wenable(ram_w4_l8192_id8_0_0_wenable),
    .ram_w4_l8192_id8_0_1_addr(ram_w4_l8192_id8_0_1_addr),
    .ram_w4_l8192_id8_0_1_rdata(ram_w4_l8192_id8_0_1_rdata),
    .ram_w4_l8192_id8_0_1_wdata(ram_w4_l8192_id8_0_1_wdata),
    .ram_w4_l8192_id8_0_1_wenable(ram_w4_l8192_id8_0_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id8_1_0_addr;
  wire [4-1:0] ram_w4_l8192_id8_1_0_rdata;
  reg [4-1:0] ram_w4_l8192_id8_1_0_wdata;
  reg ram_w4_l8192_id8_1_0_wenable;
  reg [10-1:0] ram_w4_l8192_id8_1_1_addr;
  wire [4-1:0] ram_w4_l8192_id8_1_1_rdata;
  reg [4-1:0] ram_w4_l8192_id8_1_1_wdata;
  reg ram_w4_l8192_id8_1_1_wenable;

  ram_w4_l8192_id8_1
  inst_ram_w4_l8192_id8_1
  (
    .CLK(CLK),
    .ram_w4_l8192_id8_1_0_addr(ram_w4_l8192_id8_1_0_addr),
    .ram_w4_l8192_id8_1_0_rdata(ram_w4_l8192_id8_1_0_rdata),
    .ram_w4_l8192_id8_1_0_wdata(ram_w4_l8192_id8_1_0_wdata),
    .ram_w4_l8192_id8_1_0_wenable(ram_w4_l8192_id8_1_0_wenable),
    .ram_w4_l8192_id8_1_1_addr(ram_w4_l8192_id8_1_1_addr),
    .ram_w4_l8192_id8_1_1_rdata(ram_w4_l8192_id8_1_1_rdata),
    .ram_w4_l8192_id8_1_1_wdata(ram_w4_l8192_id8_1_1_wdata),
    .ram_w4_l8192_id8_1_1_wenable(ram_w4_l8192_id8_1_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id8_2_0_addr;
  wire [4-1:0] ram_w4_l8192_id8_2_0_rdata;
  reg [4-1:0] ram_w4_l8192_id8_2_0_wdata;
  reg ram_w4_l8192_id8_2_0_wenable;
  reg [10-1:0] ram_w4_l8192_id8_2_1_addr;
  wire [4-1:0] ram_w4_l8192_id8_2_1_rdata;
  reg [4-1:0] ram_w4_l8192_id8_2_1_wdata;
  reg ram_w4_l8192_id8_2_1_wenable;

  ram_w4_l8192_id8_2
  inst_ram_w4_l8192_id8_2
  (
    .CLK(CLK),
    .ram_w4_l8192_id8_2_0_addr(ram_w4_l8192_id8_2_0_addr),
    .ram_w4_l8192_id8_2_0_rdata(ram_w4_l8192_id8_2_0_rdata),
    .ram_w4_l8192_id8_2_0_wdata(ram_w4_l8192_id8_2_0_wdata),
    .ram_w4_l8192_id8_2_0_wenable(ram_w4_l8192_id8_2_0_wenable),
    .ram_w4_l8192_id8_2_1_addr(ram_w4_l8192_id8_2_1_addr),
    .ram_w4_l8192_id8_2_1_rdata(ram_w4_l8192_id8_2_1_rdata),
    .ram_w4_l8192_id8_2_1_wdata(ram_w4_l8192_id8_2_1_wdata),
    .ram_w4_l8192_id8_2_1_wenable(ram_w4_l8192_id8_2_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id8_3_0_addr;
  wire [4-1:0] ram_w4_l8192_id8_3_0_rdata;
  reg [4-1:0] ram_w4_l8192_id8_3_0_wdata;
  reg ram_w4_l8192_id8_3_0_wenable;
  reg [10-1:0] ram_w4_l8192_id8_3_1_addr;
  wire [4-1:0] ram_w4_l8192_id8_3_1_rdata;
  reg [4-1:0] ram_w4_l8192_id8_3_1_wdata;
  reg ram_w4_l8192_id8_3_1_wenable;

  ram_w4_l8192_id8_3
  inst_ram_w4_l8192_id8_3
  (
    .CLK(CLK),
    .ram_w4_l8192_id8_3_0_addr(ram_w4_l8192_id8_3_0_addr),
    .ram_w4_l8192_id8_3_0_rdata(ram_w4_l8192_id8_3_0_rdata),
    .ram_w4_l8192_id8_3_0_wdata(ram_w4_l8192_id8_3_0_wdata),
    .ram_w4_l8192_id8_3_0_wenable(ram_w4_l8192_id8_3_0_wenable),
    .ram_w4_l8192_id8_3_1_addr(ram_w4_l8192_id8_3_1_addr),
    .ram_w4_l8192_id8_3_1_rdata(ram_w4_l8192_id8_3_1_rdata),
    .ram_w4_l8192_id8_3_1_wdata(ram_w4_l8192_id8_3_1_wdata),
    .ram_w4_l8192_id8_3_1_wenable(ram_w4_l8192_id8_3_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id8_4_0_addr;
  wire [4-1:0] ram_w4_l8192_id8_4_0_rdata;
  reg [4-1:0] ram_w4_l8192_id8_4_0_wdata;
  reg ram_w4_l8192_id8_4_0_wenable;
  reg [10-1:0] ram_w4_l8192_id8_4_1_addr;
  wire [4-1:0] ram_w4_l8192_id8_4_1_rdata;
  reg [4-1:0] ram_w4_l8192_id8_4_1_wdata;
  reg ram_w4_l8192_id8_4_1_wenable;

  ram_w4_l8192_id8_4
  inst_ram_w4_l8192_id8_4
  (
    .CLK(CLK),
    .ram_w4_l8192_id8_4_0_addr(ram_w4_l8192_id8_4_0_addr),
    .ram_w4_l8192_id8_4_0_rdata(ram_w4_l8192_id8_4_0_rdata),
    .ram_w4_l8192_id8_4_0_wdata(ram_w4_l8192_id8_4_0_wdata),
    .ram_w4_l8192_id8_4_0_wenable(ram_w4_l8192_id8_4_0_wenable),
    .ram_w4_l8192_id8_4_1_addr(ram_w4_l8192_id8_4_1_addr),
    .ram_w4_l8192_id8_4_1_rdata(ram_w4_l8192_id8_4_1_rdata),
    .ram_w4_l8192_id8_4_1_wdata(ram_w4_l8192_id8_4_1_wdata),
    .ram_w4_l8192_id8_4_1_wenable(ram_w4_l8192_id8_4_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id8_5_0_addr;
  wire [4-1:0] ram_w4_l8192_id8_5_0_rdata;
  reg [4-1:0] ram_w4_l8192_id8_5_0_wdata;
  reg ram_w4_l8192_id8_5_0_wenable;
  reg [10-1:0] ram_w4_l8192_id8_5_1_addr;
  wire [4-1:0] ram_w4_l8192_id8_5_1_rdata;
  reg [4-1:0] ram_w4_l8192_id8_5_1_wdata;
  reg ram_w4_l8192_id8_5_1_wenable;

  ram_w4_l8192_id8_5
  inst_ram_w4_l8192_id8_5
  (
    .CLK(CLK),
    .ram_w4_l8192_id8_5_0_addr(ram_w4_l8192_id8_5_0_addr),
    .ram_w4_l8192_id8_5_0_rdata(ram_w4_l8192_id8_5_0_rdata),
    .ram_w4_l8192_id8_5_0_wdata(ram_w4_l8192_id8_5_0_wdata),
    .ram_w4_l8192_id8_5_0_wenable(ram_w4_l8192_id8_5_0_wenable),
    .ram_w4_l8192_id8_5_1_addr(ram_w4_l8192_id8_5_1_addr),
    .ram_w4_l8192_id8_5_1_rdata(ram_w4_l8192_id8_5_1_rdata),
    .ram_w4_l8192_id8_5_1_wdata(ram_w4_l8192_id8_5_1_wdata),
    .ram_w4_l8192_id8_5_1_wenable(ram_w4_l8192_id8_5_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id8_6_0_addr;
  wire [4-1:0] ram_w4_l8192_id8_6_0_rdata;
  reg [4-1:0] ram_w4_l8192_id8_6_0_wdata;
  reg ram_w4_l8192_id8_6_0_wenable;
  reg [10-1:0] ram_w4_l8192_id8_6_1_addr;
  wire [4-1:0] ram_w4_l8192_id8_6_1_rdata;
  reg [4-1:0] ram_w4_l8192_id8_6_1_wdata;
  reg ram_w4_l8192_id8_6_1_wenable;

  ram_w4_l8192_id8_6
  inst_ram_w4_l8192_id8_6
  (
    .CLK(CLK),
    .ram_w4_l8192_id8_6_0_addr(ram_w4_l8192_id8_6_0_addr),
    .ram_w4_l8192_id8_6_0_rdata(ram_w4_l8192_id8_6_0_rdata),
    .ram_w4_l8192_id8_6_0_wdata(ram_w4_l8192_id8_6_0_wdata),
    .ram_w4_l8192_id8_6_0_wenable(ram_w4_l8192_id8_6_0_wenable),
    .ram_w4_l8192_id8_6_1_addr(ram_w4_l8192_id8_6_1_addr),
    .ram_w4_l8192_id8_6_1_rdata(ram_w4_l8192_id8_6_1_rdata),
    .ram_w4_l8192_id8_6_1_wdata(ram_w4_l8192_id8_6_1_wdata),
    .ram_w4_l8192_id8_6_1_wenable(ram_w4_l8192_id8_6_1_wenable)
  );

  reg [10-1:0] ram_w4_l8192_id8_7_0_addr;
  wire [4-1:0] ram_w4_l8192_id8_7_0_rdata;
  reg [4-1:0] ram_w4_l8192_id8_7_0_wdata;
  reg ram_w4_l8192_id8_7_0_wenable;
  reg [10-1:0] ram_w4_l8192_id8_7_1_addr;
  wire [4-1:0] ram_w4_l8192_id8_7_1_rdata;
  reg [4-1:0] ram_w4_l8192_id8_7_1_wdata;
  reg ram_w4_l8192_id8_7_1_wenable;

  ram_w4_l8192_id8_7
  inst_ram_w4_l8192_id8_7
  (
    .CLK(CLK),
    .ram_w4_l8192_id8_7_0_addr(ram_w4_l8192_id8_7_0_addr),
    .ram_w4_l8192_id8_7_0_rdata(ram_w4_l8192_id8_7_0_rdata),
    .ram_w4_l8192_id8_7_0_wdata(ram_w4_l8192_id8_7_0_wdata),
    .ram_w4_l8192_id8_7_0_wenable(ram_w4_l8192_id8_7_0_wenable),
    .ram_w4_l8192_id8_7_1_addr(ram_w4_l8192_id8_7_1_addr),
    .ram_w4_l8192_id8_7_1_rdata(ram_w4_l8192_id8_7_1_rdata),
    .ram_w4_l8192_id8_7_1_wdata(ram_w4_l8192_id8_7_1_wdata),
    .ram_w4_l8192_id8_7_1_wenable(ram_w4_l8192_id8_7_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id0_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id0_0_0_rdata;
  reg [8-1:0] ram_w8_l2048_id0_0_0_wdata;
  reg ram_w8_l2048_id0_0_0_wenable;
  reg [9-1:0] ram_w8_l2048_id0_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id0_0_1_rdata;
  reg [8-1:0] ram_w8_l2048_id0_0_1_wdata;
  reg ram_w8_l2048_id0_0_1_wenable;

  ram_w8_l2048_id0_0
  inst_ram_w8_l2048_id0_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id0_0_0_addr(ram_w8_l2048_id0_0_0_addr),
    .ram_w8_l2048_id0_0_0_rdata(ram_w8_l2048_id0_0_0_rdata),
    .ram_w8_l2048_id0_0_0_wdata(ram_w8_l2048_id0_0_0_wdata),
    .ram_w8_l2048_id0_0_0_wenable(ram_w8_l2048_id0_0_0_wenable),
    .ram_w8_l2048_id0_0_1_addr(ram_w8_l2048_id0_0_1_addr),
    .ram_w8_l2048_id0_0_1_rdata(ram_w8_l2048_id0_0_1_rdata),
    .ram_w8_l2048_id0_0_1_wdata(ram_w8_l2048_id0_0_1_wdata),
    .ram_w8_l2048_id0_0_1_wenable(ram_w8_l2048_id0_0_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id0_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id0_1_0_rdata;
  reg [8-1:0] ram_w8_l2048_id0_1_0_wdata;
  reg ram_w8_l2048_id0_1_0_wenable;
  reg [9-1:0] ram_w8_l2048_id0_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id0_1_1_rdata;
  reg [8-1:0] ram_w8_l2048_id0_1_1_wdata;
  reg ram_w8_l2048_id0_1_1_wenable;

  ram_w8_l2048_id0_1
  inst_ram_w8_l2048_id0_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id0_1_0_addr(ram_w8_l2048_id0_1_0_addr),
    .ram_w8_l2048_id0_1_0_rdata(ram_w8_l2048_id0_1_0_rdata),
    .ram_w8_l2048_id0_1_0_wdata(ram_w8_l2048_id0_1_0_wdata),
    .ram_w8_l2048_id0_1_0_wenable(ram_w8_l2048_id0_1_0_wenable),
    .ram_w8_l2048_id0_1_1_addr(ram_w8_l2048_id0_1_1_addr),
    .ram_w8_l2048_id0_1_1_rdata(ram_w8_l2048_id0_1_1_rdata),
    .ram_w8_l2048_id0_1_1_wdata(ram_w8_l2048_id0_1_1_wdata),
    .ram_w8_l2048_id0_1_1_wenable(ram_w8_l2048_id0_1_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id0_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id0_2_0_rdata;
  reg [8-1:0] ram_w8_l2048_id0_2_0_wdata;
  reg ram_w8_l2048_id0_2_0_wenable;
  reg [9-1:0] ram_w8_l2048_id0_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id0_2_1_rdata;
  reg [8-1:0] ram_w8_l2048_id0_2_1_wdata;
  reg ram_w8_l2048_id0_2_1_wenable;

  ram_w8_l2048_id0_2
  inst_ram_w8_l2048_id0_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id0_2_0_addr(ram_w8_l2048_id0_2_0_addr),
    .ram_w8_l2048_id0_2_0_rdata(ram_w8_l2048_id0_2_0_rdata),
    .ram_w8_l2048_id0_2_0_wdata(ram_w8_l2048_id0_2_0_wdata),
    .ram_w8_l2048_id0_2_0_wenable(ram_w8_l2048_id0_2_0_wenable),
    .ram_w8_l2048_id0_2_1_addr(ram_w8_l2048_id0_2_1_addr),
    .ram_w8_l2048_id0_2_1_rdata(ram_w8_l2048_id0_2_1_rdata),
    .ram_w8_l2048_id0_2_1_wdata(ram_w8_l2048_id0_2_1_wdata),
    .ram_w8_l2048_id0_2_1_wenable(ram_w8_l2048_id0_2_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id0_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id0_3_0_rdata;
  reg [8-1:0] ram_w8_l2048_id0_3_0_wdata;
  reg ram_w8_l2048_id0_3_0_wenable;
  reg [9-1:0] ram_w8_l2048_id0_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id0_3_1_rdata;
  reg [8-1:0] ram_w8_l2048_id0_3_1_wdata;
  reg ram_w8_l2048_id0_3_1_wenable;

  ram_w8_l2048_id0_3
  inst_ram_w8_l2048_id0_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id0_3_0_addr(ram_w8_l2048_id0_3_0_addr),
    .ram_w8_l2048_id0_3_0_rdata(ram_w8_l2048_id0_3_0_rdata),
    .ram_w8_l2048_id0_3_0_wdata(ram_w8_l2048_id0_3_0_wdata),
    .ram_w8_l2048_id0_3_0_wenable(ram_w8_l2048_id0_3_0_wenable),
    .ram_w8_l2048_id0_3_1_addr(ram_w8_l2048_id0_3_1_addr),
    .ram_w8_l2048_id0_3_1_rdata(ram_w8_l2048_id0_3_1_rdata),
    .ram_w8_l2048_id0_3_1_wdata(ram_w8_l2048_id0_3_1_wdata),
    .ram_w8_l2048_id0_3_1_wenable(ram_w8_l2048_id0_3_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id1_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id1_0_0_rdata;
  reg [8-1:0] ram_w8_l2048_id1_0_0_wdata;
  reg ram_w8_l2048_id1_0_0_wenable;
  reg [9-1:0] ram_w8_l2048_id1_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id1_0_1_rdata;
  reg [8-1:0] ram_w8_l2048_id1_0_1_wdata;
  reg ram_w8_l2048_id1_0_1_wenable;

  ram_w8_l2048_id1_0
  inst_ram_w8_l2048_id1_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id1_0_0_addr(ram_w8_l2048_id1_0_0_addr),
    .ram_w8_l2048_id1_0_0_rdata(ram_w8_l2048_id1_0_0_rdata),
    .ram_w8_l2048_id1_0_0_wdata(ram_w8_l2048_id1_0_0_wdata),
    .ram_w8_l2048_id1_0_0_wenable(ram_w8_l2048_id1_0_0_wenable),
    .ram_w8_l2048_id1_0_1_addr(ram_w8_l2048_id1_0_1_addr),
    .ram_w8_l2048_id1_0_1_rdata(ram_w8_l2048_id1_0_1_rdata),
    .ram_w8_l2048_id1_0_1_wdata(ram_w8_l2048_id1_0_1_wdata),
    .ram_w8_l2048_id1_0_1_wenable(ram_w8_l2048_id1_0_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id1_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id1_1_0_rdata;
  reg [8-1:0] ram_w8_l2048_id1_1_0_wdata;
  reg ram_w8_l2048_id1_1_0_wenable;
  reg [9-1:0] ram_w8_l2048_id1_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id1_1_1_rdata;
  reg [8-1:0] ram_w8_l2048_id1_1_1_wdata;
  reg ram_w8_l2048_id1_1_1_wenable;

  ram_w8_l2048_id1_1
  inst_ram_w8_l2048_id1_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id1_1_0_addr(ram_w8_l2048_id1_1_0_addr),
    .ram_w8_l2048_id1_1_0_rdata(ram_w8_l2048_id1_1_0_rdata),
    .ram_w8_l2048_id1_1_0_wdata(ram_w8_l2048_id1_1_0_wdata),
    .ram_w8_l2048_id1_1_0_wenable(ram_w8_l2048_id1_1_0_wenable),
    .ram_w8_l2048_id1_1_1_addr(ram_w8_l2048_id1_1_1_addr),
    .ram_w8_l2048_id1_1_1_rdata(ram_w8_l2048_id1_1_1_rdata),
    .ram_w8_l2048_id1_1_1_wdata(ram_w8_l2048_id1_1_1_wdata),
    .ram_w8_l2048_id1_1_1_wenable(ram_w8_l2048_id1_1_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id1_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id1_2_0_rdata;
  reg [8-1:0] ram_w8_l2048_id1_2_0_wdata;
  reg ram_w8_l2048_id1_2_0_wenable;
  reg [9-1:0] ram_w8_l2048_id1_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id1_2_1_rdata;
  reg [8-1:0] ram_w8_l2048_id1_2_1_wdata;
  reg ram_w8_l2048_id1_2_1_wenable;

  ram_w8_l2048_id1_2
  inst_ram_w8_l2048_id1_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id1_2_0_addr(ram_w8_l2048_id1_2_0_addr),
    .ram_w8_l2048_id1_2_0_rdata(ram_w8_l2048_id1_2_0_rdata),
    .ram_w8_l2048_id1_2_0_wdata(ram_w8_l2048_id1_2_0_wdata),
    .ram_w8_l2048_id1_2_0_wenable(ram_w8_l2048_id1_2_0_wenable),
    .ram_w8_l2048_id1_2_1_addr(ram_w8_l2048_id1_2_1_addr),
    .ram_w8_l2048_id1_2_1_rdata(ram_w8_l2048_id1_2_1_rdata),
    .ram_w8_l2048_id1_2_1_wdata(ram_w8_l2048_id1_2_1_wdata),
    .ram_w8_l2048_id1_2_1_wenable(ram_w8_l2048_id1_2_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id1_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id1_3_0_rdata;
  reg [8-1:0] ram_w8_l2048_id1_3_0_wdata;
  reg ram_w8_l2048_id1_3_0_wenable;
  reg [9-1:0] ram_w8_l2048_id1_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id1_3_1_rdata;
  reg [8-1:0] ram_w8_l2048_id1_3_1_wdata;
  reg ram_w8_l2048_id1_3_1_wenable;

  ram_w8_l2048_id1_3
  inst_ram_w8_l2048_id1_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id1_3_0_addr(ram_w8_l2048_id1_3_0_addr),
    .ram_w8_l2048_id1_3_0_rdata(ram_w8_l2048_id1_3_0_rdata),
    .ram_w8_l2048_id1_3_0_wdata(ram_w8_l2048_id1_3_0_wdata),
    .ram_w8_l2048_id1_3_0_wenable(ram_w8_l2048_id1_3_0_wenable),
    .ram_w8_l2048_id1_3_1_addr(ram_w8_l2048_id1_3_1_addr),
    .ram_w8_l2048_id1_3_1_rdata(ram_w8_l2048_id1_3_1_rdata),
    .ram_w8_l2048_id1_3_1_wdata(ram_w8_l2048_id1_3_1_wdata),
    .ram_w8_l2048_id1_3_1_wenable(ram_w8_l2048_id1_3_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id2_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id2_0_0_rdata;
  reg [8-1:0] ram_w8_l2048_id2_0_0_wdata;
  reg ram_w8_l2048_id2_0_0_wenable;
  reg [9-1:0] ram_w8_l2048_id2_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id2_0_1_rdata;
  reg [8-1:0] ram_w8_l2048_id2_0_1_wdata;
  reg ram_w8_l2048_id2_0_1_wenable;

  ram_w8_l2048_id2_0
  inst_ram_w8_l2048_id2_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id2_0_0_addr(ram_w8_l2048_id2_0_0_addr),
    .ram_w8_l2048_id2_0_0_rdata(ram_w8_l2048_id2_0_0_rdata),
    .ram_w8_l2048_id2_0_0_wdata(ram_w8_l2048_id2_0_0_wdata),
    .ram_w8_l2048_id2_0_0_wenable(ram_w8_l2048_id2_0_0_wenable),
    .ram_w8_l2048_id2_0_1_addr(ram_w8_l2048_id2_0_1_addr),
    .ram_w8_l2048_id2_0_1_rdata(ram_w8_l2048_id2_0_1_rdata),
    .ram_w8_l2048_id2_0_1_wdata(ram_w8_l2048_id2_0_1_wdata),
    .ram_w8_l2048_id2_0_1_wenable(ram_w8_l2048_id2_0_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id2_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id2_1_0_rdata;
  reg [8-1:0] ram_w8_l2048_id2_1_0_wdata;
  reg ram_w8_l2048_id2_1_0_wenable;
  reg [9-1:0] ram_w8_l2048_id2_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id2_1_1_rdata;
  reg [8-1:0] ram_w8_l2048_id2_1_1_wdata;
  reg ram_w8_l2048_id2_1_1_wenable;

  ram_w8_l2048_id2_1
  inst_ram_w8_l2048_id2_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id2_1_0_addr(ram_w8_l2048_id2_1_0_addr),
    .ram_w8_l2048_id2_1_0_rdata(ram_w8_l2048_id2_1_0_rdata),
    .ram_w8_l2048_id2_1_0_wdata(ram_w8_l2048_id2_1_0_wdata),
    .ram_w8_l2048_id2_1_0_wenable(ram_w8_l2048_id2_1_0_wenable),
    .ram_w8_l2048_id2_1_1_addr(ram_w8_l2048_id2_1_1_addr),
    .ram_w8_l2048_id2_1_1_rdata(ram_w8_l2048_id2_1_1_rdata),
    .ram_w8_l2048_id2_1_1_wdata(ram_w8_l2048_id2_1_1_wdata),
    .ram_w8_l2048_id2_1_1_wenable(ram_w8_l2048_id2_1_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id2_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id2_2_0_rdata;
  reg [8-1:0] ram_w8_l2048_id2_2_0_wdata;
  reg ram_w8_l2048_id2_2_0_wenable;
  reg [9-1:0] ram_w8_l2048_id2_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id2_2_1_rdata;
  reg [8-1:0] ram_w8_l2048_id2_2_1_wdata;
  reg ram_w8_l2048_id2_2_1_wenable;

  ram_w8_l2048_id2_2
  inst_ram_w8_l2048_id2_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id2_2_0_addr(ram_w8_l2048_id2_2_0_addr),
    .ram_w8_l2048_id2_2_0_rdata(ram_w8_l2048_id2_2_0_rdata),
    .ram_w8_l2048_id2_2_0_wdata(ram_w8_l2048_id2_2_0_wdata),
    .ram_w8_l2048_id2_2_0_wenable(ram_w8_l2048_id2_2_0_wenable),
    .ram_w8_l2048_id2_2_1_addr(ram_w8_l2048_id2_2_1_addr),
    .ram_w8_l2048_id2_2_1_rdata(ram_w8_l2048_id2_2_1_rdata),
    .ram_w8_l2048_id2_2_1_wdata(ram_w8_l2048_id2_2_1_wdata),
    .ram_w8_l2048_id2_2_1_wenable(ram_w8_l2048_id2_2_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id2_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id2_3_0_rdata;
  reg [8-1:0] ram_w8_l2048_id2_3_0_wdata;
  reg ram_w8_l2048_id2_3_0_wenable;
  reg [9-1:0] ram_w8_l2048_id2_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id2_3_1_rdata;
  reg [8-1:0] ram_w8_l2048_id2_3_1_wdata;
  reg ram_w8_l2048_id2_3_1_wenable;

  ram_w8_l2048_id2_3
  inst_ram_w8_l2048_id2_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id2_3_0_addr(ram_w8_l2048_id2_3_0_addr),
    .ram_w8_l2048_id2_3_0_rdata(ram_w8_l2048_id2_3_0_rdata),
    .ram_w8_l2048_id2_3_0_wdata(ram_w8_l2048_id2_3_0_wdata),
    .ram_w8_l2048_id2_3_0_wenable(ram_w8_l2048_id2_3_0_wenable),
    .ram_w8_l2048_id2_3_1_addr(ram_w8_l2048_id2_3_1_addr),
    .ram_w8_l2048_id2_3_1_rdata(ram_w8_l2048_id2_3_1_rdata),
    .ram_w8_l2048_id2_3_1_wdata(ram_w8_l2048_id2_3_1_wdata),
    .ram_w8_l2048_id2_3_1_wenable(ram_w8_l2048_id2_3_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id3_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id3_0_0_rdata;
  reg [8-1:0] ram_w8_l2048_id3_0_0_wdata;
  reg ram_w8_l2048_id3_0_0_wenable;
  reg [9-1:0] ram_w8_l2048_id3_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id3_0_1_rdata;
  reg [8-1:0] ram_w8_l2048_id3_0_1_wdata;
  reg ram_w8_l2048_id3_0_1_wenable;

  ram_w8_l2048_id3_0
  inst_ram_w8_l2048_id3_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id3_0_0_addr(ram_w8_l2048_id3_0_0_addr),
    .ram_w8_l2048_id3_0_0_rdata(ram_w8_l2048_id3_0_0_rdata),
    .ram_w8_l2048_id3_0_0_wdata(ram_w8_l2048_id3_0_0_wdata),
    .ram_w8_l2048_id3_0_0_wenable(ram_w8_l2048_id3_0_0_wenable),
    .ram_w8_l2048_id3_0_1_addr(ram_w8_l2048_id3_0_1_addr),
    .ram_w8_l2048_id3_0_1_rdata(ram_w8_l2048_id3_0_1_rdata),
    .ram_w8_l2048_id3_0_1_wdata(ram_w8_l2048_id3_0_1_wdata),
    .ram_w8_l2048_id3_0_1_wenable(ram_w8_l2048_id3_0_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id3_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id3_1_0_rdata;
  reg [8-1:0] ram_w8_l2048_id3_1_0_wdata;
  reg ram_w8_l2048_id3_1_0_wenable;
  reg [9-1:0] ram_w8_l2048_id3_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id3_1_1_rdata;
  reg [8-1:0] ram_w8_l2048_id3_1_1_wdata;
  reg ram_w8_l2048_id3_1_1_wenable;

  ram_w8_l2048_id3_1
  inst_ram_w8_l2048_id3_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id3_1_0_addr(ram_w8_l2048_id3_1_0_addr),
    .ram_w8_l2048_id3_1_0_rdata(ram_w8_l2048_id3_1_0_rdata),
    .ram_w8_l2048_id3_1_0_wdata(ram_w8_l2048_id3_1_0_wdata),
    .ram_w8_l2048_id3_1_0_wenable(ram_w8_l2048_id3_1_0_wenable),
    .ram_w8_l2048_id3_1_1_addr(ram_w8_l2048_id3_1_1_addr),
    .ram_w8_l2048_id3_1_1_rdata(ram_w8_l2048_id3_1_1_rdata),
    .ram_w8_l2048_id3_1_1_wdata(ram_w8_l2048_id3_1_1_wdata),
    .ram_w8_l2048_id3_1_1_wenable(ram_w8_l2048_id3_1_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id3_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id3_2_0_rdata;
  reg [8-1:0] ram_w8_l2048_id3_2_0_wdata;
  reg ram_w8_l2048_id3_2_0_wenable;
  reg [9-1:0] ram_w8_l2048_id3_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id3_2_1_rdata;
  reg [8-1:0] ram_w8_l2048_id3_2_1_wdata;
  reg ram_w8_l2048_id3_2_1_wenable;

  ram_w8_l2048_id3_2
  inst_ram_w8_l2048_id3_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id3_2_0_addr(ram_w8_l2048_id3_2_0_addr),
    .ram_w8_l2048_id3_2_0_rdata(ram_w8_l2048_id3_2_0_rdata),
    .ram_w8_l2048_id3_2_0_wdata(ram_w8_l2048_id3_2_0_wdata),
    .ram_w8_l2048_id3_2_0_wenable(ram_w8_l2048_id3_2_0_wenable),
    .ram_w8_l2048_id3_2_1_addr(ram_w8_l2048_id3_2_1_addr),
    .ram_w8_l2048_id3_2_1_rdata(ram_w8_l2048_id3_2_1_rdata),
    .ram_w8_l2048_id3_2_1_wdata(ram_w8_l2048_id3_2_1_wdata),
    .ram_w8_l2048_id3_2_1_wenable(ram_w8_l2048_id3_2_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id3_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id3_3_0_rdata;
  reg [8-1:0] ram_w8_l2048_id3_3_0_wdata;
  reg ram_w8_l2048_id3_3_0_wenable;
  reg [9-1:0] ram_w8_l2048_id3_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id3_3_1_rdata;
  reg [8-1:0] ram_w8_l2048_id3_3_1_wdata;
  reg ram_w8_l2048_id3_3_1_wenable;

  ram_w8_l2048_id3_3
  inst_ram_w8_l2048_id3_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id3_3_0_addr(ram_w8_l2048_id3_3_0_addr),
    .ram_w8_l2048_id3_3_0_rdata(ram_w8_l2048_id3_3_0_rdata),
    .ram_w8_l2048_id3_3_0_wdata(ram_w8_l2048_id3_3_0_wdata),
    .ram_w8_l2048_id3_3_0_wenable(ram_w8_l2048_id3_3_0_wenable),
    .ram_w8_l2048_id3_3_1_addr(ram_w8_l2048_id3_3_1_addr),
    .ram_w8_l2048_id3_3_1_rdata(ram_w8_l2048_id3_3_1_rdata),
    .ram_w8_l2048_id3_3_1_wdata(ram_w8_l2048_id3_3_1_wdata),
    .ram_w8_l2048_id3_3_1_wenable(ram_w8_l2048_id3_3_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id4_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id4_0_0_rdata;
  reg [8-1:0] ram_w8_l2048_id4_0_0_wdata;
  reg ram_w8_l2048_id4_0_0_wenable;
  reg [9-1:0] ram_w8_l2048_id4_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id4_0_1_rdata;
  reg [8-1:0] ram_w8_l2048_id4_0_1_wdata;
  reg ram_w8_l2048_id4_0_1_wenable;

  ram_w8_l2048_id4_0
  inst_ram_w8_l2048_id4_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id4_0_0_addr(ram_w8_l2048_id4_0_0_addr),
    .ram_w8_l2048_id4_0_0_rdata(ram_w8_l2048_id4_0_0_rdata),
    .ram_w8_l2048_id4_0_0_wdata(ram_w8_l2048_id4_0_0_wdata),
    .ram_w8_l2048_id4_0_0_wenable(ram_w8_l2048_id4_0_0_wenable),
    .ram_w8_l2048_id4_0_1_addr(ram_w8_l2048_id4_0_1_addr),
    .ram_w8_l2048_id4_0_1_rdata(ram_w8_l2048_id4_0_1_rdata),
    .ram_w8_l2048_id4_0_1_wdata(ram_w8_l2048_id4_0_1_wdata),
    .ram_w8_l2048_id4_0_1_wenable(ram_w8_l2048_id4_0_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id4_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id4_1_0_rdata;
  reg [8-1:0] ram_w8_l2048_id4_1_0_wdata;
  reg ram_w8_l2048_id4_1_0_wenable;
  reg [9-1:0] ram_w8_l2048_id4_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id4_1_1_rdata;
  reg [8-1:0] ram_w8_l2048_id4_1_1_wdata;
  reg ram_w8_l2048_id4_1_1_wenable;

  ram_w8_l2048_id4_1
  inst_ram_w8_l2048_id4_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id4_1_0_addr(ram_w8_l2048_id4_1_0_addr),
    .ram_w8_l2048_id4_1_0_rdata(ram_w8_l2048_id4_1_0_rdata),
    .ram_w8_l2048_id4_1_0_wdata(ram_w8_l2048_id4_1_0_wdata),
    .ram_w8_l2048_id4_1_0_wenable(ram_w8_l2048_id4_1_0_wenable),
    .ram_w8_l2048_id4_1_1_addr(ram_w8_l2048_id4_1_1_addr),
    .ram_w8_l2048_id4_1_1_rdata(ram_w8_l2048_id4_1_1_rdata),
    .ram_w8_l2048_id4_1_1_wdata(ram_w8_l2048_id4_1_1_wdata),
    .ram_w8_l2048_id4_1_1_wenable(ram_w8_l2048_id4_1_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id4_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id4_2_0_rdata;
  reg [8-1:0] ram_w8_l2048_id4_2_0_wdata;
  reg ram_w8_l2048_id4_2_0_wenable;
  reg [9-1:0] ram_w8_l2048_id4_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id4_2_1_rdata;
  reg [8-1:0] ram_w8_l2048_id4_2_1_wdata;
  reg ram_w8_l2048_id4_2_1_wenable;

  ram_w8_l2048_id4_2
  inst_ram_w8_l2048_id4_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id4_2_0_addr(ram_w8_l2048_id4_2_0_addr),
    .ram_w8_l2048_id4_2_0_rdata(ram_w8_l2048_id4_2_0_rdata),
    .ram_w8_l2048_id4_2_0_wdata(ram_w8_l2048_id4_2_0_wdata),
    .ram_w8_l2048_id4_2_0_wenable(ram_w8_l2048_id4_2_0_wenable),
    .ram_w8_l2048_id4_2_1_addr(ram_w8_l2048_id4_2_1_addr),
    .ram_w8_l2048_id4_2_1_rdata(ram_w8_l2048_id4_2_1_rdata),
    .ram_w8_l2048_id4_2_1_wdata(ram_w8_l2048_id4_2_1_wdata),
    .ram_w8_l2048_id4_2_1_wenable(ram_w8_l2048_id4_2_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id4_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id4_3_0_rdata;
  reg [8-1:0] ram_w8_l2048_id4_3_0_wdata;
  reg ram_w8_l2048_id4_3_0_wenable;
  reg [9-1:0] ram_w8_l2048_id4_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id4_3_1_rdata;
  reg [8-1:0] ram_w8_l2048_id4_3_1_wdata;
  reg ram_w8_l2048_id4_3_1_wenable;

  ram_w8_l2048_id4_3
  inst_ram_w8_l2048_id4_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id4_3_0_addr(ram_w8_l2048_id4_3_0_addr),
    .ram_w8_l2048_id4_3_0_rdata(ram_w8_l2048_id4_3_0_rdata),
    .ram_w8_l2048_id4_3_0_wdata(ram_w8_l2048_id4_3_0_wdata),
    .ram_w8_l2048_id4_3_0_wenable(ram_w8_l2048_id4_3_0_wenable),
    .ram_w8_l2048_id4_3_1_addr(ram_w8_l2048_id4_3_1_addr),
    .ram_w8_l2048_id4_3_1_rdata(ram_w8_l2048_id4_3_1_rdata),
    .ram_w8_l2048_id4_3_1_wdata(ram_w8_l2048_id4_3_1_wdata),
    .ram_w8_l2048_id4_3_1_wenable(ram_w8_l2048_id4_3_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id5_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id5_0_0_rdata;
  reg [8-1:0] ram_w8_l2048_id5_0_0_wdata;
  reg ram_w8_l2048_id5_0_0_wenable;
  reg [9-1:0] ram_w8_l2048_id5_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id5_0_1_rdata;
  reg [8-1:0] ram_w8_l2048_id5_0_1_wdata;
  reg ram_w8_l2048_id5_0_1_wenable;

  ram_w8_l2048_id5_0
  inst_ram_w8_l2048_id5_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id5_0_0_addr(ram_w8_l2048_id5_0_0_addr),
    .ram_w8_l2048_id5_0_0_rdata(ram_w8_l2048_id5_0_0_rdata),
    .ram_w8_l2048_id5_0_0_wdata(ram_w8_l2048_id5_0_0_wdata),
    .ram_w8_l2048_id5_0_0_wenable(ram_w8_l2048_id5_0_0_wenable),
    .ram_w8_l2048_id5_0_1_addr(ram_w8_l2048_id5_0_1_addr),
    .ram_w8_l2048_id5_0_1_rdata(ram_w8_l2048_id5_0_1_rdata),
    .ram_w8_l2048_id5_0_1_wdata(ram_w8_l2048_id5_0_1_wdata),
    .ram_w8_l2048_id5_0_1_wenable(ram_w8_l2048_id5_0_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id5_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id5_1_0_rdata;
  reg [8-1:0] ram_w8_l2048_id5_1_0_wdata;
  reg ram_w8_l2048_id5_1_0_wenable;
  reg [9-1:0] ram_w8_l2048_id5_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id5_1_1_rdata;
  reg [8-1:0] ram_w8_l2048_id5_1_1_wdata;
  reg ram_w8_l2048_id5_1_1_wenable;

  ram_w8_l2048_id5_1
  inst_ram_w8_l2048_id5_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id5_1_0_addr(ram_w8_l2048_id5_1_0_addr),
    .ram_w8_l2048_id5_1_0_rdata(ram_w8_l2048_id5_1_0_rdata),
    .ram_w8_l2048_id5_1_0_wdata(ram_w8_l2048_id5_1_0_wdata),
    .ram_w8_l2048_id5_1_0_wenable(ram_w8_l2048_id5_1_0_wenable),
    .ram_w8_l2048_id5_1_1_addr(ram_w8_l2048_id5_1_1_addr),
    .ram_w8_l2048_id5_1_1_rdata(ram_w8_l2048_id5_1_1_rdata),
    .ram_w8_l2048_id5_1_1_wdata(ram_w8_l2048_id5_1_1_wdata),
    .ram_w8_l2048_id5_1_1_wenable(ram_w8_l2048_id5_1_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id5_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id5_2_0_rdata;
  reg [8-1:0] ram_w8_l2048_id5_2_0_wdata;
  reg ram_w8_l2048_id5_2_0_wenable;
  reg [9-1:0] ram_w8_l2048_id5_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id5_2_1_rdata;
  reg [8-1:0] ram_w8_l2048_id5_2_1_wdata;
  reg ram_w8_l2048_id5_2_1_wenable;

  ram_w8_l2048_id5_2
  inst_ram_w8_l2048_id5_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id5_2_0_addr(ram_w8_l2048_id5_2_0_addr),
    .ram_w8_l2048_id5_2_0_rdata(ram_w8_l2048_id5_2_0_rdata),
    .ram_w8_l2048_id5_2_0_wdata(ram_w8_l2048_id5_2_0_wdata),
    .ram_w8_l2048_id5_2_0_wenable(ram_w8_l2048_id5_2_0_wenable),
    .ram_w8_l2048_id5_2_1_addr(ram_w8_l2048_id5_2_1_addr),
    .ram_w8_l2048_id5_2_1_rdata(ram_w8_l2048_id5_2_1_rdata),
    .ram_w8_l2048_id5_2_1_wdata(ram_w8_l2048_id5_2_1_wdata),
    .ram_w8_l2048_id5_2_1_wenable(ram_w8_l2048_id5_2_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id5_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id5_3_0_rdata;
  reg [8-1:0] ram_w8_l2048_id5_3_0_wdata;
  reg ram_w8_l2048_id5_3_0_wenable;
  reg [9-1:0] ram_w8_l2048_id5_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id5_3_1_rdata;
  reg [8-1:0] ram_w8_l2048_id5_3_1_wdata;
  reg ram_w8_l2048_id5_3_1_wenable;

  ram_w8_l2048_id5_3
  inst_ram_w8_l2048_id5_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id5_3_0_addr(ram_w8_l2048_id5_3_0_addr),
    .ram_w8_l2048_id5_3_0_rdata(ram_w8_l2048_id5_3_0_rdata),
    .ram_w8_l2048_id5_3_0_wdata(ram_w8_l2048_id5_3_0_wdata),
    .ram_w8_l2048_id5_3_0_wenable(ram_w8_l2048_id5_3_0_wenable),
    .ram_w8_l2048_id5_3_1_addr(ram_w8_l2048_id5_3_1_addr),
    .ram_w8_l2048_id5_3_1_rdata(ram_w8_l2048_id5_3_1_rdata),
    .ram_w8_l2048_id5_3_1_wdata(ram_w8_l2048_id5_3_1_wdata),
    .ram_w8_l2048_id5_3_1_wenable(ram_w8_l2048_id5_3_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id6_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id6_0_0_rdata;
  reg [8-1:0] ram_w8_l2048_id6_0_0_wdata;
  reg ram_w8_l2048_id6_0_0_wenable;
  reg [9-1:0] ram_w8_l2048_id6_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id6_0_1_rdata;
  reg [8-1:0] ram_w8_l2048_id6_0_1_wdata;
  reg ram_w8_l2048_id6_0_1_wenable;

  ram_w8_l2048_id6_0
  inst_ram_w8_l2048_id6_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id6_0_0_addr(ram_w8_l2048_id6_0_0_addr),
    .ram_w8_l2048_id6_0_0_rdata(ram_w8_l2048_id6_0_0_rdata),
    .ram_w8_l2048_id6_0_0_wdata(ram_w8_l2048_id6_0_0_wdata),
    .ram_w8_l2048_id6_0_0_wenable(ram_w8_l2048_id6_0_0_wenable),
    .ram_w8_l2048_id6_0_1_addr(ram_w8_l2048_id6_0_1_addr),
    .ram_w8_l2048_id6_0_1_rdata(ram_w8_l2048_id6_0_1_rdata),
    .ram_w8_l2048_id6_0_1_wdata(ram_w8_l2048_id6_0_1_wdata),
    .ram_w8_l2048_id6_0_1_wenable(ram_w8_l2048_id6_0_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id6_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id6_1_0_rdata;
  reg [8-1:0] ram_w8_l2048_id6_1_0_wdata;
  reg ram_w8_l2048_id6_1_0_wenable;
  reg [9-1:0] ram_w8_l2048_id6_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id6_1_1_rdata;
  reg [8-1:0] ram_w8_l2048_id6_1_1_wdata;
  reg ram_w8_l2048_id6_1_1_wenable;

  ram_w8_l2048_id6_1
  inst_ram_w8_l2048_id6_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id6_1_0_addr(ram_w8_l2048_id6_1_0_addr),
    .ram_w8_l2048_id6_1_0_rdata(ram_w8_l2048_id6_1_0_rdata),
    .ram_w8_l2048_id6_1_0_wdata(ram_w8_l2048_id6_1_0_wdata),
    .ram_w8_l2048_id6_1_0_wenable(ram_w8_l2048_id6_1_0_wenable),
    .ram_w8_l2048_id6_1_1_addr(ram_w8_l2048_id6_1_1_addr),
    .ram_w8_l2048_id6_1_1_rdata(ram_w8_l2048_id6_1_1_rdata),
    .ram_w8_l2048_id6_1_1_wdata(ram_w8_l2048_id6_1_1_wdata),
    .ram_w8_l2048_id6_1_1_wenable(ram_w8_l2048_id6_1_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id6_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id6_2_0_rdata;
  reg [8-1:0] ram_w8_l2048_id6_2_0_wdata;
  reg ram_w8_l2048_id6_2_0_wenable;
  reg [9-1:0] ram_w8_l2048_id6_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id6_2_1_rdata;
  reg [8-1:0] ram_w8_l2048_id6_2_1_wdata;
  reg ram_w8_l2048_id6_2_1_wenable;

  ram_w8_l2048_id6_2
  inst_ram_w8_l2048_id6_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id6_2_0_addr(ram_w8_l2048_id6_2_0_addr),
    .ram_w8_l2048_id6_2_0_rdata(ram_w8_l2048_id6_2_0_rdata),
    .ram_w8_l2048_id6_2_0_wdata(ram_w8_l2048_id6_2_0_wdata),
    .ram_w8_l2048_id6_2_0_wenable(ram_w8_l2048_id6_2_0_wenable),
    .ram_w8_l2048_id6_2_1_addr(ram_w8_l2048_id6_2_1_addr),
    .ram_w8_l2048_id6_2_1_rdata(ram_w8_l2048_id6_2_1_rdata),
    .ram_w8_l2048_id6_2_1_wdata(ram_w8_l2048_id6_2_1_wdata),
    .ram_w8_l2048_id6_2_1_wenable(ram_w8_l2048_id6_2_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id6_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id6_3_0_rdata;
  reg [8-1:0] ram_w8_l2048_id6_3_0_wdata;
  reg ram_w8_l2048_id6_3_0_wenable;
  reg [9-1:0] ram_w8_l2048_id6_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id6_3_1_rdata;
  reg [8-1:0] ram_w8_l2048_id6_3_1_wdata;
  reg ram_w8_l2048_id6_3_1_wenable;

  ram_w8_l2048_id6_3
  inst_ram_w8_l2048_id6_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id6_3_0_addr(ram_w8_l2048_id6_3_0_addr),
    .ram_w8_l2048_id6_3_0_rdata(ram_w8_l2048_id6_3_0_rdata),
    .ram_w8_l2048_id6_3_0_wdata(ram_w8_l2048_id6_3_0_wdata),
    .ram_w8_l2048_id6_3_0_wenable(ram_w8_l2048_id6_3_0_wenable),
    .ram_w8_l2048_id6_3_1_addr(ram_w8_l2048_id6_3_1_addr),
    .ram_w8_l2048_id6_3_1_rdata(ram_w8_l2048_id6_3_1_rdata),
    .ram_w8_l2048_id6_3_1_wdata(ram_w8_l2048_id6_3_1_wdata),
    .ram_w8_l2048_id6_3_1_wenable(ram_w8_l2048_id6_3_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id7_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id7_0_0_rdata;
  reg [8-1:0] ram_w8_l2048_id7_0_0_wdata;
  reg ram_w8_l2048_id7_0_0_wenable;
  reg [9-1:0] ram_w8_l2048_id7_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id7_0_1_rdata;
  reg [8-1:0] ram_w8_l2048_id7_0_1_wdata;
  reg ram_w8_l2048_id7_0_1_wenable;

  ram_w8_l2048_id7_0
  inst_ram_w8_l2048_id7_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id7_0_0_addr(ram_w8_l2048_id7_0_0_addr),
    .ram_w8_l2048_id7_0_0_rdata(ram_w8_l2048_id7_0_0_rdata),
    .ram_w8_l2048_id7_0_0_wdata(ram_w8_l2048_id7_0_0_wdata),
    .ram_w8_l2048_id7_0_0_wenable(ram_w8_l2048_id7_0_0_wenable),
    .ram_w8_l2048_id7_0_1_addr(ram_w8_l2048_id7_0_1_addr),
    .ram_w8_l2048_id7_0_1_rdata(ram_w8_l2048_id7_0_1_rdata),
    .ram_w8_l2048_id7_0_1_wdata(ram_w8_l2048_id7_0_1_wdata),
    .ram_w8_l2048_id7_0_1_wenable(ram_w8_l2048_id7_0_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id7_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id7_1_0_rdata;
  reg [8-1:0] ram_w8_l2048_id7_1_0_wdata;
  reg ram_w8_l2048_id7_1_0_wenable;
  reg [9-1:0] ram_w8_l2048_id7_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id7_1_1_rdata;
  reg [8-1:0] ram_w8_l2048_id7_1_1_wdata;
  reg ram_w8_l2048_id7_1_1_wenable;

  ram_w8_l2048_id7_1
  inst_ram_w8_l2048_id7_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id7_1_0_addr(ram_w8_l2048_id7_1_0_addr),
    .ram_w8_l2048_id7_1_0_rdata(ram_w8_l2048_id7_1_0_rdata),
    .ram_w8_l2048_id7_1_0_wdata(ram_w8_l2048_id7_1_0_wdata),
    .ram_w8_l2048_id7_1_0_wenable(ram_w8_l2048_id7_1_0_wenable),
    .ram_w8_l2048_id7_1_1_addr(ram_w8_l2048_id7_1_1_addr),
    .ram_w8_l2048_id7_1_1_rdata(ram_w8_l2048_id7_1_1_rdata),
    .ram_w8_l2048_id7_1_1_wdata(ram_w8_l2048_id7_1_1_wdata),
    .ram_w8_l2048_id7_1_1_wenable(ram_w8_l2048_id7_1_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id7_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id7_2_0_rdata;
  reg [8-1:0] ram_w8_l2048_id7_2_0_wdata;
  reg ram_w8_l2048_id7_2_0_wenable;
  reg [9-1:0] ram_w8_l2048_id7_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id7_2_1_rdata;
  reg [8-1:0] ram_w8_l2048_id7_2_1_wdata;
  reg ram_w8_l2048_id7_2_1_wenable;

  ram_w8_l2048_id7_2
  inst_ram_w8_l2048_id7_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id7_2_0_addr(ram_w8_l2048_id7_2_0_addr),
    .ram_w8_l2048_id7_2_0_rdata(ram_w8_l2048_id7_2_0_rdata),
    .ram_w8_l2048_id7_2_0_wdata(ram_w8_l2048_id7_2_0_wdata),
    .ram_w8_l2048_id7_2_0_wenable(ram_w8_l2048_id7_2_0_wenable),
    .ram_w8_l2048_id7_2_1_addr(ram_w8_l2048_id7_2_1_addr),
    .ram_w8_l2048_id7_2_1_rdata(ram_w8_l2048_id7_2_1_rdata),
    .ram_w8_l2048_id7_2_1_wdata(ram_w8_l2048_id7_2_1_wdata),
    .ram_w8_l2048_id7_2_1_wenable(ram_w8_l2048_id7_2_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id7_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id7_3_0_rdata;
  reg [8-1:0] ram_w8_l2048_id7_3_0_wdata;
  reg ram_w8_l2048_id7_3_0_wenable;
  reg [9-1:0] ram_w8_l2048_id7_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id7_3_1_rdata;
  reg [8-1:0] ram_w8_l2048_id7_3_1_wdata;
  reg ram_w8_l2048_id7_3_1_wenable;

  ram_w8_l2048_id7_3
  inst_ram_w8_l2048_id7_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id7_3_0_addr(ram_w8_l2048_id7_3_0_addr),
    .ram_w8_l2048_id7_3_0_rdata(ram_w8_l2048_id7_3_0_rdata),
    .ram_w8_l2048_id7_3_0_wdata(ram_w8_l2048_id7_3_0_wdata),
    .ram_w8_l2048_id7_3_0_wenable(ram_w8_l2048_id7_3_0_wenable),
    .ram_w8_l2048_id7_3_1_addr(ram_w8_l2048_id7_3_1_addr),
    .ram_w8_l2048_id7_3_1_rdata(ram_w8_l2048_id7_3_1_rdata),
    .ram_w8_l2048_id7_3_1_wdata(ram_w8_l2048_id7_3_1_wdata),
    .ram_w8_l2048_id7_3_1_wenable(ram_w8_l2048_id7_3_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id8_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id8_0_0_rdata;
  reg [8-1:0] ram_w8_l2048_id8_0_0_wdata;
  reg ram_w8_l2048_id8_0_0_wenable;
  reg [9-1:0] ram_w8_l2048_id8_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id8_0_1_rdata;
  reg [8-1:0] ram_w8_l2048_id8_0_1_wdata;
  reg ram_w8_l2048_id8_0_1_wenable;

  ram_w8_l2048_id8_0
  inst_ram_w8_l2048_id8_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id8_0_0_addr(ram_w8_l2048_id8_0_0_addr),
    .ram_w8_l2048_id8_0_0_rdata(ram_w8_l2048_id8_0_0_rdata),
    .ram_w8_l2048_id8_0_0_wdata(ram_w8_l2048_id8_0_0_wdata),
    .ram_w8_l2048_id8_0_0_wenable(ram_w8_l2048_id8_0_0_wenable),
    .ram_w8_l2048_id8_0_1_addr(ram_w8_l2048_id8_0_1_addr),
    .ram_w8_l2048_id8_0_1_rdata(ram_w8_l2048_id8_0_1_rdata),
    .ram_w8_l2048_id8_0_1_wdata(ram_w8_l2048_id8_0_1_wdata),
    .ram_w8_l2048_id8_0_1_wenable(ram_w8_l2048_id8_0_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id8_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id8_1_0_rdata;
  reg [8-1:0] ram_w8_l2048_id8_1_0_wdata;
  reg ram_w8_l2048_id8_1_0_wenable;
  reg [9-1:0] ram_w8_l2048_id8_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id8_1_1_rdata;
  reg [8-1:0] ram_w8_l2048_id8_1_1_wdata;
  reg ram_w8_l2048_id8_1_1_wenable;

  ram_w8_l2048_id8_1
  inst_ram_w8_l2048_id8_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id8_1_0_addr(ram_w8_l2048_id8_1_0_addr),
    .ram_w8_l2048_id8_1_0_rdata(ram_w8_l2048_id8_1_0_rdata),
    .ram_w8_l2048_id8_1_0_wdata(ram_w8_l2048_id8_1_0_wdata),
    .ram_w8_l2048_id8_1_0_wenable(ram_w8_l2048_id8_1_0_wenable),
    .ram_w8_l2048_id8_1_1_addr(ram_w8_l2048_id8_1_1_addr),
    .ram_w8_l2048_id8_1_1_rdata(ram_w8_l2048_id8_1_1_rdata),
    .ram_w8_l2048_id8_1_1_wdata(ram_w8_l2048_id8_1_1_wdata),
    .ram_w8_l2048_id8_1_1_wenable(ram_w8_l2048_id8_1_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id8_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id8_2_0_rdata;
  reg [8-1:0] ram_w8_l2048_id8_2_0_wdata;
  reg ram_w8_l2048_id8_2_0_wenable;
  reg [9-1:0] ram_w8_l2048_id8_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id8_2_1_rdata;
  reg [8-1:0] ram_w8_l2048_id8_2_1_wdata;
  reg ram_w8_l2048_id8_2_1_wenable;

  ram_w8_l2048_id8_2
  inst_ram_w8_l2048_id8_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id8_2_0_addr(ram_w8_l2048_id8_2_0_addr),
    .ram_w8_l2048_id8_2_0_rdata(ram_w8_l2048_id8_2_0_rdata),
    .ram_w8_l2048_id8_2_0_wdata(ram_w8_l2048_id8_2_0_wdata),
    .ram_w8_l2048_id8_2_0_wenable(ram_w8_l2048_id8_2_0_wenable),
    .ram_w8_l2048_id8_2_1_addr(ram_w8_l2048_id8_2_1_addr),
    .ram_w8_l2048_id8_2_1_rdata(ram_w8_l2048_id8_2_1_rdata),
    .ram_w8_l2048_id8_2_1_wdata(ram_w8_l2048_id8_2_1_wdata),
    .ram_w8_l2048_id8_2_1_wenable(ram_w8_l2048_id8_2_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id8_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id8_3_0_rdata;
  reg [8-1:0] ram_w8_l2048_id8_3_0_wdata;
  reg ram_w8_l2048_id8_3_0_wenable;
  reg [9-1:0] ram_w8_l2048_id8_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id8_3_1_rdata;
  reg [8-1:0] ram_w8_l2048_id8_3_1_wdata;
  reg ram_w8_l2048_id8_3_1_wenable;

  ram_w8_l2048_id8_3
  inst_ram_w8_l2048_id8_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id8_3_0_addr(ram_w8_l2048_id8_3_0_addr),
    .ram_w8_l2048_id8_3_0_rdata(ram_w8_l2048_id8_3_0_rdata),
    .ram_w8_l2048_id8_3_0_wdata(ram_w8_l2048_id8_3_0_wdata),
    .ram_w8_l2048_id8_3_0_wenable(ram_w8_l2048_id8_3_0_wenable),
    .ram_w8_l2048_id8_3_1_addr(ram_w8_l2048_id8_3_1_addr),
    .ram_w8_l2048_id8_3_1_rdata(ram_w8_l2048_id8_3_1_rdata),
    .ram_w8_l2048_id8_3_1_wdata(ram_w8_l2048_id8_3_1_wdata),
    .ram_w8_l2048_id8_3_1_wenable(ram_w8_l2048_id8_3_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id9_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id9_0_0_rdata;
  reg [8-1:0] ram_w8_l2048_id9_0_0_wdata;
  reg ram_w8_l2048_id9_0_0_wenable;
  reg [9-1:0] ram_w8_l2048_id9_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id9_0_1_rdata;
  reg [8-1:0] ram_w8_l2048_id9_0_1_wdata;
  reg ram_w8_l2048_id9_0_1_wenable;

  ram_w8_l2048_id9_0
  inst_ram_w8_l2048_id9_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id9_0_0_addr(ram_w8_l2048_id9_0_0_addr),
    .ram_w8_l2048_id9_0_0_rdata(ram_w8_l2048_id9_0_0_rdata),
    .ram_w8_l2048_id9_0_0_wdata(ram_w8_l2048_id9_0_0_wdata),
    .ram_w8_l2048_id9_0_0_wenable(ram_w8_l2048_id9_0_0_wenable),
    .ram_w8_l2048_id9_0_1_addr(ram_w8_l2048_id9_0_1_addr),
    .ram_w8_l2048_id9_0_1_rdata(ram_w8_l2048_id9_0_1_rdata),
    .ram_w8_l2048_id9_0_1_wdata(ram_w8_l2048_id9_0_1_wdata),
    .ram_w8_l2048_id9_0_1_wenable(ram_w8_l2048_id9_0_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id9_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id9_1_0_rdata;
  reg [8-1:0] ram_w8_l2048_id9_1_0_wdata;
  reg ram_w8_l2048_id9_1_0_wenable;
  reg [9-1:0] ram_w8_l2048_id9_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id9_1_1_rdata;
  reg [8-1:0] ram_w8_l2048_id9_1_1_wdata;
  reg ram_w8_l2048_id9_1_1_wenable;

  ram_w8_l2048_id9_1
  inst_ram_w8_l2048_id9_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id9_1_0_addr(ram_w8_l2048_id9_1_0_addr),
    .ram_w8_l2048_id9_1_0_rdata(ram_w8_l2048_id9_1_0_rdata),
    .ram_w8_l2048_id9_1_0_wdata(ram_w8_l2048_id9_1_0_wdata),
    .ram_w8_l2048_id9_1_0_wenable(ram_w8_l2048_id9_1_0_wenable),
    .ram_w8_l2048_id9_1_1_addr(ram_w8_l2048_id9_1_1_addr),
    .ram_w8_l2048_id9_1_1_rdata(ram_w8_l2048_id9_1_1_rdata),
    .ram_w8_l2048_id9_1_1_wdata(ram_w8_l2048_id9_1_1_wdata),
    .ram_w8_l2048_id9_1_1_wenable(ram_w8_l2048_id9_1_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id9_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id9_2_0_rdata;
  reg [8-1:0] ram_w8_l2048_id9_2_0_wdata;
  reg ram_w8_l2048_id9_2_0_wenable;
  reg [9-1:0] ram_w8_l2048_id9_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id9_2_1_rdata;
  reg [8-1:0] ram_w8_l2048_id9_2_1_wdata;
  reg ram_w8_l2048_id9_2_1_wenable;

  ram_w8_l2048_id9_2
  inst_ram_w8_l2048_id9_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id9_2_0_addr(ram_w8_l2048_id9_2_0_addr),
    .ram_w8_l2048_id9_2_0_rdata(ram_w8_l2048_id9_2_0_rdata),
    .ram_w8_l2048_id9_2_0_wdata(ram_w8_l2048_id9_2_0_wdata),
    .ram_w8_l2048_id9_2_0_wenable(ram_w8_l2048_id9_2_0_wenable),
    .ram_w8_l2048_id9_2_1_addr(ram_w8_l2048_id9_2_1_addr),
    .ram_w8_l2048_id9_2_1_rdata(ram_w8_l2048_id9_2_1_rdata),
    .ram_w8_l2048_id9_2_1_wdata(ram_w8_l2048_id9_2_1_wdata),
    .ram_w8_l2048_id9_2_1_wenable(ram_w8_l2048_id9_2_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id9_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id9_3_0_rdata;
  reg [8-1:0] ram_w8_l2048_id9_3_0_wdata;
  reg ram_w8_l2048_id9_3_0_wenable;
  reg [9-1:0] ram_w8_l2048_id9_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id9_3_1_rdata;
  reg [8-1:0] ram_w8_l2048_id9_3_1_wdata;
  reg ram_w8_l2048_id9_3_1_wenable;

  ram_w8_l2048_id9_3
  inst_ram_w8_l2048_id9_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id9_3_0_addr(ram_w8_l2048_id9_3_0_addr),
    .ram_w8_l2048_id9_3_0_rdata(ram_w8_l2048_id9_3_0_rdata),
    .ram_w8_l2048_id9_3_0_wdata(ram_w8_l2048_id9_3_0_wdata),
    .ram_w8_l2048_id9_3_0_wenable(ram_w8_l2048_id9_3_0_wenable),
    .ram_w8_l2048_id9_3_1_addr(ram_w8_l2048_id9_3_1_addr),
    .ram_w8_l2048_id9_3_1_rdata(ram_w8_l2048_id9_3_1_rdata),
    .ram_w8_l2048_id9_3_1_wdata(ram_w8_l2048_id9_3_1_wdata),
    .ram_w8_l2048_id9_3_1_wenable(ram_w8_l2048_id9_3_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id10_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id10_0_0_rdata;
  reg [8-1:0] ram_w8_l2048_id10_0_0_wdata;
  reg ram_w8_l2048_id10_0_0_wenable;
  reg [9-1:0] ram_w8_l2048_id10_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id10_0_1_rdata;
  reg [8-1:0] ram_w8_l2048_id10_0_1_wdata;
  reg ram_w8_l2048_id10_0_1_wenable;

  ram_w8_l2048_id10_0
  inst_ram_w8_l2048_id10_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id10_0_0_addr(ram_w8_l2048_id10_0_0_addr),
    .ram_w8_l2048_id10_0_0_rdata(ram_w8_l2048_id10_0_0_rdata),
    .ram_w8_l2048_id10_0_0_wdata(ram_w8_l2048_id10_0_0_wdata),
    .ram_w8_l2048_id10_0_0_wenable(ram_w8_l2048_id10_0_0_wenable),
    .ram_w8_l2048_id10_0_1_addr(ram_w8_l2048_id10_0_1_addr),
    .ram_w8_l2048_id10_0_1_rdata(ram_w8_l2048_id10_0_1_rdata),
    .ram_w8_l2048_id10_0_1_wdata(ram_w8_l2048_id10_0_1_wdata),
    .ram_w8_l2048_id10_0_1_wenable(ram_w8_l2048_id10_0_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id10_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id10_1_0_rdata;
  reg [8-1:0] ram_w8_l2048_id10_1_0_wdata;
  reg ram_w8_l2048_id10_1_0_wenable;
  reg [9-1:0] ram_w8_l2048_id10_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id10_1_1_rdata;
  reg [8-1:0] ram_w8_l2048_id10_1_1_wdata;
  reg ram_w8_l2048_id10_1_1_wenable;

  ram_w8_l2048_id10_1
  inst_ram_w8_l2048_id10_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id10_1_0_addr(ram_w8_l2048_id10_1_0_addr),
    .ram_w8_l2048_id10_1_0_rdata(ram_w8_l2048_id10_1_0_rdata),
    .ram_w8_l2048_id10_1_0_wdata(ram_w8_l2048_id10_1_0_wdata),
    .ram_w8_l2048_id10_1_0_wenable(ram_w8_l2048_id10_1_0_wenable),
    .ram_w8_l2048_id10_1_1_addr(ram_w8_l2048_id10_1_1_addr),
    .ram_w8_l2048_id10_1_1_rdata(ram_w8_l2048_id10_1_1_rdata),
    .ram_w8_l2048_id10_1_1_wdata(ram_w8_l2048_id10_1_1_wdata),
    .ram_w8_l2048_id10_1_1_wenable(ram_w8_l2048_id10_1_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id10_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id10_2_0_rdata;
  reg [8-1:0] ram_w8_l2048_id10_2_0_wdata;
  reg ram_w8_l2048_id10_2_0_wenable;
  reg [9-1:0] ram_w8_l2048_id10_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id10_2_1_rdata;
  reg [8-1:0] ram_w8_l2048_id10_2_1_wdata;
  reg ram_w8_l2048_id10_2_1_wenable;

  ram_w8_l2048_id10_2
  inst_ram_w8_l2048_id10_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id10_2_0_addr(ram_w8_l2048_id10_2_0_addr),
    .ram_w8_l2048_id10_2_0_rdata(ram_w8_l2048_id10_2_0_rdata),
    .ram_w8_l2048_id10_2_0_wdata(ram_w8_l2048_id10_2_0_wdata),
    .ram_w8_l2048_id10_2_0_wenable(ram_w8_l2048_id10_2_0_wenable),
    .ram_w8_l2048_id10_2_1_addr(ram_w8_l2048_id10_2_1_addr),
    .ram_w8_l2048_id10_2_1_rdata(ram_w8_l2048_id10_2_1_rdata),
    .ram_w8_l2048_id10_2_1_wdata(ram_w8_l2048_id10_2_1_wdata),
    .ram_w8_l2048_id10_2_1_wenable(ram_w8_l2048_id10_2_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id10_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id10_3_0_rdata;
  reg [8-1:0] ram_w8_l2048_id10_3_0_wdata;
  reg ram_w8_l2048_id10_3_0_wenable;
  reg [9-1:0] ram_w8_l2048_id10_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id10_3_1_rdata;
  reg [8-1:0] ram_w8_l2048_id10_3_1_wdata;
  reg ram_w8_l2048_id10_3_1_wenable;

  ram_w8_l2048_id10_3
  inst_ram_w8_l2048_id10_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id10_3_0_addr(ram_w8_l2048_id10_3_0_addr),
    .ram_w8_l2048_id10_3_0_rdata(ram_w8_l2048_id10_3_0_rdata),
    .ram_w8_l2048_id10_3_0_wdata(ram_w8_l2048_id10_3_0_wdata),
    .ram_w8_l2048_id10_3_0_wenable(ram_w8_l2048_id10_3_0_wenable),
    .ram_w8_l2048_id10_3_1_addr(ram_w8_l2048_id10_3_1_addr),
    .ram_w8_l2048_id10_3_1_rdata(ram_w8_l2048_id10_3_1_rdata),
    .ram_w8_l2048_id10_3_1_wdata(ram_w8_l2048_id10_3_1_wdata),
    .ram_w8_l2048_id10_3_1_wenable(ram_w8_l2048_id10_3_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id11_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id11_0_0_rdata;
  reg [8-1:0] ram_w8_l2048_id11_0_0_wdata;
  reg ram_w8_l2048_id11_0_0_wenable;
  reg [9-1:0] ram_w8_l2048_id11_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id11_0_1_rdata;
  reg [8-1:0] ram_w8_l2048_id11_0_1_wdata;
  reg ram_w8_l2048_id11_0_1_wenable;

  ram_w8_l2048_id11_0
  inst_ram_w8_l2048_id11_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id11_0_0_addr(ram_w8_l2048_id11_0_0_addr),
    .ram_w8_l2048_id11_0_0_rdata(ram_w8_l2048_id11_0_0_rdata),
    .ram_w8_l2048_id11_0_0_wdata(ram_w8_l2048_id11_0_0_wdata),
    .ram_w8_l2048_id11_0_0_wenable(ram_w8_l2048_id11_0_0_wenable),
    .ram_w8_l2048_id11_0_1_addr(ram_w8_l2048_id11_0_1_addr),
    .ram_w8_l2048_id11_0_1_rdata(ram_w8_l2048_id11_0_1_rdata),
    .ram_w8_l2048_id11_0_1_wdata(ram_w8_l2048_id11_0_1_wdata),
    .ram_w8_l2048_id11_0_1_wenable(ram_w8_l2048_id11_0_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id11_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id11_1_0_rdata;
  reg [8-1:0] ram_w8_l2048_id11_1_0_wdata;
  reg ram_w8_l2048_id11_1_0_wenable;
  reg [9-1:0] ram_w8_l2048_id11_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id11_1_1_rdata;
  reg [8-1:0] ram_w8_l2048_id11_1_1_wdata;
  reg ram_w8_l2048_id11_1_1_wenable;

  ram_w8_l2048_id11_1
  inst_ram_w8_l2048_id11_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id11_1_0_addr(ram_w8_l2048_id11_1_0_addr),
    .ram_w8_l2048_id11_1_0_rdata(ram_w8_l2048_id11_1_0_rdata),
    .ram_w8_l2048_id11_1_0_wdata(ram_w8_l2048_id11_1_0_wdata),
    .ram_w8_l2048_id11_1_0_wenable(ram_w8_l2048_id11_1_0_wenable),
    .ram_w8_l2048_id11_1_1_addr(ram_w8_l2048_id11_1_1_addr),
    .ram_w8_l2048_id11_1_1_rdata(ram_w8_l2048_id11_1_1_rdata),
    .ram_w8_l2048_id11_1_1_wdata(ram_w8_l2048_id11_1_1_wdata),
    .ram_w8_l2048_id11_1_1_wenable(ram_w8_l2048_id11_1_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id11_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id11_2_0_rdata;
  reg [8-1:0] ram_w8_l2048_id11_2_0_wdata;
  reg ram_w8_l2048_id11_2_0_wenable;
  reg [9-1:0] ram_w8_l2048_id11_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id11_2_1_rdata;
  reg [8-1:0] ram_w8_l2048_id11_2_1_wdata;
  reg ram_w8_l2048_id11_2_1_wenable;

  ram_w8_l2048_id11_2
  inst_ram_w8_l2048_id11_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id11_2_0_addr(ram_w8_l2048_id11_2_0_addr),
    .ram_w8_l2048_id11_2_0_rdata(ram_w8_l2048_id11_2_0_rdata),
    .ram_w8_l2048_id11_2_0_wdata(ram_w8_l2048_id11_2_0_wdata),
    .ram_w8_l2048_id11_2_0_wenable(ram_w8_l2048_id11_2_0_wenable),
    .ram_w8_l2048_id11_2_1_addr(ram_w8_l2048_id11_2_1_addr),
    .ram_w8_l2048_id11_2_1_rdata(ram_w8_l2048_id11_2_1_rdata),
    .ram_w8_l2048_id11_2_1_wdata(ram_w8_l2048_id11_2_1_wdata),
    .ram_w8_l2048_id11_2_1_wenable(ram_w8_l2048_id11_2_1_wenable)
  );

  reg [9-1:0] ram_w8_l2048_id11_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id11_3_0_rdata;
  reg [8-1:0] ram_w8_l2048_id11_3_0_wdata;
  reg ram_w8_l2048_id11_3_0_wenable;
  reg [9-1:0] ram_w8_l2048_id11_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id11_3_1_rdata;
  reg [8-1:0] ram_w8_l2048_id11_3_1_wdata;
  reg ram_w8_l2048_id11_3_1_wenable;

  ram_w8_l2048_id11_3
  inst_ram_w8_l2048_id11_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id11_3_0_addr(ram_w8_l2048_id11_3_0_addr),
    .ram_w8_l2048_id11_3_0_rdata(ram_w8_l2048_id11_3_0_rdata),
    .ram_w8_l2048_id11_3_0_wdata(ram_w8_l2048_id11_3_0_wdata),
    .ram_w8_l2048_id11_3_0_wenable(ram_w8_l2048_id11_3_0_wenable),
    .ram_w8_l2048_id11_3_1_addr(ram_w8_l2048_id11_3_1_addr),
    .ram_w8_l2048_id11_3_1_rdata(ram_w8_l2048_id11_3_1_rdata),
    .ram_w8_l2048_id11_3_1_wdata(ram_w8_l2048_id11_3_1_wdata),
    .ram_w8_l2048_id11_3_1_wenable(ram_w8_l2048_id11_3_1_wenable)
  );

  wire [6-1:0] cparam_conv2d_16_act_num_col;
  wire [6-1:0] cparam_conv2d_16_act_num_row;
  wire [7-1:0] cparam_conv2d_16_filter_num_och;
  wire [1-1:0] cparam_conv2d_16_bias_scala;
  wire [7-1:0] cparam_conv2d_16_bias_num;
  wire [1-1:0] cparam_conv2d_16_scale_scala;
  wire [1-1:0] cparam_conv2d_16_scale_num;
  wire [1-1:0] cparam_conv2d_16_vshamt_mul_scala;
  wire [1-1:0] cparam_conv2d_16_vshamt_mul_num;
  wire [1-1:0] cparam_conv2d_16_vshamt_sum_scala;
  wire [1-1:0] cparam_conv2d_16_vshamt_sum_num;
  wire [1-1:0] cparam_conv2d_16_vshamt_out_scala;
  wire [1-1:0] cparam_conv2d_16_vshamt_out_num;
  wire [1-1:0] cparam_conv2d_16_cshamt_mul_value;
  wire [1-1:0] cparam_conv2d_16_cshamt_sum_value;
  wire [4-1:0] cparam_conv2d_16_cshamt_out_value;
  wire [1-1:0] cparam_conv2d_16_act_func_index;
  wire [6-1:0] cparam_conv2d_16_out_num_col;
  wire [6-1:0] cparam_conv2d_16_out_num_row;
  wire [1-1:0] cparam_conv2d_16_pad_col_left;
  wire [1-1:0] cparam_conv2d_16_pad_row_top;
  wire [5-1:0] cparam_conv2d_16_max_col_count;
  wire [5-1:0] cparam_conv2d_16_max_row_count;
  wire [1-1:0] cparam_conv2d_16_max_bat_count;
  wire [1-1:0] cparam_conv2d_16_max_och_count;
  wire [8-1:0] cparam_conv2d_16_och_count_step;
  wire [1-1:0] cparam_conv2d_16_dma_flag_conds_0;
  wire [1-1:0] cparam_conv2d_16_dma_flag_conds_1;
  wire [1-1:0] cparam_conv2d_16_dma_flag_conds_2;
  wire signed [32-1:0] cparam_conv2d_16_act_offset_values_0;
  wire signed [32-1:0] cparam_conv2d_16_act_offset_values_1;
  wire signed [32-1:0] cparam_conv2d_16_act_offset_values_2;
  wire [9-1:0] cparam_conv2d_16_act_row_step;
  wire [13-1:0] cparam_conv2d_16_act_bat_step;
  wire [9-1:0] cparam_conv2d_16_act_read_size;
  wire [6-1:0] cparam_conv2d_16_act_read_block;
  wire [7-1:0] cparam_conv2d_16_act_read_step;
  wire [14-1:0] cparam_conv2d_16_filter_base_step;
  wire [15-1:0] cparam_conv2d_16_filter_read_size;
  wire [6-1:0] cparam_conv2d_16_filter_read_block;
  wire [12-1:0] cparam_conv2d_16_filter_read_step;
  wire [1-1:0] cparam_conv2d_16_out_offset_values_0;
  wire [7-1:0] cparam_conv2d_16_out_col_step;
  wire [10-1:0] cparam_conv2d_16_out_row_step;
  wire [15-1:0] cparam_conv2d_16_out_bat_step;
  wire [7-1:0] cparam_conv2d_16_out_och_step;
  wire [10-1:0] cparam_conv2d_16_out_write_size;
  wire [10-1:0] cparam_conv2d_16_out_write_size_res;
  wire [7-1:0] cparam_conv2d_16_out_write_block;
  wire [1-1:0] cparam_conv2d_16_keep_filter;
  wire [1-1:0] cparam_conv2d_16_keep_input;
  wire [1-1:0] cparam_conv2d_16_data_stationary;
  wire [7-1:0] cparam_conv2d_16_stream_num_ops;
  wire [7-1:0] cparam_conv2d_16_stream_num_ops_res;
  wire [7-1:0] cparam_conv2d_16_stream_num_ops_par;
  wire [7-1:0] cparam_conv2d_16_stream_num_ops_res_par;
  wire [6-1:0] cparam_conv2d_16_stream_reduce_size;
  wire [6-1:0] cparam_conv2d_16_stream_aligned_reduce_size;
  wire [1-1:0] cparam_conv2d_16_stream_omit_mask;
  wire [2-1:0] cparam_conv2d_16_col_select_initval;
  wire [1-1:0] cparam_conv2d_16_stride_col_par_col;
  wire [1-1:0] cparam_conv2d_16_stride_row_par_row;
  wire [1-1:0] cparam_conv2d_16_stride_col_mod_filter_num;
  wire [2-1:0] cparam_conv2d_16_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_0;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_1;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_2;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_3;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_4;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_5;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_6;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_7;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_8;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_9;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_10;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_11;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_12;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_13;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_14;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_15;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_16;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_17;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_18;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_19;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_20;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_21;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_22;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_23;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_24;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_25;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_conds_26;
  wire [1-1:0] cparam_conv2d_16_inc_act_laddr_small;
  wire [6-1:0] cparam_conv2d_16_inc_act_laddr_large;
  wire [7-1:0] cparam_conv2d_16_inc_out_laddr_col;
  wire [1-1:0] cparam_conv2d_16_stream_act_local_small_offset;
  wire signed [7-1:0] cparam_conv2d_16_stream_act_local_large_offset;
  wire [1-1:0] cparam_conv2d_16_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_conv2d_16_stream_act_local_small_flags_1;
  wire [1-1:0] cparam_conv2d_16_stream_act_local_small_flags_2;
  wire [1-1:0] cparam_conv2d_16_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_conv2d_16_stream_act_local_large_flags_1;
  wire [1-1:0] cparam_conv2d_16_stream_act_local_large_flags_2;
  wire [6-1:0] cparam_conv2d_16_inc_sync_out;
  wire [1-1:0] cparam_conv2d_16_inc_sync_out_res;
  reg [2-1:0] conv2d_16_control_param_index;
  assign cparam_conv2d_16_act_num_col = (conv2d_16_control_param_index == 0)? 32 : 
                                        (conv2d_16_control_param_index == 1)? 16 : 8;
  assign cparam_conv2d_16_act_num_row = (conv2d_16_control_param_index == 0)? 32 : 
                                        (conv2d_16_control_param_index == 1)? 16 : 8;
  assign cparam_conv2d_16_filter_num_och = (conv2d_16_control_param_index == 0)? 16 : 
                                           (conv2d_16_control_param_index == 1)? 32 : 64;
  assign cparam_conv2d_16_bias_scala = (conv2d_16_control_param_index == 0)? 0 : 
                                       (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_bias_num = (conv2d_16_control_param_index == 0)? 16 : 
                                     (conv2d_16_control_param_index == 1)? 32 : 64;
  assign cparam_conv2d_16_scale_scala = (conv2d_16_control_param_index == 0)? 1 : 
                                        (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_scale_num = (conv2d_16_control_param_index == 0)? 1 : 
                                      (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_vshamt_mul_scala = (conv2d_16_control_param_index == 0)? 0 : 
                                             (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_vshamt_mul_num = (conv2d_16_control_param_index == 0)? 0 : 
                                           (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_vshamt_sum_scala = (conv2d_16_control_param_index == 0)? 0 : 
                                             (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_vshamt_sum_num = (conv2d_16_control_param_index == 0)? 0 : 
                                           (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_vshamt_out_scala = (conv2d_16_control_param_index == 0)? 0 : 
                                             (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_vshamt_out_num = (conv2d_16_control_param_index == 0)? 0 : 
                                           (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_cshamt_mul_value = (conv2d_16_control_param_index == 0)? 0 : 
                                             (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_cshamt_sum_value = (conv2d_16_control_param_index == 0)? 0 : 
                                             (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_cshamt_out_value = (conv2d_16_control_param_index == 0)? 12 : 
                                             (conv2d_16_control_param_index == 1)? 10 : 11;
  assign cparam_conv2d_16_act_func_index = (conv2d_16_control_param_index == 0)? 0 : 
                                           (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_out_num_col = (conv2d_16_control_param_index == 0)? 32 : 
                                        (conv2d_16_control_param_index == 1)? 16 : 8;
  assign cparam_conv2d_16_out_num_row = (conv2d_16_control_param_index == 0)? 32 : 
                                        (conv2d_16_control_param_index == 1)? 16 : 8;
  assign cparam_conv2d_16_pad_col_left = (conv2d_16_control_param_index == 0)? 1 : 
                                         (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_pad_row_top = (conv2d_16_control_param_index == 0)? 1 : 
                                        (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_max_col_count = (conv2d_16_control_param_index == 0)? 31 : 
                                          (conv2d_16_control_param_index == 1)? 15 : 7;
  assign cparam_conv2d_16_max_row_count = (conv2d_16_control_param_index == 0)? 31 : 
                                          (conv2d_16_control_param_index == 1)? 15 : 7;
  assign cparam_conv2d_16_max_bat_count = (conv2d_16_control_param_index == 0)? 0 : 
                                          (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_max_och_count = (conv2d_16_control_param_index == 0)? 0 : 
                                          (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_och_count_step = (conv2d_16_control_param_index == 0)? 32 : 
                                           (conv2d_16_control_param_index == 1)? 64 : 128;
  assign cparam_conv2d_16_dma_flag_conds_0 = (conv2d_16_control_param_index == 0)? 1 : 
                                             (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_dma_flag_conds_1 = (conv2d_16_control_param_index == 0)? 0 : 
                                             (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_dma_flag_conds_2 = (conv2d_16_control_param_index == 0)? 0 : 
                                             (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_act_offset_values_0 = (conv2d_16_control_param_index == 0)? -128 : 
                                                (conv2d_16_control_param_index == 1)? -256 : -256;
  assign cparam_conv2d_16_act_offset_values_1 = (conv2d_16_control_param_index == 0)? 0 : 
                                                (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_act_offset_values_2 = (conv2d_16_control_param_index == 0)? 128 : 
                                                (conv2d_16_control_param_index == 1)? 256 : 256;
  assign cparam_conv2d_16_act_row_step = (conv2d_16_control_param_index == 0)? 128 : 
                                         (conv2d_16_control_param_index == 1)? 256 : 256;
  assign cparam_conv2d_16_act_bat_step = (conv2d_16_control_param_index == 0)? 4096 : 
                                         (conv2d_16_control_param_index == 1)? 4096 : 2048;
  assign cparam_conv2d_16_act_read_size = (conv2d_16_control_param_index == 0)? 128 : 
                                          (conv2d_16_control_param_index == 1)? 256 : 256;
  assign cparam_conv2d_16_act_read_block = (conv2d_16_control_param_index == 0)? 4 : 
                                           (conv2d_16_control_param_index == 1)? 16 : 32;
  assign cparam_conv2d_16_act_read_step = (conv2d_16_control_param_index == 0)? 44 : 
                                          (conv2d_16_control_param_index == 1)? 96 : 96;
  assign cparam_conv2d_16_filter_base_step = (conv2d_16_control_param_index == 0)? 576 : 
                                             (conv2d_16_control_param_index == 1)? 2304 : 9216;
  assign cparam_conv2d_16_filter_read_size = (conv2d_16_control_param_index == 0)? 1152 : 
                                             (conv2d_16_control_param_index == 1)? 4608 : 18432;
  assign cparam_conv2d_16_filter_read_block = (conv2d_16_control_param_index == 0)? 8 : 
                                              (conv2d_16_control_param_index == 1)? 16 : 32;
  assign cparam_conv2d_16_filter_read_step = (conv2d_16_control_param_index == 0)? 128 : 
                                             (conv2d_16_control_param_index == 1)? 512 : 2048;
  assign cparam_conv2d_16_out_offset_values_0 = (conv2d_16_control_param_index == 0)? 0 : 
                                                (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_out_col_step = (conv2d_16_control_param_index == 0)? 16 : 
                                         (conv2d_16_control_param_index == 1)? 32 : 64;
  assign cparam_conv2d_16_out_row_step = (conv2d_16_control_param_index == 0)? 512 : 
                                         (conv2d_16_control_param_index == 1)? 512 : 512;
  assign cparam_conv2d_16_out_bat_step = (conv2d_16_control_param_index == 0)? 16384 : 
                                         (conv2d_16_control_param_index == 1)? 8192 : 4096;
  assign cparam_conv2d_16_out_och_step = (conv2d_16_control_param_index == 0)? 16 : 
                                         (conv2d_16_control_param_index == 1)? 32 : 64;
  assign cparam_conv2d_16_out_write_size = (conv2d_16_control_param_index == 0)? 512 : 
                                           (conv2d_16_control_param_index == 1)? 512 : 512;
  assign cparam_conv2d_16_out_write_size_res = (conv2d_16_control_param_index == 0)? 512 : 
                                               (conv2d_16_control_param_index == 1)? 512 : 512;
  assign cparam_conv2d_16_out_write_block = (conv2d_16_control_param_index == 0)? 16 : 
                                            (conv2d_16_control_param_index == 1)? 32 : 64;
  assign cparam_conv2d_16_keep_filter = (conv2d_16_control_param_index == 0)? 1 : 
                                        (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_keep_input = (conv2d_16_control_param_index == 0)? 1 : 
                                       (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_data_stationary = (conv2d_16_control_param_index == 0)? 0 : 
                                            (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_stream_num_ops = (conv2d_16_control_param_index == 0)? 16 : 
                                           (conv2d_16_control_param_index == 1)? 32 : 64;
  assign cparam_conv2d_16_stream_num_ops_res = (conv2d_16_control_param_index == 0)? 16 : 
                                               (conv2d_16_control_param_index == 1)? 32 : 64;
  assign cparam_conv2d_16_stream_num_ops_par = (conv2d_16_control_param_index == 0)? 16 : 
                                               (conv2d_16_control_param_index == 1)? 32 : 64;
  assign cparam_conv2d_16_stream_num_ops_res_par = (conv2d_16_control_param_index == 0)? 16 : 
                                                   (conv2d_16_control_param_index == 1)? 32 : 64;
  assign cparam_conv2d_16_stream_reduce_size = (conv2d_16_control_param_index == 0)? 3 : 
                                               (conv2d_16_control_param_index == 1)? 16 : 32;
  assign cparam_conv2d_16_stream_aligned_reduce_size = (conv2d_16_control_param_index == 0)? 8 : 
                                                       (conv2d_16_control_param_index == 1)? 16 : 32;
  assign cparam_conv2d_16_stream_omit_mask = (conv2d_16_control_param_index == 0)? 0 : 
                                             (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_col_select_initval = (conv2d_16_control_param_index == 0)? 2 : 
                                               (conv2d_16_control_param_index == 1)? 2 : 2;
  assign cparam_conv2d_16_stride_col_par_col = (conv2d_16_control_param_index == 0)? 1 : 
                                               (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_stride_row_par_row = (conv2d_16_control_param_index == 0)? 1 : 
                                               (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_stride_col_mod_filter_num = (conv2d_16_control_param_index == 0)? 1 : 
                                                      (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_filter_num_col_minus_stride_col_mod = (conv2d_16_control_param_index == 0)? 2 : 
                                                                (conv2d_16_control_param_index == 1)? 2 : 2;
  assign cparam_conv2d_16_inc_act_laddr_conds_0 = (conv2d_16_control_param_index == 0)? 1 : 
                                                  (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_inc_act_laddr_conds_1 = (conv2d_16_control_param_index == 0)? 0 : 
                                                  (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_2 = (conv2d_16_control_param_index == 0)? 0 : 
                                                  (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_3 = (conv2d_16_control_param_index == 0)? 0 : 
                                                  (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_4 = (conv2d_16_control_param_index == 0)? 1 : 
                                                  (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_inc_act_laddr_conds_5 = (conv2d_16_control_param_index == 0)? 0 : 
                                                  (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_6 = (conv2d_16_control_param_index == 0)? 0 : 
                                                  (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_7 = (conv2d_16_control_param_index == 0)? 0 : 
                                                  (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_8 = (conv2d_16_control_param_index == 0)? 1 : 
                                                  (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_inc_act_laddr_conds_9 = (conv2d_16_control_param_index == 0)? 1 : 
                                                  (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_inc_act_laddr_conds_10 = (conv2d_16_control_param_index == 0)? 0 : 
                                                   (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_11 = (conv2d_16_control_param_index == 0)? 0 : 
                                                   (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_12 = (conv2d_16_control_param_index == 0)? 0 : 
                                                   (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_13 = (conv2d_16_control_param_index == 0)? 1 : 
                                                   (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_inc_act_laddr_conds_14 = (conv2d_16_control_param_index == 0)? 0 : 
                                                   (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_15 = (conv2d_16_control_param_index == 0)? 0 : 
                                                   (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_16 = (conv2d_16_control_param_index == 0)? 0 : 
                                                   (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_17 = (conv2d_16_control_param_index == 0)? 1 : 
                                                   (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_inc_act_laddr_conds_18 = (conv2d_16_control_param_index == 0)? 1 : 
                                                   (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_inc_act_laddr_conds_19 = (conv2d_16_control_param_index == 0)? 0 : 
                                                   (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_20 = (conv2d_16_control_param_index == 0)? 0 : 
                                                   (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_21 = (conv2d_16_control_param_index == 0)? 0 : 
                                                   (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_22 = (conv2d_16_control_param_index == 0)? 1 : 
                                                   (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_inc_act_laddr_conds_23 = (conv2d_16_control_param_index == 0)? 0 : 
                                                   (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_24 = (conv2d_16_control_param_index == 0)? 0 : 
                                                   (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_25 = (conv2d_16_control_param_index == 0)? 0 : 
                                                   (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_conds_26 = (conv2d_16_control_param_index == 0)? 1 : 
                                                   (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_inc_act_laddr_small = (conv2d_16_control_param_index == 0)? 0 : 
                                                (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_inc_act_laddr_large = (conv2d_16_control_param_index == 0)? 4 : 
                                                (conv2d_16_control_param_index == 1)? 16 : 32;
  assign cparam_conv2d_16_inc_out_laddr_col = (conv2d_16_control_param_index == 0)? 16 : 
                                              (conv2d_16_control_param_index == 1)? 32 : 64;
  assign cparam_conv2d_16_stream_act_local_small_offset = (conv2d_16_control_param_index == 0)? 0 : 
                                                          (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_stream_act_local_large_offset = (conv2d_16_control_param_index == 0)? -4 : 
                                                          (conv2d_16_control_param_index == 1)? -16 : -32;
  assign cparam_conv2d_16_stream_act_local_small_flags_0 = (conv2d_16_control_param_index == 0)? 0 : 
                                                           (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_stream_act_local_small_flags_1 = (conv2d_16_control_param_index == 0)? 0 : 
                                                           (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_stream_act_local_small_flags_2 = (conv2d_16_control_param_index == 0)? 1 : 
                                                           (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_stream_act_local_large_flags_0 = (conv2d_16_control_param_index == 0)? 0 : 
                                                           (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_stream_act_local_large_flags_1 = (conv2d_16_control_param_index == 0)? 0 : 
                                                           (conv2d_16_control_param_index == 1)? 0 : 0;
  assign cparam_conv2d_16_stream_act_local_large_flags_2 = (conv2d_16_control_param_index == 0)? 1 : 
                                                           (conv2d_16_control_param_index == 1)? 1 : 1;
  assign cparam_conv2d_16_inc_sync_out = (conv2d_16_control_param_index == 0)? 32 : 
                                         (conv2d_16_control_param_index == 1)? 16 : 8;
  assign cparam_conv2d_16_inc_sync_out_res = (conv2d_16_control_param_index == 0)? 0 : 
                                             (conv2d_16_control_param_index == 1)? 0 : 0;
  wire [6-1:0] cparam_max_pool_serial_18_act_num_col;
  wire [6-1:0] cparam_max_pool_serial_18_act_num_row;
  wire [2-1:0] cparam_max_pool_serial_18_stride_col;
  wire [2-1:0] cparam_max_pool_serial_18_stride_row;
  wire [5-1:0] cparam_max_pool_serial_18_out_num_col;
  wire [5-1:0] cparam_max_pool_serial_18_out_num_row;
  wire [1-1:0] cparam_max_pool_serial_18_pad_col_left;
  wire [1-1:0] cparam_max_pool_serial_18_pad_row_top;
  wire [5-1:0] cparam_max_pool_serial_18_max_col_count;
  wire [5-1:0] cparam_max_pool_serial_18_max_row_count;
  wire [1-1:0] cparam_max_pool_serial_18_max_bat_count;
  wire signed [32-1:0] cparam_max_pool_serial_18_act_offset_values_0;
  wire signed [32-1:0] cparam_max_pool_serial_18_act_offset_values_1;
  wire [11-1:0] cparam_max_pool_serial_18_act_row_step;
  wire [15-1:0] cparam_max_pool_serial_18_act_bat_step;
  wire [10-1:0] cparam_max_pool_serial_18_act_read_size;
  wire [7-1:0] cparam_max_pool_serial_18_act_read_block;
  wire [9-1:0] cparam_max_pool_serial_18_out_row_step;
  wire [13-1:0] cparam_max_pool_serial_18_out_bat_step;
  wire [9-1:0] cparam_max_pool_serial_18_out_write_size;
  wire [7-1:0] cparam_max_pool_serial_18_stream_size;
  wire [1-1:0] cparam_max_pool_serial_18_col_select_initval;
  wire [1-1:0] cparam_max_pool_serial_18_stride_col_mod_ksize;
  wire [2-1:0] cparam_max_pool_serial_18_ksize_col_minus_stride_col_mod;
  wire [1-1:0] cparam_max_pool_serial_18_local_pad_offset;
  wire [8-1:0] cparam_max_pool_serial_18_inc_act_laddr;
  wire [7-1:0] cparam_max_pool_serial_18_inc_out_laddr;
  reg [2-1:0] max_pool_serial_18_control_param_index;
  assign cparam_max_pool_serial_18_act_num_col = (max_pool_serial_18_control_param_index == 0)? 32 : 
                                                 (max_pool_serial_18_control_param_index == 1)? 16 : 8;
  assign cparam_max_pool_serial_18_act_num_row = (max_pool_serial_18_control_param_index == 0)? 32 : 
                                                 (max_pool_serial_18_control_param_index == 1)? 16 : 8;
  assign cparam_max_pool_serial_18_stride_col = (max_pool_serial_18_control_param_index == 0)? 2 : 
                                                (max_pool_serial_18_control_param_index == 1)? 2 : 2;
  assign cparam_max_pool_serial_18_stride_row = (max_pool_serial_18_control_param_index == 0)? 2 : 
                                                (max_pool_serial_18_control_param_index == 1)? 2 : 2;
  assign cparam_max_pool_serial_18_out_num_col = (max_pool_serial_18_control_param_index == 0)? 16 : 
                                                 (max_pool_serial_18_control_param_index == 1)? 8 : 4;
  assign cparam_max_pool_serial_18_out_num_row = (max_pool_serial_18_control_param_index == 0)? 16 : 
                                                 (max_pool_serial_18_control_param_index == 1)? 8 : 4;
  assign cparam_max_pool_serial_18_pad_col_left = (max_pool_serial_18_control_param_index == 0)? 0 : 
                                                  (max_pool_serial_18_control_param_index == 1)? 0 : 0;
  assign cparam_max_pool_serial_18_pad_row_top = (max_pool_serial_18_control_param_index == 0)? 0 : 
                                                 (max_pool_serial_18_control_param_index == 1)? 0 : 0;
  assign cparam_max_pool_serial_18_max_col_count = (max_pool_serial_18_control_param_index == 0)? 29 : 
                                                   (max_pool_serial_18_control_param_index == 1)? 13 : 5;
  assign cparam_max_pool_serial_18_max_row_count = (max_pool_serial_18_control_param_index == 0)? 29 : 
                                                   (max_pool_serial_18_control_param_index == 1)? 13 : 5;
  assign cparam_max_pool_serial_18_max_bat_count = (max_pool_serial_18_control_param_index == 0)? 0 : 
                                                   (max_pool_serial_18_control_param_index == 1)? 0 : 0;
  assign cparam_max_pool_serial_18_act_offset_values_0 = (max_pool_serial_18_control_param_index == 0)? 0 : 
                                                         (max_pool_serial_18_control_param_index == 1)? 0 : 0;
  assign cparam_max_pool_serial_18_act_offset_values_1 = (max_pool_serial_18_control_param_index == 0)? 512 : 
                                                         (max_pool_serial_18_control_param_index == 1)? 512 : 512;
  assign cparam_max_pool_serial_18_act_row_step = (max_pool_serial_18_control_param_index == 0)? 1024 : 
                                                  (max_pool_serial_18_control_param_index == 1)? 1024 : 1024;
  assign cparam_max_pool_serial_18_act_bat_step = (max_pool_serial_18_control_param_index == 0)? 16384 : 
                                                  (max_pool_serial_18_control_param_index == 1)? 8192 : 4096;
  assign cparam_max_pool_serial_18_act_read_size = (max_pool_serial_18_control_param_index == 0)? 512 : 
                                                   (max_pool_serial_18_control_param_index == 1)? 512 : 512;
  assign cparam_max_pool_serial_18_act_read_block = (max_pool_serial_18_control_param_index == 0)? 16 : 
                                                    (max_pool_serial_18_control_param_index == 1)? 32 : 64;
  assign cparam_max_pool_serial_18_out_row_step = (max_pool_serial_18_control_param_index == 0)? 256 : 
                                                  (max_pool_serial_18_control_param_index == 1)? 256 : 256;
  assign cparam_max_pool_serial_18_out_bat_step = (max_pool_serial_18_control_param_index == 0)? 4096 : 
                                                  (max_pool_serial_18_control_param_index == 1)? 2048 : 1024;
  assign cparam_max_pool_serial_18_out_write_size = (max_pool_serial_18_control_param_index == 0)? 256 : 
                                                    (max_pool_serial_18_control_param_index == 1)? 256 : 256;
  assign cparam_max_pool_serial_18_stream_size = (max_pool_serial_18_control_param_index == 0)? 16 : 
                                                 (max_pool_serial_18_control_param_index == 1)? 32 : 64;
  assign cparam_max_pool_serial_18_col_select_initval = (max_pool_serial_18_control_param_index == 0)? 0 : 
                                                        (max_pool_serial_18_control_param_index == 1)? 0 : 0;
  assign cparam_max_pool_serial_18_stride_col_mod_ksize = (max_pool_serial_18_control_param_index == 0)? 0 : 
                                                          (max_pool_serial_18_control_param_index == 1)? 0 : 0;
  assign cparam_max_pool_serial_18_ksize_col_minus_stride_col_mod = (max_pool_serial_18_control_param_index == 0)? 2 : 
                                                                    (max_pool_serial_18_control_param_index == 1)? 2 : 2;
  assign cparam_max_pool_serial_18_local_pad_offset = (max_pool_serial_18_control_param_index == 0)? 0 : 
                                                      (max_pool_serial_18_control_param_index == 1)? 0 : 0;
  assign cparam_max_pool_serial_18_inc_act_laddr = (max_pool_serial_18_control_param_index == 0)? 32 : 
                                                   (max_pool_serial_18_control_param_index == 1)? 64 : 128;
  assign cparam_max_pool_serial_18_inc_out_laddr = (max_pool_serial_18_control_param_index == 0)? 16 : 
                                                   (max_pool_serial_18_control_param_index == 1)? 32 : 64;
  wire [1-1:0] cparam_matmul_29_act_num_col;
  wire [1-1:0] cparam_matmul_29_act_num_row;
  wire [9-1:0] cparam_matmul_29_filter_num_och;
  wire [1-1:0] cparam_matmul_29_bias_scala;
  wire [9-1:0] cparam_matmul_29_bias_num;
  wire [1-1:0] cparam_matmul_29_scale_scala;
  wire [1-1:0] cparam_matmul_29_scale_num;
  wire [1-1:0] cparam_matmul_29_vshamt_mul_scala;
  wire [1-1:0] cparam_matmul_29_vshamt_mul_num;
  wire [1-1:0] cparam_matmul_29_vshamt_sum_scala;
  wire [1-1:0] cparam_matmul_29_vshamt_sum_num;
  wire [1-1:0] cparam_matmul_29_vshamt_out_scala;
  wire [1-1:0] cparam_matmul_29_vshamt_out_num;
  wire [1-1:0] cparam_matmul_29_cshamt_mul_value;
  wire [1-1:0] cparam_matmul_29_cshamt_sum_value;
  wire [4-1:0] cparam_matmul_29_cshamt_out_value;
  wire [1-1:0] cparam_matmul_29_act_func_index;
  wire [1-1:0] cparam_matmul_29_out_num_col;
  wire [1-1:0] cparam_matmul_29_out_num_row;
  wire [1-1:0] cparam_matmul_29_pad_col_left;
  wire [1-1:0] cparam_matmul_29_pad_row_top;
  wire [1-1:0] cparam_matmul_29_max_col_count;
  wire [1-1:0] cparam_matmul_29_max_row_count;
  wire [1-1:0] cparam_matmul_29_max_bat_count;
  wire [8-1:0] cparam_matmul_29_max_och_count;
  wire [6-1:0] cparam_matmul_29_och_count_step;
  wire [1-1:0] cparam_matmul_29_dma_flag_conds_0;
  wire signed [32-1:0] cparam_matmul_29_act_offset_values_0;
  wire [11-1:0] cparam_matmul_29_act_row_step;
  wire [11-1:0] cparam_matmul_29_act_bat_step;
  wire [11-1:0] cparam_matmul_29_act_read_size;
  wire [11-1:0] cparam_matmul_29_act_read_block;
  wire [11-1:0] cparam_matmul_29_act_read_step;
  wire [12-1:0] cparam_matmul_29_filter_base_step;
  wire [13-1:0] cparam_matmul_29_filter_read_size;
  wire [11-1:0] cparam_matmul_29_filter_read_block;
  wire [13-1:0] cparam_matmul_29_filter_read_step;
  wire [1-1:0] cparam_matmul_29_out_offset_values_0;
  wire [9-1:0] cparam_matmul_29_out_col_step;
  wire [9-1:0] cparam_matmul_29_out_row_step;
  wire [9-1:0] cparam_matmul_29_out_bat_step;
  wire [5-1:0] cparam_matmul_29_out_och_step;
  wire [5-1:0] cparam_matmul_29_out_write_size;
  wire [5-1:0] cparam_matmul_29_out_write_size_res;
  wire [4-1:0] cparam_matmul_29_out_write_block;
  wire [1-1:0] cparam_matmul_29_keep_filter;
  wire [1-1:0] cparam_matmul_29_keep_input;
  wire [1-1:0] cparam_matmul_29_data_stationary;
  wire [5-1:0] cparam_matmul_29_stream_num_ops;
  wire [5-1:0] cparam_matmul_29_stream_num_ops_res;
  wire [5-1:0] cparam_matmul_29_stream_num_ops_par;
  wire [5-1:0] cparam_matmul_29_stream_num_ops_res_par;
  wire [11-1:0] cparam_matmul_29_stream_reduce_size;
  wire [11-1:0] cparam_matmul_29_stream_aligned_reduce_size;
  wire [1-1:0] cparam_matmul_29_stream_omit_mask;
  wire [1-1:0] cparam_matmul_29_col_select_initval;
  wire [1-1:0] cparam_matmul_29_stride_col_par_col;
  wire [1-1:0] cparam_matmul_29_stride_row_par_row;
  wire [1-1:0] cparam_matmul_29_stride_col_mod_filter_num;
  wire [1-1:0] cparam_matmul_29_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_matmul_29_inc_act_laddr_conds_0;
  wire [11-1:0] cparam_matmul_29_inc_act_laddr_small;
  wire [11-1:0] cparam_matmul_29_inc_act_laddr_large;
  wire [9-1:0] cparam_matmul_29_inc_out_laddr_col;
  wire [1-1:0] cparam_matmul_29_stream_act_local_small_offset;
  wire [1-1:0] cparam_matmul_29_stream_act_local_large_offset;
  wire [1-1:0] cparam_matmul_29_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_matmul_29_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_matmul_29_inc_sync_out;
  wire [1-1:0] cparam_matmul_29_inc_sync_out_res;
  reg [2-1:0] matmul_29_control_param_index;
  assign cparam_matmul_29_act_num_col = (matmul_29_control_param_index == 0)? 1 : 
                                        (matmul_29_control_param_index == 1)? 1 : 1;
  assign cparam_matmul_29_act_num_row = (matmul_29_control_param_index == 0)? 1 : 
                                        (matmul_29_control_param_index == 1)? 1 : 1;
  assign cparam_matmul_29_filter_num_och = (matmul_29_control_param_index == 0)? 256 : 
                                           (matmul_29_control_param_index == 1)? 128 : 10;
  assign cparam_matmul_29_bias_scala = (matmul_29_control_param_index == 0)? 0 : 
                                       (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_bias_num = (matmul_29_control_param_index == 0)? 256 : 
                                     (matmul_29_control_param_index == 1)? 128 : 10;
  assign cparam_matmul_29_scale_scala = (matmul_29_control_param_index == 0)? 1 : 
                                        (matmul_29_control_param_index == 1)? 1 : 1;
  assign cparam_matmul_29_scale_num = (matmul_29_control_param_index == 0)? 1 : 
                                      (matmul_29_control_param_index == 1)? 1 : 1;
  assign cparam_matmul_29_vshamt_mul_scala = (matmul_29_control_param_index == 0)? 0 : 
                                             (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_vshamt_mul_num = (matmul_29_control_param_index == 0)? 0 : 
                                           (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_vshamt_sum_scala = (matmul_29_control_param_index == 0)? 0 : 
                                             (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_vshamt_sum_num = (matmul_29_control_param_index == 0)? 0 : 
                                           (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_vshamt_out_scala = (matmul_29_control_param_index == 0)? 0 : 
                                             (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_vshamt_out_num = (matmul_29_control_param_index == 0)? 0 : 
                                           (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_cshamt_mul_value = (matmul_29_control_param_index == 0)? 0 : 
                                             (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_cshamt_sum_value = (matmul_29_control_param_index == 0)? 0 : 
                                             (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_cshamt_out_value = (matmul_29_control_param_index == 0)? 12 : 
                                             (matmul_29_control_param_index == 1)? 10 : 13;
  assign cparam_matmul_29_act_func_index = (matmul_29_control_param_index == 0)? 0 : 
                                           (matmul_29_control_param_index == 1)? 0 : 1;
  assign cparam_matmul_29_out_num_col = (matmul_29_control_param_index == 0)? 1 : 
                                        (matmul_29_control_param_index == 1)? 1 : 1;
  assign cparam_matmul_29_out_num_row = (matmul_29_control_param_index == 0)? 1 : 
                                        (matmul_29_control_param_index == 1)? 1 : 1;
  assign cparam_matmul_29_pad_col_left = (matmul_29_control_param_index == 0)? 0 : 
                                         (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_pad_row_top = (matmul_29_control_param_index == 0)? 0 : 
                                        (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_max_col_count = (matmul_29_control_param_index == 0)? 0 : 
                                          (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_max_row_count = (matmul_29_control_param_index == 0)? 0 : 
                                          (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_max_bat_count = (matmul_29_control_param_index == 0)? 0 : 
                                          (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_max_och_count = (matmul_29_control_param_index == 0)? 252 : 
                                          (matmul_29_control_param_index == 1)? 112 : 0;
  assign cparam_matmul_29_och_count_step = (matmul_29_control_param_index == 0)? 4 : 
                                           (matmul_29_control_param_index == 1)? 16 : 32;
  assign cparam_matmul_29_dma_flag_conds_0 = (matmul_29_control_param_index == 0)? 1 : 
                                             (matmul_29_control_param_index == 1)? 1 : 1;
  assign cparam_matmul_29_act_offset_values_0 = (matmul_29_control_param_index == 0)? 0 : 
                                                (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_act_row_step = (matmul_29_control_param_index == 0)? 1024 : 
                                         (matmul_29_control_param_index == 1)? 256 : 128;
  assign cparam_matmul_29_act_bat_step = (matmul_29_control_param_index == 0)? 1024 : 
                                         (matmul_29_control_param_index == 1)? 256 : 128;
  assign cparam_matmul_29_act_read_size = (matmul_29_control_param_index == 0)? 1024 : 
                                          (matmul_29_control_param_index == 1)? 256 : 128;
  assign cparam_matmul_29_act_read_block = (matmul_29_control_param_index == 0)? 1024 : 
                                           (matmul_29_control_param_index == 1)? 256 : 128;
  assign cparam_matmul_29_act_read_step = (matmul_29_control_param_index == 0)? 1024 : 
                                          (matmul_29_control_param_index == 1)? 256 : 128;
  assign cparam_matmul_29_filter_base_step = (matmul_29_control_param_index == 0)? 2048 : 
                                             (matmul_29_control_param_index == 1)? 2048 : 640;
  assign cparam_matmul_29_filter_read_size = (matmul_29_control_param_index == 0)? 4096 : 
                                             (matmul_29_control_param_index == 1)? 4096 : 1280;
  assign cparam_matmul_29_filter_read_block = (matmul_29_control_param_index == 0)? 1024 : 
                                              (matmul_29_control_param_index == 1)? 256 : 128;
  assign cparam_matmul_29_filter_read_step = (matmul_29_control_param_index == 0)? 4096 : 
                                             (matmul_29_control_param_index == 1)? 4096 : 1280;
  assign cparam_matmul_29_out_offset_values_0 = (matmul_29_control_param_index == 0)? 0 : 
                                                (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_out_col_step = (matmul_29_control_param_index == 0)? 256 : 
                                         (matmul_29_control_param_index == 1)? 128 : 12;
  assign cparam_matmul_29_out_row_step = (matmul_29_control_param_index == 0)? 256 : 
                                         (matmul_29_control_param_index == 1)? 128 : 12;
  assign cparam_matmul_29_out_bat_step = (matmul_29_control_param_index == 0)? 256 : 
                                         (matmul_29_control_param_index == 1)? 128 : 12;
  assign cparam_matmul_29_out_och_step = (matmul_29_control_param_index == 0)? 4 : 
                                         (matmul_29_control_param_index == 1)? 16 : 10;
  assign cparam_matmul_29_out_write_size = (matmul_29_control_param_index == 0)? 4 : 
                                           (matmul_29_control_param_index == 1)? 16 : 12;
  assign cparam_matmul_29_out_write_size_res = (matmul_29_control_param_index == 0)? 4 : 
                                               (matmul_29_control_param_index == 1)? 16 : 12;
  assign cparam_matmul_29_out_write_block = (matmul_29_control_param_index == 0)? 0 : 
                                            (matmul_29_control_param_index == 1)? 0 : 12;
  assign cparam_matmul_29_keep_filter = (matmul_29_control_param_index == 0)? 0 : 
                                        (matmul_29_control_param_index == 1)? 0 : 1;
  assign cparam_matmul_29_keep_input = (matmul_29_control_param_index == 0)? 1 : 
                                       (matmul_29_control_param_index == 1)? 1 : 1;
  assign cparam_matmul_29_data_stationary = (matmul_29_control_param_index == 0)? 0 : 
                                            (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_stream_num_ops = (matmul_29_control_param_index == 0)? 4 : 
                                           (matmul_29_control_param_index == 1)? 16 : 12;
  assign cparam_matmul_29_stream_num_ops_res = (matmul_29_control_param_index == 0)? 4 : 
                                               (matmul_29_control_param_index == 1)? 16 : 12;
  assign cparam_matmul_29_stream_num_ops_par = (matmul_29_control_param_index == 0)? 4 : 
                                               (matmul_29_control_param_index == 1)? 16 : 12;
  assign cparam_matmul_29_stream_num_ops_res_par = (matmul_29_control_param_index == 0)? 4 : 
                                                   (matmul_29_control_param_index == 1)? 16 : 12;
  assign cparam_matmul_29_stream_reduce_size = (matmul_29_control_param_index == 0)? 1024 : 
                                               (matmul_29_control_param_index == 1)? 256 : 128;
  assign cparam_matmul_29_stream_aligned_reduce_size = (matmul_29_control_param_index == 0)? 1024 : 
                                                       (matmul_29_control_param_index == 1)? 256 : 128;
  assign cparam_matmul_29_stream_omit_mask = (matmul_29_control_param_index == 0)? 0 : 
                                             (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_col_select_initval = (matmul_29_control_param_index == 0)? 0 : 
                                               (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_stride_col_par_col = (matmul_29_control_param_index == 0)? 1 : 
                                               (matmul_29_control_param_index == 1)? 1 : 1;
  assign cparam_matmul_29_stride_row_par_row = (matmul_29_control_param_index == 0)? 1 : 
                                               (matmul_29_control_param_index == 1)? 1 : 1;
  assign cparam_matmul_29_stride_col_mod_filter_num = (matmul_29_control_param_index == 0)? 0 : 
                                                      (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_filter_num_col_minus_stride_col_mod = (matmul_29_control_param_index == 0)? 1 : 
                                                                (matmul_29_control_param_index == 1)? 1 : 1;
  assign cparam_matmul_29_inc_act_laddr_conds_0 = (matmul_29_control_param_index == 0)? 0 : 
                                                  (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_inc_act_laddr_small = (matmul_29_control_param_index == 0)? 1024 : 
                                                (matmul_29_control_param_index == 1)? 256 : 128;
  assign cparam_matmul_29_inc_act_laddr_large = (matmul_29_control_param_index == 0)? 1024 : 
                                                (matmul_29_control_param_index == 1)? 256 : 128;
  assign cparam_matmul_29_inc_out_laddr_col = (matmul_29_control_param_index == 0)? 256 : 
                                              (matmul_29_control_param_index == 1)? 128 : 10;
  assign cparam_matmul_29_stream_act_local_small_offset = (matmul_29_control_param_index == 0)? 0 : 
                                                          (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_stream_act_local_large_offset = (matmul_29_control_param_index == 0)? 0 : 
                                                          (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_stream_act_local_small_flags_0 = (matmul_29_control_param_index == 0)? 0 : 
                                                           (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_stream_act_local_large_flags_0 = (matmul_29_control_param_index == 0)? 0 : 
                                                           (matmul_29_control_param_index == 1)? 0 : 0;
  assign cparam_matmul_29_inc_sync_out = (matmul_29_control_param_index == 0)? 1 : 
                                         (matmul_29_control_param_index == 1)? 1 : 1;
  assign cparam_matmul_29_inc_sync_out_res = (matmul_29_control_param_index == 0)? 0 : 
                                             (matmul_29_control_param_index == 1)? 0 : 0;
  reg [32-1:0] _acc_0_fsm;
  localparam _acc_0_fsm_init = 0;
  wire _acc_0_start_flag;
  reg _acc_0_start;
  reg _acc_0_end_flag;
  reg _acc_0_term_sink;
  reg _acc_0_source_busy;
  reg _acc_0_sink_busy;
  reg _acc_0_x_idle;
  reg [3-1:0] _acc_0_x_source_mode;
  reg [32-1:0] _acc_0_x_source_offset;
  reg [33-1:0] _acc_0_x_source_size;
  reg [32-1:0] _acc_0_x_source_stride;
  reg [33-1:0] _acc_0_x_source_count;
  reg [32-1:0] _acc_0_x_source_offset_buf;
  reg [32-1:0] _acc_0_x_source_stride_buf;
  reg [8-1:0] _acc_0_x_source_ram_sel;
  reg [32-1:0] _acc_0_x_source_ram_raddr;
  reg _acc_0_x_source_ram_renable;
  wire [32-1:0] _acc_0_x_source_ram_rdata;
  reg _acc_0_x_source_ram_rvalid;
  reg [32-1:0] _acc_0_x_source_empty_data;
  reg _acc_0_rshift_idle;
  reg [3-1:0] _acc_0_rshift_source_mode;
  reg [32-1:0] _acc_0_rshift_source_offset;
  reg [33-1:0] _acc_0_rshift_source_size;
  reg [32-1:0] _acc_0_rshift_source_stride;
  reg [33-1:0] _acc_0_rshift_source_count;
  reg [32-1:0] _acc_0_rshift_source_offset_buf;
  reg [32-1:0] _acc_0_rshift_source_stride_buf;
  reg [8-1:0] _acc_0_rshift_source_ram_sel;
  reg [32-1:0] _acc_0_rshift_source_ram_raddr;
  reg _acc_0_rshift_source_ram_renable;
  wire [32-1:0] _acc_0_rshift_source_ram_rdata;
  reg _acc_0_rshift_source_ram_rvalid;
  reg [32-1:0] _acc_0_rshift_source_empty_data;
  reg [32-1:0] _acc_0_size_next_constant_data;
  reg _acc_0_reduce_reset;
  reg [3-1:0] _acc_0_sum_sink_mode;
  reg [32-1:0] _acc_0_sum_sink_offset;
  reg [33-1:0] _acc_0_sum_sink_size;
  reg [32-1:0] _acc_0_sum_sink_stride;
  reg [33-1:0] _acc_0_sum_sink_count;
  reg [32-1:0] _acc_0_sum_sink_offset_buf;
  reg [32-1:0] _acc_0_sum_sink_stride_buf;
  reg [8-1:0] _acc_0_sum_sink_ram_sel;
  reg [32-1:0] _acc_0_sum_sink_waddr;
  reg _acc_0_sum_sink_wenable;
  reg [32-1:0] _acc_0_sum_sink_wdata;
  reg [3-1:0] _acc_0_valid_sink_mode;
  reg [32-1:0] _acc_0_valid_sink_offset;
  reg [33-1:0] _acc_0_valid_sink_size;
  reg [32-1:0] _acc_0_valid_sink_stride;
  reg [33-1:0] _acc_0_valid_sink_count;
  reg [32-1:0] _acc_0_valid_sink_offset_buf;
  reg [32-1:0] _acc_0_valid_sink_stride_buf;
  reg [8-1:0] _acc_0_valid_sink_ram_sel;
  reg [32-1:0] _acc_0_valid_sink_waddr;
  reg _acc_0_valid_sink_wenable;
  reg [1-1:0] _acc_0_valid_sink_wdata;
  reg [32-1:0] _add_tree_1_fsm;
  localparam _add_tree_1_fsm_init = 0;
  wire _add_tree_1_start_flag;
  reg _add_tree_1_start;
  reg _add_tree_1_end_flag;
  reg _add_tree_1_term_sink;
  reg _add_tree_1_source_busy;
  reg _add_tree_1_sink_busy;
  reg _add_tree_1_var0_idle;
  reg [3-1:0] _add_tree_1_var0_source_mode;
  reg [32-1:0] _add_tree_1_var0_source_offset;
  reg [33-1:0] _add_tree_1_var0_source_size;
  reg [32-1:0] _add_tree_1_var0_source_stride;
  reg [33-1:0] _add_tree_1_var0_source_count;
  reg [32-1:0] _add_tree_1_var0_source_offset_buf;
  reg [32-1:0] _add_tree_1_var0_source_stride_buf;
  reg [8-1:0] _add_tree_1_var0_source_ram_sel;
  reg [32-1:0] _add_tree_1_var0_source_ram_raddr;
  reg _add_tree_1_var0_source_ram_renable;
  wire [32-1:0] _add_tree_1_var0_source_ram_rdata;
  reg _add_tree_1_var0_source_ram_rvalid;
  reg [32-1:0] _add_tree_1_var0_source_empty_data;
  reg [3-1:0] _add_tree_1_sum_sink_mode;
  reg [32-1:0] _add_tree_1_sum_sink_offset;
  reg [33-1:0] _add_tree_1_sum_sink_size;
  reg [32-1:0] _add_tree_1_sum_sink_stride;
  reg [33-1:0] _add_tree_1_sum_sink_count;
  reg [32-1:0] _add_tree_1_sum_sink_offset_buf;
  reg [32-1:0] _add_tree_1_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_1_sum_sink_ram_sel;
  reg [32-1:0] _add_tree_1_sum_sink_waddr;
  reg _add_tree_1_sum_sink_wenable;
  reg [32-1:0] _add_tree_1_sum_sink_wdata;
  reg [32-1:0] _add_tree_2_fsm;
  localparam _add_tree_2_fsm_init = 0;
  wire _add_tree_2_start_flag;
  reg _add_tree_2_start;
  reg _add_tree_2_end_flag;
  reg _add_tree_2_term_sink;
  reg _add_tree_2_source_busy;
  reg _add_tree_2_sink_busy;
  reg _add_tree_2_var0_idle;
  reg [3-1:0] _add_tree_2_var0_source_mode;
  reg [32-1:0] _add_tree_2_var0_source_offset;
  reg [33-1:0] _add_tree_2_var0_source_size;
  reg [32-1:0] _add_tree_2_var0_source_stride;
  reg [33-1:0] _add_tree_2_var0_source_count;
  reg [32-1:0] _add_tree_2_var0_source_offset_buf;
  reg [32-1:0] _add_tree_2_var0_source_stride_buf;
  reg [8-1:0] _add_tree_2_var0_source_ram_sel;
  reg [32-1:0] _add_tree_2_var0_source_ram_raddr;
  reg _add_tree_2_var0_source_ram_renable;
  wire [32-1:0] _add_tree_2_var0_source_ram_rdata;
  reg _add_tree_2_var0_source_ram_rvalid;
  reg [32-1:0] _add_tree_2_var0_source_empty_data;
  reg _add_tree_2_var1_idle;
  reg [3-1:0] _add_tree_2_var1_source_mode;
  reg [32-1:0] _add_tree_2_var1_source_offset;
  reg [33-1:0] _add_tree_2_var1_source_size;
  reg [32-1:0] _add_tree_2_var1_source_stride;
  reg [33-1:0] _add_tree_2_var1_source_count;
  reg [32-1:0] _add_tree_2_var1_source_offset_buf;
  reg [32-1:0] _add_tree_2_var1_source_stride_buf;
  reg [8-1:0] _add_tree_2_var1_source_ram_sel;
  reg [32-1:0] _add_tree_2_var1_source_ram_raddr;
  reg _add_tree_2_var1_source_ram_renable;
  wire [32-1:0] _add_tree_2_var1_source_ram_rdata;
  reg _add_tree_2_var1_source_ram_rvalid;
  reg [32-1:0] _add_tree_2_var1_source_empty_data;
  reg _add_tree_2_var2_idle;
  reg [3-1:0] _add_tree_2_var2_source_mode;
  reg [32-1:0] _add_tree_2_var2_source_offset;
  reg [33-1:0] _add_tree_2_var2_source_size;
  reg [32-1:0] _add_tree_2_var2_source_stride;
  reg [33-1:0] _add_tree_2_var2_source_count;
  reg [32-1:0] _add_tree_2_var2_source_offset_buf;
  reg [32-1:0] _add_tree_2_var2_source_stride_buf;
  reg [8-1:0] _add_tree_2_var2_source_ram_sel;
  reg [32-1:0] _add_tree_2_var2_source_ram_raddr;
  reg _add_tree_2_var2_source_ram_renable;
  wire [32-1:0] _add_tree_2_var2_source_ram_rdata;
  reg _add_tree_2_var2_source_ram_rvalid;
  reg [32-1:0] _add_tree_2_var2_source_empty_data;
  reg _add_tree_2_var3_idle;
  reg [3-1:0] _add_tree_2_var3_source_mode;
  reg [32-1:0] _add_tree_2_var3_source_offset;
  reg [33-1:0] _add_tree_2_var3_source_size;
  reg [32-1:0] _add_tree_2_var3_source_stride;
  reg [33-1:0] _add_tree_2_var3_source_count;
  reg [32-1:0] _add_tree_2_var3_source_offset_buf;
  reg [32-1:0] _add_tree_2_var3_source_stride_buf;
  reg [8-1:0] _add_tree_2_var3_source_ram_sel;
  reg [32-1:0] _add_tree_2_var3_source_ram_raddr;
  reg _add_tree_2_var3_source_ram_renable;
  wire [32-1:0] _add_tree_2_var3_source_ram_rdata;
  reg _add_tree_2_var3_source_ram_rvalid;
  reg [32-1:0] _add_tree_2_var3_source_empty_data;
  reg _add_tree_2_var4_idle;
  reg [3-1:0] _add_tree_2_var4_source_mode;
  reg [32-1:0] _add_tree_2_var4_source_offset;
  reg [33-1:0] _add_tree_2_var4_source_size;
  reg [32-1:0] _add_tree_2_var4_source_stride;
  reg [33-1:0] _add_tree_2_var4_source_count;
  reg [32-1:0] _add_tree_2_var4_source_offset_buf;
  reg [32-1:0] _add_tree_2_var4_source_stride_buf;
  reg [8-1:0] _add_tree_2_var4_source_ram_sel;
  reg [32-1:0] _add_tree_2_var4_source_ram_raddr;
  reg _add_tree_2_var4_source_ram_renable;
  wire [32-1:0] _add_tree_2_var4_source_ram_rdata;
  reg _add_tree_2_var4_source_ram_rvalid;
  reg [32-1:0] _add_tree_2_var4_source_empty_data;
  reg _add_tree_2_var5_idle;
  reg [3-1:0] _add_tree_2_var5_source_mode;
  reg [32-1:0] _add_tree_2_var5_source_offset;
  reg [33-1:0] _add_tree_2_var5_source_size;
  reg [32-1:0] _add_tree_2_var5_source_stride;
  reg [33-1:0] _add_tree_2_var5_source_count;
  reg [32-1:0] _add_tree_2_var5_source_offset_buf;
  reg [32-1:0] _add_tree_2_var5_source_stride_buf;
  reg [8-1:0] _add_tree_2_var5_source_ram_sel;
  reg [32-1:0] _add_tree_2_var5_source_ram_raddr;
  reg _add_tree_2_var5_source_ram_renable;
  wire [32-1:0] _add_tree_2_var5_source_ram_rdata;
  reg _add_tree_2_var5_source_ram_rvalid;
  reg [32-1:0] _add_tree_2_var5_source_empty_data;
  reg _add_tree_2_var6_idle;
  reg [3-1:0] _add_tree_2_var6_source_mode;
  reg [32-1:0] _add_tree_2_var6_source_offset;
  reg [33-1:0] _add_tree_2_var6_source_size;
  reg [32-1:0] _add_tree_2_var6_source_stride;
  reg [33-1:0] _add_tree_2_var6_source_count;
  reg [32-1:0] _add_tree_2_var6_source_offset_buf;
  reg [32-1:0] _add_tree_2_var6_source_stride_buf;
  reg [8-1:0] _add_tree_2_var6_source_ram_sel;
  reg [32-1:0] _add_tree_2_var6_source_ram_raddr;
  reg _add_tree_2_var6_source_ram_renable;
  wire [32-1:0] _add_tree_2_var6_source_ram_rdata;
  reg _add_tree_2_var6_source_ram_rvalid;
  reg [32-1:0] _add_tree_2_var6_source_empty_data;
  reg _add_tree_2_var7_idle;
  reg [3-1:0] _add_tree_2_var7_source_mode;
  reg [32-1:0] _add_tree_2_var7_source_offset;
  reg [33-1:0] _add_tree_2_var7_source_size;
  reg [32-1:0] _add_tree_2_var7_source_stride;
  reg [33-1:0] _add_tree_2_var7_source_count;
  reg [32-1:0] _add_tree_2_var7_source_offset_buf;
  reg [32-1:0] _add_tree_2_var7_source_stride_buf;
  reg [8-1:0] _add_tree_2_var7_source_ram_sel;
  reg [32-1:0] _add_tree_2_var7_source_ram_raddr;
  reg _add_tree_2_var7_source_ram_renable;
  wire [32-1:0] _add_tree_2_var7_source_ram_rdata;
  reg _add_tree_2_var7_source_ram_rvalid;
  reg [32-1:0] _add_tree_2_var7_source_empty_data;
  reg _add_tree_2_var8_idle;
  reg [3-1:0] _add_tree_2_var8_source_mode;
  reg [32-1:0] _add_tree_2_var8_source_offset;
  reg [33-1:0] _add_tree_2_var8_source_size;
  reg [32-1:0] _add_tree_2_var8_source_stride;
  reg [33-1:0] _add_tree_2_var8_source_count;
  reg [32-1:0] _add_tree_2_var8_source_offset_buf;
  reg [32-1:0] _add_tree_2_var8_source_stride_buf;
  reg [8-1:0] _add_tree_2_var8_source_ram_sel;
  reg [32-1:0] _add_tree_2_var8_source_ram_raddr;
  reg _add_tree_2_var8_source_ram_renable;
  wire [32-1:0] _add_tree_2_var8_source_ram_rdata;
  reg _add_tree_2_var8_source_ram_rvalid;
  reg [32-1:0] _add_tree_2_var8_source_empty_data;
  reg [3-1:0] _add_tree_2_sum_sink_mode;
  reg [32-1:0] _add_tree_2_sum_sink_offset;
  reg [33-1:0] _add_tree_2_sum_sink_size;
  reg [32-1:0] _add_tree_2_sum_sink_stride;
  reg [33-1:0] _add_tree_2_sum_sink_count;
  reg [32-1:0] _add_tree_2_sum_sink_offset_buf;
  reg [32-1:0] _add_tree_2_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_2_sum_sink_ram_sel;
  reg [32-1:0] _add_tree_2_sum_sink_waddr;
  reg _add_tree_2_sum_sink_wenable;
  reg [32-1:0] _add_tree_2_sum_sink_wdata;
  reg [32-1:0] _mul_rshift_clip_3_fsm;
  localparam _mul_rshift_clip_3_fsm_init = 0;
  wire _mul_rshift_clip_3_start_flag;
  reg _mul_rshift_clip_3_start;
  reg _mul_rshift_clip_3_end_flag;
  reg _mul_rshift_clip_3_term_sink;
  reg _mul_rshift_clip_3_source_busy;
  reg _mul_rshift_clip_3_sink_busy;
  reg _mul_rshift_clip_3_x_idle;
  reg [3-1:0] _mul_rshift_clip_3_x_source_mode;
  reg [32-1:0] _mul_rshift_clip_3_x_source_offset;
  reg [33-1:0] _mul_rshift_clip_3_x_source_size;
  reg [32-1:0] _mul_rshift_clip_3_x_source_stride;
  reg [33-1:0] _mul_rshift_clip_3_x_source_count;
  reg [32-1:0] _mul_rshift_clip_3_x_source_offset_buf;
  reg [32-1:0] _mul_rshift_clip_3_x_source_stride_buf;
  reg [8-1:0] _mul_rshift_clip_3_x_source_ram_sel;
  reg [32-1:0] _mul_rshift_clip_3_x_source_ram_raddr;
  reg _mul_rshift_clip_3_x_source_ram_renable;
  wire [32-1:0] _mul_rshift_clip_3_x_source_ram_rdata;
  reg _mul_rshift_clip_3_x_source_ram_rvalid;
  reg [32-1:0] _mul_rshift_clip_3_x_source_empty_data;
  reg _mul_rshift_clip_3_y_idle;
  reg [3-1:0] _mul_rshift_clip_3_y_source_mode;
  reg [32-1:0] _mul_rshift_clip_3_y_source_offset;
  reg [33-1:0] _mul_rshift_clip_3_y_source_size;
  reg [32-1:0] _mul_rshift_clip_3_y_source_stride;
  reg [33-1:0] _mul_rshift_clip_3_y_source_count;
  reg [32-1:0] _mul_rshift_clip_3_y_source_offset_buf;
  reg [32-1:0] _mul_rshift_clip_3_y_source_stride_buf;
  reg [8-1:0] _mul_rshift_clip_3_y_source_ram_sel;
  reg [32-1:0] _mul_rshift_clip_3_y_source_ram_raddr;
  reg _mul_rshift_clip_3_y_source_ram_renable;
  wire [8-1:0] _mul_rshift_clip_3_y_source_ram_rdata;
  reg _mul_rshift_clip_3_y_source_ram_rvalid;
  reg [8-1:0] _mul_rshift_clip_3_y_source_empty_data;
  reg _mul_rshift_clip_3_rshift_idle;
  reg [3-1:0] _mul_rshift_clip_3_rshift_source_mode;
  reg [32-1:0] _mul_rshift_clip_3_rshift_source_offset;
  reg [33-1:0] _mul_rshift_clip_3_rshift_source_size;
  reg [32-1:0] _mul_rshift_clip_3_rshift_source_stride;
  reg [33-1:0] _mul_rshift_clip_3_rshift_source_count;
  reg [32-1:0] _mul_rshift_clip_3_rshift_source_offset_buf;
  reg [32-1:0] _mul_rshift_clip_3_rshift_source_stride_buf;
  reg [8-1:0] _mul_rshift_clip_3_rshift_source_ram_sel;
  reg [32-1:0] _mul_rshift_clip_3_rshift_source_ram_raddr;
  reg _mul_rshift_clip_3_rshift_source_ram_renable;
  wire [32-1:0] _mul_rshift_clip_3_rshift_source_ram_rdata;
  reg _mul_rshift_clip_3_rshift_source_ram_rvalid;
  reg [32-1:0] _mul_rshift_clip_3_rshift_source_empty_data;
  reg [3-1:0] _mul_rshift_clip_3_z_sink_mode;
  reg [32-1:0] _mul_rshift_clip_3_z_sink_offset;
  reg [33-1:0] _mul_rshift_clip_3_z_sink_size;
  reg [32-1:0] _mul_rshift_clip_3_z_sink_stride;
  reg [33-1:0] _mul_rshift_clip_3_z_sink_count;
  reg [32-1:0] _mul_rshift_clip_3_z_sink_offset_buf;
  reg [32-1:0] _mul_rshift_clip_3_z_sink_stride_buf;
  reg [8-1:0] _mul_rshift_clip_3_z_sink_ram_sel;
  reg [32-1:0] _mul_rshift_clip_3_z_sink_waddr;
  reg _mul_rshift_clip_3_z_sink_wenable;
  reg [8-1:0] _mul_rshift_clip_3_z_sink_wdata;
  reg [32-1:0] _mul_4_fsm;
  localparam _mul_4_fsm_init = 0;
  wire _mul_4_start_flag;
  reg _mul_4_start;
  reg _mul_4_end_flag;
  reg _mul_4_term_sink;
  reg _mul_4_source_busy;
  reg _mul_4_sink_busy;
  reg _mul_4_x_idle;
  reg [3-1:0] _mul_4_x_source_mode;
  reg [32-1:0] _mul_4_x_source_offset;
  reg [33-1:0] _mul_4_x_source_size;
  reg [32-1:0] _mul_4_x_source_stride;
  reg [33-1:0] _mul_4_x_source_count;
  reg [32-1:0] _mul_4_x_source_offset_buf;
  reg [32-1:0] _mul_4_x_source_stride_buf;
  reg [8-1:0] _mul_4_x_source_ram_sel;
  reg [32-1:0] _mul_4_x_source_ram_raddr;
  reg _mul_4_x_source_ram_renable;
  wire [8-1:0] _mul_4_x_source_ram_rdata;
  reg _mul_4_x_source_ram_rvalid;
  reg [8-1:0] _mul_4_x_source_empty_data;
  reg _mul_4_y_idle;
  reg [3-1:0] _mul_4_y_source_mode;
  reg [32-1:0] _mul_4_y_source_offset;
  reg [33-1:0] _mul_4_y_source_size;
  reg [32-1:0] _mul_4_y_source_stride;
  reg [33-1:0] _mul_4_y_source_count;
  reg [32-1:0] _mul_4_y_source_offset_buf;
  reg [32-1:0] _mul_4_y_source_stride_buf;
  reg [8-1:0] _mul_4_y_source_ram_sel;
  reg [32-1:0] _mul_4_y_source_ram_raddr;
  reg _mul_4_y_source_ram_renable;
  wire [4-1:0] _mul_4_y_source_ram_rdata;
  reg _mul_4_y_source_ram_rvalid;
  reg [4-1:0] _mul_4_y_source_empty_data;
  reg _mul_4_rshift_idle;
  reg [3-1:0] _mul_4_rshift_source_mode;
  reg [32-1:0] _mul_4_rshift_source_offset;
  reg [33-1:0] _mul_4_rshift_source_size;
  reg [32-1:0] _mul_4_rshift_source_stride;
  reg [33-1:0] _mul_4_rshift_source_count;
  reg [32-1:0] _mul_4_rshift_source_offset_buf;
  reg [32-1:0] _mul_4_rshift_source_stride_buf;
  reg [8-1:0] _mul_4_rshift_source_ram_sel;
  reg [32-1:0] _mul_4_rshift_source_ram_raddr;
  reg _mul_4_rshift_source_ram_renable;
  wire [8-1:0] _mul_4_rshift_source_ram_rdata;
  reg _mul_4_rshift_source_ram_rvalid;
  reg [8-1:0] _mul_4_rshift_source_empty_data;
  reg [3-1:0] _mul_4_z_sink_mode;
  reg [32-1:0] _mul_4_z_sink_offset;
  reg [33-1:0] _mul_4_z_sink_size;
  reg [32-1:0] _mul_4_z_sink_stride;
  reg [33-1:0] _mul_4_z_sink_count;
  reg [32-1:0] _mul_4_z_sink_offset_buf;
  reg [32-1:0] _mul_4_z_sink_stride_buf;
  reg [8-1:0] _mul_4_z_sink_ram_sel;
  reg [32-1:0] _mul_4_z_sink_waddr;
  reg _mul_4_z_sink_wenable;
  reg [12-1:0] _mul_4_z_sink_wdata;
  reg [32-1:0] _mul_5_fsm;
  localparam _mul_5_fsm_init = 0;
  wire _mul_5_start_flag;
  reg _mul_5_start;
  reg _mul_5_end_flag;
  reg _mul_5_term_sink;
  reg _mul_5_source_busy;
  reg _mul_5_sink_busy;
  reg _mul_5_x_idle;
  reg [3-1:0] _mul_5_x_source_mode;
  reg [32-1:0] _mul_5_x_source_offset;
  reg [33-1:0] _mul_5_x_source_size;
  reg [32-1:0] _mul_5_x_source_stride;
  reg [33-1:0] _mul_5_x_source_count;
  reg [32-1:0] _mul_5_x_source_offset_buf;
  reg [32-1:0] _mul_5_x_source_stride_buf;
  reg [8-1:0] _mul_5_x_source_ram_sel;
  reg [32-1:0] _mul_5_x_source_ram_raddr;
  reg _mul_5_x_source_ram_renable;
  wire [8-1:0] _mul_5_x_source_ram_rdata;
  reg _mul_5_x_source_ram_rvalid;
  reg [8-1:0] _mul_5_x_source_empty_data;
  reg _mul_5_y_idle;
  reg [3-1:0] _mul_5_y_source_mode;
  reg [32-1:0] _mul_5_y_source_offset;
  reg [33-1:0] _mul_5_y_source_size;
  reg [32-1:0] _mul_5_y_source_stride;
  reg [33-1:0] _mul_5_y_source_count;
  reg [32-1:0] _mul_5_y_source_offset_buf;
  reg [32-1:0] _mul_5_y_source_stride_buf;
  reg [8-1:0] _mul_5_y_source_ram_sel;
  reg [32-1:0] _mul_5_y_source_ram_raddr;
  reg _mul_5_y_source_ram_renable;
  wire [4-1:0] _mul_5_y_source_ram_rdata;
  reg _mul_5_y_source_ram_rvalid;
  reg [4-1:0] _mul_5_y_source_empty_data;
  reg _mul_5_rshift_idle;
  reg [3-1:0] _mul_5_rshift_source_mode;
  reg [32-1:0] _mul_5_rshift_source_offset;
  reg [33-1:0] _mul_5_rshift_source_size;
  reg [32-1:0] _mul_5_rshift_source_stride;
  reg [33-1:0] _mul_5_rshift_source_count;
  reg [32-1:0] _mul_5_rshift_source_offset_buf;
  reg [32-1:0] _mul_5_rshift_source_stride_buf;
  reg [8-1:0] _mul_5_rshift_source_ram_sel;
  reg [32-1:0] _mul_5_rshift_source_ram_raddr;
  reg _mul_5_rshift_source_ram_renable;
  wire [8-1:0] _mul_5_rshift_source_ram_rdata;
  reg _mul_5_rshift_source_ram_rvalid;
  reg [8-1:0] _mul_5_rshift_source_empty_data;
  reg [3-1:0] _mul_5_z_sink_mode;
  reg [32-1:0] _mul_5_z_sink_offset;
  reg [33-1:0] _mul_5_z_sink_size;
  reg [32-1:0] _mul_5_z_sink_stride;
  reg [33-1:0] _mul_5_z_sink_count;
  reg [32-1:0] _mul_5_z_sink_offset_buf;
  reg [32-1:0] _mul_5_z_sink_stride_buf;
  reg [8-1:0] _mul_5_z_sink_ram_sel;
  reg [32-1:0] _mul_5_z_sink_waddr;
  reg _mul_5_z_sink_wenable;
  reg [12-1:0] _mul_5_z_sink_wdata;
  reg [32-1:0] _mul_6_fsm;
  localparam _mul_6_fsm_init = 0;
  wire _mul_6_start_flag;
  reg _mul_6_start;
  reg _mul_6_end_flag;
  reg _mul_6_term_sink;
  reg _mul_6_source_busy;
  reg _mul_6_sink_busy;
  reg _mul_6_x_idle;
  reg [3-1:0] _mul_6_x_source_mode;
  reg [32-1:0] _mul_6_x_source_offset;
  reg [33-1:0] _mul_6_x_source_size;
  reg [32-1:0] _mul_6_x_source_stride;
  reg [33-1:0] _mul_6_x_source_count;
  reg [32-1:0] _mul_6_x_source_offset_buf;
  reg [32-1:0] _mul_6_x_source_stride_buf;
  reg [8-1:0] _mul_6_x_source_ram_sel;
  reg [32-1:0] _mul_6_x_source_ram_raddr;
  reg _mul_6_x_source_ram_renable;
  wire [8-1:0] _mul_6_x_source_ram_rdata;
  reg _mul_6_x_source_ram_rvalid;
  reg [8-1:0] _mul_6_x_source_empty_data;
  reg _mul_6_y_idle;
  reg [3-1:0] _mul_6_y_source_mode;
  reg [32-1:0] _mul_6_y_source_offset;
  reg [33-1:0] _mul_6_y_source_size;
  reg [32-1:0] _mul_6_y_source_stride;
  reg [33-1:0] _mul_6_y_source_count;
  reg [32-1:0] _mul_6_y_source_offset_buf;
  reg [32-1:0] _mul_6_y_source_stride_buf;
  reg [8-1:0] _mul_6_y_source_ram_sel;
  reg [32-1:0] _mul_6_y_source_ram_raddr;
  reg _mul_6_y_source_ram_renable;
  wire [4-1:0] _mul_6_y_source_ram_rdata;
  reg _mul_6_y_source_ram_rvalid;
  reg [4-1:0] _mul_6_y_source_empty_data;
  reg _mul_6_rshift_idle;
  reg [3-1:0] _mul_6_rshift_source_mode;
  reg [32-1:0] _mul_6_rshift_source_offset;
  reg [33-1:0] _mul_6_rshift_source_size;
  reg [32-1:0] _mul_6_rshift_source_stride;
  reg [33-1:0] _mul_6_rshift_source_count;
  reg [32-1:0] _mul_6_rshift_source_offset_buf;
  reg [32-1:0] _mul_6_rshift_source_stride_buf;
  reg [8-1:0] _mul_6_rshift_source_ram_sel;
  reg [32-1:0] _mul_6_rshift_source_ram_raddr;
  reg _mul_6_rshift_source_ram_renable;
  wire [8-1:0] _mul_6_rshift_source_ram_rdata;
  reg _mul_6_rshift_source_ram_rvalid;
  reg [8-1:0] _mul_6_rshift_source_empty_data;
  reg [3-1:0] _mul_6_z_sink_mode;
  reg [32-1:0] _mul_6_z_sink_offset;
  reg [33-1:0] _mul_6_z_sink_size;
  reg [32-1:0] _mul_6_z_sink_stride;
  reg [33-1:0] _mul_6_z_sink_count;
  reg [32-1:0] _mul_6_z_sink_offset_buf;
  reg [32-1:0] _mul_6_z_sink_stride_buf;
  reg [8-1:0] _mul_6_z_sink_ram_sel;
  reg [32-1:0] _mul_6_z_sink_waddr;
  reg _mul_6_z_sink_wenable;
  reg [12-1:0] _mul_6_z_sink_wdata;
  reg [32-1:0] _mul_7_fsm;
  localparam _mul_7_fsm_init = 0;
  wire _mul_7_start_flag;
  reg _mul_7_start;
  reg _mul_7_end_flag;
  reg _mul_7_term_sink;
  reg _mul_7_source_busy;
  reg _mul_7_sink_busy;
  reg _mul_7_x_idle;
  reg [3-1:0] _mul_7_x_source_mode;
  reg [32-1:0] _mul_7_x_source_offset;
  reg [33-1:0] _mul_7_x_source_size;
  reg [32-1:0] _mul_7_x_source_stride;
  reg [33-1:0] _mul_7_x_source_count;
  reg [32-1:0] _mul_7_x_source_offset_buf;
  reg [32-1:0] _mul_7_x_source_stride_buf;
  reg [8-1:0] _mul_7_x_source_ram_sel;
  reg [32-1:0] _mul_7_x_source_ram_raddr;
  reg _mul_7_x_source_ram_renable;
  wire [8-1:0] _mul_7_x_source_ram_rdata;
  reg _mul_7_x_source_ram_rvalid;
  reg [8-1:0] _mul_7_x_source_empty_data;
  reg _mul_7_y_idle;
  reg [3-1:0] _mul_7_y_source_mode;
  reg [32-1:0] _mul_7_y_source_offset;
  reg [33-1:0] _mul_7_y_source_size;
  reg [32-1:0] _mul_7_y_source_stride;
  reg [33-1:0] _mul_7_y_source_count;
  reg [32-1:0] _mul_7_y_source_offset_buf;
  reg [32-1:0] _mul_7_y_source_stride_buf;
  reg [8-1:0] _mul_7_y_source_ram_sel;
  reg [32-1:0] _mul_7_y_source_ram_raddr;
  reg _mul_7_y_source_ram_renable;
  wire [4-1:0] _mul_7_y_source_ram_rdata;
  reg _mul_7_y_source_ram_rvalid;
  reg [4-1:0] _mul_7_y_source_empty_data;
  reg _mul_7_rshift_idle;
  reg [3-1:0] _mul_7_rshift_source_mode;
  reg [32-1:0] _mul_7_rshift_source_offset;
  reg [33-1:0] _mul_7_rshift_source_size;
  reg [32-1:0] _mul_7_rshift_source_stride;
  reg [33-1:0] _mul_7_rshift_source_count;
  reg [32-1:0] _mul_7_rshift_source_offset_buf;
  reg [32-1:0] _mul_7_rshift_source_stride_buf;
  reg [8-1:0] _mul_7_rshift_source_ram_sel;
  reg [32-1:0] _mul_7_rshift_source_ram_raddr;
  reg _mul_7_rshift_source_ram_renable;
  wire [8-1:0] _mul_7_rshift_source_ram_rdata;
  reg _mul_7_rshift_source_ram_rvalid;
  reg [8-1:0] _mul_7_rshift_source_empty_data;
  reg [3-1:0] _mul_7_z_sink_mode;
  reg [32-1:0] _mul_7_z_sink_offset;
  reg [33-1:0] _mul_7_z_sink_size;
  reg [32-1:0] _mul_7_z_sink_stride;
  reg [33-1:0] _mul_7_z_sink_count;
  reg [32-1:0] _mul_7_z_sink_offset_buf;
  reg [32-1:0] _mul_7_z_sink_stride_buf;
  reg [8-1:0] _mul_7_z_sink_ram_sel;
  reg [32-1:0] _mul_7_z_sink_waddr;
  reg _mul_7_z_sink_wenable;
  reg [12-1:0] _mul_7_z_sink_wdata;
  reg [32-1:0] _mul_8_fsm;
  localparam _mul_8_fsm_init = 0;
  wire _mul_8_start_flag;
  reg _mul_8_start;
  reg _mul_8_end_flag;
  reg _mul_8_term_sink;
  reg _mul_8_source_busy;
  reg _mul_8_sink_busy;
  reg _mul_8_x_idle;
  reg [3-1:0] _mul_8_x_source_mode;
  reg [32-1:0] _mul_8_x_source_offset;
  reg [33-1:0] _mul_8_x_source_size;
  reg [32-1:0] _mul_8_x_source_stride;
  reg [33-1:0] _mul_8_x_source_count;
  reg [32-1:0] _mul_8_x_source_offset_buf;
  reg [32-1:0] _mul_8_x_source_stride_buf;
  reg [8-1:0] _mul_8_x_source_ram_sel;
  reg [32-1:0] _mul_8_x_source_ram_raddr;
  reg _mul_8_x_source_ram_renable;
  wire [8-1:0] _mul_8_x_source_ram_rdata;
  reg _mul_8_x_source_ram_rvalid;
  reg [8-1:0] _mul_8_x_source_empty_data;
  reg _mul_8_y_idle;
  reg [3-1:0] _mul_8_y_source_mode;
  reg [32-1:0] _mul_8_y_source_offset;
  reg [33-1:0] _mul_8_y_source_size;
  reg [32-1:0] _mul_8_y_source_stride;
  reg [33-1:0] _mul_8_y_source_count;
  reg [32-1:0] _mul_8_y_source_offset_buf;
  reg [32-1:0] _mul_8_y_source_stride_buf;
  reg [8-1:0] _mul_8_y_source_ram_sel;
  reg [32-1:0] _mul_8_y_source_ram_raddr;
  reg _mul_8_y_source_ram_renable;
  wire [4-1:0] _mul_8_y_source_ram_rdata;
  reg _mul_8_y_source_ram_rvalid;
  reg [4-1:0] _mul_8_y_source_empty_data;
  reg _mul_8_rshift_idle;
  reg [3-1:0] _mul_8_rshift_source_mode;
  reg [32-1:0] _mul_8_rshift_source_offset;
  reg [33-1:0] _mul_8_rshift_source_size;
  reg [32-1:0] _mul_8_rshift_source_stride;
  reg [33-1:0] _mul_8_rshift_source_count;
  reg [32-1:0] _mul_8_rshift_source_offset_buf;
  reg [32-1:0] _mul_8_rshift_source_stride_buf;
  reg [8-1:0] _mul_8_rshift_source_ram_sel;
  reg [32-1:0] _mul_8_rshift_source_ram_raddr;
  reg _mul_8_rshift_source_ram_renable;
  wire [8-1:0] _mul_8_rshift_source_ram_rdata;
  reg _mul_8_rshift_source_ram_rvalid;
  reg [8-1:0] _mul_8_rshift_source_empty_data;
  reg [3-1:0] _mul_8_z_sink_mode;
  reg [32-1:0] _mul_8_z_sink_offset;
  reg [33-1:0] _mul_8_z_sink_size;
  reg [32-1:0] _mul_8_z_sink_stride;
  reg [33-1:0] _mul_8_z_sink_count;
  reg [32-1:0] _mul_8_z_sink_offset_buf;
  reg [32-1:0] _mul_8_z_sink_stride_buf;
  reg [8-1:0] _mul_8_z_sink_ram_sel;
  reg [32-1:0] _mul_8_z_sink_waddr;
  reg _mul_8_z_sink_wenable;
  reg [12-1:0] _mul_8_z_sink_wdata;
  reg [32-1:0] _mul_9_fsm;
  localparam _mul_9_fsm_init = 0;
  wire _mul_9_start_flag;
  reg _mul_9_start;
  reg _mul_9_end_flag;
  reg _mul_9_term_sink;
  reg _mul_9_source_busy;
  reg _mul_9_sink_busy;
  reg _mul_9_x_idle;
  reg [3-1:0] _mul_9_x_source_mode;
  reg [32-1:0] _mul_9_x_source_offset;
  reg [33-1:0] _mul_9_x_source_size;
  reg [32-1:0] _mul_9_x_source_stride;
  reg [33-1:0] _mul_9_x_source_count;
  reg [32-1:0] _mul_9_x_source_offset_buf;
  reg [32-1:0] _mul_9_x_source_stride_buf;
  reg [8-1:0] _mul_9_x_source_ram_sel;
  reg [32-1:0] _mul_9_x_source_ram_raddr;
  reg _mul_9_x_source_ram_renable;
  wire [8-1:0] _mul_9_x_source_ram_rdata;
  reg _mul_9_x_source_ram_rvalid;
  reg [8-1:0] _mul_9_x_source_empty_data;
  reg _mul_9_y_idle;
  reg [3-1:0] _mul_9_y_source_mode;
  reg [32-1:0] _mul_9_y_source_offset;
  reg [33-1:0] _mul_9_y_source_size;
  reg [32-1:0] _mul_9_y_source_stride;
  reg [33-1:0] _mul_9_y_source_count;
  reg [32-1:0] _mul_9_y_source_offset_buf;
  reg [32-1:0] _mul_9_y_source_stride_buf;
  reg [8-1:0] _mul_9_y_source_ram_sel;
  reg [32-1:0] _mul_9_y_source_ram_raddr;
  reg _mul_9_y_source_ram_renable;
  wire [4-1:0] _mul_9_y_source_ram_rdata;
  reg _mul_9_y_source_ram_rvalid;
  reg [4-1:0] _mul_9_y_source_empty_data;
  reg _mul_9_rshift_idle;
  reg [3-1:0] _mul_9_rshift_source_mode;
  reg [32-1:0] _mul_9_rshift_source_offset;
  reg [33-1:0] _mul_9_rshift_source_size;
  reg [32-1:0] _mul_9_rshift_source_stride;
  reg [33-1:0] _mul_9_rshift_source_count;
  reg [32-1:0] _mul_9_rshift_source_offset_buf;
  reg [32-1:0] _mul_9_rshift_source_stride_buf;
  reg [8-1:0] _mul_9_rshift_source_ram_sel;
  reg [32-1:0] _mul_9_rshift_source_ram_raddr;
  reg _mul_9_rshift_source_ram_renable;
  wire [8-1:0] _mul_9_rshift_source_ram_rdata;
  reg _mul_9_rshift_source_ram_rvalid;
  reg [8-1:0] _mul_9_rshift_source_empty_data;
  reg [3-1:0] _mul_9_z_sink_mode;
  reg [32-1:0] _mul_9_z_sink_offset;
  reg [33-1:0] _mul_9_z_sink_size;
  reg [32-1:0] _mul_9_z_sink_stride;
  reg [33-1:0] _mul_9_z_sink_count;
  reg [32-1:0] _mul_9_z_sink_offset_buf;
  reg [32-1:0] _mul_9_z_sink_stride_buf;
  reg [8-1:0] _mul_9_z_sink_ram_sel;
  reg [32-1:0] _mul_9_z_sink_waddr;
  reg _mul_9_z_sink_wenable;
  reg [12-1:0] _mul_9_z_sink_wdata;
  reg [32-1:0] _mul_10_fsm;
  localparam _mul_10_fsm_init = 0;
  wire _mul_10_start_flag;
  reg _mul_10_start;
  reg _mul_10_end_flag;
  reg _mul_10_term_sink;
  reg _mul_10_source_busy;
  reg _mul_10_sink_busy;
  reg _mul_10_x_idle;
  reg [3-1:0] _mul_10_x_source_mode;
  reg [32-1:0] _mul_10_x_source_offset;
  reg [33-1:0] _mul_10_x_source_size;
  reg [32-1:0] _mul_10_x_source_stride;
  reg [33-1:0] _mul_10_x_source_count;
  reg [32-1:0] _mul_10_x_source_offset_buf;
  reg [32-1:0] _mul_10_x_source_stride_buf;
  reg [8-1:0] _mul_10_x_source_ram_sel;
  reg [32-1:0] _mul_10_x_source_ram_raddr;
  reg _mul_10_x_source_ram_renable;
  wire [8-1:0] _mul_10_x_source_ram_rdata;
  reg _mul_10_x_source_ram_rvalid;
  reg [8-1:0] _mul_10_x_source_empty_data;
  reg _mul_10_y_idle;
  reg [3-1:0] _mul_10_y_source_mode;
  reg [32-1:0] _mul_10_y_source_offset;
  reg [33-1:0] _mul_10_y_source_size;
  reg [32-1:0] _mul_10_y_source_stride;
  reg [33-1:0] _mul_10_y_source_count;
  reg [32-1:0] _mul_10_y_source_offset_buf;
  reg [32-1:0] _mul_10_y_source_stride_buf;
  reg [8-1:0] _mul_10_y_source_ram_sel;
  reg [32-1:0] _mul_10_y_source_ram_raddr;
  reg _mul_10_y_source_ram_renable;
  wire [4-1:0] _mul_10_y_source_ram_rdata;
  reg _mul_10_y_source_ram_rvalid;
  reg [4-1:0] _mul_10_y_source_empty_data;
  reg _mul_10_rshift_idle;
  reg [3-1:0] _mul_10_rshift_source_mode;
  reg [32-1:0] _mul_10_rshift_source_offset;
  reg [33-1:0] _mul_10_rshift_source_size;
  reg [32-1:0] _mul_10_rshift_source_stride;
  reg [33-1:0] _mul_10_rshift_source_count;
  reg [32-1:0] _mul_10_rshift_source_offset_buf;
  reg [32-1:0] _mul_10_rshift_source_stride_buf;
  reg [8-1:0] _mul_10_rshift_source_ram_sel;
  reg [32-1:0] _mul_10_rshift_source_ram_raddr;
  reg _mul_10_rshift_source_ram_renable;
  wire [8-1:0] _mul_10_rshift_source_ram_rdata;
  reg _mul_10_rshift_source_ram_rvalid;
  reg [8-1:0] _mul_10_rshift_source_empty_data;
  reg [3-1:0] _mul_10_z_sink_mode;
  reg [32-1:0] _mul_10_z_sink_offset;
  reg [33-1:0] _mul_10_z_sink_size;
  reg [32-1:0] _mul_10_z_sink_stride;
  reg [33-1:0] _mul_10_z_sink_count;
  reg [32-1:0] _mul_10_z_sink_offset_buf;
  reg [32-1:0] _mul_10_z_sink_stride_buf;
  reg [8-1:0] _mul_10_z_sink_ram_sel;
  reg [32-1:0] _mul_10_z_sink_waddr;
  reg _mul_10_z_sink_wenable;
  reg [12-1:0] _mul_10_z_sink_wdata;
  reg [32-1:0] _mul_11_fsm;
  localparam _mul_11_fsm_init = 0;
  wire _mul_11_start_flag;
  reg _mul_11_start;
  reg _mul_11_end_flag;
  reg _mul_11_term_sink;
  reg _mul_11_source_busy;
  reg _mul_11_sink_busy;
  reg _mul_11_x_idle;
  reg [3-1:0] _mul_11_x_source_mode;
  reg [32-1:0] _mul_11_x_source_offset;
  reg [33-1:0] _mul_11_x_source_size;
  reg [32-1:0] _mul_11_x_source_stride;
  reg [33-1:0] _mul_11_x_source_count;
  reg [32-1:0] _mul_11_x_source_offset_buf;
  reg [32-1:0] _mul_11_x_source_stride_buf;
  reg [8-1:0] _mul_11_x_source_ram_sel;
  reg [32-1:0] _mul_11_x_source_ram_raddr;
  reg _mul_11_x_source_ram_renable;
  wire [8-1:0] _mul_11_x_source_ram_rdata;
  reg _mul_11_x_source_ram_rvalid;
  reg [8-1:0] _mul_11_x_source_empty_data;
  reg _mul_11_y_idle;
  reg [3-1:0] _mul_11_y_source_mode;
  reg [32-1:0] _mul_11_y_source_offset;
  reg [33-1:0] _mul_11_y_source_size;
  reg [32-1:0] _mul_11_y_source_stride;
  reg [33-1:0] _mul_11_y_source_count;
  reg [32-1:0] _mul_11_y_source_offset_buf;
  reg [32-1:0] _mul_11_y_source_stride_buf;
  reg [8-1:0] _mul_11_y_source_ram_sel;
  reg [32-1:0] _mul_11_y_source_ram_raddr;
  reg _mul_11_y_source_ram_renable;
  wire [4-1:0] _mul_11_y_source_ram_rdata;
  reg _mul_11_y_source_ram_rvalid;
  reg [4-1:0] _mul_11_y_source_empty_data;
  reg _mul_11_rshift_idle;
  reg [3-1:0] _mul_11_rshift_source_mode;
  reg [32-1:0] _mul_11_rshift_source_offset;
  reg [33-1:0] _mul_11_rshift_source_size;
  reg [32-1:0] _mul_11_rshift_source_stride;
  reg [33-1:0] _mul_11_rshift_source_count;
  reg [32-1:0] _mul_11_rshift_source_offset_buf;
  reg [32-1:0] _mul_11_rshift_source_stride_buf;
  reg [8-1:0] _mul_11_rshift_source_ram_sel;
  reg [32-1:0] _mul_11_rshift_source_ram_raddr;
  reg _mul_11_rshift_source_ram_renable;
  wire [8-1:0] _mul_11_rshift_source_ram_rdata;
  reg _mul_11_rshift_source_ram_rvalid;
  reg [8-1:0] _mul_11_rshift_source_empty_data;
  reg [3-1:0] _mul_11_z_sink_mode;
  reg [32-1:0] _mul_11_z_sink_offset;
  reg [33-1:0] _mul_11_z_sink_size;
  reg [32-1:0] _mul_11_z_sink_stride;
  reg [33-1:0] _mul_11_z_sink_count;
  reg [32-1:0] _mul_11_z_sink_offset_buf;
  reg [32-1:0] _mul_11_z_sink_stride_buf;
  reg [8-1:0] _mul_11_z_sink_ram_sel;
  reg [32-1:0] _mul_11_z_sink_waddr;
  reg _mul_11_z_sink_wenable;
  reg [12-1:0] _mul_11_z_sink_wdata;
  reg [32-1:0] _mul_12_fsm;
  localparam _mul_12_fsm_init = 0;
  wire _mul_12_start_flag;
  reg _mul_12_start;
  reg _mul_12_end_flag;
  reg _mul_12_term_sink;
  reg _mul_12_source_busy;
  reg _mul_12_sink_busy;
  reg _mul_12_x_idle;
  reg [3-1:0] _mul_12_x_source_mode;
  reg [32-1:0] _mul_12_x_source_offset;
  reg [33-1:0] _mul_12_x_source_size;
  reg [32-1:0] _mul_12_x_source_stride;
  reg [33-1:0] _mul_12_x_source_count;
  reg [32-1:0] _mul_12_x_source_offset_buf;
  reg [32-1:0] _mul_12_x_source_stride_buf;
  reg [8-1:0] _mul_12_x_source_ram_sel;
  reg [32-1:0] _mul_12_x_source_ram_raddr;
  reg _mul_12_x_source_ram_renable;
  wire [8-1:0] _mul_12_x_source_ram_rdata;
  reg _mul_12_x_source_ram_rvalid;
  reg [8-1:0] _mul_12_x_source_empty_data;
  reg _mul_12_y_idle;
  reg [3-1:0] _mul_12_y_source_mode;
  reg [32-1:0] _mul_12_y_source_offset;
  reg [33-1:0] _mul_12_y_source_size;
  reg [32-1:0] _mul_12_y_source_stride;
  reg [33-1:0] _mul_12_y_source_count;
  reg [32-1:0] _mul_12_y_source_offset_buf;
  reg [32-1:0] _mul_12_y_source_stride_buf;
  reg [8-1:0] _mul_12_y_source_ram_sel;
  reg [32-1:0] _mul_12_y_source_ram_raddr;
  reg _mul_12_y_source_ram_renable;
  wire [4-1:0] _mul_12_y_source_ram_rdata;
  reg _mul_12_y_source_ram_rvalid;
  reg [4-1:0] _mul_12_y_source_empty_data;
  reg _mul_12_rshift_idle;
  reg [3-1:0] _mul_12_rshift_source_mode;
  reg [32-1:0] _mul_12_rshift_source_offset;
  reg [33-1:0] _mul_12_rshift_source_size;
  reg [32-1:0] _mul_12_rshift_source_stride;
  reg [33-1:0] _mul_12_rshift_source_count;
  reg [32-1:0] _mul_12_rshift_source_offset_buf;
  reg [32-1:0] _mul_12_rshift_source_stride_buf;
  reg [8-1:0] _mul_12_rshift_source_ram_sel;
  reg [32-1:0] _mul_12_rshift_source_ram_raddr;
  reg _mul_12_rshift_source_ram_renable;
  wire [8-1:0] _mul_12_rshift_source_ram_rdata;
  reg _mul_12_rshift_source_ram_rvalid;
  reg [8-1:0] _mul_12_rshift_source_empty_data;
  reg [3-1:0] _mul_12_z_sink_mode;
  reg [32-1:0] _mul_12_z_sink_offset;
  reg [33-1:0] _mul_12_z_sink_size;
  reg [32-1:0] _mul_12_z_sink_stride;
  reg [33-1:0] _mul_12_z_sink_count;
  reg [32-1:0] _mul_12_z_sink_offset_buf;
  reg [32-1:0] _mul_12_z_sink_stride_buf;
  reg [8-1:0] _mul_12_z_sink_ram_sel;
  reg [32-1:0] _mul_12_z_sink_waddr;
  reg _mul_12_z_sink_wenable;
  reg [12-1:0] _mul_12_z_sink_wdata;
  reg [32-1:0] __reduce_max_13_fsm;
  localparam __reduce_max_13_fsm_init = 0;
  wire __reduce_max_13_start_flag;
  reg __reduce_max_13_start;
  reg __reduce_max_13_end_flag;
  reg __reduce_max_13_term_sink;
  reg __reduce_max_13_source_busy;
  reg __reduce_max_13_sink_busy;
  reg __reduce_max_13_x_idle;
  reg [3-1:0] __reduce_max_13_x_source_mode;
  reg [32-1:0] __reduce_max_13_x_source_offset;
  reg [33-1:0] __reduce_max_13_x_source_size;
  reg [32-1:0] __reduce_max_13_x_source_stride;
  reg [33-1:0] __reduce_max_13_x_source_count;
  reg [32-1:0] __reduce_max_13_x_source_offset_buf;
  reg [32-1:0] __reduce_max_13_x_source_stride_buf;
  reg [8-1:0] __reduce_max_13_x_source_ram_sel;
  reg [32-1:0] __reduce_max_13_x_source_ram_raddr;
  reg __reduce_max_13_x_source_ram_renable;
  wire [8-1:0] __reduce_max_13_x_source_ram_rdata;
  reg __reduce_max_13_x_source_ram_rvalid;
  reg [8-1:0] __reduce_max_13_x_source_empty_data;
  reg [8-1:0] __reduce_max_13_size_next_constant_data;
  reg __reduce_max_13_reduce_reset;
  reg [3-1:0] __reduce_max_13_data_sink_mode;
  reg [32-1:0] __reduce_max_13_data_sink_offset;
  reg [33-1:0] __reduce_max_13_data_sink_size;
  reg [32-1:0] __reduce_max_13_data_sink_stride;
  reg [33-1:0] __reduce_max_13_data_sink_count;
  reg [32-1:0] __reduce_max_13_data_sink_offset_buf;
  reg [32-1:0] __reduce_max_13_data_sink_stride_buf;
  reg [8-1:0] __reduce_max_13_data_sink_ram_sel;
  reg [32-1:0] __reduce_max_13_data_sink_waddr;
  reg __reduce_max_13_data_sink_wenable;
  reg [8-1:0] __reduce_max_13_data_sink_wdata;
  reg [3-1:0] __reduce_max_13_valid_sink_mode;
  reg [32-1:0] __reduce_max_13_valid_sink_offset;
  reg [33-1:0] __reduce_max_13_valid_sink_size;
  reg [32-1:0] __reduce_max_13_valid_sink_stride;
  reg [33-1:0] __reduce_max_13_valid_sink_count;
  reg [32-1:0] __reduce_max_13_valid_sink_offset_buf;
  reg [32-1:0] __reduce_max_13_valid_sink_stride_buf;
  reg [8-1:0] __reduce_max_13_valid_sink_ram_sel;
  reg [32-1:0] __reduce_max_13_valid_sink_waddr;
  reg __reduce_max_13_valid_sink_wenable;
  reg [1-1:0] __reduce_max_13_valid_sink_wdata;
  reg [32-1:0] _stream_conv2d_16_fsm;
  localparam _stream_conv2d_16_fsm_init = 0;
  wire _stream_conv2d_16_start_flag;
  reg _stream_conv2d_16_start;
  reg _stream_conv2d_16_end_flag;
  reg _stream_conv2d_16_term_sink;
  reg _stream_conv2d_16_source_busy;
  reg _stream_conv2d_16_sink_busy;
  reg [6-1:0] _stream_conv2d_16_constant_0_next_constant_data;
  reg [2-1:0] _stream_conv2d_16_constant_1_next_constant_data;
  reg [2-1:0] _stream_conv2d_16_constant_2_next_constant_data;
  reg [9-1:0] _stream_conv2d_16_constant_3_next_constant_data;
  reg [1-1:0] _stream_conv2d_16_constant_4_next_constant_data;
  reg _stream_conv2d_16_reduce_reset;
  reg [1-1:0] _stream_conv2d_16_constant_5_next_constant_data;
  reg _stream_conv2d_16_source_6_idle;
  reg [3-1:0] _stream_conv2d_16_source_6_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_6_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_6_source_size;
  reg [32-1:0] _stream_conv2d_16_source_6_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_6_source_count;
  reg [32-1:0] _stream_conv2d_16_source_6_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_6_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_6_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_6_source_ram_raddr;
  reg _stream_conv2d_16_source_6_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_6_source_ram_rdata;
  reg _stream_conv2d_16_source_6_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_6_source_empty_data;
  reg [1-1:0] _stream_conv2d_16_constant_7_next_constant_data;
  reg _stream_conv2d_16_source_8_idle;
  reg [3-1:0] _stream_conv2d_16_source_8_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_8_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_8_source_size;
  reg [32-1:0] _stream_conv2d_16_source_8_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_8_source_count;
  reg [32-1:0] _stream_conv2d_16_source_8_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_8_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_8_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_8_source_ram_raddr;
  reg _stream_conv2d_16_source_8_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_8_source_ram_rdata;
  reg _stream_conv2d_16_source_8_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_8_source_empty_data;
  reg [1-1:0] _stream_conv2d_16_constant_9_next_constant_data;
  reg _stream_conv2d_16_source_10_idle;
  reg [3-1:0] _stream_conv2d_16_source_10_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_10_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_10_source_size;
  reg [32-1:0] _stream_conv2d_16_source_10_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_10_source_count;
  reg [32-1:0] _stream_conv2d_16_source_10_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_10_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_10_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_10_source_ram_raddr;
  reg _stream_conv2d_16_source_10_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_10_source_ram_rdata;
  reg _stream_conv2d_16_source_10_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_10_source_empty_data;
  reg [1-1:0] _stream_conv2d_16_constant_11_next_constant_data;
  reg _stream_conv2d_16_source_12_idle;
  reg [3-1:0] _stream_conv2d_16_source_12_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_12_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_12_source_size;
  reg [32-1:0] _stream_conv2d_16_source_12_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_12_source_count;
  reg [32-1:0] _stream_conv2d_16_source_12_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_12_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_12_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_12_source_ram_raddr;
  reg _stream_conv2d_16_source_12_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_12_source_ram_rdata;
  reg _stream_conv2d_16_source_12_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_12_source_empty_data;
  reg [1-1:0] _stream_conv2d_16_constant_13_next_constant_data;
  reg _stream_conv2d_16_source_14_idle;
  reg [3-1:0] _stream_conv2d_16_source_14_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_14_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_14_source_size;
  reg [32-1:0] _stream_conv2d_16_source_14_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_14_source_count;
  reg [32-1:0] _stream_conv2d_16_source_14_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_14_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_14_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_14_source_ram_raddr;
  reg _stream_conv2d_16_source_14_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_14_source_ram_rdata;
  reg _stream_conv2d_16_source_14_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_14_source_empty_data;
  reg [1-1:0] _stream_conv2d_16_constant_15_next_constant_data;
  reg [1-1:0] _stream_conv2d_16_constant_16_next_constant_data;
  reg [4-1:0] _stream_conv2d_16_constant_17_next_constant_data;
  reg [1-1:0] _stream_conv2d_16_constant_18_next_constant_data;
  reg _stream_conv2d_16_source_19_idle;
  reg [3-1:0] _stream_conv2d_16_source_19_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_19_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_19_source_size;
  reg [32-1:0] _stream_conv2d_16_source_19_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_19_source_count;
  reg [32-1:0] _stream_conv2d_16_source_19_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_19_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_19_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_19_source_ram_raddr;
  reg _stream_conv2d_16_source_19_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_19_source_ram_rdata;
  reg _stream_conv2d_16_source_19_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_19_source_empty_data;
  reg _stream_conv2d_16_source_20_idle;
  reg [3-1:0] _stream_conv2d_16_source_20_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_20_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_20_source_size;
  reg [32-1:0] _stream_conv2d_16_source_20_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_20_source_count;
  reg [32-1:0] _stream_conv2d_16_source_20_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_20_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_20_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_20_source_ram_raddr;
  reg _stream_conv2d_16_source_20_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_20_source_ram_rdata;
  reg _stream_conv2d_16_source_20_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_20_source_empty_data;
  reg _stream_conv2d_16_source_21_idle;
  reg [3-1:0] _stream_conv2d_16_source_21_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_21_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_21_source_size;
  reg [32-1:0] _stream_conv2d_16_source_21_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_21_source_count;
  reg [32-1:0] _stream_conv2d_16_source_21_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_21_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_21_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_21_source_ram_raddr;
  reg _stream_conv2d_16_source_21_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_21_source_ram_rdata;
  reg _stream_conv2d_16_source_21_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_21_source_empty_data;
  reg _stream_conv2d_16_source_22_idle;
  reg [3-1:0] _stream_conv2d_16_source_22_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_22_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_22_source_size;
  reg [32-1:0] _stream_conv2d_16_source_22_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_22_source_count;
  reg [32-1:0] _stream_conv2d_16_source_22_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_22_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_22_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_22_source_ram_raddr;
  reg _stream_conv2d_16_source_22_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_22_source_ram_rdata;
  reg _stream_conv2d_16_source_22_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_22_source_empty_data;
  reg _stream_conv2d_16_source_23_idle;
  reg [3-1:0] _stream_conv2d_16_source_23_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_23_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_23_source_size;
  reg [32-1:0] _stream_conv2d_16_source_23_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_23_source_count;
  reg [32-1:0] _stream_conv2d_16_source_23_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_23_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_23_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_23_source_ram_raddr;
  reg _stream_conv2d_16_source_23_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_23_source_ram_rdata;
  reg _stream_conv2d_16_source_23_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_23_source_empty_data;
  reg _stream_conv2d_16_source_24_idle;
  reg [3-1:0] _stream_conv2d_16_source_24_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_24_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_24_source_size;
  reg [32-1:0] _stream_conv2d_16_source_24_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_24_source_count;
  reg [32-1:0] _stream_conv2d_16_source_24_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_24_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_24_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_24_source_ram_raddr;
  reg _stream_conv2d_16_source_24_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_24_source_ram_rdata;
  reg _stream_conv2d_16_source_24_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_24_source_empty_data;
  reg _stream_conv2d_16_source_25_idle;
  reg [3-1:0] _stream_conv2d_16_source_25_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_25_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_25_source_size;
  reg [32-1:0] _stream_conv2d_16_source_25_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_25_source_count;
  reg [32-1:0] _stream_conv2d_16_source_25_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_25_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_25_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_25_source_ram_raddr;
  reg _stream_conv2d_16_source_25_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_25_source_ram_rdata;
  reg _stream_conv2d_16_source_25_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_25_source_empty_data;
  reg _stream_conv2d_16_source_26_idle;
  reg [3-1:0] _stream_conv2d_16_source_26_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_26_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_26_source_size;
  reg [32-1:0] _stream_conv2d_16_source_26_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_26_source_count;
  reg [32-1:0] _stream_conv2d_16_source_26_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_26_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_26_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_26_source_ram_raddr;
  reg _stream_conv2d_16_source_26_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_26_source_ram_rdata;
  reg _stream_conv2d_16_source_26_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_26_source_empty_data;
  reg _stream_conv2d_16_source_27_idle;
  reg [3-1:0] _stream_conv2d_16_source_27_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_27_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_27_source_size;
  reg [32-1:0] _stream_conv2d_16_source_27_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_27_source_count;
  reg [32-1:0] _stream_conv2d_16_source_27_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_27_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_27_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_27_source_ram_raddr;
  reg _stream_conv2d_16_source_27_source_ram_renable;
  wire [8-1:0] _stream_conv2d_16_source_27_source_ram_rdata;
  reg _stream_conv2d_16_source_27_source_ram_rvalid;
  reg [8-1:0] _stream_conv2d_16_source_27_source_empty_data;
  reg _stream_conv2d_16_source_28_idle;
  reg [3-1:0] _stream_conv2d_16_source_28_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_28_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_28_source_size;
  reg [32-1:0] _stream_conv2d_16_source_28_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_28_source_count;
  reg [32-1:0] _stream_conv2d_16_source_28_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_28_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_28_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_28_source_ram_raddr;
  reg _stream_conv2d_16_source_28_source_ram_renable;
  wire [4-1:0] _stream_conv2d_16_source_28_source_ram_rdata;
  reg _stream_conv2d_16_source_28_source_ram_rvalid;
  reg [4-1:0] _stream_conv2d_16_source_28_source_empty_data;
  reg _stream_conv2d_16_source_29_idle;
  reg [3-1:0] _stream_conv2d_16_source_29_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_29_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_29_source_size;
  reg [32-1:0] _stream_conv2d_16_source_29_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_29_source_count;
  reg [32-1:0] _stream_conv2d_16_source_29_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_29_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_29_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_29_source_ram_raddr;
  reg _stream_conv2d_16_source_29_source_ram_renable;
  wire [4-1:0] _stream_conv2d_16_source_29_source_ram_rdata;
  reg _stream_conv2d_16_source_29_source_ram_rvalid;
  reg [4-1:0] _stream_conv2d_16_source_29_source_empty_data;
  reg _stream_conv2d_16_source_30_idle;
  reg [3-1:0] _stream_conv2d_16_source_30_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_30_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_30_source_size;
  reg [32-1:0] _stream_conv2d_16_source_30_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_30_source_count;
  reg [32-1:0] _stream_conv2d_16_source_30_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_30_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_30_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_30_source_ram_raddr;
  reg _stream_conv2d_16_source_30_source_ram_renable;
  wire [4-1:0] _stream_conv2d_16_source_30_source_ram_rdata;
  reg _stream_conv2d_16_source_30_source_ram_rvalid;
  reg [4-1:0] _stream_conv2d_16_source_30_source_empty_data;
  reg _stream_conv2d_16_source_31_idle;
  reg [3-1:0] _stream_conv2d_16_source_31_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_31_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_31_source_size;
  reg [32-1:0] _stream_conv2d_16_source_31_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_31_source_count;
  reg [32-1:0] _stream_conv2d_16_source_31_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_31_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_31_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_31_source_ram_raddr;
  reg _stream_conv2d_16_source_31_source_ram_renable;
  wire [4-1:0] _stream_conv2d_16_source_31_source_ram_rdata;
  reg _stream_conv2d_16_source_31_source_ram_rvalid;
  reg [4-1:0] _stream_conv2d_16_source_31_source_empty_data;
  reg _stream_conv2d_16_source_32_idle;
  reg [3-1:0] _stream_conv2d_16_source_32_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_32_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_32_source_size;
  reg [32-1:0] _stream_conv2d_16_source_32_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_32_source_count;
  reg [32-1:0] _stream_conv2d_16_source_32_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_32_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_32_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_32_source_ram_raddr;
  reg _stream_conv2d_16_source_32_source_ram_renable;
  wire [4-1:0] _stream_conv2d_16_source_32_source_ram_rdata;
  reg _stream_conv2d_16_source_32_source_ram_rvalid;
  reg [4-1:0] _stream_conv2d_16_source_32_source_empty_data;
  reg _stream_conv2d_16_source_33_idle;
  reg [3-1:0] _stream_conv2d_16_source_33_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_33_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_33_source_size;
  reg [32-1:0] _stream_conv2d_16_source_33_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_33_source_count;
  reg [32-1:0] _stream_conv2d_16_source_33_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_33_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_33_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_33_source_ram_raddr;
  reg _stream_conv2d_16_source_33_source_ram_renable;
  wire [4-1:0] _stream_conv2d_16_source_33_source_ram_rdata;
  reg _stream_conv2d_16_source_33_source_ram_rvalid;
  reg [4-1:0] _stream_conv2d_16_source_33_source_empty_data;
  reg _stream_conv2d_16_source_34_idle;
  reg [3-1:0] _stream_conv2d_16_source_34_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_34_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_34_source_size;
  reg [32-1:0] _stream_conv2d_16_source_34_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_34_source_count;
  reg [32-1:0] _stream_conv2d_16_source_34_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_34_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_34_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_34_source_ram_raddr;
  reg _stream_conv2d_16_source_34_source_ram_renable;
  wire [4-1:0] _stream_conv2d_16_source_34_source_ram_rdata;
  reg _stream_conv2d_16_source_34_source_ram_rvalid;
  reg [4-1:0] _stream_conv2d_16_source_34_source_empty_data;
  reg _stream_conv2d_16_source_35_idle;
  reg [3-1:0] _stream_conv2d_16_source_35_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_35_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_35_source_size;
  reg [32-1:0] _stream_conv2d_16_source_35_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_35_source_count;
  reg [32-1:0] _stream_conv2d_16_source_35_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_35_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_35_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_35_source_ram_raddr;
  reg _stream_conv2d_16_source_35_source_ram_renable;
  wire [4-1:0] _stream_conv2d_16_source_35_source_ram_rdata;
  reg _stream_conv2d_16_source_35_source_ram_rvalid;
  reg [4-1:0] _stream_conv2d_16_source_35_source_empty_data;
  reg _stream_conv2d_16_source_36_idle;
  reg [3-1:0] _stream_conv2d_16_source_36_source_mode;
  reg [32-1:0] _stream_conv2d_16_source_36_source_offset;
  reg [33-1:0] _stream_conv2d_16_source_36_source_size;
  reg [32-1:0] _stream_conv2d_16_source_36_source_stride;
  reg [33-1:0] _stream_conv2d_16_source_36_source_count;
  reg [32-1:0] _stream_conv2d_16_source_36_source_offset_buf;
  reg [32-1:0] _stream_conv2d_16_source_36_source_stride_buf;
  reg [8-1:0] _stream_conv2d_16_source_36_source_ram_sel;
  reg [32-1:0] _stream_conv2d_16_source_36_source_ram_raddr;
  reg _stream_conv2d_16_source_36_source_ram_renable;
  wire [4-1:0] _stream_conv2d_16_source_36_source_ram_rdata;
  reg _stream_conv2d_16_source_36_source_ram_rvalid;
  reg [4-1:0] _stream_conv2d_16_source_36_source_empty_data;
  wire signed [8-1:0] mul_4_x_data;
  wire signed [4-1:0] mul_4_y_data;
  wire [4-1:0] mul_4_rshift_data;
  reg [1-1:0] _greaterthan_data_57;
  reg [4-1:0] _minus_data_59;
  reg signed [8-1:0] __delay_data_594;
  reg signed [4-1:0] __delay_data_597;
  reg [4-1:0] __delay_data_600;
  reg signed [18-1:0] _sll_data_61;
  reg [1-1:0] __delay_data_593;
  reg signed [8-1:0] __delay_data_595;
  reg signed [4-1:0] __delay_data_598;
  reg [4-1:0] __delay_data_601;
  reg signed [12-1:0] _cond_data_67;
  reg signed [8-1:0] __delay_data_596;
  reg signed [4-1:0] __delay_data_599;
  reg [4-1:0] __delay_data_602;
  wire signed [12-1:0] __muladd_madd_odata_69;
  reg signed [12-1:0] __muladd_madd_odata_reg_69;
  wire signed [12-1:0] __muladd_data_69;
  assign __muladd_data_69 = __muladd_madd_odata_reg_69;
  wire __muladd_madd_update_69;
  assign __muladd_madd_update_69 = 1'd1;

  madd_0
  __muladd_madd_69
  (
    .CLK(CLK),
    .update(__muladd_madd_update_69),
    .a(__delay_data_596),
    .b(__delay_data_599),
    .c(_cond_data_67),
    .d(__muladd_madd_odata_69)
  );

  reg [4-1:0] __delay_data_603;
  reg [4-1:0] __delay_data_604;
  reg [4-1:0] __delay_data_605;
  reg [4-1:0] __delay_data_606;
  reg signed [12-1:0] _sra_data_70;
  wire signed [12-1:0] mul_4_z_data;
  assign mul_4_z_data = _sra_data_70;
  reg _substream_mul_4_x_data_cond_592_0;
  reg _substream_mul_4_y_data_cond_592_1;
  reg _substream_mul_4_rshift_data_cond_592_2;
  wire signed [8-1:0] mul_5_x_data;
  wire signed [4-1:0] mul_5_y_data;
  wire [4-1:0] mul_5_rshift_data;
  reg [1-1:0] _greaterthan_data_74;
  reg [4-1:0] _minus_data_76;
  reg signed [8-1:0] __delay_data_611;
  reg signed [4-1:0] __delay_data_614;
  reg [4-1:0] __delay_data_617;
  reg signed [18-1:0] _sll_data_78;
  reg [1-1:0] __delay_data_610;
  reg signed [8-1:0] __delay_data_612;
  reg signed [4-1:0] __delay_data_615;
  reg [4-1:0] __delay_data_618;
  reg signed [12-1:0] _cond_data_84;
  reg signed [8-1:0] __delay_data_613;
  reg signed [4-1:0] __delay_data_616;
  reg [4-1:0] __delay_data_619;
  wire signed [12-1:0] __muladd_madd_odata_86;
  reg signed [12-1:0] __muladd_madd_odata_reg_86;
  wire signed [12-1:0] __muladd_data_86;
  assign __muladd_data_86 = __muladd_madd_odata_reg_86;
  wire __muladd_madd_update_86;
  assign __muladd_madd_update_86 = 1'd1;

  madd_1
  __muladd_madd_86
  (
    .CLK(CLK),
    .update(__muladd_madd_update_86),
    .a(__delay_data_613),
    .b(__delay_data_616),
    .c(_cond_data_84),
    .d(__muladd_madd_odata_86)
  );

  reg [4-1:0] __delay_data_620;
  reg [4-1:0] __delay_data_621;
  reg [4-1:0] __delay_data_622;
  reg [4-1:0] __delay_data_623;
  reg signed [12-1:0] _sra_data_87;
  wire signed [12-1:0] mul_5_z_data;
  assign mul_5_z_data = _sra_data_87;
  reg _substream_mul_5_x_data_cond_609_3;
  reg _substream_mul_5_y_data_cond_609_4;
  reg _substream_mul_5_rshift_data_cond_609_5;
  wire signed [8-1:0] mul_6_x_data;
  wire signed [4-1:0] mul_6_y_data;
  wire [4-1:0] mul_6_rshift_data;
  reg [1-1:0] _greaterthan_data_91;
  reg [4-1:0] _minus_data_93;
  reg signed [8-1:0] __delay_data_628;
  reg signed [4-1:0] __delay_data_631;
  reg [4-1:0] __delay_data_634;
  reg signed [18-1:0] _sll_data_95;
  reg [1-1:0] __delay_data_627;
  reg signed [8-1:0] __delay_data_629;
  reg signed [4-1:0] __delay_data_632;
  reg [4-1:0] __delay_data_635;
  reg signed [12-1:0] _cond_data_101;
  reg signed [8-1:0] __delay_data_630;
  reg signed [4-1:0] __delay_data_633;
  reg [4-1:0] __delay_data_636;
  wire signed [12-1:0] __muladd_madd_odata_103;
  reg signed [12-1:0] __muladd_madd_odata_reg_103;
  wire signed [12-1:0] __muladd_data_103;
  assign __muladd_data_103 = __muladd_madd_odata_reg_103;
  wire __muladd_madd_update_103;
  assign __muladd_madd_update_103 = 1'd1;

  madd_2
  __muladd_madd_103
  (
    .CLK(CLK),
    .update(__muladd_madd_update_103),
    .a(__delay_data_630),
    .b(__delay_data_633),
    .c(_cond_data_101),
    .d(__muladd_madd_odata_103)
  );

  reg [4-1:0] __delay_data_637;
  reg [4-1:0] __delay_data_638;
  reg [4-1:0] __delay_data_639;
  reg [4-1:0] __delay_data_640;
  reg signed [12-1:0] _sra_data_104;
  wire signed [12-1:0] mul_6_z_data;
  assign mul_6_z_data = _sra_data_104;
  reg _substream_mul_6_x_data_cond_626_6;
  reg _substream_mul_6_y_data_cond_626_7;
  reg _substream_mul_6_rshift_data_cond_626_8;
  wire signed [8-1:0] mul_7_x_data;
  wire signed [4-1:0] mul_7_y_data;
  wire [4-1:0] mul_7_rshift_data;
  reg [1-1:0] _greaterthan_data_108;
  reg [4-1:0] _minus_data_110;
  reg signed [8-1:0] __delay_data_645;
  reg signed [4-1:0] __delay_data_648;
  reg [4-1:0] __delay_data_651;
  reg signed [18-1:0] _sll_data_112;
  reg [1-1:0] __delay_data_644;
  reg signed [8-1:0] __delay_data_646;
  reg signed [4-1:0] __delay_data_649;
  reg [4-1:0] __delay_data_652;
  reg signed [12-1:0] _cond_data_118;
  reg signed [8-1:0] __delay_data_647;
  reg signed [4-1:0] __delay_data_650;
  reg [4-1:0] __delay_data_653;
  wire signed [12-1:0] __muladd_madd_odata_120;
  reg signed [12-1:0] __muladd_madd_odata_reg_120;
  wire signed [12-1:0] __muladd_data_120;
  assign __muladd_data_120 = __muladd_madd_odata_reg_120;
  wire __muladd_madd_update_120;
  assign __muladd_madd_update_120 = 1'd1;

  madd_3
  __muladd_madd_120
  (
    .CLK(CLK),
    .update(__muladd_madd_update_120),
    .a(__delay_data_647),
    .b(__delay_data_650),
    .c(_cond_data_118),
    .d(__muladd_madd_odata_120)
  );

  reg [4-1:0] __delay_data_654;
  reg [4-1:0] __delay_data_655;
  reg [4-1:0] __delay_data_656;
  reg [4-1:0] __delay_data_657;
  reg signed [12-1:0] _sra_data_121;
  wire signed [12-1:0] mul_7_z_data;
  assign mul_7_z_data = _sra_data_121;
  reg _substream_mul_7_x_data_cond_643_9;
  reg _substream_mul_7_y_data_cond_643_10;
  reg _substream_mul_7_rshift_data_cond_643_11;
  wire signed [8-1:0] mul_8_x_data;
  wire signed [4-1:0] mul_8_y_data;
  wire [4-1:0] mul_8_rshift_data;
  reg [1-1:0] _greaterthan_data_125;
  reg [4-1:0] _minus_data_127;
  reg signed [8-1:0] __delay_data_662;
  reg signed [4-1:0] __delay_data_665;
  reg [4-1:0] __delay_data_668;
  reg signed [18-1:0] _sll_data_129;
  reg [1-1:0] __delay_data_661;
  reg signed [8-1:0] __delay_data_663;
  reg signed [4-1:0] __delay_data_666;
  reg [4-1:0] __delay_data_669;
  reg signed [12-1:0] _cond_data_135;
  reg signed [8-1:0] __delay_data_664;
  reg signed [4-1:0] __delay_data_667;
  reg [4-1:0] __delay_data_670;
  wire signed [12-1:0] __muladd_madd_odata_137;
  reg signed [12-1:0] __muladd_madd_odata_reg_137;
  wire signed [12-1:0] __muladd_data_137;
  assign __muladd_data_137 = __muladd_madd_odata_reg_137;
  wire __muladd_madd_update_137;
  assign __muladd_madd_update_137 = 1'd1;

  madd_4
  __muladd_madd_137
  (
    .CLK(CLK),
    .update(__muladd_madd_update_137),
    .a(__delay_data_664),
    .b(__delay_data_667),
    .c(_cond_data_135),
    .d(__muladd_madd_odata_137)
  );

  reg [4-1:0] __delay_data_671;
  reg [4-1:0] __delay_data_672;
  reg [4-1:0] __delay_data_673;
  reg [4-1:0] __delay_data_674;
  reg signed [12-1:0] _sra_data_138;
  wire signed [12-1:0] mul_8_z_data;
  assign mul_8_z_data = _sra_data_138;
  reg _substream_mul_8_x_data_cond_660_12;
  reg _substream_mul_8_y_data_cond_660_13;
  reg _substream_mul_8_rshift_data_cond_660_14;
  wire signed [8-1:0] mul_9_x_data;
  wire signed [4-1:0] mul_9_y_data;
  wire [4-1:0] mul_9_rshift_data;
  reg [1-1:0] _greaterthan_data_142;
  reg [4-1:0] _minus_data_144;
  reg signed [8-1:0] __delay_data_679;
  reg signed [4-1:0] __delay_data_682;
  reg [4-1:0] __delay_data_685;
  reg signed [18-1:0] _sll_data_146;
  reg [1-1:0] __delay_data_678;
  reg signed [8-1:0] __delay_data_680;
  reg signed [4-1:0] __delay_data_683;
  reg [4-1:0] __delay_data_686;
  reg signed [12-1:0] _cond_data_152;
  reg signed [8-1:0] __delay_data_681;
  reg signed [4-1:0] __delay_data_684;
  reg [4-1:0] __delay_data_687;
  wire signed [12-1:0] __muladd_madd_odata_154;
  reg signed [12-1:0] __muladd_madd_odata_reg_154;
  wire signed [12-1:0] __muladd_data_154;
  assign __muladd_data_154 = __muladd_madd_odata_reg_154;
  wire __muladd_madd_update_154;
  assign __muladd_madd_update_154 = 1'd1;

  madd_5
  __muladd_madd_154
  (
    .CLK(CLK),
    .update(__muladd_madd_update_154),
    .a(__delay_data_681),
    .b(__delay_data_684),
    .c(_cond_data_152),
    .d(__muladd_madd_odata_154)
  );

  reg [4-1:0] __delay_data_688;
  reg [4-1:0] __delay_data_689;
  reg [4-1:0] __delay_data_690;
  reg [4-1:0] __delay_data_691;
  reg signed [12-1:0] _sra_data_155;
  wire signed [12-1:0] mul_9_z_data;
  assign mul_9_z_data = _sra_data_155;
  reg _substream_mul_9_x_data_cond_677_15;
  reg _substream_mul_9_y_data_cond_677_16;
  reg _substream_mul_9_rshift_data_cond_677_17;
  wire signed [8-1:0] mul_10_x_data;
  wire signed [4-1:0] mul_10_y_data;
  wire [4-1:0] mul_10_rshift_data;
  reg [1-1:0] _greaterthan_data_159;
  reg [4-1:0] _minus_data_161;
  reg signed [8-1:0] __delay_data_696;
  reg signed [4-1:0] __delay_data_699;
  reg [4-1:0] __delay_data_702;
  reg signed [18-1:0] _sll_data_163;
  reg [1-1:0] __delay_data_695;
  reg signed [8-1:0] __delay_data_697;
  reg signed [4-1:0] __delay_data_700;
  reg [4-1:0] __delay_data_703;
  reg signed [12-1:0] _cond_data_169;
  reg signed [8-1:0] __delay_data_698;
  reg signed [4-1:0] __delay_data_701;
  reg [4-1:0] __delay_data_704;
  wire signed [12-1:0] __muladd_madd_odata_171;
  reg signed [12-1:0] __muladd_madd_odata_reg_171;
  wire signed [12-1:0] __muladd_data_171;
  assign __muladd_data_171 = __muladd_madd_odata_reg_171;
  wire __muladd_madd_update_171;
  assign __muladd_madd_update_171 = 1'd1;

  madd_6
  __muladd_madd_171
  (
    .CLK(CLK),
    .update(__muladd_madd_update_171),
    .a(__delay_data_698),
    .b(__delay_data_701),
    .c(_cond_data_169),
    .d(__muladd_madd_odata_171)
  );

  reg [4-1:0] __delay_data_705;
  reg [4-1:0] __delay_data_706;
  reg [4-1:0] __delay_data_707;
  reg [4-1:0] __delay_data_708;
  reg signed [12-1:0] _sra_data_172;
  wire signed [12-1:0] mul_10_z_data;
  assign mul_10_z_data = _sra_data_172;
  reg _substream_mul_10_x_data_cond_694_18;
  reg _substream_mul_10_y_data_cond_694_19;
  reg _substream_mul_10_rshift_data_cond_694_20;
  wire signed [8-1:0] mul_11_x_data;
  wire signed [4-1:0] mul_11_y_data;
  wire [4-1:0] mul_11_rshift_data;
  reg [1-1:0] _greaterthan_data_176;
  reg [4-1:0] _minus_data_178;
  reg signed [8-1:0] __delay_data_713;
  reg signed [4-1:0] __delay_data_716;
  reg [4-1:0] __delay_data_719;
  reg signed [18-1:0] _sll_data_180;
  reg [1-1:0] __delay_data_712;
  reg signed [8-1:0] __delay_data_714;
  reg signed [4-1:0] __delay_data_717;
  reg [4-1:0] __delay_data_720;
  reg signed [12-1:0] _cond_data_186;
  reg signed [8-1:0] __delay_data_715;
  reg signed [4-1:0] __delay_data_718;
  reg [4-1:0] __delay_data_721;
  wire signed [12-1:0] __muladd_madd_odata_188;
  reg signed [12-1:0] __muladd_madd_odata_reg_188;
  wire signed [12-1:0] __muladd_data_188;
  assign __muladd_data_188 = __muladd_madd_odata_reg_188;
  wire __muladd_madd_update_188;
  assign __muladd_madd_update_188 = 1'd1;

  madd_7
  __muladd_madd_188
  (
    .CLK(CLK),
    .update(__muladd_madd_update_188),
    .a(__delay_data_715),
    .b(__delay_data_718),
    .c(_cond_data_186),
    .d(__muladd_madd_odata_188)
  );

  reg [4-1:0] __delay_data_722;
  reg [4-1:0] __delay_data_723;
  reg [4-1:0] __delay_data_724;
  reg [4-1:0] __delay_data_725;
  reg signed [12-1:0] _sra_data_189;
  wire signed [12-1:0] mul_11_z_data;
  assign mul_11_z_data = _sra_data_189;
  reg _substream_mul_11_x_data_cond_711_21;
  reg _substream_mul_11_y_data_cond_711_22;
  reg _substream_mul_11_rshift_data_cond_711_23;
  wire signed [8-1:0] mul_12_x_data;
  wire signed [4-1:0] mul_12_y_data;
  wire [4-1:0] mul_12_rshift_data;
  reg [1-1:0] _greaterthan_data_193;
  reg [4-1:0] _minus_data_195;
  reg signed [8-1:0] __delay_data_730;
  reg signed [4-1:0] __delay_data_733;
  reg [4-1:0] __delay_data_736;
  reg signed [18-1:0] _sll_data_197;
  reg [1-1:0] __delay_data_729;
  reg signed [8-1:0] __delay_data_731;
  reg signed [4-1:0] __delay_data_734;
  reg [4-1:0] __delay_data_737;
  reg signed [12-1:0] _cond_data_203;
  reg signed [8-1:0] __delay_data_732;
  reg signed [4-1:0] __delay_data_735;
  reg [4-1:0] __delay_data_738;
  wire signed [12-1:0] __muladd_madd_odata_205;
  reg signed [12-1:0] __muladd_madd_odata_reg_205;
  wire signed [12-1:0] __muladd_data_205;
  assign __muladd_data_205 = __muladd_madd_odata_reg_205;
  wire __muladd_madd_update_205;
  assign __muladd_madd_update_205 = 1'd1;

  madd_8
  __muladd_madd_205
  (
    .CLK(CLK),
    .update(__muladd_madd_update_205),
    .a(__delay_data_732),
    .b(__delay_data_735),
    .c(_cond_data_203),
    .d(__muladd_madd_odata_205)
  );

  reg [4-1:0] __delay_data_739;
  reg [4-1:0] __delay_data_740;
  reg [4-1:0] __delay_data_741;
  reg [4-1:0] __delay_data_742;
  reg signed [12-1:0] _sra_data_206;
  wire signed [12-1:0] mul_12_z_data;
  assign mul_12_z_data = _sra_data_206;
  reg _substream_mul_12_x_data_cond_728_24;
  reg _substream_mul_12_y_data_cond_728_25;
  reg _substream_mul_12_rshift_data_cond_728_26;
  wire signed [32-1:0] add_tree_2_var0_data;
  wire signed [32-1:0] add_tree_2_var1_data;
  wire signed [32-1:0] add_tree_2_var2_data;
  wire signed [32-1:0] add_tree_2_var3_data;
  wire signed [32-1:0] add_tree_2_var4_data;
  wire signed [32-1:0] add_tree_2_var5_data;
  wire signed [32-1:0] add_tree_2_var6_data;
  wire signed [32-1:0] add_tree_2_var7_data;
  wire signed [32-1:0] add_tree_2_var8_data;
  reg signed [32-1:0] __plusn_data_34;
  reg signed [32-1:0] __plusn_data_35;
  reg signed [32-1:0] __plusn_data_36;
  reg signed [32-1:0] __plusn_data_37;
  wire signed [32-1:0] add_tree_2_sum_data;
  assign add_tree_2_sum_data = __plusn_data_37;
  reg _substream_add_tree_2_var0_data_cond_745_27;
  reg _substream_add_tree_2_var1_data_cond_745_28;
  reg _substream_add_tree_2_var2_data_cond_745_29;
  reg _substream_add_tree_2_var3_data_cond_745_30;
  reg _substream_add_tree_2_var4_data_cond_745_31;
  reg _substream_add_tree_2_var5_data_cond_745_32;
  reg _substream_add_tree_2_var6_data_cond_745_33;
  reg _substream_add_tree_2_var7_data_cond_745_34;
  reg _substream_add_tree_2_var8_data_cond_745_35;
  wire signed [32-1:0] acc_0_x_data;
  wire [6-1:0] acc_0_rshift_data;
  wire [32-1:0] acc_0_size_data;
  reg [1-1:0] _greaterthan_data_3;
  reg [6-1:0] _minus_data_5;
  reg signed [32-1:0] _reduceadd_data_17;
  reg [33-1:0] _reduceadd_count_17;
  reg [1-1:0] _pulse_data_19;
  reg [33-1:0] _pulse_count_19;
  reg [6-1:0] __delay_data_751;
  reg signed [66-1:0] _sll_data_7;
  reg [1-1:0] __delay_data_748;
  reg signed [32-1:0] __delay_data_749;
  reg [6-1:0] __delay_data_752;
  reg [1-1:0] __delay_data_755;
  reg signed [32-1:0] _cond_data_13;
  reg signed [32-1:0] __delay_data_750;
  reg [6-1:0] __delay_data_753;
  reg [1-1:0] __delay_data_756;
  reg signed [32-1:0] _plus_data_20;
  reg [6-1:0] __delay_data_754;
  reg [1-1:0] __delay_data_757;
  reg signed [32-1:0] _sra_data_21;
  reg [1-1:0] __delay_data_758;
  wire signed [32-1:0] acc_0_sum_data;
  assign acc_0_sum_data = _sra_data_21;
  wire [1-1:0] acc_0_valid_data;
  assign acc_0_valid_data = __delay_data_758;
  reg _substream_acc_0_x_data_cond_747_36;
  reg _substream_acc_0_rshift_data_cond_747_37;
  reg _substream_acc_0_size_data_cond_747_38;
  wire signed [32-1:0] mul_rshift_clip_3_x_data;
  wire signed [8-1:0] mul_rshift_clip_3_y_data;
  wire [6-1:0] mul_rshift_clip_3_rshift_data;
  wire signed [40-1:0] _times_mul_odata_41;
  reg signed [40-1:0] _times_mul_odata_reg_41;
  wire signed [40-1:0] _times_data_41;
  assign _times_data_41 = _times_mul_odata_reg_41;
  wire _times_mul_update_41;
  assign _times_mul_update_41 = 1'd1;

  multiplier_0
  _times_mul_41
  (
    .CLK(CLK),
    .update(_times_mul_update_41),
    .a(mul_rshift_clip_3_x_data),
    .b(mul_rshift_clip_3_y_data),
    .c(_times_mul_odata_41)
  );

  reg [6-1:0] __delay_data_764;
  reg [6-1:0] __delay_data_765;
  reg [6-1:0] __delay_data_766;
  reg [6-1:0] __delay_data_767;
  reg signed [40-1:0] _sra_data_42;
  reg [1-1:0] _greaterthan_data_43;
  reg [1-1:0] _lessthan_data_47;
  reg [1-1:0] _greatereq_data_51;
  reg signed [40-1:0] __delay_data_768;
  reg signed [40-1:0] _cond_data_45;
  reg signed [40-1:0] _cond_data_49;
  reg [1-1:0] __delay_data_769;
  reg signed [8-1:0] _cond_data_53;
  wire signed [8-1:0] mul_rshift_clip_3_z_data;
  assign mul_rshift_clip_3_z_data = _cond_data_53;
  reg _substream_mul_rshift_clip_3_x_data_cond_763_39;
  reg _substream_mul_rshift_clip_3_y_data_cond_763_40;
  reg _substream_mul_rshift_clip_3_rshift_data_cond_763_41;
  reg [3-1:0] _stream_conv2d_16_sink_37_sink_mode;
  reg [32-1:0] _stream_conv2d_16_sink_37_sink_offset;
  reg [33-1:0] _stream_conv2d_16_sink_37_sink_size;
  reg [32-1:0] _stream_conv2d_16_sink_37_sink_stride;
  reg [33-1:0] _stream_conv2d_16_sink_37_sink_count;
  reg [32-1:0] _stream_conv2d_16_sink_37_sink_offset_buf;
  reg [32-1:0] _stream_conv2d_16_sink_37_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_16_sink_37_sink_ram_sel;
  reg [32-1:0] _stream_conv2d_16_sink_37_sink_waddr;
  reg _stream_conv2d_16_sink_37_sink_wenable;
  reg [8-1:0] _stream_conv2d_16_sink_37_sink_wdata;
  reg [3-1:0] _stream_conv2d_16_sink_38_sink_mode;
  reg [32-1:0] _stream_conv2d_16_sink_38_sink_offset;
  reg [33-1:0] _stream_conv2d_16_sink_38_sink_size;
  reg [32-1:0] _stream_conv2d_16_sink_38_sink_stride;
  reg [33-1:0] _stream_conv2d_16_sink_38_sink_count;
  reg [32-1:0] _stream_conv2d_16_sink_38_sink_offset_buf;
  reg [32-1:0] _stream_conv2d_16_sink_38_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_16_sink_38_sink_ram_sel;
  reg [32-1:0] _stream_conv2d_16_sink_38_sink_waddr;
  reg _stream_conv2d_16_sink_38_sink_wenable;
  reg [1-1:0] _stream_conv2d_16_sink_38_sink_wdata;
  reg [32-1:0] _stream_max_pool_serial_18_fsm;
  localparam _stream_max_pool_serial_18_fsm_init = 0;
  wire _stream_max_pool_serial_18_start_flag;
  reg _stream_max_pool_serial_18_start;
  reg _stream_max_pool_serial_18_end_flag;
  reg _stream_max_pool_serial_18_term_sink;
  reg _stream_max_pool_serial_18_source_busy;
  reg _stream_max_pool_serial_18_sink_busy;
  reg [3-1:0] _stream_max_pool_serial_18_constant_0_next_constant_data;
  reg _stream_max_pool_serial_18_source_1_idle;
  reg [3-1:0] _stream_max_pool_serial_18_source_1_source_mode;
  reg [32-1:0] _stream_max_pool_serial_18_source_1_source_offset;
  reg [33-1:0] _stream_max_pool_serial_18_source_1_source_size;
  reg [32-1:0] _stream_max_pool_serial_18_source_1_source_stride;
  reg [33-1:0] _stream_max_pool_serial_18_source_1_source_count;
  reg [32-1:0] _stream_max_pool_serial_18_source_1_source_offset_buf;
  reg [32-1:0] _stream_max_pool_serial_18_source_1_source_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_18_source_1_source_ram_sel;
  reg [32-1:0] _stream_max_pool_serial_18_source_1_source_ram_raddr;
  reg _stream_max_pool_serial_18_source_1_source_ram_renable;
  wire [8-1:0] _stream_max_pool_serial_18_source_1_source_ram_rdata;
  reg _stream_max_pool_serial_18_source_1_source_ram_rvalid;
  reg [8-1:0] _stream_max_pool_serial_18_source_1_source_empty_data;
  reg [4-1:0] _stream_max_pool_serial_18_constant_2_next_constant_data;
  reg _stream_max_pool_serial_18_reduce_reset;
  wire signed [8-1:0] _reduce_max_13_x_data;
  wire [8-1:0] _reduce_max_13_size_data;
  reg signed [8-1:0] _reducemax_data_211;
  reg [9-1:0] _reducemax_count_211;
  reg [1-1:0] _pulse_data_213;
  reg [9-1:0] _pulse_count_213;
  wire signed [8-1:0] _reduce_max_13_data_data;
  assign _reduce_max_13_data_data = _reducemax_data_211;
  wire [1-1:0] _reduce_max_13_valid_data;
  assign _reduce_max_13_valid_data = _pulse_data_213;
  reg _substream__reduce_max_13_x_data_cond_792_42;
  reg _substream__reduce_max_13_size_data_cond_792_43;
  reg [3-1:0] _stream_max_pool_serial_18_sink_3_sink_mode;
  reg [32-1:0] _stream_max_pool_serial_18_sink_3_sink_offset;
  reg [33-1:0] _stream_max_pool_serial_18_sink_3_sink_size;
  reg [32-1:0] _stream_max_pool_serial_18_sink_3_sink_stride;
  reg [33-1:0] _stream_max_pool_serial_18_sink_3_sink_count;
  reg [32-1:0] _stream_max_pool_serial_18_sink_3_sink_offset_buf;
  reg [32-1:0] _stream_max_pool_serial_18_sink_3_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_18_sink_3_sink_ram_sel;
  reg [32-1:0] _stream_max_pool_serial_18_sink_3_sink_waddr;
  reg _stream_max_pool_serial_18_sink_3_sink_wenable;
  reg [8-1:0] _stream_max_pool_serial_18_sink_3_sink_wdata;
  reg [3-1:0] _stream_max_pool_serial_18_sink_4_sink_mode;
  reg [32-1:0] _stream_max_pool_serial_18_sink_4_sink_offset;
  reg [33-1:0] _stream_max_pool_serial_18_sink_4_sink_size;
  reg [32-1:0] _stream_max_pool_serial_18_sink_4_sink_stride;
  reg [33-1:0] _stream_max_pool_serial_18_sink_4_sink_count;
  reg [32-1:0] _stream_max_pool_serial_18_sink_4_sink_offset_buf;
  reg [32-1:0] _stream_max_pool_serial_18_sink_4_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_18_sink_4_sink_ram_sel;
  reg [32-1:0] _stream_max_pool_serial_18_sink_4_sink_waddr;
  reg _stream_max_pool_serial_18_sink_4_sink_wenable;
  reg [1-1:0] _stream_max_pool_serial_18_sink_4_sink_wdata;
  reg [32-1:0] _stream_matmul_29_fsm;
  localparam _stream_matmul_29_fsm_init = 0;
  wire _stream_matmul_29_start_flag;
  reg _stream_matmul_29_start;
  reg _stream_matmul_29_end_flag;
  reg _stream_matmul_29_term_sink;
  reg _stream_matmul_29_source_busy;
  reg _stream_matmul_29_sink_busy;
  reg [11-1:0] _stream_matmul_29_constant_0_next_constant_data;
  reg [1-1:0] _stream_matmul_29_constant_1_next_constant_data;
  reg [1-1:0] _stream_matmul_29_constant_2_next_constant_data;
  reg [1-1:0] _stream_matmul_29_constant_3_next_constant_data;
  reg [1-1:0] _stream_matmul_29_constant_4_next_constant_data;
  reg _stream_matmul_29_reduce_reset;
  reg [1-1:0] _stream_matmul_29_constant_5_next_constant_data;
  reg _stream_matmul_29_source_6_idle;
  reg [3-1:0] _stream_matmul_29_source_6_source_mode;
  reg [32-1:0] _stream_matmul_29_source_6_source_offset;
  reg [33-1:0] _stream_matmul_29_source_6_source_size;
  reg [32-1:0] _stream_matmul_29_source_6_source_stride;
  reg [33-1:0] _stream_matmul_29_source_6_source_count;
  reg [32-1:0] _stream_matmul_29_source_6_source_offset_buf;
  reg [32-1:0] _stream_matmul_29_source_6_source_stride_buf;
  reg [8-1:0] _stream_matmul_29_source_6_source_ram_sel;
  reg [32-1:0] _stream_matmul_29_source_6_source_ram_raddr;
  reg _stream_matmul_29_source_6_source_ram_renable;
  wire [8-1:0] _stream_matmul_29_source_6_source_ram_rdata;
  reg _stream_matmul_29_source_6_source_ram_rvalid;
  reg [8-1:0] _stream_matmul_29_source_6_source_empty_data;
  reg [1-1:0] _stream_matmul_29_constant_7_next_constant_data;
  reg _stream_matmul_29_source_8_idle;
  reg [3-1:0] _stream_matmul_29_source_8_source_mode;
  reg [32-1:0] _stream_matmul_29_source_8_source_offset;
  reg [33-1:0] _stream_matmul_29_source_8_source_size;
  reg [32-1:0] _stream_matmul_29_source_8_source_stride;
  reg [33-1:0] _stream_matmul_29_source_8_source_count;
  reg [32-1:0] _stream_matmul_29_source_8_source_offset_buf;
  reg [32-1:0] _stream_matmul_29_source_8_source_stride_buf;
  reg [8-1:0] _stream_matmul_29_source_8_source_ram_sel;
  reg [32-1:0] _stream_matmul_29_source_8_source_ram_raddr;
  reg _stream_matmul_29_source_8_source_ram_renable;
  wire [8-1:0] _stream_matmul_29_source_8_source_ram_rdata;
  reg _stream_matmul_29_source_8_source_ram_rvalid;
  reg [8-1:0] _stream_matmul_29_source_8_source_empty_data;
  reg [1-1:0] _stream_matmul_29_constant_9_next_constant_data;
  reg _stream_matmul_29_source_10_idle;
  reg [3-1:0] _stream_matmul_29_source_10_source_mode;
  reg [32-1:0] _stream_matmul_29_source_10_source_offset;
  reg [33-1:0] _stream_matmul_29_source_10_source_size;
  reg [32-1:0] _stream_matmul_29_source_10_source_stride;
  reg [33-1:0] _stream_matmul_29_source_10_source_count;
  reg [32-1:0] _stream_matmul_29_source_10_source_offset_buf;
  reg [32-1:0] _stream_matmul_29_source_10_source_stride_buf;
  reg [8-1:0] _stream_matmul_29_source_10_source_ram_sel;
  reg [32-1:0] _stream_matmul_29_source_10_source_ram_raddr;
  reg _stream_matmul_29_source_10_source_ram_renable;
  wire [8-1:0] _stream_matmul_29_source_10_source_ram_rdata;
  reg _stream_matmul_29_source_10_source_ram_rvalid;
  reg [8-1:0] _stream_matmul_29_source_10_source_empty_data;
  reg [1-1:0] _stream_matmul_29_constant_11_next_constant_data;
  reg _stream_matmul_29_source_12_idle;
  reg [3-1:0] _stream_matmul_29_source_12_source_mode;
  reg [32-1:0] _stream_matmul_29_source_12_source_offset;
  reg [33-1:0] _stream_matmul_29_source_12_source_size;
  reg [32-1:0] _stream_matmul_29_source_12_source_stride;
  reg [33-1:0] _stream_matmul_29_source_12_source_count;
  reg [32-1:0] _stream_matmul_29_source_12_source_offset_buf;
  reg [32-1:0] _stream_matmul_29_source_12_source_stride_buf;
  reg [8-1:0] _stream_matmul_29_source_12_source_ram_sel;
  reg [32-1:0] _stream_matmul_29_source_12_source_ram_raddr;
  reg _stream_matmul_29_source_12_source_ram_renable;
  wire [8-1:0] _stream_matmul_29_source_12_source_ram_rdata;
  reg _stream_matmul_29_source_12_source_ram_rvalid;
  reg [8-1:0] _stream_matmul_29_source_12_source_empty_data;
  reg [1-1:0] _stream_matmul_29_constant_13_next_constant_data;
  reg _stream_matmul_29_source_14_idle;
  reg [3-1:0] _stream_matmul_29_source_14_source_mode;
  reg [32-1:0] _stream_matmul_29_source_14_source_offset;
  reg [33-1:0] _stream_matmul_29_source_14_source_size;
  reg [32-1:0] _stream_matmul_29_source_14_source_stride;
  reg [33-1:0] _stream_matmul_29_source_14_source_count;
  reg [32-1:0] _stream_matmul_29_source_14_source_offset_buf;
  reg [32-1:0] _stream_matmul_29_source_14_source_stride_buf;
  reg [8-1:0] _stream_matmul_29_source_14_source_ram_sel;
  reg [32-1:0] _stream_matmul_29_source_14_source_ram_raddr;
  reg _stream_matmul_29_source_14_source_ram_renable;
  wire [8-1:0] _stream_matmul_29_source_14_source_ram_rdata;
  reg _stream_matmul_29_source_14_source_ram_rvalid;
  reg [8-1:0] _stream_matmul_29_source_14_source_empty_data;
  reg [1-1:0] _stream_matmul_29_constant_15_next_constant_data;
  reg [1-1:0] _stream_matmul_29_constant_16_next_constant_data;
  reg [4-1:0] _stream_matmul_29_constant_17_next_constant_data;
  reg [2-1:0] _stream_matmul_29_constant_18_next_constant_data;
  reg _stream_matmul_29_source_19_idle;
  reg [3-1:0] _stream_matmul_29_source_19_source_mode;
  reg [32-1:0] _stream_matmul_29_source_19_source_offset;
  reg [33-1:0] _stream_matmul_29_source_19_source_size;
  reg [32-1:0] _stream_matmul_29_source_19_source_stride;
  reg [33-1:0] _stream_matmul_29_source_19_source_count;
  reg [32-1:0] _stream_matmul_29_source_19_source_offset_buf;
  reg [32-1:0] _stream_matmul_29_source_19_source_stride_buf;
  reg [8-1:0] _stream_matmul_29_source_19_source_ram_sel;
  reg [32-1:0] _stream_matmul_29_source_19_source_ram_raddr;
  reg _stream_matmul_29_source_19_source_ram_renable;
  wire [8-1:0] _stream_matmul_29_source_19_source_ram_rdata;
  reg _stream_matmul_29_source_19_source_ram_rvalid;
  reg [8-1:0] _stream_matmul_29_source_19_source_empty_data;
  reg _stream_matmul_29_source_20_idle;
  reg [3-1:0] _stream_matmul_29_source_20_source_mode;
  reg [32-1:0] _stream_matmul_29_source_20_source_offset;
  reg [33-1:0] _stream_matmul_29_source_20_source_size;
  reg [32-1:0] _stream_matmul_29_source_20_source_stride;
  reg [33-1:0] _stream_matmul_29_source_20_source_count;
  reg [32-1:0] _stream_matmul_29_source_20_source_offset_buf;
  reg [32-1:0] _stream_matmul_29_source_20_source_stride_buf;
  reg [8-1:0] _stream_matmul_29_source_20_source_ram_sel;
  reg [32-1:0] _stream_matmul_29_source_20_source_ram_raddr;
  reg _stream_matmul_29_source_20_source_ram_renable;
  wire [4-1:0] _stream_matmul_29_source_20_source_ram_rdata;
  reg _stream_matmul_29_source_20_source_ram_rvalid;
  reg [4-1:0] _stream_matmul_29_source_20_source_empty_data;
  reg _substream_mul_4_x_data_cond_874_44;
  reg _substream_mul_4_y_data_cond_874_45;
  reg _substream_mul_4_rshift_data_cond_874_46;
  wire signed [32-1:0] add_tree_1_var0_data;
  wire signed [32-1:0] _cast_src_23;
  assign _cast_src_23 = add_tree_1_var0_data;
  wire signed [32-1:0] _cast_data_23;
  assign _cast_data_23 = _cast_src_23;
  wire signed [32-1:0] add_tree_1_sum_data;
  assign add_tree_1_sum_data = _cast_data_23;
  reg _substream_add_tree_1_var0_data_cond_877_47;
  reg _substream_acc_0_x_data_cond_879_48;
  reg _substream_acc_0_rshift_data_cond_879_49;
  reg _substream_acc_0_size_data_cond_879_50;
  reg _substream_mul_rshift_clip_3_x_data_cond_884_51;
  reg _substream_mul_rshift_clip_3_y_data_cond_884_52;
  reg _substream_mul_rshift_clip_3_rshift_data_cond_884_53;
  reg [3-1:0] _stream_matmul_29_sink_21_sink_mode;
  reg [32-1:0] _stream_matmul_29_sink_21_sink_offset;
  reg [33-1:0] _stream_matmul_29_sink_21_sink_size;
  reg [32-1:0] _stream_matmul_29_sink_21_sink_stride;
  reg [33-1:0] _stream_matmul_29_sink_21_sink_count;
  reg [32-1:0] _stream_matmul_29_sink_21_sink_offset_buf;
  reg [32-1:0] _stream_matmul_29_sink_21_sink_stride_buf;
  reg [8-1:0] _stream_matmul_29_sink_21_sink_ram_sel;
  reg [32-1:0] _stream_matmul_29_sink_21_sink_waddr;
  reg _stream_matmul_29_sink_21_sink_wenable;
  reg [8-1:0] _stream_matmul_29_sink_21_sink_wdata;
  reg [3-1:0] _stream_matmul_29_sink_22_sink_mode;
  reg [32-1:0] _stream_matmul_29_sink_22_sink_offset;
  reg [33-1:0] _stream_matmul_29_sink_22_sink_size;
  reg [32-1:0] _stream_matmul_29_sink_22_sink_stride;
  reg [33-1:0] _stream_matmul_29_sink_22_sink_count;
  reg [32-1:0] _stream_matmul_29_sink_22_sink_offset_buf;
  reg [32-1:0] _stream_matmul_29_sink_22_sink_stride_buf;
  reg [8-1:0] _stream_matmul_29_sink_22_sink_ram_sel;
  reg [32-1:0] _stream_matmul_29_sink_22_sink_waddr;
  reg _stream_matmul_29_sink_22_sink_wenable;
  reg [1-1:0] _stream_matmul_29_sink_22_sink_wdata;
  reg [32-1:0] main_fsm;
  localparam main_fsm_init = 0;
  reg [32-1:0] conv2d_16_objaddr;
  reg [32-1:0] conv2d_16_arg_objaddr_0;
  reg [32-1:0] conv2d_16_arg_objaddr_1;
  reg [32-1:0] conv2d_16_arg_objaddr_2;
  reg [32-1:0] conv2d_16_arg_objaddr_3;
  reg [32-1:0] control_conv2d_16;
  localparam control_conv2d_16_init = 0;
  reg _control_conv2d_16_called;
  wire signed [32-1:0] conv2d_16_act_base_offset;
  reg signed [32-1:0] conv2d_16_act_base_offset_row;
  reg signed [32-1:0] conv2d_16_act_base_offset_bat;
  assign conv2d_16_act_base_offset = conv2d_16_act_base_offset_row + conv2d_16_act_base_offset_bat;
  reg signed [32-1:0] conv2d_16_filter_base_offset;
  reg [32-1:0] conv2d_16_next_stream_num_ops;
  wire signed [32-1:0] conv2d_16_out_base_offset;
  reg signed [32-1:0] conv2d_16_out_base_offset_val;
  reg signed [32-1:0] conv2d_16_out_base_offset_col;
  reg signed [32-1:0] conv2d_16_out_base_offset_row;
  reg signed [32-1:0] conv2d_16_out_base_offset_bat;
  reg signed [32-1:0] conv2d_16_out_base_offset_och;
  assign conv2d_16_out_base_offset = conv2d_16_out_base_offset_val + conv2d_16_out_base_offset_col + conv2d_16_out_base_offset_row + conv2d_16_out_base_offset_bat + conv2d_16_out_base_offset_och;
  reg conv2d_16_dma_flag_0;
  reg conv2d_16_dma_flag_1;
  reg conv2d_16_dma_flag_2;
  reg [32-1:0] conv2d_16_sync_comp_count;
  reg [32-1:0] conv2d_16_sync_out_count;
  reg [32-1:0] conv2d_16_write_count;
  reg [32-1:0] conv2d_16_next_out_write_size;
  reg [32-1:0] conv2d_16_col_count;
  reg [32-1:0] conv2d_16_row_count;
  reg [32-1:0] conv2d_16_bat_count;
  reg [32-1:0] conv2d_16_och_count;
  reg [2-1:0] conv2d_16_col_select;
  reg [2-1:0] conv2d_16_row_select;
  reg [32-1:0] conv2d_16_out_col_count;
  reg [32-1:0] conv2d_16_out_row_count;
  reg [32-1:0] conv2d_16_out_ram_select;
  reg [32-1:0] conv2d_16_prev_col_count;
  reg [32-1:0] conv2d_16_prev_row_count;
  reg [32-1:0] conv2d_16_prev_bat_count;
  reg [32-1:0] conv2d_16_prev_och_count;
  reg [2-1:0] conv2d_16_prev_row_select;
  reg [32-1:0] conv2d_16_stream_act_local_0;
  reg [32-1:0] conv2d_16_stream_act_local_1;
  reg [32-1:0] conv2d_16_stream_act_local_2;
  reg [32-1:0] conv2d_16_stream_act_local_3;
  reg [32-1:0] conv2d_16_stream_act_local_4;
  reg [32-1:0] conv2d_16_stream_act_local_5;
  reg [32-1:0] conv2d_16_stream_act_local_6;
  reg [32-1:0] conv2d_16_stream_act_local_7;
  reg [32-1:0] conv2d_16_stream_act_local_8;
  reg [32-1:0] conv2d_16_stream_out_local_val;
  reg [32-1:0] conv2d_16_stream_out_local_col;
  wire [32-1:0] conv2d_16_stream_out_local;
  assign conv2d_16_stream_out_local = conv2d_16_stream_out_local_val + conv2d_16_stream_out_local_col;
  reg [32-1:0] conv2d_16_act_page_comp_offset_0;
  reg [32-1:0] conv2d_16_act_page_comp_offset_1;
  reg [32-1:0] conv2d_16_act_page_comp_offset_2;
  reg [32-1:0] conv2d_16_act_page_dma_offset_0;
  reg [32-1:0] conv2d_16_act_page_dma_offset_1;
  reg [32-1:0] conv2d_16_act_page_dma_offset_2;
  reg [32-1:0] conv2d_16_filter_page_comp_offset;
  reg [32-1:0] conv2d_16_filter_page_dma_offset;
  reg conv2d_16_out_page;
  reg [32-1:0] conv2d_16_out_page_comp_offset;
  reg [32-1:0] conv2d_16_out_page_dma_offset;
  reg [32-1:0] conv2d_16_out_laddr_offset;
  reg conv2d_16_skip_read_filter;
  reg conv2d_16_skip_read_act;
  reg conv2d_16_skip_comp;
  reg conv2d_16_skip_write_out;
  reg axim_flag_9;
  reg [32-1:0] _d1_control_conv2d_16;
  reg _control_conv2d_16_cond_3_0_1;
  reg _maxi_ram_w8_l2048_id1_1_read_start;
  reg [8-1:0] _maxi_ram_w8_l2048_id1_1_read_op_sel;
  reg [32-1:0] _maxi_ram_w8_l2048_id1_1_read_local_addr;
  reg [32-1:0] _maxi_ram_w8_l2048_id1_1_read_global_addr;
  reg [33-1:0] _maxi_ram_w8_l2048_id1_1_read_size;
  reg [32-1:0] _maxi_ram_w8_l2048_id1_1_read_local_stride;
  reg [32-1:0] _maxi_read_fsm;
  localparam _maxi_read_fsm_init = 0;
  reg [32-1:0] _maxi_read_cur_global_addr;
  reg [33-1:0] _maxi_read_cur_size;
  reg [33-1:0] _maxi_read_rest_size;
  reg [32-1:0] _wdata_10;
  reg _wvalid_11;
  reg [34-1:0] _tmp_12;
  reg _tmp_13;
  wire [8-1:0] _dataflow_slice_odata_3;
  wire _dataflow_slice_ovalid_3;
  wire _dataflow_slice_oready_3;
  assign _dataflow_slice_oready_3 = (_tmp_12 > 0) && !_tmp_13;
  reg _ram_w8_l2048_id1_0_cond_0_1;
  reg [34-1:0] _tmp_14;
  reg _tmp_15;
  wire [8-1:0] _dataflow_slice_odata_6;
  wire _dataflow_slice_ovalid_6;
  wire _dataflow_slice_oready_6;
  assign _dataflow_slice_oready_6 = (_tmp_14 > 0) && !_tmp_15;
  reg _ram_w8_l2048_id1_1_cond_0_1;
  reg [34-1:0] _tmp_16;
  reg _tmp_17;
  wire [8-1:0] _dataflow_slice_odata_9;
  wire _dataflow_slice_ovalid_9;
  wire _dataflow_slice_oready_9;
  assign _dataflow_slice_oready_9 = (_tmp_16 > 0) && !_tmp_17;
  reg _ram_w8_l2048_id1_2_cond_0_1;
  reg [34-1:0] _tmp_18;
  reg _tmp_19;
  wire [8-1:0] _dataflow_slice_odata_12;
  wire _dataflow_slice_ovalid_12;
  wire _dataflow_slice_oready_12;
  assign _dataflow_slice_oready_12 = (_tmp_18 > 0) && !_tmp_19;
  reg _ram_w8_l2048_id1_3_cond_0_1;
  reg [9-1:0] _tmp_20;
  reg _maxi_cond_0_1;
  assign maxi_rready = _maxi_read_fsm == 3;
  reg [32-1:0] _d1__maxi_read_fsm;
  reg __maxi_read_fsm_cond_3_0_1;
  reg axim_flag_21;
  reg __maxi_read_fsm_cond_4_1_1;
  reg axim_flag_22;
  reg _control_conv2d_16_cond_8_1_1;
  reg _maxi_ram_w8_l2048_id0_1_read_start;
  reg [8-1:0] _maxi_ram_w8_l2048_id0_1_read_op_sel;
  reg [32-1:0] _maxi_ram_w8_l2048_id0_1_read_local_addr;
  reg [32-1:0] _maxi_ram_w8_l2048_id0_1_read_global_addr;
  reg [33-1:0] _maxi_ram_w8_l2048_id0_1_read_size;
  reg [32-1:0] _maxi_ram_w8_l2048_id0_1_read_local_stride;
  reg [32-1:0] _wdata_23;
  reg _wvalid_24;
  reg [34-1:0] _tmp_25;
  reg _tmp_26;
  wire [8-1:0] _dataflow_slice_odata_16;
  wire _dataflow_slice_ovalid_16;
  wire _dataflow_slice_oready_16;
  assign _dataflow_slice_oready_16 = (_tmp_25 > 0) && !_tmp_26;
  reg _ram_w8_l2048_id0_0_cond_0_1;
  reg [34-1:0] _tmp_27;
  reg _tmp_28;
  wire [8-1:0] _dataflow_slice_odata_19;
  wire _dataflow_slice_ovalid_19;
  wire _dataflow_slice_oready_19;
  assign _dataflow_slice_oready_19 = (_tmp_27 > 0) && !_tmp_28;
  reg _ram_w8_l2048_id0_1_cond_0_1;
  reg [34-1:0] _tmp_29;
  reg _tmp_30;
  wire [8-1:0] _dataflow_slice_odata_22;
  wire _dataflow_slice_ovalid_22;
  wire _dataflow_slice_oready_22;
  assign _dataflow_slice_oready_22 = (_tmp_29 > 0) && !_tmp_30;
  reg _ram_w8_l2048_id0_2_cond_0_1;
  reg [34-1:0] _tmp_31;
  reg _tmp_32;
  wire [8-1:0] _dataflow_slice_odata_25;
  wire _dataflow_slice_ovalid_25;
  wire _dataflow_slice_oready_25;
  assign _dataflow_slice_oready_25 = (_tmp_31 > 0) && !_tmp_32;
  reg _ram_w8_l2048_id0_3_cond_0_1;
  reg __maxi_read_fsm_cond_3_2_1;
  reg [10-1:0] req_block_size_33;
  reg set_req_34;
  reg _control_conv2d_16_cond_14_2_1;
  reg axim_flag_35;
  reg _control_conv2d_16_cond_15_3_1;
  reg _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start;
  reg [8-1:0] _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_op_sel;
  reg [32-1:0] _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_addr;
  reg [32-1:0] _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_global_addr;
  reg [33-1:0] _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_size;
  reg [32-1:0] _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_stride;
  reg [32-1:0] _wdata_36;
  reg _wvalid_37;
  reg [11-1:0] _tmp_38;
  reg [34-1:0] _tmp_39;
  reg _tmp_40;
  wire [4-1:0] _dataflow_slice_odata_29;
  wire _dataflow_slice_ovalid_29;
  wire _dataflow_slice_oready_29;
  assign _dataflow_slice_oready_29 = (_tmp_39 > 0) && !_tmp_40;
  reg [10-1:0] _tmp_41;
  reg [10-1:0] _tmp_42;
  reg [10-1:0] _tmp_43;
  reg [10-1:0] _tmp_44;
  reg [10-1:0] _tmp_45;
  reg [10-1:0] _tmp_46;
  reg [10-1:0] _tmp_47;
  reg [10-1:0] _tmp_48;
  reg [10-1:0] _tmp_49;
  wire [10-1:0] _tmp_50;
  wire [10-1:0] _tmp_51;
  wire [10-1:0] _tmp_52;
  wire [10-1:0] _tmp_53;
  wire [10-1:0] _tmp_54;
  wire [10-1:0] _tmp_55;
  wire [10-1:0] _tmp_56;
  wire [10-1:0] _tmp_57;
  wire [10-1:0] _tmp_58;
  assign _tmp_50 = _tmp_41 + _maxi_read_local_stride;
  assign _tmp_51 = _tmp_42 + _maxi_read_local_stride;
  assign _tmp_52 = _tmp_43 + _maxi_read_local_stride;
  assign _tmp_53 = _tmp_44 + _maxi_read_local_stride;
  assign _tmp_54 = _tmp_45 + _maxi_read_local_stride;
  assign _tmp_55 = _tmp_46 + _maxi_read_local_stride;
  assign _tmp_56 = _tmp_47 + _maxi_read_local_stride;
  assign _tmp_57 = _tmp_48 + _maxi_read_local_stride;
  assign _tmp_58 = _tmp_49 + _maxi_read_local_stride;
  wire [10-1:0] _tmp_59;
  wire [10-1:0] _tmp_60;
  wire [10-1:0] _tmp_61;
  wire [10-1:0] _tmp_62;
  wire [10-1:0] _tmp_63;
  wire [10-1:0] _tmp_64;
  wire [10-1:0] _tmp_65;
  wire [10-1:0] _tmp_66;
  wire [10-1:0] _tmp_67;
  assign _tmp_59 = _tmp_50;
  assign _tmp_60 = _tmp_51;
  assign _tmp_61 = _tmp_52;
  assign _tmp_62 = _tmp_53;
  assign _tmp_63 = _tmp_54;
  assign _tmp_64 = _tmp_55;
  assign _tmp_65 = _tmp_56;
  assign _tmp_66 = _tmp_57;
  assign _tmp_67 = _tmp_58;
  reg [4-1:0] _tmp_68;
  reg _ram_w4_l8192_id0_0_cond_0_1;
  reg _ram_w4_l8192_id0_0_cond_1_1;
  reg _ram_w4_l8192_id1_0_cond_0_1;
  reg _ram_w4_l8192_id2_0_cond_0_1;
  reg _ram_w4_l8192_id3_0_cond_0_1;
  reg _ram_w4_l8192_id4_0_cond_0_1;
  reg _ram_w4_l8192_id5_0_cond_0_1;
  reg _ram_w4_l8192_id6_0_cond_0_1;
  reg _ram_w4_l8192_id7_0_cond_0_1;
  reg _ram_w4_l8192_id8_0_cond_0_1;
  reg [11-1:0] _tmp_69;
  reg [34-1:0] _tmp_70;
  reg _tmp_71;
  wire [4-1:0] _dataflow_slice_odata_32;
  wire _dataflow_slice_ovalid_32;
  wire _dataflow_slice_oready_32;
  assign _dataflow_slice_oready_32 = (_tmp_70 > 0) && !_tmp_71;
  reg [10-1:0] _tmp_72;
  reg [10-1:0] _tmp_73;
  reg [10-1:0] _tmp_74;
  reg [10-1:0] _tmp_75;
  reg [10-1:0] _tmp_76;
  reg [10-1:0] _tmp_77;
  reg [10-1:0] _tmp_78;
  reg [10-1:0] _tmp_79;
  reg [10-1:0] _tmp_80;
  wire [10-1:0] _tmp_81;
  wire [10-1:0] _tmp_82;
  wire [10-1:0] _tmp_83;
  wire [10-1:0] _tmp_84;
  wire [10-1:0] _tmp_85;
  wire [10-1:0] _tmp_86;
  wire [10-1:0] _tmp_87;
  wire [10-1:0] _tmp_88;
  wire [10-1:0] _tmp_89;
  assign _tmp_81 = _tmp_72 + _maxi_read_local_stride;
  assign _tmp_82 = _tmp_73 + _maxi_read_local_stride;
  assign _tmp_83 = _tmp_74 + _maxi_read_local_stride;
  assign _tmp_84 = _tmp_75 + _maxi_read_local_stride;
  assign _tmp_85 = _tmp_76 + _maxi_read_local_stride;
  assign _tmp_86 = _tmp_77 + _maxi_read_local_stride;
  assign _tmp_87 = _tmp_78 + _maxi_read_local_stride;
  assign _tmp_88 = _tmp_79 + _maxi_read_local_stride;
  assign _tmp_89 = _tmp_80 + _maxi_read_local_stride;
  wire [10-1:0] _tmp_90;
  wire [10-1:0] _tmp_91;
  wire [10-1:0] _tmp_92;
  wire [10-1:0] _tmp_93;
  wire [10-1:0] _tmp_94;
  wire [10-1:0] _tmp_95;
  wire [10-1:0] _tmp_96;
  wire [10-1:0] _tmp_97;
  wire [10-1:0] _tmp_98;
  assign _tmp_90 = _tmp_81;
  assign _tmp_91 = _tmp_82;
  assign _tmp_92 = _tmp_83;
  assign _tmp_93 = _tmp_84;
  assign _tmp_94 = _tmp_85;
  assign _tmp_95 = _tmp_86;
  assign _tmp_96 = _tmp_87;
  assign _tmp_97 = _tmp_88;
  assign _tmp_98 = _tmp_89;
  reg [4-1:0] _tmp_99;
  reg _ram_w4_l8192_id0_1_cond_0_1;
  reg _ram_w4_l8192_id0_1_cond_1_1;
  reg _ram_w4_l8192_id1_1_cond_0_1;
  reg _ram_w4_l8192_id2_1_cond_0_1;
  reg _ram_w4_l8192_id3_1_cond_0_1;
  reg _ram_w4_l8192_id4_1_cond_0_1;
  reg _ram_w4_l8192_id5_1_cond_0_1;
  reg _ram_w4_l8192_id6_1_cond_0_1;
  reg _ram_w4_l8192_id7_1_cond_0_1;
  reg _ram_w4_l8192_id8_1_cond_0_1;
  reg [11-1:0] _tmp_100;
  reg [34-1:0] _tmp_101;
  reg _tmp_102;
  wire [4-1:0] _dataflow_slice_odata_35;
  wire _dataflow_slice_ovalid_35;
  wire _dataflow_slice_oready_35;
  assign _dataflow_slice_oready_35 = (_tmp_101 > 0) && !_tmp_102;
  reg [10-1:0] _tmp_103;
  reg [10-1:0] _tmp_104;
  reg [10-1:0] _tmp_105;
  reg [10-1:0] _tmp_106;
  reg [10-1:0] _tmp_107;
  reg [10-1:0] _tmp_108;
  reg [10-1:0] _tmp_109;
  reg [10-1:0] _tmp_110;
  reg [10-1:0] _tmp_111;
  wire [10-1:0] _tmp_112;
  wire [10-1:0] _tmp_113;
  wire [10-1:0] _tmp_114;
  wire [10-1:0] _tmp_115;
  wire [10-1:0] _tmp_116;
  wire [10-1:0] _tmp_117;
  wire [10-1:0] _tmp_118;
  wire [10-1:0] _tmp_119;
  wire [10-1:0] _tmp_120;
  assign _tmp_112 = _tmp_103 + _maxi_read_local_stride;
  assign _tmp_113 = _tmp_104 + _maxi_read_local_stride;
  assign _tmp_114 = _tmp_105 + _maxi_read_local_stride;
  assign _tmp_115 = _tmp_106 + _maxi_read_local_stride;
  assign _tmp_116 = _tmp_107 + _maxi_read_local_stride;
  assign _tmp_117 = _tmp_108 + _maxi_read_local_stride;
  assign _tmp_118 = _tmp_109 + _maxi_read_local_stride;
  assign _tmp_119 = _tmp_110 + _maxi_read_local_stride;
  assign _tmp_120 = _tmp_111 + _maxi_read_local_stride;
  wire [10-1:0] _tmp_121;
  wire [10-1:0] _tmp_122;
  wire [10-1:0] _tmp_123;
  wire [10-1:0] _tmp_124;
  wire [10-1:0] _tmp_125;
  wire [10-1:0] _tmp_126;
  wire [10-1:0] _tmp_127;
  wire [10-1:0] _tmp_128;
  wire [10-1:0] _tmp_129;
  assign _tmp_121 = _tmp_112;
  assign _tmp_122 = _tmp_113;
  assign _tmp_123 = _tmp_114;
  assign _tmp_124 = _tmp_115;
  assign _tmp_125 = _tmp_116;
  assign _tmp_126 = _tmp_117;
  assign _tmp_127 = _tmp_118;
  assign _tmp_128 = _tmp_119;
  assign _tmp_129 = _tmp_120;
  reg [4-1:0] _tmp_130;
  reg _ram_w4_l8192_id0_2_cond_0_1;
  reg _ram_w4_l8192_id0_2_cond_1_1;
  reg _ram_w4_l8192_id1_2_cond_0_1;
  reg _ram_w4_l8192_id2_2_cond_0_1;
  reg _ram_w4_l8192_id3_2_cond_0_1;
  reg _ram_w4_l8192_id4_2_cond_0_1;
  reg _ram_w4_l8192_id5_2_cond_0_1;
  reg _ram_w4_l8192_id6_2_cond_0_1;
  reg _ram_w4_l8192_id7_2_cond_0_1;
  reg _ram_w4_l8192_id8_2_cond_0_1;
  reg [11-1:0] _tmp_131;
  reg [34-1:0] _tmp_132;
  reg _tmp_133;
  wire [4-1:0] _dataflow_slice_odata_38;
  wire _dataflow_slice_ovalid_38;
  wire _dataflow_slice_oready_38;
  assign _dataflow_slice_oready_38 = (_tmp_132 > 0) && !_tmp_133;
  reg [10-1:0] _tmp_134;
  reg [10-1:0] _tmp_135;
  reg [10-1:0] _tmp_136;
  reg [10-1:0] _tmp_137;
  reg [10-1:0] _tmp_138;
  reg [10-1:0] _tmp_139;
  reg [10-1:0] _tmp_140;
  reg [10-1:0] _tmp_141;
  reg [10-1:0] _tmp_142;
  wire [10-1:0] _tmp_143;
  wire [10-1:0] _tmp_144;
  wire [10-1:0] _tmp_145;
  wire [10-1:0] _tmp_146;
  wire [10-1:0] _tmp_147;
  wire [10-1:0] _tmp_148;
  wire [10-1:0] _tmp_149;
  wire [10-1:0] _tmp_150;
  wire [10-1:0] _tmp_151;
  assign _tmp_143 = _tmp_134 + _maxi_read_local_stride;
  assign _tmp_144 = _tmp_135 + _maxi_read_local_stride;
  assign _tmp_145 = _tmp_136 + _maxi_read_local_stride;
  assign _tmp_146 = _tmp_137 + _maxi_read_local_stride;
  assign _tmp_147 = _tmp_138 + _maxi_read_local_stride;
  assign _tmp_148 = _tmp_139 + _maxi_read_local_stride;
  assign _tmp_149 = _tmp_140 + _maxi_read_local_stride;
  assign _tmp_150 = _tmp_141 + _maxi_read_local_stride;
  assign _tmp_151 = _tmp_142 + _maxi_read_local_stride;
  wire [10-1:0] _tmp_152;
  wire [10-1:0] _tmp_153;
  wire [10-1:0] _tmp_154;
  wire [10-1:0] _tmp_155;
  wire [10-1:0] _tmp_156;
  wire [10-1:0] _tmp_157;
  wire [10-1:0] _tmp_158;
  wire [10-1:0] _tmp_159;
  wire [10-1:0] _tmp_160;
  assign _tmp_152 = _tmp_143;
  assign _tmp_153 = _tmp_144;
  assign _tmp_154 = _tmp_145;
  assign _tmp_155 = _tmp_146;
  assign _tmp_156 = _tmp_147;
  assign _tmp_157 = _tmp_148;
  assign _tmp_158 = _tmp_149;
  assign _tmp_159 = _tmp_150;
  assign _tmp_160 = _tmp_151;
  reg [4-1:0] _tmp_161;
  reg _ram_w4_l8192_id0_3_cond_0_1;
  reg _ram_w4_l8192_id0_3_cond_1_1;
  reg _ram_w4_l8192_id1_3_cond_0_1;
  reg _ram_w4_l8192_id2_3_cond_0_1;
  reg _ram_w4_l8192_id3_3_cond_0_1;
  reg _ram_w4_l8192_id4_3_cond_0_1;
  reg _ram_w4_l8192_id5_3_cond_0_1;
  reg _ram_w4_l8192_id6_3_cond_0_1;
  reg _ram_w4_l8192_id7_3_cond_0_1;
  reg _ram_w4_l8192_id8_3_cond_0_1;
  reg [11-1:0] _tmp_162;
  reg [34-1:0] _tmp_163;
  reg _tmp_164;
  wire [4-1:0] _dataflow_slice_odata_41;
  wire _dataflow_slice_ovalid_41;
  wire _dataflow_slice_oready_41;
  assign _dataflow_slice_oready_41 = (_tmp_163 > 0) && !_tmp_164;
  reg [10-1:0] _tmp_165;
  reg [10-1:0] _tmp_166;
  reg [10-1:0] _tmp_167;
  reg [10-1:0] _tmp_168;
  reg [10-1:0] _tmp_169;
  reg [10-1:0] _tmp_170;
  reg [10-1:0] _tmp_171;
  reg [10-1:0] _tmp_172;
  reg [10-1:0] _tmp_173;
  wire [10-1:0] _tmp_174;
  wire [10-1:0] _tmp_175;
  wire [10-1:0] _tmp_176;
  wire [10-1:0] _tmp_177;
  wire [10-1:0] _tmp_178;
  wire [10-1:0] _tmp_179;
  wire [10-1:0] _tmp_180;
  wire [10-1:0] _tmp_181;
  wire [10-1:0] _tmp_182;
  assign _tmp_174 = _tmp_165 + _maxi_read_local_stride;
  assign _tmp_175 = _tmp_166 + _maxi_read_local_stride;
  assign _tmp_176 = _tmp_167 + _maxi_read_local_stride;
  assign _tmp_177 = _tmp_168 + _maxi_read_local_stride;
  assign _tmp_178 = _tmp_169 + _maxi_read_local_stride;
  assign _tmp_179 = _tmp_170 + _maxi_read_local_stride;
  assign _tmp_180 = _tmp_171 + _maxi_read_local_stride;
  assign _tmp_181 = _tmp_172 + _maxi_read_local_stride;
  assign _tmp_182 = _tmp_173 + _maxi_read_local_stride;
  wire [10-1:0] _tmp_183;
  wire [10-1:0] _tmp_184;
  wire [10-1:0] _tmp_185;
  wire [10-1:0] _tmp_186;
  wire [10-1:0] _tmp_187;
  wire [10-1:0] _tmp_188;
  wire [10-1:0] _tmp_189;
  wire [10-1:0] _tmp_190;
  wire [10-1:0] _tmp_191;
  assign _tmp_183 = _tmp_174;
  assign _tmp_184 = _tmp_175;
  assign _tmp_185 = _tmp_176;
  assign _tmp_186 = _tmp_177;
  assign _tmp_187 = _tmp_178;
  assign _tmp_188 = _tmp_179;
  assign _tmp_189 = _tmp_180;
  assign _tmp_190 = _tmp_181;
  assign _tmp_191 = _tmp_182;
  reg [4-1:0] _tmp_192;
  reg _ram_w4_l8192_id0_4_cond_0_1;
  reg _ram_w4_l8192_id0_4_cond_1_1;
  reg _ram_w4_l8192_id1_4_cond_0_1;
  reg _ram_w4_l8192_id2_4_cond_0_1;
  reg _ram_w4_l8192_id3_4_cond_0_1;
  reg _ram_w4_l8192_id4_4_cond_0_1;
  reg _ram_w4_l8192_id5_4_cond_0_1;
  reg _ram_w4_l8192_id6_4_cond_0_1;
  reg _ram_w4_l8192_id7_4_cond_0_1;
  reg _ram_w4_l8192_id8_4_cond_0_1;
  reg [11-1:0] _tmp_193;
  reg [34-1:0] _tmp_194;
  reg _tmp_195;
  wire [4-1:0] _dataflow_slice_odata_44;
  wire _dataflow_slice_ovalid_44;
  wire _dataflow_slice_oready_44;
  assign _dataflow_slice_oready_44 = (_tmp_194 > 0) && !_tmp_195;
  reg [10-1:0] _tmp_196;
  reg [10-1:0] _tmp_197;
  reg [10-1:0] _tmp_198;
  reg [10-1:0] _tmp_199;
  reg [10-1:0] _tmp_200;
  reg [10-1:0] _tmp_201;
  reg [10-1:0] _tmp_202;
  reg [10-1:0] _tmp_203;
  reg [10-1:0] _tmp_204;
  wire [10-1:0] _tmp_205;
  wire [10-1:0] _tmp_206;
  wire [10-1:0] _tmp_207;
  wire [10-1:0] _tmp_208;
  wire [10-1:0] _tmp_209;
  wire [10-1:0] _tmp_210;
  wire [10-1:0] _tmp_211;
  wire [10-1:0] _tmp_212;
  wire [10-1:0] _tmp_213;
  assign _tmp_205 = _tmp_196 + _maxi_read_local_stride;
  assign _tmp_206 = _tmp_197 + _maxi_read_local_stride;
  assign _tmp_207 = _tmp_198 + _maxi_read_local_stride;
  assign _tmp_208 = _tmp_199 + _maxi_read_local_stride;
  assign _tmp_209 = _tmp_200 + _maxi_read_local_stride;
  assign _tmp_210 = _tmp_201 + _maxi_read_local_stride;
  assign _tmp_211 = _tmp_202 + _maxi_read_local_stride;
  assign _tmp_212 = _tmp_203 + _maxi_read_local_stride;
  assign _tmp_213 = _tmp_204 + _maxi_read_local_stride;
  wire [10-1:0] _tmp_214;
  wire [10-1:0] _tmp_215;
  wire [10-1:0] _tmp_216;
  wire [10-1:0] _tmp_217;
  wire [10-1:0] _tmp_218;
  wire [10-1:0] _tmp_219;
  wire [10-1:0] _tmp_220;
  wire [10-1:0] _tmp_221;
  wire [10-1:0] _tmp_222;
  assign _tmp_214 = _tmp_205;
  assign _tmp_215 = _tmp_206;
  assign _tmp_216 = _tmp_207;
  assign _tmp_217 = _tmp_208;
  assign _tmp_218 = _tmp_209;
  assign _tmp_219 = _tmp_210;
  assign _tmp_220 = _tmp_211;
  assign _tmp_221 = _tmp_212;
  assign _tmp_222 = _tmp_213;
  reg [4-1:0] _tmp_223;
  reg _ram_w4_l8192_id0_5_cond_0_1;
  reg _ram_w4_l8192_id0_5_cond_1_1;
  reg _ram_w4_l8192_id1_5_cond_0_1;
  reg _ram_w4_l8192_id2_5_cond_0_1;
  reg _ram_w4_l8192_id3_5_cond_0_1;
  reg _ram_w4_l8192_id4_5_cond_0_1;
  reg _ram_w4_l8192_id5_5_cond_0_1;
  reg _ram_w4_l8192_id6_5_cond_0_1;
  reg _ram_w4_l8192_id7_5_cond_0_1;
  reg _ram_w4_l8192_id8_5_cond_0_1;
  reg [11-1:0] _tmp_224;
  reg [34-1:0] _tmp_225;
  reg _tmp_226;
  wire [4-1:0] _dataflow_slice_odata_47;
  wire _dataflow_slice_ovalid_47;
  wire _dataflow_slice_oready_47;
  assign _dataflow_slice_oready_47 = (_tmp_225 > 0) && !_tmp_226;
  reg [10-1:0] _tmp_227;
  reg [10-1:0] _tmp_228;
  reg [10-1:0] _tmp_229;
  reg [10-1:0] _tmp_230;
  reg [10-1:0] _tmp_231;
  reg [10-1:0] _tmp_232;
  reg [10-1:0] _tmp_233;
  reg [10-1:0] _tmp_234;
  reg [10-1:0] _tmp_235;
  wire [10-1:0] _tmp_236;
  wire [10-1:0] _tmp_237;
  wire [10-1:0] _tmp_238;
  wire [10-1:0] _tmp_239;
  wire [10-1:0] _tmp_240;
  wire [10-1:0] _tmp_241;
  wire [10-1:0] _tmp_242;
  wire [10-1:0] _tmp_243;
  wire [10-1:0] _tmp_244;
  assign _tmp_236 = _tmp_227 + _maxi_read_local_stride;
  assign _tmp_237 = _tmp_228 + _maxi_read_local_stride;
  assign _tmp_238 = _tmp_229 + _maxi_read_local_stride;
  assign _tmp_239 = _tmp_230 + _maxi_read_local_stride;
  assign _tmp_240 = _tmp_231 + _maxi_read_local_stride;
  assign _tmp_241 = _tmp_232 + _maxi_read_local_stride;
  assign _tmp_242 = _tmp_233 + _maxi_read_local_stride;
  assign _tmp_243 = _tmp_234 + _maxi_read_local_stride;
  assign _tmp_244 = _tmp_235 + _maxi_read_local_stride;
  wire [10-1:0] _tmp_245;
  wire [10-1:0] _tmp_246;
  wire [10-1:0] _tmp_247;
  wire [10-1:0] _tmp_248;
  wire [10-1:0] _tmp_249;
  wire [10-1:0] _tmp_250;
  wire [10-1:0] _tmp_251;
  wire [10-1:0] _tmp_252;
  wire [10-1:0] _tmp_253;
  assign _tmp_245 = _tmp_236;
  assign _tmp_246 = _tmp_237;
  assign _tmp_247 = _tmp_238;
  assign _tmp_248 = _tmp_239;
  assign _tmp_249 = _tmp_240;
  assign _tmp_250 = _tmp_241;
  assign _tmp_251 = _tmp_242;
  assign _tmp_252 = _tmp_243;
  assign _tmp_253 = _tmp_244;
  reg [4-1:0] _tmp_254;
  reg _ram_w4_l8192_id0_6_cond_0_1;
  reg _ram_w4_l8192_id0_6_cond_1_1;
  reg _ram_w4_l8192_id1_6_cond_0_1;
  reg _ram_w4_l8192_id2_6_cond_0_1;
  reg _ram_w4_l8192_id3_6_cond_0_1;
  reg _ram_w4_l8192_id4_6_cond_0_1;
  reg _ram_w4_l8192_id5_6_cond_0_1;
  reg _ram_w4_l8192_id6_6_cond_0_1;
  reg _ram_w4_l8192_id7_6_cond_0_1;
  reg _ram_w4_l8192_id8_6_cond_0_1;
  reg [11-1:0] _tmp_255;
  reg [34-1:0] _tmp_256;
  reg _tmp_257;
  wire [4-1:0] _dataflow_slice_odata_50;
  wire _dataflow_slice_ovalid_50;
  wire _dataflow_slice_oready_50;
  assign _dataflow_slice_oready_50 = (_tmp_256 > 0) && !_tmp_257;
  reg [10-1:0] _tmp_258;
  reg [10-1:0] _tmp_259;
  reg [10-1:0] _tmp_260;
  reg [10-1:0] _tmp_261;
  reg [10-1:0] _tmp_262;
  reg [10-1:0] _tmp_263;
  reg [10-1:0] _tmp_264;
  reg [10-1:0] _tmp_265;
  reg [10-1:0] _tmp_266;
  wire [10-1:0] _tmp_267;
  wire [10-1:0] _tmp_268;
  wire [10-1:0] _tmp_269;
  wire [10-1:0] _tmp_270;
  wire [10-1:0] _tmp_271;
  wire [10-1:0] _tmp_272;
  wire [10-1:0] _tmp_273;
  wire [10-1:0] _tmp_274;
  wire [10-1:0] _tmp_275;
  assign _tmp_267 = _tmp_258 + _maxi_read_local_stride;
  assign _tmp_268 = _tmp_259 + _maxi_read_local_stride;
  assign _tmp_269 = _tmp_260 + _maxi_read_local_stride;
  assign _tmp_270 = _tmp_261 + _maxi_read_local_stride;
  assign _tmp_271 = _tmp_262 + _maxi_read_local_stride;
  assign _tmp_272 = _tmp_263 + _maxi_read_local_stride;
  assign _tmp_273 = _tmp_264 + _maxi_read_local_stride;
  assign _tmp_274 = _tmp_265 + _maxi_read_local_stride;
  assign _tmp_275 = _tmp_266 + _maxi_read_local_stride;
  wire [10-1:0] _tmp_276;
  wire [10-1:0] _tmp_277;
  wire [10-1:0] _tmp_278;
  wire [10-1:0] _tmp_279;
  wire [10-1:0] _tmp_280;
  wire [10-1:0] _tmp_281;
  wire [10-1:0] _tmp_282;
  wire [10-1:0] _tmp_283;
  wire [10-1:0] _tmp_284;
  assign _tmp_276 = _tmp_267;
  assign _tmp_277 = _tmp_268;
  assign _tmp_278 = _tmp_269;
  assign _tmp_279 = _tmp_270;
  assign _tmp_280 = _tmp_271;
  assign _tmp_281 = _tmp_272;
  assign _tmp_282 = _tmp_273;
  assign _tmp_283 = _tmp_274;
  assign _tmp_284 = _tmp_275;
  reg [4-1:0] _tmp_285;
  reg _ram_w4_l8192_id0_7_cond_0_1;
  reg _ram_w4_l8192_id0_7_cond_1_1;
  reg _ram_w4_l8192_id1_7_cond_0_1;
  reg _ram_w4_l8192_id2_7_cond_0_1;
  reg _ram_w4_l8192_id3_7_cond_0_1;
  reg _ram_w4_l8192_id4_7_cond_0_1;
  reg _ram_w4_l8192_id5_7_cond_0_1;
  reg _ram_w4_l8192_id6_7_cond_0_1;
  reg _ram_w4_l8192_id7_7_cond_0_1;
  reg _ram_w4_l8192_id8_7_cond_0_1;
  reg __maxi_read_fsm_cond_3_3_1;
  wire [32-1:0] conv2d_16_mux_act_gaddr_0;
  assign conv2d_16_mux_act_gaddr_0 = (conv2d_16_row_select == 0)? conv2d_16_arg_objaddr_0 + (conv2d_16_act_base_offset + cparam_conv2d_16_act_offset_values_0) : 
                                     (conv2d_16_row_select == 1)? conv2d_16_arg_objaddr_0 + (conv2d_16_act_base_offset + cparam_conv2d_16_act_offset_values_2) : 
                                     (conv2d_16_row_select == 2)? conv2d_16_arg_objaddr_0 + (conv2d_16_act_base_offset + cparam_conv2d_16_act_offset_values_1) : 1'd0;
  wire [32-1:0] conv2d_16_mux_act_gaddr_1;
  assign conv2d_16_mux_act_gaddr_1 = (conv2d_16_row_select == 0)? conv2d_16_arg_objaddr_0 + (conv2d_16_act_base_offset + cparam_conv2d_16_act_offset_values_1) : 
                                     (conv2d_16_row_select == 1)? conv2d_16_arg_objaddr_0 + (conv2d_16_act_base_offset + cparam_conv2d_16_act_offset_values_0) : 
                                     (conv2d_16_row_select == 2)? conv2d_16_arg_objaddr_0 + (conv2d_16_act_base_offset + cparam_conv2d_16_act_offset_values_2) : 1'd0;
  wire [32-1:0] conv2d_16_mux_act_gaddr_2;
  assign conv2d_16_mux_act_gaddr_2 = (conv2d_16_row_select == 0)? conv2d_16_arg_objaddr_0 + (conv2d_16_act_base_offset + cparam_conv2d_16_act_offset_values_2) : 
                                     (conv2d_16_row_select == 1)? conv2d_16_arg_objaddr_0 + (conv2d_16_act_base_offset + cparam_conv2d_16_act_offset_values_1) : 
                                     (conv2d_16_row_select == 2)? conv2d_16_arg_objaddr_0 + (conv2d_16_act_base_offset + cparam_conv2d_16_act_offset_values_0) : 1'd0;
  wire conv2d_16_dma_pad_mask_0;
  assign conv2d_16_dma_pad_mask_0 = (conv2d_16_row_count + 0 < cparam_conv2d_16_pad_row_top) || (conv2d_16_row_count + 0 >= cparam_conv2d_16_act_num_row + cparam_conv2d_16_pad_row_top);
  wire conv2d_16_dma_pad_mask_1;
  assign conv2d_16_dma_pad_mask_1 = (conv2d_16_row_count + 1 < cparam_conv2d_16_pad_row_top) || (conv2d_16_row_count + 1 >= cparam_conv2d_16_act_num_row + cparam_conv2d_16_pad_row_top);
  wire conv2d_16_dma_pad_mask_2;
  assign conv2d_16_dma_pad_mask_2 = (conv2d_16_row_count + 2 < cparam_conv2d_16_pad_row_top) || (conv2d_16_row_count + 2 >= cparam_conv2d_16_act_num_row + cparam_conv2d_16_pad_row_top);
  wire conv2d_16_mux_dma_pad_mask_0;
  assign conv2d_16_mux_dma_pad_mask_0 = (conv2d_16_row_select == 0)? conv2d_16_dma_pad_mask_0 : 
                                        (conv2d_16_row_select == 1)? conv2d_16_dma_pad_mask_2 : 
                                        (conv2d_16_row_select == 2)? conv2d_16_dma_pad_mask_1 : 1'd0;
  wire conv2d_16_mux_dma_pad_mask_1;
  assign conv2d_16_mux_dma_pad_mask_1 = (conv2d_16_row_select == 0)? conv2d_16_dma_pad_mask_1 : 
                                        (conv2d_16_row_select == 1)? conv2d_16_dma_pad_mask_0 : 
                                        (conv2d_16_row_select == 2)? conv2d_16_dma_pad_mask_2 : 1'd0;
  wire conv2d_16_mux_dma_pad_mask_2;
  assign conv2d_16_mux_dma_pad_mask_2 = (conv2d_16_row_select == 0)? conv2d_16_dma_pad_mask_2 : 
                                        (conv2d_16_row_select == 1)? conv2d_16_dma_pad_mask_1 : 
                                        (conv2d_16_row_select == 2)? conv2d_16_dma_pad_mask_0 : 1'd0;
  wire conv2d_16_mux_dma_flag_0;
  assign conv2d_16_mux_dma_flag_0 = (conv2d_16_prev_row_select == 0)? conv2d_16_dma_flag_0 : 
                                    (conv2d_16_prev_row_select == 1)? conv2d_16_dma_flag_2 : 
                                    (conv2d_16_prev_row_select == 2)? conv2d_16_dma_flag_1 : 1'd0;
  wire conv2d_16_mux_dma_flag_1;
  assign conv2d_16_mux_dma_flag_1 = (conv2d_16_prev_row_select == 0)? conv2d_16_dma_flag_1 : 
                                    (conv2d_16_prev_row_select == 1)? conv2d_16_dma_flag_0 : 
                                    (conv2d_16_prev_row_select == 2)? conv2d_16_dma_flag_2 : 1'd0;
  wire conv2d_16_mux_dma_flag_2;
  assign conv2d_16_mux_dma_flag_2 = (conv2d_16_prev_row_select == 0)? conv2d_16_dma_flag_2 : 
                                    (conv2d_16_prev_row_select == 1)? conv2d_16_dma_flag_1 : 
                                    (conv2d_16_prev_row_select == 2)? conv2d_16_dma_flag_0 : 1'd0;
  reg [9-1:0] req_block_size_286;
  reg set_req_287;
  reg _control_conv2d_16_cond_23_4_1;
  reg axim_flag_288;
  reg _control_conv2d_16_cond_24_5_1;
  reg _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start;
  reg [8-1:0] _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_op_sel;
  reg [32-1:0] _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_addr;
  reg [32-1:0] _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_global_addr;
  reg [33-1:0] _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_size;
  reg [32-1:0] _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_stride;
  reg [32-1:0] _wdata_289;
  reg _wvalid_290;
  reg [10-1:0] _tmp_291;
  reg [34-1:0] _tmp_292;
  reg _tmp_293;
  wire [8-1:0] _dataflow_slice_odata_54;
  wire _dataflow_slice_ovalid_54;
  wire _dataflow_slice_oready_54;
  assign _dataflow_slice_oready_54 = (_tmp_292 > 0) && !_tmp_293;
  reg [9-1:0] _tmp_294;
  reg [9-1:0] _tmp_295;
  reg [9-1:0] _tmp_296;
  wire [9-1:0] _tmp_297;
  wire [9-1:0] _tmp_298;
  wire [9-1:0] _tmp_299;
  assign _tmp_297 = _tmp_294 + _maxi_read_local_stride;
  assign _tmp_298 = _tmp_295 + _maxi_read_local_stride;
  assign _tmp_299 = _tmp_296 + _maxi_read_local_stride;
  wire [9-1:0] _tmp_300;
  wire [9-1:0] _tmp_301;
  wire [9-1:0] _tmp_302;
  assign _tmp_300 = _tmp_297;
  assign _tmp_301 = _tmp_298;
  assign _tmp_302 = _tmp_299;
  reg [2-1:0] _tmp_303;
  reg _ram_w8_l2048_id2_0_cond_0_1;
  reg _ram_w8_l2048_id2_0_cond_1_1;
  reg _ram_w8_l2048_id3_0_cond_0_1;
  reg _ram_w8_l2048_id4_0_cond_0_1;
  reg [10-1:0] _tmp_304;
  reg [34-1:0] _tmp_305;
  reg _tmp_306;
  wire [8-1:0] _dataflow_slice_odata_57;
  wire _dataflow_slice_ovalid_57;
  wire _dataflow_slice_oready_57;
  assign _dataflow_slice_oready_57 = (_tmp_305 > 0) && !_tmp_306;
  reg [9-1:0] _tmp_307;
  reg [9-1:0] _tmp_308;
  reg [9-1:0] _tmp_309;
  wire [9-1:0] _tmp_310;
  wire [9-1:0] _tmp_311;
  wire [9-1:0] _tmp_312;
  assign _tmp_310 = _tmp_307 + _maxi_read_local_stride;
  assign _tmp_311 = _tmp_308 + _maxi_read_local_stride;
  assign _tmp_312 = _tmp_309 + _maxi_read_local_stride;
  wire [9-1:0] _tmp_313;
  wire [9-1:0] _tmp_314;
  wire [9-1:0] _tmp_315;
  assign _tmp_313 = _tmp_310;
  assign _tmp_314 = _tmp_311;
  assign _tmp_315 = _tmp_312;
  reg [2-1:0] _tmp_316;
  reg _ram_w8_l2048_id2_1_cond_0_1;
  reg _ram_w8_l2048_id2_1_cond_1_1;
  reg _ram_w8_l2048_id3_1_cond_0_1;
  reg _ram_w8_l2048_id4_1_cond_0_1;
  reg [10-1:0] _tmp_317;
  reg [34-1:0] _tmp_318;
  reg _tmp_319;
  wire [8-1:0] _dataflow_slice_odata_60;
  wire _dataflow_slice_ovalid_60;
  wire _dataflow_slice_oready_60;
  assign _dataflow_slice_oready_60 = (_tmp_318 > 0) && !_tmp_319;
  reg [9-1:0] _tmp_320;
  reg [9-1:0] _tmp_321;
  reg [9-1:0] _tmp_322;
  wire [9-1:0] _tmp_323;
  wire [9-1:0] _tmp_324;
  wire [9-1:0] _tmp_325;
  assign _tmp_323 = _tmp_320 + _maxi_read_local_stride;
  assign _tmp_324 = _tmp_321 + _maxi_read_local_stride;
  assign _tmp_325 = _tmp_322 + _maxi_read_local_stride;
  wire [9-1:0] _tmp_326;
  wire [9-1:0] _tmp_327;
  wire [9-1:0] _tmp_328;
  assign _tmp_326 = _tmp_323;
  assign _tmp_327 = _tmp_324;
  assign _tmp_328 = _tmp_325;
  reg [2-1:0] _tmp_329;
  reg _ram_w8_l2048_id2_2_cond_0_1;
  reg _ram_w8_l2048_id2_2_cond_1_1;
  reg _ram_w8_l2048_id3_2_cond_0_1;
  reg _ram_w8_l2048_id4_2_cond_0_1;
  reg [10-1:0] _tmp_330;
  reg [34-1:0] _tmp_331;
  reg _tmp_332;
  wire [8-1:0] _dataflow_slice_odata_63;
  wire _dataflow_slice_ovalid_63;
  wire _dataflow_slice_oready_63;
  assign _dataflow_slice_oready_63 = (_tmp_331 > 0) && !_tmp_332;
  reg [9-1:0] _tmp_333;
  reg [9-1:0] _tmp_334;
  reg [9-1:0] _tmp_335;
  wire [9-1:0] _tmp_336;
  wire [9-1:0] _tmp_337;
  wire [9-1:0] _tmp_338;
  assign _tmp_336 = _tmp_333 + _maxi_read_local_stride;
  assign _tmp_337 = _tmp_334 + _maxi_read_local_stride;
  assign _tmp_338 = _tmp_335 + _maxi_read_local_stride;
  wire [9-1:0] _tmp_339;
  wire [9-1:0] _tmp_340;
  wire [9-1:0] _tmp_341;
  assign _tmp_339 = _tmp_336;
  assign _tmp_340 = _tmp_337;
  assign _tmp_341 = _tmp_338;
  reg [2-1:0] _tmp_342;
  reg _ram_w8_l2048_id2_3_cond_0_1;
  reg _ram_w8_l2048_id2_3_cond_1_1;
  reg _ram_w8_l2048_id3_3_cond_0_1;
  reg _ram_w8_l2048_id4_3_cond_0_1;
  reg __maxi_read_fsm_cond_3_4_1;
  reg [9-1:0] req_block_size_343;
  reg set_req_344;
  reg _control_conv2d_16_cond_30_6_1;
  reg axim_flag_345;
  reg _control_conv2d_16_cond_31_7_1;
  reg _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start;
  reg [8-1:0] _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_op_sel;
  reg [32-1:0] _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_addr;
  reg [32-1:0] _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_global_addr;
  reg [33-1:0] _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_size;
  reg [32-1:0] _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_stride;
  reg [32-1:0] _wdata_346;
  reg _wvalid_347;
  reg [10-1:0] _tmp_348;
  reg [34-1:0] _tmp_349;
  reg _tmp_350;
  wire [8-1:0] _dataflow_slice_odata_67;
  wire _dataflow_slice_ovalid_67;
  wire _dataflow_slice_oready_67;
  assign _dataflow_slice_oready_67 = (_tmp_349 > 0) && !_tmp_350;
  reg [9-1:0] _tmp_351;
  reg [9-1:0] _tmp_352;
  reg [9-1:0] _tmp_353;
  wire [9-1:0] _tmp_354;
  wire [9-1:0] _tmp_355;
  wire [9-1:0] _tmp_356;
  assign _tmp_354 = _tmp_351 + _maxi_read_local_stride;
  assign _tmp_355 = _tmp_352 + _maxi_read_local_stride;
  assign _tmp_356 = _tmp_353 + _maxi_read_local_stride;
  wire [9-1:0] _tmp_357;
  wire [9-1:0] _tmp_358;
  wire [9-1:0] _tmp_359;
  assign _tmp_357 = _tmp_354;
  assign _tmp_358 = _tmp_355;
  assign _tmp_359 = _tmp_356;
  reg [2-1:0] _tmp_360;
  reg _ram_w8_l2048_id5_0_cond_0_1;
  reg _ram_w8_l2048_id5_0_cond_1_1;
  reg _ram_w8_l2048_id6_0_cond_0_1;
  reg _ram_w8_l2048_id7_0_cond_0_1;
  reg [10-1:0] _tmp_361;
  reg [34-1:0] _tmp_362;
  reg _tmp_363;
  wire [8-1:0] _dataflow_slice_odata_70;
  wire _dataflow_slice_ovalid_70;
  wire _dataflow_slice_oready_70;
  assign _dataflow_slice_oready_70 = (_tmp_362 > 0) && !_tmp_363;
  reg [9-1:0] _tmp_364;
  reg [9-1:0] _tmp_365;
  reg [9-1:0] _tmp_366;
  wire [9-1:0] _tmp_367;
  wire [9-1:0] _tmp_368;
  wire [9-1:0] _tmp_369;
  assign _tmp_367 = _tmp_364 + _maxi_read_local_stride;
  assign _tmp_368 = _tmp_365 + _maxi_read_local_stride;
  assign _tmp_369 = _tmp_366 + _maxi_read_local_stride;
  wire [9-1:0] _tmp_370;
  wire [9-1:0] _tmp_371;
  wire [9-1:0] _tmp_372;
  assign _tmp_370 = _tmp_367;
  assign _tmp_371 = _tmp_368;
  assign _tmp_372 = _tmp_369;
  reg [2-1:0] _tmp_373;
  reg _ram_w8_l2048_id5_1_cond_0_1;
  reg _ram_w8_l2048_id5_1_cond_1_1;
  reg _ram_w8_l2048_id6_1_cond_0_1;
  reg _ram_w8_l2048_id7_1_cond_0_1;
  reg [10-1:0] _tmp_374;
  reg [34-1:0] _tmp_375;
  reg _tmp_376;
  wire [8-1:0] _dataflow_slice_odata_73;
  wire _dataflow_slice_ovalid_73;
  wire _dataflow_slice_oready_73;
  assign _dataflow_slice_oready_73 = (_tmp_375 > 0) && !_tmp_376;
  reg [9-1:0] _tmp_377;
  reg [9-1:0] _tmp_378;
  reg [9-1:0] _tmp_379;
  wire [9-1:0] _tmp_380;
  wire [9-1:0] _tmp_381;
  wire [9-1:0] _tmp_382;
  assign _tmp_380 = _tmp_377 + _maxi_read_local_stride;
  assign _tmp_381 = _tmp_378 + _maxi_read_local_stride;
  assign _tmp_382 = _tmp_379 + _maxi_read_local_stride;
  wire [9-1:0] _tmp_383;
  wire [9-1:0] _tmp_384;
  wire [9-1:0] _tmp_385;
  assign _tmp_383 = _tmp_380;
  assign _tmp_384 = _tmp_381;
  assign _tmp_385 = _tmp_382;
  reg [2-1:0] _tmp_386;
  reg _ram_w8_l2048_id5_2_cond_0_1;
  reg _ram_w8_l2048_id5_2_cond_1_1;
  reg _ram_w8_l2048_id6_2_cond_0_1;
  reg _ram_w8_l2048_id7_2_cond_0_1;
  reg [10-1:0] _tmp_387;
  reg [34-1:0] _tmp_388;
  reg _tmp_389;
  wire [8-1:0] _dataflow_slice_odata_76;
  wire _dataflow_slice_ovalid_76;
  wire _dataflow_slice_oready_76;
  assign _dataflow_slice_oready_76 = (_tmp_388 > 0) && !_tmp_389;
  reg [9-1:0] _tmp_390;
  reg [9-1:0] _tmp_391;
  reg [9-1:0] _tmp_392;
  wire [9-1:0] _tmp_393;
  wire [9-1:0] _tmp_394;
  wire [9-1:0] _tmp_395;
  assign _tmp_393 = _tmp_390 + _maxi_read_local_stride;
  assign _tmp_394 = _tmp_391 + _maxi_read_local_stride;
  assign _tmp_395 = _tmp_392 + _maxi_read_local_stride;
  wire [9-1:0] _tmp_396;
  wire [9-1:0] _tmp_397;
  wire [9-1:0] _tmp_398;
  assign _tmp_396 = _tmp_393;
  assign _tmp_397 = _tmp_394;
  assign _tmp_398 = _tmp_395;
  reg [2-1:0] _tmp_399;
  reg _ram_w8_l2048_id5_3_cond_0_1;
  reg _ram_w8_l2048_id5_3_cond_1_1;
  reg _ram_w8_l2048_id6_3_cond_0_1;
  reg _ram_w8_l2048_id7_3_cond_0_1;
  reg __maxi_read_fsm_cond_3_5_1;
  reg [9-1:0] req_block_size_400;
  reg set_req_401;
  reg _control_conv2d_16_cond_37_8_1;
  reg axim_flag_402;
  reg _control_conv2d_16_cond_38_9_1;
  reg _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start;
  reg [8-1:0] _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_op_sel;
  reg [32-1:0] _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_addr;
  reg [32-1:0] _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_global_addr;
  reg [33-1:0] _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_size;
  reg [32-1:0] _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_stride;
  reg [32-1:0] _wdata_403;
  reg _wvalid_404;
  reg [10-1:0] _tmp_405;
  reg [34-1:0] _tmp_406;
  reg _tmp_407;
  wire [8-1:0] _dataflow_slice_odata_80;
  wire _dataflow_slice_ovalid_80;
  wire _dataflow_slice_oready_80;
  assign _dataflow_slice_oready_80 = (_tmp_406 > 0) && !_tmp_407;
  reg [9-1:0] _tmp_408;
  reg [9-1:0] _tmp_409;
  reg [9-1:0] _tmp_410;
  wire [9-1:0] _tmp_411;
  wire [9-1:0] _tmp_412;
  wire [9-1:0] _tmp_413;
  assign _tmp_411 = _tmp_408 + _maxi_read_local_stride;
  assign _tmp_412 = _tmp_409 + _maxi_read_local_stride;
  assign _tmp_413 = _tmp_410 + _maxi_read_local_stride;
  wire [9-1:0] _tmp_414;
  wire [9-1:0] _tmp_415;
  wire [9-1:0] _tmp_416;
  assign _tmp_414 = _tmp_411;
  assign _tmp_415 = _tmp_412;
  assign _tmp_416 = _tmp_413;
  reg [2-1:0] _tmp_417;
  reg _ram_w8_l2048_id8_0_cond_0_1;
  reg _ram_w8_l2048_id8_0_cond_1_1;
  reg _ram_w8_l2048_id9_0_cond_0_1;
  reg _ram_w8_l2048_id10_0_cond_0_1;
  reg [10-1:0] _tmp_418;
  reg [34-1:0] _tmp_419;
  reg _tmp_420;
  wire [8-1:0] _dataflow_slice_odata_83;
  wire _dataflow_slice_ovalid_83;
  wire _dataflow_slice_oready_83;
  assign _dataflow_slice_oready_83 = (_tmp_419 > 0) && !_tmp_420;
  reg [9-1:0] _tmp_421;
  reg [9-1:0] _tmp_422;
  reg [9-1:0] _tmp_423;
  wire [9-1:0] _tmp_424;
  wire [9-1:0] _tmp_425;
  wire [9-1:0] _tmp_426;
  assign _tmp_424 = _tmp_421 + _maxi_read_local_stride;
  assign _tmp_425 = _tmp_422 + _maxi_read_local_stride;
  assign _tmp_426 = _tmp_423 + _maxi_read_local_stride;
  wire [9-1:0] _tmp_427;
  wire [9-1:0] _tmp_428;
  wire [9-1:0] _tmp_429;
  assign _tmp_427 = _tmp_424;
  assign _tmp_428 = _tmp_425;
  assign _tmp_429 = _tmp_426;
  reg [2-1:0] _tmp_430;
  reg _ram_w8_l2048_id8_1_cond_0_1;
  reg _ram_w8_l2048_id8_1_cond_1_1;
  reg _ram_w8_l2048_id9_1_cond_0_1;
  reg _ram_w8_l2048_id10_1_cond_0_1;
  reg [10-1:0] _tmp_431;
  reg [34-1:0] _tmp_432;
  reg _tmp_433;
  wire [8-1:0] _dataflow_slice_odata_86;
  wire _dataflow_slice_ovalid_86;
  wire _dataflow_slice_oready_86;
  assign _dataflow_slice_oready_86 = (_tmp_432 > 0) && !_tmp_433;
  reg [9-1:0] _tmp_434;
  reg [9-1:0] _tmp_435;
  reg [9-1:0] _tmp_436;
  wire [9-1:0] _tmp_437;
  wire [9-1:0] _tmp_438;
  wire [9-1:0] _tmp_439;
  assign _tmp_437 = _tmp_434 + _maxi_read_local_stride;
  assign _tmp_438 = _tmp_435 + _maxi_read_local_stride;
  assign _tmp_439 = _tmp_436 + _maxi_read_local_stride;
  wire [9-1:0] _tmp_440;
  wire [9-1:0] _tmp_441;
  wire [9-1:0] _tmp_442;
  assign _tmp_440 = _tmp_437;
  assign _tmp_441 = _tmp_438;
  assign _tmp_442 = _tmp_439;
  reg [2-1:0] _tmp_443;
  reg _ram_w8_l2048_id8_2_cond_0_1;
  reg _ram_w8_l2048_id8_2_cond_1_1;
  reg _ram_w8_l2048_id9_2_cond_0_1;
  reg _ram_w8_l2048_id10_2_cond_0_1;
  reg [10-1:0] _tmp_444;
  reg [34-1:0] _tmp_445;
  reg _tmp_446;
  wire [8-1:0] _dataflow_slice_odata_89;
  wire _dataflow_slice_ovalid_89;
  wire _dataflow_slice_oready_89;
  assign _dataflow_slice_oready_89 = (_tmp_445 > 0) && !_tmp_446;
  reg [9-1:0] _tmp_447;
  reg [9-1:0] _tmp_448;
  reg [9-1:0] _tmp_449;
  wire [9-1:0] _tmp_450;
  wire [9-1:0] _tmp_451;
  wire [9-1:0] _tmp_452;
  assign _tmp_450 = _tmp_447 + _maxi_read_local_stride;
  assign _tmp_451 = _tmp_448 + _maxi_read_local_stride;
  assign _tmp_452 = _tmp_449 + _maxi_read_local_stride;
  wire [9-1:0] _tmp_453;
  wire [9-1:0] _tmp_454;
  wire [9-1:0] _tmp_455;
  assign _tmp_453 = _tmp_450;
  assign _tmp_454 = _tmp_451;
  assign _tmp_455 = _tmp_452;
  reg [2-1:0] _tmp_456;
  reg _ram_w8_l2048_id8_3_cond_0_1;
  reg _ram_w8_l2048_id8_3_cond_1_1;
  reg _ram_w8_l2048_id9_3_cond_0_1;
  reg _ram_w8_l2048_id10_3_cond_0_1;
  reg __maxi_read_fsm_cond_3_6_1;
  reg [32-1:0] conv2d_16_comp_fsm;
  localparam conv2d_16_comp_fsm_init = 0;
  reg [32-1:0] conv2d_16_filter_page_comp_offset_buf;
  reg [32-1:0] conv2d_16_act_page_comp_offset_buf_0;
  reg [32-1:0] conv2d_16_act_page_comp_offset_buf_1;
  reg [32-1:0] conv2d_16_act_page_comp_offset_buf_2;
  reg [32-1:0] conv2d_16_out_page_comp_offset_buf;
  reg [32-1:0] conv2d_16_row_count_buf;
  reg [2-1:0] conv2d_16_row_select_buf;
  reg [32-1:0] conv2d_16_och_count_buf;
  wire conv2d_16_stream_pad_mask_0_0;
  assign conv2d_16_stream_pad_mask_0_0 = (conv2d_16_col_count + 0 < cparam_conv2d_16_pad_col_left) || (conv2d_16_col_count + 0 >= cparam_conv2d_16_act_num_col + cparam_conv2d_16_pad_col_left) || (conv2d_16_row_count_buf + 0 < cparam_conv2d_16_pad_row_top) || (conv2d_16_row_count_buf + 0 >= cparam_conv2d_16_act_num_row + cparam_conv2d_16_pad_row_top);
  wire conv2d_16_stream_pad_mask_0_1;
  assign conv2d_16_stream_pad_mask_0_1 = (conv2d_16_col_count + 1 < cparam_conv2d_16_pad_col_left) || (conv2d_16_col_count + 1 >= cparam_conv2d_16_act_num_col + cparam_conv2d_16_pad_col_left) || (conv2d_16_row_count_buf + 0 < cparam_conv2d_16_pad_row_top) || (conv2d_16_row_count_buf + 0 >= cparam_conv2d_16_act_num_row + cparam_conv2d_16_pad_row_top);
  wire conv2d_16_stream_pad_mask_0_2;
  assign conv2d_16_stream_pad_mask_0_2 = (conv2d_16_col_count + 2 < cparam_conv2d_16_pad_col_left) || (conv2d_16_col_count + 2 >= cparam_conv2d_16_act_num_col + cparam_conv2d_16_pad_col_left) || (conv2d_16_row_count_buf + 0 < cparam_conv2d_16_pad_row_top) || (conv2d_16_row_count_buf + 0 >= cparam_conv2d_16_act_num_row + cparam_conv2d_16_pad_row_top);
  wire conv2d_16_stream_pad_mask_1_0;
  assign conv2d_16_stream_pad_mask_1_0 = (conv2d_16_col_count + 0 < cparam_conv2d_16_pad_col_left) || (conv2d_16_col_count + 0 >= cparam_conv2d_16_act_num_col + cparam_conv2d_16_pad_col_left) || (conv2d_16_row_count_buf + 1 < cparam_conv2d_16_pad_row_top) || (conv2d_16_row_count_buf + 1 >= cparam_conv2d_16_act_num_row + cparam_conv2d_16_pad_row_top);
  wire conv2d_16_stream_pad_mask_1_1;
  assign conv2d_16_stream_pad_mask_1_1 = (conv2d_16_col_count + 1 < cparam_conv2d_16_pad_col_left) || (conv2d_16_col_count + 1 >= cparam_conv2d_16_act_num_col + cparam_conv2d_16_pad_col_left) || (conv2d_16_row_count_buf + 1 < cparam_conv2d_16_pad_row_top) || (conv2d_16_row_count_buf + 1 >= cparam_conv2d_16_act_num_row + cparam_conv2d_16_pad_row_top);
  wire conv2d_16_stream_pad_mask_1_2;
  assign conv2d_16_stream_pad_mask_1_2 = (conv2d_16_col_count + 2 < cparam_conv2d_16_pad_col_left) || (conv2d_16_col_count + 2 >= cparam_conv2d_16_act_num_col + cparam_conv2d_16_pad_col_left) || (conv2d_16_row_count_buf + 1 < cparam_conv2d_16_pad_row_top) || (conv2d_16_row_count_buf + 1 >= cparam_conv2d_16_act_num_row + cparam_conv2d_16_pad_row_top);
  wire conv2d_16_stream_pad_mask_2_0;
  assign conv2d_16_stream_pad_mask_2_0 = (conv2d_16_col_count + 0 < cparam_conv2d_16_pad_col_left) || (conv2d_16_col_count + 0 >= cparam_conv2d_16_act_num_col + cparam_conv2d_16_pad_col_left) || (conv2d_16_row_count_buf + 2 < cparam_conv2d_16_pad_row_top) || (conv2d_16_row_count_buf + 2 >= cparam_conv2d_16_act_num_row + cparam_conv2d_16_pad_row_top);
  wire conv2d_16_stream_pad_mask_2_1;
  assign conv2d_16_stream_pad_mask_2_1 = (conv2d_16_col_count + 1 < cparam_conv2d_16_pad_col_left) || (conv2d_16_col_count + 1 >= cparam_conv2d_16_act_num_col + cparam_conv2d_16_pad_col_left) || (conv2d_16_row_count_buf + 2 < cparam_conv2d_16_pad_row_top) || (conv2d_16_row_count_buf + 2 >= cparam_conv2d_16_act_num_row + cparam_conv2d_16_pad_row_top);
  wire conv2d_16_stream_pad_mask_2_2;
  assign conv2d_16_stream_pad_mask_2_2 = (conv2d_16_col_count + 2 < cparam_conv2d_16_pad_col_left) || (conv2d_16_col_count + 2 >= cparam_conv2d_16_act_num_col + cparam_conv2d_16_pad_col_left) || (conv2d_16_row_count_buf + 2 < cparam_conv2d_16_pad_row_top) || (conv2d_16_row_count_buf + 2 >= cparam_conv2d_16_act_num_row + cparam_conv2d_16_pad_row_top);
  reg [9-1:0] conv2d_16_stream_pad_masks;
  wire [6-1:0] stream_conv2d_16_constant_0_data;
  wire [2-1:0] stream_conv2d_16_constant_1_data;
  wire [2-1:0] stream_conv2d_16_constant_2_data;
  wire [9-1:0] stream_conv2d_16_constant_3_data;
  wire [1-1:0] stream_conv2d_16_constant_4_data;
  wire [1-1:0] stream_conv2d_16_constant_5_data;
  wire [8-1:0] stream_conv2d_16_source_6_data;
  wire [1-1:0] stream_conv2d_16_constant_7_data;
  wire [8-1:0] stream_conv2d_16_source_8_data;
  wire [1-1:0] stream_conv2d_16_constant_9_data;
  wire [8-1:0] stream_conv2d_16_source_10_data;
  wire [1-1:0] stream_conv2d_16_constant_11_data;
  wire [8-1:0] stream_conv2d_16_source_12_data;
  wire [1-1:0] stream_conv2d_16_constant_13_data;
  wire [8-1:0] stream_conv2d_16_source_14_data;
  wire [1-1:0] stream_conv2d_16_constant_15_data;
  wire [1-1:0] stream_conv2d_16_constant_16_data;
  wire [4-1:0] stream_conv2d_16_constant_17_data;
  wire [1-1:0] stream_conv2d_16_constant_18_data;
  wire [8-1:0] stream_conv2d_16_source_19_data;
  wire [8-1:0] stream_conv2d_16_source_20_data;
  wire [8-1:0] stream_conv2d_16_source_21_data;
  wire [8-1:0] stream_conv2d_16_source_22_data;
  wire [8-1:0] stream_conv2d_16_source_23_data;
  wire [8-1:0] stream_conv2d_16_source_24_data;
  wire [8-1:0] stream_conv2d_16_source_25_data;
  wire [8-1:0] stream_conv2d_16_source_26_data;
  wire [8-1:0] stream_conv2d_16_source_27_data;
  wire [4-1:0] stream_conv2d_16_source_28_data;
  wire [4-1:0] stream_conv2d_16_source_29_data;
  wire [4-1:0] stream_conv2d_16_source_30_data;
  wire [4-1:0] stream_conv2d_16_source_31_data;
  wire [4-1:0] stream_conv2d_16_source_32_data;
  wire [4-1:0] stream_conv2d_16_source_33_data;
  wire [4-1:0] stream_conv2d_16_source_34_data;
  wire [4-1:0] stream_conv2d_16_source_35_data;
  wire [4-1:0] stream_conv2d_16_source_36_data;
  wire [8-1:0] _slice_data_233;
  assign _slice_data_233 = stream_conv2d_16_source_6_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_234;
  assign _reinterpretcast_src_234 = _slice_data_233;
  wire signed [8-1:0] _reinterpretcast_data_234;
  assign _reinterpretcast_data_234 = _reinterpretcast_src_234;
  reg signed [8-1:0] _cond_data_235;
  wire [8-1:0] _slice_data_240;
  assign _slice_data_240 = stream_conv2d_16_source_8_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_241;
  assign _reinterpretcast_src_241 = _slice_data_240;
  wire signed [8-1:0] _reinterpretcast_data_241;
  assign _reinterpretcast_data_241 = _reinterpretcast_src_241;
  reg signed [8-1:0] _cond_data_242;
  wire [8-1:0] _slice_data_247;
  assign _slice_data_247 = stream_conv2d_16_source_10_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_248;
  assign _reinterpretcast_src_248 = _slice_data_247;
  wire [8-1:0] _reinterpretcast_data_248;
  assign _reinterpretcast_data_248 = _reinterpretcast_src_248;
  reg [8-1:0] _cond_data_249;
  wire [8-1:0] _slice_data_254;
  assign _slice_data_254 = stream_conv2d_16_source_12_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_255;
  assign _reinterpretcast_src_255 = _slice_data_254;
  wire [8-1:0] _reinterpretcast_data_255;
  assign _reinterpretcast_data_255 = _reinterpretcast_src_255;
  reg [8-1:0] _cond_data_256;
  wire [8-1:0] _slice_data_261;
  assign _slice_data_261 = stream_conv2d_16_source_14_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_262;
  assign _reinterpretcast_src_262 = _slice_data_261;
  wire [8-1:0] _reinterpretcast_data_262;
  assign _reinterpretcast_data_262 = _reinterpretcast_src_262;
  reg [8-1:0] _cond_data_263;
  reg [1-1:0] _eq_data_277;
  reg [1-1:0] _eq_data_281;
  reg [1-1:0] _eq_data_284;
  reg [1-1:0] _eq_data_287;
  reg [1-1:0] _eq_data_291;
  reg [1-1:0] _eq_data_294;
  reg [1-1:0] _eq_data_297;
  reg [1-1:0] _eq_data_301;
  reg [1-1:0] _eq_data_304;
  reg [1-1:0] _eq_data_307;
  reg [1-1:0] _eq_data_311;
  reg [1-1:0] _eq_data_314;
  reg [1-1:0] _eq_data_317;
  reg [1-1:0] _eq_data_321;
  reg [1-1:0] _eq_data_324;
  reg [1-1:0] _eq_data_327;
  reg [1-1:0] _eq_data_331;
  reg [1-1:0] _eq_data_334;
  reg [1-1:0] _eq_data_337;
  reg [1-1:0] _eq_data_341;
  reg [1-1:0] _eq_data_344;
  reg [1-1:0] _eq_data_347;
  reg [1-1:0] _eq_data_351;
  reg [1-1:0] _eq_data_354;
  reg [1-1:0] _eq_data_357;
  reg [1-1:0] _eq_data_361;
  reg [1-1:0] _eq_data_364;
  reg [1-1:0] _eq_data_367;
  reg [1-1:0] _eq_data_371;
  reg [1-1:0] _eq_data_374;
  reg [1-1:0] _eq_data_377;
  reg [1-1:0] _eq_data_381;
  reg [1-1:0] _eq_data_384;
  reg [1-1:0] _eq_data_387;
  reg [1-1:0] _eq_data_391;
  reg [1-1:0] _eq_data_394;
  reg [1-1:0] _eq_data_397;
  reg [1-1:0] _eq_data_401;
  reg [1-1:0] _eq_data_404;
  reg [1-1:0] _eq_data_407;
  reg [1-1:0] _eq_data_411;
  reg [1-1:0] _eq_data_414;
  reg [1-1:0] _eq_data_417;
  reg [1-1:0] _eq_data_421;
  reg [1-1:0] _eq_data_424;
  reg [1-1:0] _eq_data_427;
  reg [1-1:0] _eq_data_431;
  reg [1-1:0] _eq_data_434;
  reg [1-1:0] _eq_data_437;
  reg [1-1:0] _eq_data_441;
  reg [1-1:0] _eq_data_444;
  reg [1-1:0] _eq_data_447;
  reg [1-1:0] _eq_data_451;
  reg [1-1:0] _eq_data_454;
  wire [4-1:0] _reinterpretcast_src_547;
  assign _reinterpretcast_src_547 = stream_conv2d_16_source_28_data;
  wire signed [4-1:0] _reinterpretcast_data_547;
  assign _reinterpretcast_data_547 = _reinterpretcast_src_547;
  wire [4-1:0] _reinterpretcast_src_548;
  assign _reinterpretcast_src_548 = stream_conv2d_16_source_29_data;
  wire signed [4-1:0] _reinterpretcast_data_548;
  assign _reinterpretcast_data_548 = _reinterpretcast_src_548;
  wire [4-1:0] _reinterpretcast_src_549;
  assign _reinterpretcast_src_549 = stream_conv2d_16_source_30_data;
  wire signed [4-1:0] _reinterpretcast_data_549;
  assign _reinterpretcast_data_549 = _reinterpretcast_src_549;
  wire [4-1:0] _reinterpretcast_src_550;
  assign _reinterpretcast_src_550 = stream_conv2d_16_source_31_data;
  wire signed [4-1:0] _reinterpretcast_data_550;
  assign _reinterpretcast_data_550 = _reinterpretcast_src_550;
  wire [4-1:0] _reinterpretcast_src_551;
  assign _reinterpretcast_src_551 = stream_conv2d_16_source_32_data;
  wire signed [4-1:0] _reinterpretcast_data_551;
  assign _reinterpretcast_data_551 = _reinterpretcast_src_551;
  wire [4-1:0] _reinterpretcast_src_552;
  assign _reinterpretcast_src_552 = stream_conv2d_16_source_33_data;
  wire signed [4-1:0] _reinterpretcast_data_552;
  assign _reinterpretcast_data_552 = _reinterpretcast_src_552;
  wire [4-1:0] _reinterpretcast_src_553;
  assign _reinterpretcast_src_553 = stream_conv2d_16_source_34_data;
  wire signed [4-1:0] _reinterpretcast_data_553;
  assign _reinterpretcast_data_553 = _reinterpretcast_src_553;
  wire [4-1:0] _reinterpretcast_src_554;
  assign _reinterpretcast_src_554 = stream_conv2d_16_source_35_data;
  wire signed [4-1:0] _reinterpretcast_data_554;
  assign _reinterpretcast_data_554 = _reinterpretcast_src_554;
  wire [4-1:0] _reinterpretcast_src_555;
  assign _reinterpretcast_src_555 = stream_conv2d_16_source_36_data;
  wire signed [4-1:0] _reinterpretcast_data_555;
  assign _reinterpretcast_data_555 = _reinterpretcast_src_555;
  wire [1-1:0] _pointer_data_556;
  assign _pointer_data_556 = stream_conv2d_16_constant_3_data[1'sd0];
  wire [1-1:0] _pointer_data_558;
  assign _pointer_data_558 = stream_conv2d_16_constant_3_data[2'sd1];
  wire [1-1:0] _pointer_data_560;
  assign _pointer_data_560 = stream_conv2d_16_constant_3_data[3'sd2];
  wire [1-1:0] _pointer_data_562;
  assign _pointer_data_562 = stream_conv2d_16_constant_3_data[3'sd3];
  wire [1-1:0] _pointer_data_564;
  assign _pointer_data_564 = stream_conv2d_16_constant_3_data[4'sd4];
  wire [1-1:0] _pointer_data_566;
  assign _pointer_data_566 = stream_conv2d_16_constant_3_data[4'sd5];
  wire [1-1:0] _pointer_data_568;
  assign _pointer_data_568 = stream_conv2d_16_constant_3_data[4'sd6];
  wire [1-1:0] _pointer_data_570;
  assign _pointer_data_570 = stream_conv2d_16_constant_3_data[4'sd7];
  wire [1-1:0] _pointer_data_572;
  assign _pointer_data_572 = stream_conv2d_16_constant_3_data[5'sd8];
  reg [8-1:0] __delay_data_898;
  reg [8-1:0] __delay_data_900;
  reg [8-1:0] __delay_data_904;
  reg [8-1:0] __delay_data_907;
  reg [8-1:0] __delay_data_909;
  reg [8-1:0] __delay_data_913;
  reg [8-1:0] __delay_data_916;
  reg [8-1:0] __delay_data_918;
  reg [8-1:0] __delay_data_922;
  reg [1-1:0] __delay_data_940;
  reg [1-1:0] __delay_data_947;
  reg signed [4-1:0] __delay_data_948;
  reg [1-1:0] __delay_data_992;
  reg signed [4-1:0] __delay_data_999;
  reg [1-1:0] __delay_data_1040;
  reg signed [4-1:0] __delay_data_1047;
  reg [1-1:0] __delay_data_1075;
  reg signed [4-1:0] __delay_data_1082;
  reg [1-1:0] __delay_data_1110;
  reg signed [4-1:0] __delay_data_1117;
  reg [1-1:0] __delay_data_1145;
  reg signed [4-1:0] __delay_data_1152;
  reg [1-1:0] __delay_data_1179;
  reg signed [4-1:0] __delay_data_1186;
  reg [1-1:0] __delay_data_1213;
  reg signed [4-1:0] __delay_data_1220;
  reg [1-1:0] __delay_data_1247;
  reg signed [4-1:0] __delay_data_1254;
  reg [1-1:0] __delay_data_1268;
  reg [6-1:0] __delay_data_1289;
  reg [4-1:0] __delay_data_1339;
  reg signed [8-1:0] _cond_data_279;
  reg signed [8-1:0] _cond_data_289;
  reg signed [8-1:0] _cond_data_299;
  reg signed [8-1:0] _cond_data_309;
  reg signed [8-1:0] _cond_data_319;
  reg signed [8-1:0] _cond_data_329;
  reg signed [8-1:0] _cond_data_339;
  reg signed [8-1:0] _cond_data_349;
  reg signed [8-1:0] _cond_data_359;
  reg [8-1:0] _plus_data_607;
  reg [8-1:0] _plus_data_624;
  reg [8-1:0] _plus_data_641;
  reg [8-1:0] _plus_data_658;
  reg [8-1:0] _plus_data_675;
  reg [8-1:0] _plus_data_692;
  reg [8-1:0] _plus_data_709;
  reg [8-1:0] _plus_data_726;
  reg [8-1:0] _plus_data_743;
  reg [8-1:0] _plus_data_759;
  reg [8-1:0] _plus_data_770;
  reg [1-1:0] __delay_data_899;
  reg [8-1:0] __delay_data_901;
  reg [1-1:0] __delay_data_902;
  reg [8-1:0] __delay_data_905;
  reg [1-1:0] __delay_data_908;
  reg [8-1:0] __delay_data_910;
  reg [1-1:0] __delay_data_911;
  reg [8-1:0] __delay_data_914;
  reg [1-1:0] __delay_data_917;
  reg [8-1:0] __delay_data_919;
  reg [1-1:0] __delay_data_920;
  reg [8-1:0] __delay_data_923;
  reg [1-1:0] __delay_data_925;
  reg [1-1:0] __delay_data_928;
  reg [1-1:0] __delay_data_933;
  reg [1-1:0] __delay_data_941;
  reg signed [4-1:0] __delay_data_949;
  reg [1-1:0] __delay_data_962;
  reg [8-1:0] __delay_data_963;
  reg [1-1:0] __delay_data_964;
  reg [1-1:0] __delay_data_967;
  reg [8-1:0] __delay_data_968;
  reg [1-1:0] __delay_data_969;
  reg [1-1:0] __delay_data_972;
  reg [8-1:0] __delay_data_973;
  reg [1-1:0] __delay_data_974;
  reg [1-1:0] __delay_data_977;
  reg [1-1:0] __delay_data_980;
  reg [1-1:0] __delay_data_985;
  reg [1-1:0] __delay_data_993;
  reg signed [4-1:0] __delay_data_1000;
  reg [1-1:0] __delay_data_1013;
  reg [1-1:0] __delay_data_1014;
  reg [1-1:0] __delay_data_1017;
  reg [1-1:0] __delay_data_1018;
  reg [1-1:0] __delay_data_1021;
  reg [1-1:0] __delay_data_1022;
  reg [1-1:0] __delay_data_1025;
  reg [1-1:0] __delay_data_1028;
  reg [1-1:0] __delay_data_1033;
  reg [1-1:0] __delay_data_1041;
  reg signed [4-1:0] __delay_data_1048;
  reg [1-1:0] __delay_data_1061;
  reg [1-1:0] __delay_data_1064;
  reg [1-1:0] __delay_data_1069;
  reg [1-1:0] __delay_data_1076;
  reg signed [4-1:0] __delay_data_1083;
  reg [1-1:0] __delay_data_1096;
  reg [1-1:0] __delay_data_1099;
  reg [1-1:0] __delay_data_1104;
  reg [1-1:0] __delay_data_1111;
  reg signed [4-1:0] __delay_data_1118;
  reg [1-1:0] __delay_data_1131;
  reg [1-1:0] __delay_data_1134;
  reg [1-1:0] __delay_data_1139;
  reg [1-1:0] __delay_data_1146;
  reg signed [4-1:0] __delay_data_1153;
  reg [1-1:0] __delay_data_1166;
  reg [1-1:0] __delay_data_1169;
  reg [1-1:0] __delay_data_1173;
  reg [1-1:0] __delay_data_1180;
  reg signed [4-1:0] __delay_data_1187;
  reg [1-1:0] __delay_data_1200;
  reg [1-1:0] __delay_data_1203;
  reg [1-1:0] __delay_data_1207;
  reg [1-1:0] __delay_data_1214;
  reg signed [4-1:0] __delay_data_1221;
  reg [1-1:0] __delay_data_1234;
  reg [1-1:0] __delay_data_1237;
  reg [1-1:0] __delay_data_1241;
  reg [1-1:0] __delay_data_1248;
  reg signed [4-1:0] __delay_data_1255;
  reg [6-1:0] __delay_data_1290;
  reg signed [8-1:0] __delay_data_1311;
  reg signed [8-1:0] __delay_data_1340;
  reg signed [8-1:0] _cond_data_283;
  reg signed [8-1:0] _cond_data_293;
  reg signed [8-1:0] _cond_data_303;
  reg signed [8-1:0] _cond_data_313;
  reg signed [8-1:0] _cond_data_323;
  reg signed [8-1:0] _cond_data_333;
  reg signed [8-1:0] _cond_data_343;
  reg signed [8-1:0] _cond_data_353;
  reg signed [8-1:0] _cond_data_363;
  reg [1-1:0] __delay_data_903;
  reg [8-1:0] __delay_data_906;
  reg [1-1:0] __delay_data_912;
  reg [8-1:0] __delay_data_915;
  reg [1-1:0] __delay_data_921;
  reg [8-1:0] __delay_data_924;
  reg [1-1:0] __delay_data_926;
  reg [1-1:0] __delay_data_929;
  reg [1-1:0] __delay_data_934;
  reg [1-1:0] __delay_data_942;
  reg signed [4-1:0] __delay_data_950;
  reg [8-1:0] __delay_data_956;
  reg [1-1:0] __delay_data_965;
  reg [8-1:0] __delay_data_966;
  reg [1-1:0] __delay_data_970;
  reg [8-1:0] __delay_data_971;
  reg [1-1:0] __delay_data_975;
  reg [8-1:0] __delay_data_976;
  reg [1-1:0] __delay_data_978;
  reg [1-1:0] __delay_data_981;
  reg [1-1:0] __delay_data_986;
  reg [1-1:0] __delay_data_994;
  reg signed [4-1:0] __delay_data_1001;
  reg [8-1:0] __delay_data_1007;
  reg [1-1:0] __delay_data_1015;
  reg [8-1:0] __delay_data_1016;
  reg [1-1:0] __delay_data_1019;
  reg [8-1:0] __delay_data_1020;
  reg [1-1:0] __delay_data_1023;
  reg [8-1:0] __delay_data_1024;
  reg [1-1:0] __delay_data_1026;
  reg [1-1:0] __delay_data_1029;
  reg [1-1:0] __delay_data_1034;
  reg [1-1:0] __delay_data_1042;
  reg signed [4-1:0] __delay_data_1049;
  reg [8-1:0] __delay_data_1055;
  reg [1-1:0] __delay_data_1062;
  reg [1-1:0] __delay_data_1065;
  reg [1-1:0] __delay_data_1070;
  reg [1-1:0] __delay_data_1077;
  reg signed [4-1:0] __delay_data_1084;
  reg [8-1:0] __delay_data_1090;
  reg [1-1:0] __delay_data_1097;
  reg [1-1:0] __delay_data_1100;
  reg [1-1:0] __delay_data_1105;
  reg [1-1:0] __delay_data_1112;
  reg signed [4-1:0] __delay_data_1119;
  reg [8-1:0] __delay_data_1125;
  reg [1-1:0] __delay_data_1132;
  reg [1-1:0] __delay_data_1135;
  reg [1-1:0] __delay_data_1140;
  reg [1-1:0] __delay_data_1147;
  reg signed [4-1:0] __delay_data_1154;
  reg [8-1:0] __delay_data_1160;
  reg [1-1:0] __delay_data_1167;
  reg [1-1:0] __delay_data_1170;
  reg [1-1:0] __delay_data_1174;
  reg [1-1:0] __delay_data_1181;
  reg signed [4-1:0] __delay_data_1188;
  reg [8-1:0] __delay_data_1194;
  reg [1-1:0] __delay_data_1201;
  reg [1-1:0] __delay_data_1204;
  reg [1-1:0] __delay_data_1208;
  reg [1-1:0] __delay_data_1215;
  reg signed [4-1:0] __delay_data_1222;
  reg [8-1:0] __delay_data_1228;
  reg [1-1:0] __delay_data_1235;
  reg [1-1:0] __delay_data_1238;
  reg [1-1:0] __delay_data_1242;
  reg [1-1:0] __delay_data_1249;
  reg signed [4-1:0] __delay_data_1256;
  reg [8-1:0] __delay_data_1262;
  reg [8-1:0] __delay_data_1269;
  reg [6-1:0] __delay_data_1291;
  reg signed [8-1:0] __delay_data_1312;
  reg signed [8-1:0] __delay_data_1341;
  reg [8-1:0] __delay_data_1369;
  reg signed [8-1:0] _cond_data_286;
  reg signed [8-1:0] _cond_data_296;
  reg signed [8-1:0] _cond_data_306;
  reg signed [8-1:0] _cond_data_316;
  reg signed [8-1:0] _cond_data_326;
  reg signed [8-1:0] _cond_data_336;
  reg signed [8-1:0] _cond_data_346;
  reg signed [8-1:0] _cond_data_356;
  reg signed [8-1:0] _cond_data_366;
  reg [1-1:0] __delay_data_927;
  reg [1-1:0] __delay_data_930;
  reg [1-1:0] __delay_data_935;
  reg [1-1:0] __delay_data_943;
  reg signed [4-1:0] __delay_data_951;
  reg [8-1:0] __delay_data_957;
  reg [1-1:0] __delay_data_979;
  reg [1-1:0] __delay_data_982;
  reg [1-1:0] __delay_data_987;
  reg [1-1:0] __delay_data_995;
  reg signed [4-1:0] __delay_data_1002;
  reg [8-1:0] __delay_data_1008;
  reg [1-1:0] __delay_data_1027;
  reg [1-1:0] __delay_data_1030;
  reg [1-1:0] __delay_data_1035;
  reg [1-1:0] __delay_data_1043;
  reg signed [4-1:0] __delay_data_1050;
  reg [8-1:0] __delay_data_1056;
  reg [1-1:0] __delay_data_1063;
  reg [1-1:0] __delay_data_1066;
  reg [1-1:0] __delay_data_1071;
  reg [1-1:0] __delay_data_1078;
  reg signed [4-1:0] __delay_data_1085;
  reg [8-1:0] __delay_data_1091;
  reg [1-1:0] __delay_data_1098;
  reg [1-1:0] __delay_data_1101;
  reg [1-1:0] __delay_data_1106;
  reg [1-1:0] __delay_data_1113;
  reg signed [4-1:0] __delay_data_1120;
  reg [8-1:0] __delay_data_1126;
  reg [1-1:0] __delay_data_1133;
  reg [1-1:0] __delay_data_1136;
  reg [1-1:0] __delay_data_1141;
  reg [1-1:0] __delay_data_1148;
  reg signed [4-1:0] __delay_data_1155;
  reg [8-1:0] __delay_data_1161;
  reg [1-1:0] __delay_data_1168;
  reg [1-1:0] __delay_data_1171;
  reg [1-1:0] __delay_data_1175;
  reg [1-1:0] __delay_data_1182;
  reg signed [4-1:0] __delay_data_1189;
  reg [8-1:0] __delay_data_1195;
  reg [1-1:0] __delay_data_1202;
  reg [1-1:0] __delay_data_1205;
  reg [1-1:0] __delay_data_1209;
  reg [1-1:0] __delay_data_1216;
  reg signed [4-1:0] __delay_data_1223;
  reg [8-1:0] __delay_data_1229;
  reg [1-1:0] __delay_data_1236;
  reg [1-1:0] __delay_data_1239;
  reg [1-1:0] __delay_data_1243;
  reg [1-1:0] __delay_data_1250;
  reg signed [4-1:0] __delay_data_1257;
  reg [8-1:0] __delay_data_1263;
  reg [8-1:0] __delay_data_1270;
  reg [6-1:0] __delay_data_1292;
  reg signed [8-1:0] __delay_data_1313;
  reg signed [8-1:0] __delay_data_1342;
  reg [8-1:0] __delay_data_1370;
  reg signed [8-1:0] _cond_data_369;
  reg signed [8-1:0] _cond_data_379;
  reg signed [8-1:0] _cond_data_389;
  reg signed [8-1:0] _cond_data_399;
  reg signed [8-1:0] _cond_data_409;
  reg signed [8-1:0] _cond_data_419;
  reg signed [8-1:0] _cond_data_429;
  reg signed [8-1:0] _cond_data_439;
  reg signed [8-1:0] _cond_data_449;
  reg [1-1:0] __delay_data_931;
  reg signed [8-1:0] __delay_data_932;
  reg [1-1:0] __delay_data_936;
  reg signed [8-1:0] __delay_data_938;
  reg [1-1:0] __delay_data_944;
  reg signed [4-1:0] __delay_data_952;
  reg [8-1:0] __delay_data_958;
  reg [1-1:0] __delay_data_983;
  reg signed [8-1:0] __delay_data_984;
  reg [1-1:0] __delay_data_988;
  reg signed [8-1:0] __delay_data_990;
  reg [1-1:0] __delay_data_996;
  reg signed [4-1:0] __delay_data_1003;
  reg [8-1:0] __delay_data_1009;
  reg [1-1:0] __delay_data_1031;
  reg signed [8-1:0] __delay_data_1032;
  reg [1-1:0] __delay_data_1036;
  reg signed [8-1:0] __delay_data_1038;
  reg [1-1:0] __delay_data_1044;
  reg signed [4-1:0] __delay_data_1051;
  reg [8-1:0] __delay_data_1057;
  reg [1-1:0] __delay_data_1067;
  reg signed [8-1:0] __delay_data_1068;
  reg [1-1:0] __delay_data_1072;
  reg [1-1:0] __delay_data_1079;
  reg signed [4-1:0] __delay_data_1086;
  reg [8-1:0] __delay_data_1092;
  reg [1-1:0] __delay_data_1102;
  reg signed [8-1:0] __delay_data_1103;
  reg [1-1:0] __delay_data_1107;
  reg [1-1:0] __delay_data_1114;
  reg signed [4-1:0] __delay_data_1121;
  reg [8-1:0] __delay_data_1127;
  reg [1-1:0] __delay_data_1137;
  reg signed [8-1:0] __delay_data_1138;
  reg [1-1:0] __delay_data_1142;
  reg [1-1:0] __delay_data_1149;
  reg signed [4-1:0] __delay_data_1156;
  reg [8-1:0] __delay_data_1162;
  reg [1-1:0] __delay_data_1172;
  reg [1-1:0] __delay_data_1176;
  reg [1-1:0] __delay_data_1183;
  reg signed [4-1:0] __delay_data_1190;
  reg [8-1:0] __delay_data_1196;
  reg [1-1:0] __delay_data_1206;
  reg [1-1:0] __delay_data_1210;
  reg [1-1:0] __delay_data_1217;
  reg signed [4-1:0] __delay_data_1224;
  reg [8-1:0] __delay_data_1230;
  reg [1-1:0] __delay_data_1240;
  reg [1-1:0] __delay_data_1244;
  reg [1-1:0] __delay_data_1251;
  reg signed [4-1:0] __delay_data_1258;
  reg [8-1:0] __delay_data_1264;
  reg [8-1:0] __delay_data_1271;
  reg [6-1:0] __delay_data_1293;
  reg signed [8-1:0] __delay_data_1314;
  reg signed [8-1:0] __delay_data_1343;
  reg [8-1:0] __delay_data_1371;
  reg signed [8-1:0] _cond_data_373;
  reg signed [8-1:0] _cond_data_383;
  reg signed [8-1:0] _cond_data_393;
  reg signed [8-1:0] _cond_data_403;
  reg signed [8-1:0] _cond_data_413;
  reg signed [8-1:0] _cond_data_423;
  reg signed [8-1:0] _cond_data_433;
  reg signed [8-1:0] _cond_data_443;
  reg signed [8-1:0] _cond_data_453;
  reg [1-1:0] __delay_data_937;
  reg signed [8-1:0] __delay_data_939;
  reg [1-1:0] __delay_data_945;
  reg signed [4-1:0] __delay_data_953;
  reg [8-1:0] __delay_data_959;
  reg [1-1:0] __delay_data_989;
  reg signed [8-1:0] __delay_data_991;
  reg [1-1:0] __delay_data_997;
  reg signed [4-1:0] __delay_data_1004;
  reg [8-1:0] __delay_data_1010;
  reg [1-1:0] __delay_data_1037;
  reg signed [8-1:0] __delay_data_1039;
  reg [1-1:0] __delay_data_1045;
  reg signed [4-1:0] __delay_data_1052;
  reg [8-1:0] __delay_data_1058;
  reg [1-1:0] __delay_data_1073;
  reg signed [8-1:0] __delay_data_1074;
  reg [1-1:0] __delay_data_1080;
  reg signed [4-1:0] __delay_data_1087;
  reg [8-1:0] __delay_data_1093;
  reg [1-1:0] __delay_data_1108;
  reg signed [8-1:0] __delay_data_1109;
  reg [1-1:0] __delay_data_1115;
  reg signed [4-1:0] __delay_data_1122;
  reg [8-1:0] __delay_data_1128;
  reg [1-1:0] __delay_data_1143;
  reg signed [8-1:0] __delay_data_1144;
  reg [1-1:0] __delay_data_1150;
  reg signed [4-1:0] __delay_data_1157;
  reg [8-1:0] __delay_data_1163;
  reg [1-1:0] __delay_data_1177;
  reg signed [8-1:0] __delay_data_1178;
  reg [1-1:0] __delay_data_1184;
  reg signed [4-1:0] __delay_data_1191;
  reg [8-1:0] __delay_data_1197;
  reg [1-1:0] __delay_data_1211;
  reg signed [8-1:0] __delay_data_1212;
  reg [1-1:0] __delay_data_1218;
  reg signed [4-1:0] __delay_data_1225;
  reg [8-1:0] __delay_data_1231;
  reg [1-1:0] __delay_data_1245;
  reg signed [8-1:0] __delay_data_1246;
  reg [1-1:0] __delay_data_1252;
  reg signed [4-1:0] __delay_data_1259;
  reg [8-1:0] __delay_data_1265;
  reg [8-1:0] __delay_data_1272;
  reg [6-1:0] __delay_data_1294;
  reg signed [8-1:0] __delay_data_1315;
  reg signed [8-1:0] __delay_data_1344;
  reg [8-1:0] __delay_data_1372;
  reg signed [8-1:0] _cond_data_376;
  reg signed [8-1:0] _cond_data_386;
  reg signed [8-1:0] _cond_data_396;
  reg signed [8-1:0] _cond_data_406;
  reg signed [8-1:0] _cond_data_416;
  reg signed [8-1:0] _cond_data_426;
  reg signed [8-1:0] _cond_data_436;
  reg signed [8-1:0] _cond_data_446;
  reg signed [8-1:0] _cond_data_456;
  reg [1-1:0] __delay_data_946;
  reg signed [4-1:0] __delay_data_954;
  reg [8-1:0] __delay_data_960;
  reg [1-1:0] __delay_data_998;
  reg signed [4-1:0] __delay_data_1005;
  reg [8-1:0] __delay_data_1011;
  reg [1-1:0] __delay_data_1046;
  reg signed [4-1:0] __delay_data_1053;
  reg [8-1:0] __delay_data_1059;
  reg [1-1:0] __delay_data_1081;
  reg signed [4-1:0] __delay_data_1088;
  reg [8-1:0] __delay_data_1094;
  reg [1-1:0] __delay_data_1116;
  reg signed [4-1:0] __delay_data_1123;
  reg [8-1:0] __delay_data_1129;
  reg [1-1:0] __delay_data_1151;
  reg signed [4-1:0] __delay_data_1158;
  reg [8-1:0] __delay_data_1164;
  reg [1-1:0] __delay_data_1185;
  reg signed [4-1:0] __delay_data_1192;
  reg [8-1:0] __delay_data_1198;
  reg [1-1:0] __delay_data_1219;
  reg signed [4-1:0] __delay_data_1226;
  reg [8-1:0] __delay_data_1232;
  reg [1-1:0] __delay_data_1253;
  reg signed [4-1:0] __delay_data_1260;
  reg [8-1:0] __delay_data_1266;
  reg [8-1:0] __delay_data_1273;
  reg [6-1:0] __delay_data_1295;
  reg signed [8-1:0] __delay_data_1316;
  reg signed [8-1:0] __delay_data_1345;
  reg [8-1:0] __delay_data_1373;
  wire signed [8-1:0] _reinterpretcast_src_493;
  assign _reinterpretcast_src_493 = _cond_data_376;
  wire signed [8-1:0] _reinterpretcast_data_493;
  assign _reinterpretcast_data_493 = _reinterpretcast_src_493;
  wire signed [8-1:0] _reinterpretcast_src_494;
  assign _reinterpretcast_src_494 = _cond_data_406;
  wire signed [8-1:0] _reinterpretcast_data_494;
  assign _reinterpretcast_data_494 = _reinterpretcast_src_494;
  wire signed [8-1:0] _reinterpretcast_src_495;
  assign _reinterpretcast_src_495 = _cond_data_436;
  wire signed [8-1:0] _reinterpretcast_data_495;
  assign _reinterpretcast_data_495 = _reinterpretcast_src_495;
  wire signed [8-1:0] _reinterpretcast_src_496;
  assign _reinterpretcast_src_496 = _cond_data_386;
  wire signed [8-1:0] _reinterpretcast_data_496;
  assign _reinterpretcast_data_496 = _reinterpretcast_src_496;
  wire signed [8-1:0] _reinterpretcast_src_497;
  assign _reinterpretcast_src_497 = _cond_data_416;
  wire signed [8-1:0] _reinterpretcast_data_497;
  assign _reinterpretcast_data_497 = _reinterpretcast_src_497;
  wire signed [8-1:0] _reinterpretcast_src_498;
  assign _reinterpretcast_src_498 = _cond_data_446;
  wire signed [8-1:0] _reinterpretcast_data_498;
  assign _reinterpretcast_data_498 = _reinterpretcast_src_498;
  wire signed [8-1:0] _reinterpretcast_src_499;
  assign _reinterpretcast_src_499 = _cond_data_396;
  wire signed [8-1:0] _reinterpretcast_data_499;
  assign _reinterpretcast_data_499 = _reinterpretcast_src_499;
  wire signed [8-1:0] _reinterpretcast_src_500;
  assign _reinterpretcast_src_500 = _cond_data_426;
  wire signed [8-1:0] _reinterpretcast_data_500;
  assign _reinterpretcast_data_500 = _reinterpretcast_src_500;
  wire signed [8-1:0] _reinterpretcast_src_501;
  assign _reinterpretcast_src_501 = _cond_data_456;
  wire signed [8-1:0] _reinterpretcast_data_501;
  assign _reinterpretcast_data_501 = _reinterpretcast_src_501;
  reg signed [8-1:0] _cond_data_575;
  reg signed [8-1:0] _cond_data_577;
  reg signed [8-1:0] _cond_data_579;
  reg signed [8-1:0] _cond_data_581;
  reg signed [8-1:0] _cond_data_583;
  reg signed [8-1:0] _cond_data_585;
  reg signed [8-1:0] _cond_data_587;
  reg signed [8-1:0] _cond_data_589;
  reg signed [8-1:0] _cond_data_591;
  reg signed [4-1:0] __delay_data_955;
  reg [8-1:0] __delay_data_961;
  reg signed [4-1:0] __delay_data_1006;
  reg [8-1:0] __delay_data_1012;
  reg signed [4-1:0] __delay_data_1054;
  reg [8-1:0] __delay_data_1060;
  reg signed [4-1:0] __delay_data_1089;
  reg [8-1:0] __delay_data_1095;
  reg signed [4-1:0] __delay_data_1124;
  reg [8-1:0] __delay_data_1130;
  reg signed [4-1:0] __delay_data_1159;
  reg [8-1:0] __delay_data_1165;
  reg signed [4-1:0] __delay_data_1193;
  reg [8-1:0] __delay_data_1199;
  reg signed [4-1:0] __delay_data_1227;
  reg [8-1:0] __delay_data_1233;
  reg signed [4-1:0] __delay_data_1261;
  reg [8-1:0] __delay_data_1267;
  reg [8-1:0] __delay_data_1274;
  reg [6-1:0] __delay_data_1296;
  reg signed [8-1:0] __delay_data_1317;
  reg signed [8-1:0] __delay_data_1346;
  reg [8-1:0] __delay_data_1374;
  reg signed [8-1:0] __variable_wdata_54;
  assign mul_4_x_data = __variable_wdata_54;
  reg signed [4-1:0] __variable_wdata_55;
  assign mul_4_y_data = __variable_wdata_55;
  reg [4-1:0] __variable_wdata_56;
  assign mul_4_rshift_data = __variable_wdata_56;
  reg signed [8-1:0] __variable_wdata_71;
  assign mul_5_x_data = __variable_wdata_71;
  reg signed [4-1:0] __variable_wdata_72;
  assign mul_5_y_data = __variable_wdata_72;
  reg [4-1:0] __variable_wdata_73;
  assign mul_5_rshift_data = __variable_wdata_73;
  reg signed [8-1:0] __variable_wdata_88;
  assign mul_6_x_data = __variable_wdata_88;
  reg signed [4-1:0] __variable_wdata_89;
  assign mul_6_y_data = __variable_wdata_89;
  reg [4-1:0] __variable_wdata_90;
  assign mul_6_rshift_data = __variable_wdata_90;
  reg signed [8-1:0] __variable_wdata_105;
  assign mul_7_x_data = __variable_wdata_105;
  reg signed [4-1:0] __variable_wdata_106;
  assign mul_7_y_data = __variable_wdata_106;
  reg [4-1:0] __variable_wdata_107;
  assign mul_7_rshift_data = __variable_wdata_107;
  reg signed [8-1:0] __variable_wdata_122;
  assign mul_8_x_data = __variable_wdata_122;
  reg signed [4-1:0] __variable_wdata_123;
  assign mul_8_y_data = __variable_wdata_123;
  reg [4-1:0] __variable_wdata_124;
  assign mul_8_rshift_data = __variable_wdata_124;
  reg signed [8-1:0] __variable_wdata_139;
  assign mul_9_x_data = __variable_wdata_139;
  reg signed [4-1:0] __variable_wdata_140;
  assign mul_9_y_data = __variable_wdata_140;
  reg [4-1:0] __variable_wdata_141;
  assign mul_9_rshift_data = __variable_wdata_141;
  reg signed [8-1:0] __variable_wdata_156;
  assign mul_10_x_data = __variable_wdata_156;
  reg signed [4-1:0] __variable_wdata_157;
  assign mul_10_y_data = __variable_wdata_157;
  reg [4-1:0] __variable_wdata_158;
  assign mul_10_rshift_data = __variable_wdata_158;
  reg signed [8-1:0] __variable_wdata_173;
  assign mul_11_x_data = __variable_wdata_173;
  reg signed [4-1:0] __variable_wdata_174;
  assign mul_11_y_data = __variable_wdata_174;
  reg [4-1:0] __variable_wdata_175;
  assign mul_11_rshift_data = __variable_wdata_175;
  reg signed [8-1:0] __variable_wdata_190;
  assign mul_12_x_data = __variable_wdata_190;
  reg signed [4-1:0] __variable_wdata_191;
  assign mul_12_y_data = __variable_wdata_191;
  reg [4-1:0] __variable_wdata_192;
  assign mul_12_rshift_data = __variable_wdata_192;
  reg [8-1:0] __delay_data_1275;
  reg [6-1:0] __delay_data_1297;
  reg signed [8-1:0] __delay_data_1318;
  reg signed [8-1:0] __delay_data_1347;
  reg [8-1:0] __delay_data_1375;
  reg [8-1:0] __delay_data_1276;
  reg [6-1:0] __delay_data_1298;
  reg signed [8-1:0] __delay_data_1319;
  reg signed [8-1:0] __delay_data_1348;
  reg [8-1:0] __delay_data_1376;
  reg [8-1:0] __delay_data_1277;
  reg [6-1:0] __delay_data_1299;
  reg signed [8-1:0] __delay_data_1320;
  reg signed [8-1:0] __delay_data_1349;
  reg [8-1:0] __delay_data_1377;
  reg [8-1:0] __delay_data_1278;
  reg [6-1:0] __delay_data_1300;
  reg signed [8-1:0] __delay_data_1321;
  reg signed [8-1:0] __delay_data_1350;
  reg [8-1:0] __delay_data_1378;
  reg [8-1:0] __delay_data_1279;
  reg [6-1:0] __delay_data_1301;
  reg signed [8-1:0] __delay_data_1322;
  reg signed [8-1:0] __delay_data_1351;
  reg [8-1:0] __delay_data_1379;
  reg [8-1:0] __delay_data_1280;
  reg [6-1:0] __delay_data_1302;
  reg signed [8-1:0] __delay_data_1323;
  reg signed [8-1:0] __delay_data_1352;
  reg [8-1:0] __delay_data_1380;
  reg [8-1:0] __delay_data_1281;
  reg [6-1:0] __delay_data_1303;
  reg signed [8-1:0] __delay_data_1324;
  reg signed [8-1:0] __delay_data_1353;
  reg [8-1:0] __delay_data_1381;
  reg [8-1:0] __delay_data_1282;
  reg [6-1:0] __delay_data_1304;
  reg signed [8-1:0] __delay_data_1325;
  reg signed [8-1:0] __delay_data_1354;
  reg [8-1:0] __delay_data_1382;
  reg [8-1:0] __delay_data_1283;
  reg [6-1:0] __delay_data_1305;
  reg signed [8-1:0] __delay_data_1326;
  reg signed [8-1:0] __delay_data_1355;
  reg [8-1:0] __delay_data_1383;
  reg signed [12-1:0] __substreamoutput_data_608;
  reg signed [12-1:0] __substreamoutput_data_625;
  reg signed [12-1:0] __substreamoutput_data_642;
  reg signed [12-1:0] __substreamoutput_data_659;
  reg signed [12-1:0] __substreamoutput_data_676;
  reg signed [12-1:0] __substreamoutput_data_693;
  reg signed [12-1:0] __substreamoutput_data_710;
  reg signed [12-1:0] __substreamoutput_data_727;
  reg signed [12-1:0] __substreamoutput_data_744;
  reg [8-1:0] __delay_data_1284;
  reg [6-1:0] __delay_data_1306;
  reg signed [8-1:0] __delay_data_1327;
  reg signed [8-1:0] __delay_data_1356;
  reg [8-1:0] __delay_data_1384;
  reg signed [32-1:0] __variable_wdata_24;
  assign add_tree_2_var0_data = __variable_wdata_24;
  reg signed [32-1:0] __variable_wdata_25;
  assign add_tree_2_var1_data = __variable_wdata_25;
  reg signed [32-1:0] __variable_wdata_26;
  assign add_tree_2_var2_data = __variable_wdata_26;
  reg signed [32-1:0] __variable_wdata_27;
  assign add_tree_2_var3_data = __variable_wdata_27;
  reg signed [32-1:0] __variable_wdata_28;
  assign add_tree_2_var4_data = __variable_wdata_28;
  reg signed [32-1:0] __variable_wdata_29;
  assign add_tree_2_var5_data = __variable_wdata_29;
  reg signed [32-1:0] __variable_wdata_30;
  assign add_tree_2_var6_data = __variable_wdata_30;
  reg signed [32-1:0] __variable_wdata_31;
  assign add_tree_2_var7_data = __variable_wdata_31;
  reg signed [32-1:0] __variable_wdata_32;
  assign add_tree_2_var8_data = __variable_wdata_32;
  reg [8-1:0] __delay_data_1285;
  reg [6-1:0] __delay_data_1307;
  reg signed [8-1:0] __delay_data_1328;
  reg signed [8-1:0] __delay_data_1357;
  reg [8-1:0] __delay_data_1385;
  reg [8-1:0] __delay_data_1286;
  reg [6-1:0] __delay_data_1308;
  reg signed [8-1:0] __delay_data_1329;
  reg signed [8-1:0] __delay_data_1358;
  reg [8-1:0] __delay_data_1386;
  reg [8-1:0] __delay_data_1287;
  reg [6-1:0] __delay_data_1309;
  reg signed [8-1:0] __delay_data_1330;
  reg signed [8-1:0] __delay_data_1359;
  reg [8-1:0] __delay_data_1387;
  reg signed [32-1:0] __substreamoutput_data_746;
  reg [8-1:0] __delay_data_1288;
  reg [6-1:0] __delay_data_1310;
  reg signed [8-1:0] __delay_data_1331;
  reg signed [8-1:0] __delay_data_1360;
  reg [8-1:0] __delay_data_1388;
  reg signed [32-1:0] __variable_wdata_0;
  assign acc_0_x_data = __variable_wdata_0;
  reg [6-1:0] __variable_wdata_1;
  assign acc_0_rshift_data = __variable_wdata_1;
  reg [32-1:0] __variable_wdata_2;
  assign acc_0_size_data = __variable_wdata_2;
  reg signed [8-1:0] __delay_data_1332;
  reg signed [8-1:0] __delay_data_1361;
  reg [8-1:0] __delay_data_1389;
  reg signed [8-1:0] __delay_data_1333;
  reg signed [8-1:0] __delay_data_1362;
  reg [8-1:0] __delay_data_1390;
  reg signed [8-1:0] __delay_data_1334;
  reg signed [8-1:0] __delay_data_1363;
  reg [8-1:0] __delay_data_1391;
  reg signed [8-1:0] __delay_data_1335;
  reg signed [8-1:0] __delay_data_1364;
  reg [8-1:0] __delay_data_1392;
  reg signed [8-1:0] __delay_data_1336;
  reg signed [8-1:0] __delay_data_1365;
  reg [8-1:0] __delay_data_1393;
  reg signed [8-1:0] __delay_data_1337;
  reg signed [8-1:0] __delay_data_1366;
  reg [8-1:0] __delay_data_1394;
  reg signed [32-1:0] __substreamoutput_data_760;
  reg [1-1:0] __substreamoutput_data_761;
  reg signed [8-1:0] __delay_data_1338;
  reg signed [8-1:0] __delay_data_1367;
  reg [8-1:0] __delay_data_1395;
  reg signed [32-1:0] _plus_data_762;
  reg signed [8-1:0] __delay_data_1368;
  reg [8-1:0] __delay_data_1396;
  reg [1-1:0] __delay_data_1398;
  reg signed [32-1:0] __variable_wdata_38;
  assign mul_rshift_clip_3_x_data = __variable_wdata_38;
  reg signed [8-1:0] __variable_wdata_39;
  assign mul_rshift_clip_3_y_data = __variable_wdata_39;
  reg [6-1:0] __variable_wdata_40;
  assign mul_rshift_clip_3_rshift_data = __variable_wdata_40;
  reg [1-1:0] __delay_data_1399;
  reg [1-1:0] __delay_data_1400;
  reg [1-1:0] __delay_data_1401;
  reg [1-1:0] __delay_data_1402;
  reg [1-1:0] __delay_data_1403;
  reg [1-1:0] __delay_data_1404;
  reg [1-1:0] __delay_data_1405;
  reg [1-1:0] __delay_data_1406;
  reg [1-1:0] __delay_data_1407;
  reg signed [8-1:0] __substreamoutput_data_771;
  reg [1-1:0] __delay_data_1408;
  reg [1-1:0] _greaterthan_data_773;
  reg signed [8-1:0] __delay_data_1397;
  reg [1-1:0] __delay_data_1409;
  reg signed [8-1:0] _cond_data_775;
  reg [1-1:0] __delay_data_1410;
  wire signed [8-1:0] _reinterpretcast_src_776;
  assign _reinterpretcast_src_776 = _cond_data_775;
  wire signed [8-1:0] _reinterpretcast_data_776;
  assign _reinterpretcast_data_776 = _reinterpretcast_src_776;
  wire signed [8-1:0] stream_conv2d_16_sink_37_data;
  assign stream_conv2d_16_sink_37_data = _reinterpretcast_data_776;
  wire [1-1:0] stream_conv2d_16_sink_38_data;
  assign stream_conv2d_16_sink_38_data = __delay_data_1410;
  reg _set_flag_457;
  reg [6-1:0] __variable_wdata_214;
  assign stream_conv2d_16_constant_0_data = __variable_wdata_214;
  reg _set_flag_458;
  reg [2-1:0] __variable_wdata_215;
  assign stream_conv2d_16_constant_1_data = __variable_wdata_215;
  reg _set_flag_459;
  reg [2-1:0] __variable_wdata_216;
  assign stream_conv2d_16_constant_2_data = __variable_wdata_216;
  reg _set_flag_460;
  reg [9-1:0] __variable_wdata_217;
  assign stream_conv2d_16_constant_3_data = __variable_wdata_217;
  reg _set_flag_461;
  reg [1-1:0] __variable_wdata_218;
  assign stream_conv2d_16_constant_4_data = __variable_wdata_218;
  reg _set_flag_462;
  reg [1-1:0] __variable_wdata_229;
  assign stream_conv2d_16_constant_5_data = __variable_wdata_229;
  reg [32-1:0] _source_stream_conv2d_16_source_6_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_6_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_6_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_6_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_6_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_6_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_6_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_6_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_6_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_6_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_6_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_6_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_6_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_6_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_6_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_6_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_6_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_6_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_6_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_6_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_6_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_6_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_6_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_6_pat_stride_buf_3;
  reg _set_flag_463;
  wire [2-1:0] _tmp_464;
  assign _tmp_464 = _stream_conv2d_16_source_6_source_ram_raddr;
  reg [2-1:0] __tmp_464_1;
  reg [2-1:0] __tmp_464_2;
  reg _tmp_465;
  reg _ram_w8_l2048_id1_0_cond_1_1;
  reg _ram_w8_l2048_id1_0_cond_2_1;
  reg _ram_w8_l2048_id1_0_cond_2_2;
  reg _tmp_466;
  reg _ram_w8_l2048_id1_1_cond_1_1;
  reg _ram_w8_l2048_id1_1_cond_2_1;
  reg _ram_w8_l2048_id1_1_cond_2_2;
  reg _tmp_467;
  reg _ram_w8_l2048_id1_2_cond_1_1;
  reg _ram_w8_l2048_id1_2_cond_2_1;
  reg _ram_w8_l2048_id1_2_cond_2_2;
  reg _tmp_468;
  reg _ram_w8_l2048_id1_3_cond_1_1;
  reg _ram_w8_l2048_id1_3_cond_2_1;
  reg _ram_w8_l2048_id1_3_cond_2_2;
  wire signed [8-1:0] _tmp_469;
  wire _tmp_470;
  assign _tmp_469 = (__tmp_464_2 == 0)? ram_w8_l2048_id1_0_0_rdata : 
                    (__tmp_464_2 == 1)? ram_w8_l2048_id1_1_0_rdata : 
                    (__tmp_464_2 == 2)? ram_w8_l2048_id1_2_0_rdata : 
                    (__tmp_464_2 == 3)? ram_w8_l2048_id1_3_0_rdata : 0;
  assign _tmp_470 = _tmp_465;
  assign _stream_conv2d_16_source_6_source_ram_rdata = (_stream_conv2d_16_source_6_source_ram_sel == 1)? _tmp_469 : 0;
  localparam _tmp_471 = 1;
  wire [_tmp_471-1:0] _tmp_472;
  assign _tmp_472 = _stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1);
  reg [_tmp_471-1:0] __tmp_472_1;
  reg [8-1:0] __variable_wdata_230;
  assign stream_conv2d_16_source_6_data = __variable_wdata_230;
  reg [32-1:0] _stream_conv2d_16_source_6_source_pat_fsm_0;
  localparam _stream_conv2d_16_source_6_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_6_source_pat_all_offset;
  assign _stream_conv2d_16_source_6_source_pat_all_offset = _stream_conv2d_16_source_6_source_offset_buf + _source_stream_conv2d_16_source_6_pat_cur_offset_0 + _source_stream_conv2d_16_source_6_pat_cur_offset_1 + _source_stream_conv2d_16_source_6_pat_cur_offset_2 + _source_stream_conv2d_16_source_6_pat_cur_offset_3;
  reg _set_flag_473;
  reg [1-1:0] __variable_wdata_236;
  assign stream_conv2d_16_constant_7_data = __variable_wdata_236;
  reg [32-1:0] _source_stream_conv2d_16_source_8_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_8_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_8_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_8_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_8_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_8_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_8_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_8_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_8_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_8_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_8_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_8_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_8_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_8_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_8_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_8_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_8_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_8_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_8_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_8_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_8_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_8_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_8_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_8_pat_stride_buf_3;
  reg _set_flag_474;
  wire [2-1:0] _tmp_475;
  assign _tmp_475 = _stream_conv2d_16_source_8_source_ram_raddr;
  reg [2-1:0] __tmp_475_1;
  reg [2-1:0] __tmp_475_2;
  reg _tmp_476;
  reg _ram_w8_l2048_id0_0_cond_1_1;
  reg _ram_w8_l2048_id0_0_cond_2_1;
  reg _ram_w8_l2048_id0_0_cond_2_2;
  reg _tmp_477;
  reg _ram_w8_l2048_id0_1_cond_1_1;
  reg _ram_w8_l2048_id0_1_cond_2_1;
  reg _ram_w8_l2048_id0_1_cond_2_2;
  reg _tmp_478;
  reg _ram_w8_l2048_id0_2_cond_1_1;
  reg _ram_w8_l2048_id0_2_cond_2_1;
  reg _ram_w8_l2048_id0_2_cond_2_2;
  reg _tmp_479;
  reg _ram_w8_l2048_id0_3_cond_1_1;
  reg _ram_w8_l2048_id0_3_cond_2_1;
  reg _ram_w8_l2048_id0_3_cond_2_2;
  wire signed [8-1:0] _tmp_480;
  wire _tmp_481;
  assign _tmp_480 = (__tmp_475_2 == 0)? ram_w8_l2048_id0_0_0_rdata : 
                    (__tmp_475_2 == 1)? ram_w8_l2048_id0_1_0_rdata : 
                    (__tmp_475_2 == 2)? ram_w8_l2048_id0_2_0_rdata : 
                    (__tmp_475_2 == 3)? ram_w8_l2048_id0_3_0_rdata : 0;
  assign _tmp_481 = _tmp_476;
  assign _stream_conv2d_16_source_8_source_ram_rdata = (_stream_conv2d_16_source_8_source_ram_sel == 2)? _tmp_480 : 0;
  localparam _tmp_482 = 1;
  wire [_tmp_482-1:0] _tmp_483;
  assign _tmp_483 = _stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2);
  reg [_tmp_482-1:0] __tmp_483_1;
  reg [8-1:0] __variable_wdata_237;
  assign stream_conv2d_16_source_8_data = __variable_wdata_237;
  reg [32-1:0] _stream_conv2d_16_source_8_source_pat_fsm_1;
  localparam _stream_conv2d_16_source_8_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_8_source_pat_all_offset;
  assign _stream_conv2d_16_source_8_source_pat_all_offset = _stream_conv2d_16_source_8_source_offset_buf + _source_stream_conv2d_16_source_8_pat_cur_offset_0 + _source_stream_conv2d_16_source_8_pat_cur_offset_1 + _source_stream_conv2d_16_source_8_pat_cur_offset_2 + _source_stream_conv2d_16_source_8_pat_cur_offset_3;
  reg _set_flag_484;
  reg [1-1:0] __variable_wdata_243;
  assign stream_conv2d_16_constant_9_data = __variable_wdata_243;
  reg _set_flag_485;
  reg [8-1:0] __variable_wdata_244;
  assign stream_conv2d_16_source_10_data = __variable_wdata_244;
  reg _set_flag_486;
  reg [1-1:0] __variable_wdata_250;
  assign stream_conv2d_16_constant_11_data = __variable_wdata_250;
  reg _set_flag_487;
  reg [8-1:0] __variable_wdata_251;
  assign stream_conv2d_16_source_12_data = __variable_wdata_251;
  reg _set_flag_488;
  reg [1-1:0] __variable_wdata_257;
  assign stream_conv2d_16_constant_13_data = __variable_wdata_257;
  reg _set_flag_489;
  reg [8-1:0] __variable_wdata_258;
  assign stream_conv2d_16_source_14_data = __variable_wdata_258;
  reg _set_flag_490;
  reg [1-1:0] __variable_wdata_264;
  assign stream_conv2d_16_constant_15_data = __variable_wdata_264;
  reg _set_flag_491;
  reg [1-1:0] __variable_wdata_265;
  assign stream_conv2d_16_constant_16_data = __variable_wdata_265;
  reg _set_flag_492;
  reg [4-1:0] __variable_wdata_266;
  assign stream_conv2d_16_constant_17_data = __variable_wdata_266;
  reg _set_flag_493;
  reg [1-1:0] __variable_wdata_267;
  assign stream_conv2d_16_constant_18_data = __variable_wdata_267;
  reg [32-1:0] _source_stream_conv2d_16_source_19_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_19_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_19_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_19_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_19_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_19_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_19_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_19_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_19_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_19_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_19_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_19_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_19_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_19_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_19_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_19_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_19_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_19_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_19_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_19_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_19_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_19_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_19_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_19_pat_stride_buf_3;
  reg _set_flag_494;
  wire [2-1:0] _tmp_495;
  assign _tmp_495 = _stream_conv2d_16_source_19_source_ram_raddr;
  reg [2-1:0] __tmp_495_1;
  reg [2-1:0] __tmp_495_2;
  reg _tmp_496;
  reg _ram_w8_l2048_id2_0_cond_2_1;
  reg _ram_w8_l2048_id2_0_cond_3_1;
  reg _ram_w8_l2048_id2_0_cond_3_2;
  reg _tmp_497;
  reg _ram_w8_l2048_id2_1_cond_2_1;
  reg _ram_w8_l2048_id2_1_cond_3_1;
  reg _ram_w8_l2048_id2_1_cond_3_2;
  reg _tmp_498;
  reg _ram_w8_l2048_id2_2_cond_2_1;
  reg _ram_w8_l2048_id2_2_cond_3_1;
  reg _ram_w8_l2048_id2_2_cond_3_2;
  reg _tmp_499;
  reg _ram_w8_l2048_id2_3_cond_2_1;
  reg _ram_w8_l2048_id2_3_cond_3_1;
  reg _ram_w8_l2048_id2_3_cond_3_2;
  wire signed [8-1:0] _tmp_500;
  wire _tmp_501;
  assign _tmp_500 = (__tmp_495_2 == 0)? ram_w8_l2048_id2_0_0_rdata : 
                    (__tmp_495_2 == 1)? ram_w8_l2048_id2_1_0_rdata : 
                    (__tmp_495_2 == 2)? ram_w8_l2048_id2_2_0_rdata : 
                    (__tmp_495_2 == 3)? ram_w8_l2048_id2_3_0_rdata : 0;
  assign _tmp_501 = _tmp_496;
  assign _stream_conv2d_16_source_19_source_ram_rdata = (_stream_conv2d_16_source_19_source_ram_sel == 3)? _tmp_500 : 0;
  localparam _tmp_502 = 1;
  wire [_tmp_502-1:0] _tmp_503;
  assign _tmp_503 = _stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3);
  reg [_tmp_502-1:0] __tmp_503_1;
  reg [8-1:0] __variable_wdata_268;
  assign stream_conv2d_16_source_19_data = __variable_wdata_268;
  reg [32-1:0] _stream_conv2d_16_source_19_source_pat_fsm_2;
  localparam _stream_conv2d_16_source_19_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_19_source_pat_all_offset;
  assign _stream_conv2d_16_source_19_source_pat_all_offset = _stream_conv2d_16_source_19_source_offset_buf + _source_stream_conv2d_16_source_19_pat_cur_offset_0 + _source_stream_conv2d_16_source_19_pat_cur_offset_1 + _source_stream_conv2d_16_source_19_pat_cur_offset_2 + _source_stream_conv2d_16_source_19_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_20_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_20_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_20_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_20_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_20_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_20_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_20_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_20_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_20_pat_stride_buf_3;
  reg _set_flag_504;
  wire [2-1:0] _tmp_505;
  assign _tmp_505 = _stream_conv2d_16_source_20_source_ram_raddr;
  reg [2-1:0] __tmp_505_1;
  reg [2-1:0] __tmp_505_2;
  reg _tmp_506;
  reg _ram_w8_l2048_id3_0_cond_1_1;
  reg _ram_w8_l2048_id3_0_cond_2_1;
  reg _ram_w8_l2048_id3_0_cond_2_2;
  reg _tmp_507;
  reg _ram_w8_l2048_id3_1_cond_1_1;
  reg _ram_w8_l2048_id3_1_cond_2_1;
  reg _ram_w8_l2048_id3_1_cond_2_2;
  reg _tmp_508;
  reg _ram_w8_l2048_id3_2_cond_1_1;
  reg _ram_w8_l2048_id3_2_cond_2_1;
  reg _ram_w8_l2048_id3_2_cond_2_2;
  reg _tmp_509;
  reg _ram_w8_l2048_id3_3_cond_1_1;
  reg _ram_w8_l2048_id3_3_cond_2_1;
  reg _ram_w8_l2048_id3_3_cond_2_2;
  wire signed [8-1:0] _tmp_510;
  wire _tmp_511;
  assign _tmp_510 = (__tmp_505_2 == 0)? ram_w8_l2048_id3_0_0_rdata : 
                    (__tmp_505_2 == 1)? ram_w8_l2048_id3_1_0_rdata : 
                    (__tmp_505_2 == 2)? ram_w8_l2048_id3_2_0_rdata : 
                    (__tmp_505_2 == 3)? ram_w8_l2048_id3_3_0_rdata : 0;
  assign _tmp_511 = _tmp_506;
  assign _stream_conv2d_16_source_20_source_ram_rdata = (_stream_conv2d_16_source_20_source_ram_sel == 4)? _tmp_510 : 0;
  localparam _tmp_512 = 1;
  wire [_tmp_512-1:0] _tmp_513;
  assign _tmp_513 = _stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4);
  reg [_tmp_512-1:0] __tmp_513_1;
  reg [8-1:0] __variable_wdata_269;
  assign stream_conv2d_16_source_20_data = __variable_wdata_269;
  reg [32-1:0] _stream_conv2d_16_source_20_source_pat_fsm_3;
  localparam _stream_conv2d_16_source_20_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_20_source_pat_all_offset;
  assign _stream_conv2d_16_source_20_source_pat_all_offset = _stream_conv2d_16_source_20_source_offset_buf + _source_stream_conv2d_16_source_20_pat_cur_offset_0 + _source_stream_conv2d_16_source_20_pat_cur_offset_1 + _source_stream_conv2d_16_source_20_pat_cur_offset_2 + _source_stream_conv2d_16_source_20_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_21_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_21_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_21_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_21_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_21_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_21_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_21_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_21_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_21_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_21_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_21_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_21_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_21_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_21_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_21_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_21_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_21_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_21_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_21_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_21_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_21_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_21_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_21_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_21_pat_stride_buf_3;
  reg _set_flag_514;
  wire [2-1:0] _tmp_515;
  assign _tmp_515 = _stream_conv2d_16_source_21_source_ram_raddr;
  reg [2-1:0] __tmp_515_1;
  reg [2-1:0] __tmp_515_2;
  reg _tmp_516;
  reg _ram_w8_l2048_id4_0_cond_1_1;
  reg _ram_w8_l2048_id4_0_cond_2_1;
  reg _ram_w8_l2048_id4_0_cond_2_2;
  reg _tmp_517;
  reg _ram_w8_l2048_id4_1_cond_1_1;
  reg _ram_w8_l2048_id4_1_cond_2_1;
  reg _ram_w8_l2048_id4_1_cond_2_2;
  reg _tmp_518;
  reg _ram_w8_l2048_id4_2_cond_1_1;
  reg _ram_w8_l2048_id4_2_cond_2_1;
  reg _ram_w8_l2048_id4_2_cond_2_2;
  reg _tmp_519;
  reg _ram_w8_l2048_id4_3_cond_1_1;
  reg _ram_w8_l2048_id4_3_cond_2_1;
  reg _ram_w8_l2048_id4_3_cond_2_2;
  wire signed [8-1:0] _tmp_520;
  wire _tmp_521;
  assign _tmp_520 = (__tmp_515_2 == 0)? ram_w8_l2048_id4_0_0_rdata : 
                    (__tmp_515_2 == 1)? ram_w8_l2048_id4_1_0_rdata : 
                    (__tmp_515_2 == 2)? ram_w8_l2048_id4_2_0_rdata : 
                    (__tmp_515_2 == 3)? ram_w8_l2048_id4_3_0_rdata : 0;
  assign _tmp_521 = _tmp_516;
  assign _stream_conv2d_16_source_21_source_ram_rdata = (_stream_conv2d_16_source_21_source_ram_sel == 5)? _tmp_520 : 0;
  localparam _tmp_522 = 1;
  wire [_tmp_522-1:0] _tmp_523;
  assign _tmp_523 = _stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5);
  reg [_tmp_522-1:0] __tmp_523_1;
  reg [8-1:0] __variable_wdata_270;
  assign stream_conv2d_16_source_21_data = __variable_wdata_270;
  reg [32-1:0] _stream_conv2d_16_source_21_source_pat_fsm_4;
  localparam _stream_conv2d_16_source_21_source_pat_fsm_4_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_21_source_pat_all_offset;
  assign _stream_conv2d_16_source_21_source_pat_all_offset = _stream_conv2d_16_source_21_source_offset_buf + _source_stream_conv2d_16_source_21_pat_cur_offset_0 + _source_stream_conv2d_16_source_21_pat_cur_offset_1 + _source_stream_conv2d_16_source_21_pat_cur_offset_2 + _source_stream_conv2d_16_source_21_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_22_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_22_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_22_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_22_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_22_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_22_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_22_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_22_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_22_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_22_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_22_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_22_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_22_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_22_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_22_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_22_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_22_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_22_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_22_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_22_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_22_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_22_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_22_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_22_pat_stride_buf_3;
  reg _set_flag_524;
  wire [2-1:0] _tmp_525;
  assign _tmp_525 = _stream_conv2d_16_source_22_source_ram_raddr;
  reg [2-1:0] __tmp_525_1;
  reg [2-1:0] __tmp_525_2;
  reg _tmp_526;
  reg _ram_w8_l2048_id5_0_cond_2_1;
  reg _ram_w8_l2048_id5_0_cond_3_1;
  reg _ram_w8_l2048_id5_0_cond_3_2;
  reg _tmp_527;
  reg _ram_w8_l2048_id5_1_cond_2_1;
  reg _ram_w8_l2048_id5_1_cond_3_1;
  reg _ram_w8_l2048_id5_1_cond_3_2;
  reg _tmp_528;
  reg _ram_w8_l2048_id5_2_cond_2_1;
  reg _ram_w8_l2048_id5_2_cond_3_1;
  reg _ram_w8_l2048_id5_2_cond_3_2;
  reg _tmp_529;
  reg _ram_w8_l2048_id5_3_cond_2_1;
  reg _ram_w8_l2048_id5_3_cond_3_1;
  reg _ram_w8_l2048_id5_3_cond_3_2;
  wire signed [8-1:0] _tmp_530;
  wire _tmp_531;
  assign _tmp_530 = (__tmp_525_2 == 0)? ram_w8_l2048_id5_0_0_rdata : 
                    (__tmp_525_2 == 1)? ram_w8_l2048_id5_1_0_rdata : 
                    (__tmp_525_2 == 2)? ram_w8_l2048_id5_2_0_rdata : 
                    (__tmp_525_2 == 3)? ram_w8_l2048_id5_3_0_rdata : 0;
  assign _tmp_531 = _tmp_526;
  assign _stream_conv2d_16_source_22_source_ram_rdata = (_stream_conv2d_16_source_22_source_ram_sel == 6)? _tmp_530 : 0;
  localparam _tmp_532 = 1;
  wire [_tmp_532-1:0] _tmp_533;
  assign _tmp_533 = _stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6);
  reg [_tmp_532-1:0] __tmp_533_1;
  reg [8-1:0] __variable_wdata_271;
  assign stream_conv2d_16_source_22_data = __variable_wdata_271;
  reg [32-1:0] _stream_conv2d_16_source_22_source_pat_fsm_5;
  localparam _stream_conv2d_16_source_22_source_pat_fsm_5_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_22_source_pat_all_offset;
  assign _stream_conv2d_16_source_22_source_pat_all_offset = _stream_conv2d_16_source_22_source_offset_buf + _source_stream_conv2d_16_source_22_pat_cur_offset_0 + _source_stream_conv2d_16_source_22_pat_cur_offset_1 + _source_stream_conv2d_16_source_22_pat_cur_offset_2 + _source_stream_conv2d_16_source_22_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_23_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_23_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_23_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_23_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_23_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_23_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_23_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_23_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_23_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_23_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_23_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_23_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_23_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_23_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_23_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_23_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_23_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_23_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_23_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_23_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_23_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_23_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_23_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_23_pat_stride_buf_3;
  reg _set_flag_534;
  wire [2-1:0] _tmp_535;
  assign _tmp_535 = _stream_conv2d_16_source_23_source_ram_raddr;
  reg [2-1:0] __tmp_535_1;
  reg [2-1:0] __tmp_535_2;
  reg _tmp_536;
  reg _ram_w8_l2048_id6_0_cond_1_1;
  reg _ram_w8_l2048_id6_0_cond_2_1;
  reg _ram_w8_l2048_id6_0_cond_2_2;
  reg _tmp_537;
  reg _ram_w8_l2048_id6_1_cond_1_1;
  reg _ram_w8_l2048_id6_1_cond_2_1;
  reg _ram_w8_l2048_id6_1_cond_2_2;
  reg _tmp_538;
  reg _ram_w8_l2048_id6_2_cond_1_1;
  reg _ram_w8_l2048_id6_2_cond_2_1;
  reg _ram_w8_l2048_id6_2_cond_2_2;
  reg _tmp_539;
  reg _ram_w8_l2048_id6_3_cond_1_1;
  reg _ram_w8_l2048_id6_3_cond_2_1;
  reg _ram_w8_l2048_id6_3_cond_2_2;
  wire signed [8-1:0] _tmp_540;
  wire _tmp_541;
  assign _tmp_540 = (__tmp_535_2 == 0)? ram_w8_l2048_id6_0_0_rdata : 
                    (__tmp_535_2 == 1)? ram_w8_l2048_id6_1_0_rdata : 
                    (__tmp_535_2 == 2)? ram_w8_l2048_id6_2_0_rdata : 
                    (__tmp_535_2 == 3)? ram_w8_l2048_id6_3_0_rdata : 0;
  assign _tmp_541 = _tmp_536;
  assign _stream_conv2d_16_source_23_source_ram_rdata = (_stream_conv2d_16_source_23_source_ram_sel == 7)? _tmp_540 : 0;
  localparam _tmp_542 = 1;
  wire [_tmp_542-1:0] _tmp_543;
  assign _tmp_543 = _stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7);
  reg [_tmp_542-1:0] __tmp_543_1;
  reg [8-1:0] __variable_wdata_272;
  assign stream_conv2d_16_source_23_data = __variable_wdata_272;
  reg [32-1:0] _stream_conv2d_16_source_23_source_pat_fsm_6;
  localparam _stream_conv2d_16_source_23_source_pat_fsm_6_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_23_source_pat_all_offset;
  assign _stream_conv2d_16_source_23_source_pat_all_offset = _stream_conv2d_16_source_23_source_offset_buf + _source_stream_conv2d_16_source_23_pat_cur_offset_0 + _source_stream_conv2d_16_source_23_pat_cur_offset_1 + _source_stream_conv2d_16_source_23_pat_cur_offset_2 + _source_stream_conv2d_16_source_23_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_24_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_24_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_24_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_24_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_24_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_24_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_24_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_24_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_24_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_24_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_24_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_24_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_24_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_24_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_24_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_24_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_24_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_24_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_24_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_24_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_24_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_24_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_24_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_24_pat_stride_buf_3;
  reg _set_flag_544;
  wire [2-1:0] _tmp_545;
  assign _tmp_545 = _stream_conv2d_16_source_24_source_ram_raddr;
  reg [2-1:0] __tmp_545_1;
  reg [2-1:0] __tmp_545_2;
  reg _tmp_546;
  reg _ram_w8_l2048_id7_0_cond_1_1;
  reg _ram_w8_l2048_id7_0_cond_2_1;
  reg _ram_w8_l2048_id7_0_cond_2_2;
  reg _tmp_547;
  reg _ram_w8_l2048_id7_1_cond_1_1;
  reg _ram_w8_l2048_id7_1_cond_2_1;
  reg _ram_w8_l2048_id7_1_cond_2_2;
  reg _tmp_548;
  reg _ram_w8_l2048_id7_2_cond_1_1;
  reg _ram_w8_l2048_id7_2_cond_2_1;
  reg _ram_w8_l2048_id7_2_cond_2_2;
  reg _tmp_549;
  reg _ram_w8_l2048_id7_3_cond_1_1;
  reg _ram_w8_l2048_id7_3_cond_2_1;
  reg _ram_w8_l2048_id7_3_cond_2_2;
  wire signed [8-1:0] _tmp_550;
  wire _tmp_551;
  assign _tmp_550 = (__tmp_545_2 == 0)? ram_w8_l2048_id7_0_0_rdata : 
                    (__tmp_545_2 == 1)? ram_w8_l2048_id7_1_0_rdata : 
                    (__tmp_545_2 == 2)? ram_w8_l2048_id7_2_0_rdata : 
                    (__tmp_545_2 == 3)? ram_w8_l2048_id7_3_0_rdata : 0;
  assign _tmp_551 = _tmp_546;
  assign _stream_conv2d_16_source_24_source_ram_rdata = (_stream_conv2d_16_source_24_source_ram_sel == 8)? _tmp_550 : 0;
  localparam _tmp_552 = 1;
  wire [_tmp_552-1:0] _tmp_553;
  assign _tmp_553 = _stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8);
  reg [_tmp_552-1:0] __tmp_553_1;
  reg [8-1:0] __variable_wdata_273;
  assign stream_conv2d_16_source_24_data = __variable_wdata_273;
  reg [32-1:0] _stream_conv2d_16_source_24_source_pat_fsm_7;
  localparam _stream_conv2d_16_source_24_source_pat_fsm_7_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_24_source_pat_all_offset;
  assign _stream_conv2d_16_source_24_source_pat_all_offset = _stream_conv2d_16_source_24_source_offset_buf + _source_stream_conv2d_16_source_24_pat_cur_offset_0 + _source_stream_conv2d_16_source_24_pat_cur_offset_1 + _source_stream_conv2d_16_source_24_pat_cur_offset_2 + _source_stream_conv2d_16_source_24_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_25_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_25_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_25_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_25_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_25_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_25_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_25_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_25_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_25_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_25_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_25_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_25_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_25_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_25_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_25_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_25_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_25_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_25_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_25_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_25_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_25_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_25_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_25_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_25_pat_stride_buf_3;
  reg _set_flag_554;
  wire [2-1:0] _tmp_555;
  assign _tmp_555 = _stream_conv2d_16_source_25_source_ram_raddr;
  reg [2-1:0] __tmp_555_1;
  reg [2-1:0] __tmp_555_2;
  reg _tmp_556;
  reg _ram_w8_l2048_id8_0_cond_2_1;
  reg _ram_w8_l2048_id8_0_cond_3_1;
  reg _ram_w8_l2048_id8_0_cond_3_2;
  reg _tmp_557;
  reg _ram_w8_l2048_id8_1_cond_2_1;
  reg _ram_w8_l2048_id8_1_cond_3_1;
  reg _ram_w8_l2048_id8_1_cond_3_2;
  reg _tmp_558;
  reg _ram_w8_l2048_id8_2_cond_2_1;
  reg _ram_w8_l2048_id8_2_cond_3_1;
  reg _ram_w8_l2048_id8_2_cond_3_2;
  reg _tmp_559;
  reg _ram_w8_l2048_id8_3_cond_2_1;
  reg _ram_w8_l2048_id8_3_cond_3_1;
  reg _ram_w8_l2048_id8_3_cond_3_2;
  wire signed [8-1:0] _tmp_560;
  wire _tmp_561;
  assign _tmp_560 = (__tmp_555_2 == 0)? ram_w8_l2048_id8_0_0_rdata : 
                    (__tmp_555_2 == 1)? ram_w8_l2048_id8_1_0_rdata : 
                    (__tmp_555_2 == 2)? ram_w8_l2048_id8_2_0_rdata : 
                    (__tmp_555_2 == 3)? ram_w8_l2048_id8_3_0_rdata : 0;
  assign _tmp_561 = _tmp_556;
  assign _stream_conv2d_16_source_25_source_ram_rdata = (_stream_conv2d_16_source_25_source_ram_sel == 9)? _tmp_560 : 0;
  localparam _tmp_562 = 1;
  wire [_tmp_562-1:0] _tmp_563;
  assign _tmp_563 = _stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9);
  reg [_tmp_562-1:0] __tmp_563_1;
  reg [8-1:0] __variable_wdata_274;
  assign stream_conv2d_16_source_25_data = __variable_wdata_274;
  reg [32-1:0] _stream_conv2d_16_source_25_source_pat_fsm_8;
  localparam _stream_conv2d_16_source_25_source_pat_fsm_8_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_25_source_pat_all_offset;
  assign _stream_conv2d_16_source_25_source_pat_all_offset = _stream_conv2d_16_source_25_source_offset_buf + _source_stream_conv2d_16_source_25_pat_cur_offset_0 + _source_stream_conv2d_16_source_25_pat_cur_offset_1 + _source_stream_conv2d_16_source_25_pat_cur_offset_2 + _source_stream_conv2d_16_source_25_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_26_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_26_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_26_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_26_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_26_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_26_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_26_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_26_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_26_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_26_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_26_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_26_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_26_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_26_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_26_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_26_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_26_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_26_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_26_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_26_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_26_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_26_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_26_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_26_pat_stride_buf_3;
  reg _set_flag_564;
  wire [2-1:0] _tmp_565;
  assign _tmp_565 = _stream_conv2d_16_source_26_source_ram_raddr;
  reg [2-1:0] __tmp_565_1;
  reg [2-1:0] __tmp_565_2;
  reg _tmp_566;
  reg _ram_w8_l2048_id9_0_cond_1_1;
  reg _ram_w8_l2048_id9_0_cond_2_1;
  reg _ram_w8_l2048_id9_0_cond_2_2;
  reg _tmp_567;
  reg _ram_w8_l2048_id9_1_cond_1_1;
  reg _ram_w8_l2048_id9_1_cond_2_1;
  reg _ram_w8_l2048_id9_1_cond_2_2;
  reg _tmp_568;
  reg _ram_w8_l2048_id9_2_cond_1_1;
  reg _ram_w8_l2048_id9_2_cond_2_1;
  reg _ram_w8_l2048_id9_2_cond_2_2;
  reg _tmp_569;
  reg _ram_w8_l2048_id9_3_cond_1_1;
  reg _ram_w8_l2048_id9_3_cond_2_1;
  reg _ram_w8_l2048_id9_3_cond_2_2;
  wire signed [8-1:0] _tmp_570;
  wire _tmp_571;
  assign _tmp_570 = (__tmp_565_2 == 0)? ram_w8_l2048_id9_0_0_rdata : 
                    (__tmp_565_2 == 1)? ram_w8_l2048_id9_1_0_rdata : 
                    (__tmp_565_2 == 2)? ram_w8_l2048_id9_2_0_rdata : 
                    (__tmp_565_2 == 3)? ram_w8_l2048_id9_3_0_rdata : 0;
  assign _tmp_571 = _tmp_566;
  assign _stream_conv2d_16_source_26_source_ram_rdata = (_stream_conv2d_16_source_26_source_ram_sel == 10)? _tmp_570 : 0;
  localparam _tmp_572 = 1;
  wire [_tmp_572-1:0] _tmp_573;
  assign _tmp_573 = _stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10);
  reg [_tmp_572-1:0] __tmp_573_1;
  reg [8-1:0] __variable_wdata_275;
  assign stream_conv2d_16_source_26_data = __variable_wdata_275;
  reg [32-1:0] _stream_conv2d_16_source_26_source_pat_fsm_9;
  localparam _stream_conv2d_16_source_26_source_pat_fsm_9_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_26_source_pat_all_offset;
  assign _stream_conv2d_16_source_26_source_pat_all_offset = _stream_conv2d_16_source_26_source_offset_buf + _source_stream_conv2d_16_source_26_pat_cur_offset_0 + _source_stream_conv2d_16_source_26_pat_cur_offset_1 + _source_stream_conv2d_16_source_26_pat_cur_offset_2 + _source_stream_conv2d_16_source_26_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_27_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_27_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_27_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_27_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_27_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_27_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_27_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_27_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_27_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_27_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_27_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_27_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_27_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_27_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_27_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_27_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_27_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_27_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_27_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_27_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_27_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_27_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_27_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_27_pat_stride_buf_3;
  reg _set_flag_574;
  wire [2-1:0] _tmp_575;
  assign _tmp_575 = _stream_conv2d_16_source_27_source_ram_raddr;
  reg [2-1:0] __tmp_575_1;
  reg [2-1:0] __tmp_575_2;
  reg _tmp_576;
  reg _ram_w8_l2048_id10_0_cond_1_1;
  reg _ram_w8_l2048_id10_0_cond_2_1;
  reg _ram_w8_l2048_id10_0_cond_2_2;
  reg _tmp_577;
  reg _ram_w8_l2048_id10_1_cond_1_1;
  reg _ram_w8_l2048_id10_1_cond_2_1;
  reg _ram_w8_l2048_id10_1_cond_2_2;
  reg _tmp_578;
  reg _ram_w8_l2048_id10_2_cond_1_1;
  reg _ram_w8_l2048_id10_2_cond_2_1;
  reg _ram_w8_l2048_id10_2_cond_2_2;
  reg _tmp_579;
  reg _ram_w8_l2048_id10_3_cond_1_1;
  reg _ram_w8_l2048_id10_3_cond_2_1;
  reg _ram_w8_l2048_id10_3_cond_2_2;
  wire signed [8-1:0] _tmp_580;
  wire _tmp_581;
  assign _tmp_580 = (__tmp_575_2 == 0)? ram_w8_l2048_id10_0_0_rdata : 
                    (__tmp_575_2 == 1)? ram_w8_l2048_id10_1_0_rdata : 
                    (__tmp_575_2 == 2)? ram_w8_l2048_id10_2_0_rdata : 
                    (__tmp_575_2 == 3)? ram_w8_l2048_id10_3_0_rdata : 0;
  assign _tmp_581 = _tmp_576;
  assign _stream_conv2d_16_source_27_source_ram_rdata = (_stream_conv2d_16_source_27_source_ram_sel == 11)? _tmp_580 : 0;
  localparam _tmp_582 = 1;
  wire [_tmp_582-1:0] _tmp_583;
  assign _tmp_583 = _stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11);
  reg [_tmp_582-1:0] __tmp_583_1;
  reg [8-1:0] __variable_wdata_276;
  assign stream_conv2d_16_source_27_data = __variable_wdata_276;
  reg [32-1:0] _stream_conv2d_16_source_27_source_pat_fsm_10;
  localparam _stream_conv2d_16_source_27_source_pat_fsm_10_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_27_source_pat_all_offset;
  assign _stream_conv2d_16_source_27_source_pat_all_offset = _stream_conv2d_16_source_27_source_offset_buf + _source_stream_conv2d_16_source_27_pat_cur_offset_0 + _source_stream_conv2d_16_source_27_pat_cur_offset_1 + _source_stream_conv2d_16_source_27_pat_cur_offset_2 + _source_stream_conv2d_16_source_27_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_28_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_28_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_28_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_28_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_28_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_28_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_28_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_28_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_28_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_28_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_28_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_28_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_28_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_28_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_28_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_28_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_28_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_28_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_28_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_28_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_28_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_28_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_28_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_28_pat_stride_buf_3;
  reg _set_flag_584;
  wire [3-1:0] _tmp_585;
  assign _tmp_585 = _stream_conv2d_16_source_28_source_ram_raddr;
  reg [3-1:0] __tmp_585_1;
  reg [3-1:0] __tmp_585_2;
  reg _tmp_586;
  reg _ram_w4_l8192_id0_0_cond_2_1;
  reg _ram_w4_l8192_id0_0_cond_3_1;
  reg _ram_w4_l8192_id0_0_cond_3_2;
  reg _tmp_587;
  reg _ram_w4_l8192_id0_1_cond_2_1;
  reg _ram_w4_l8192_id0_1_cond_3_1;
  reg _ram_w4_l8192_id0_1_cond_3_2;
  reg _tmp_588;
  reg _ram_w4_l8192_id0_2_cond_2_1;
  reg _ram_w4_l8192_id0_2_cond_3_1;
  reg _ram_w4_l8192_id0_2_cond_3_2;
  reg _tmp_589;
  reg _ram_w4_l8192_id0_3_cond_2_1;
  reg _ram_w4_l8192_id0_3_cond_3_1;
  reg _ram_w4_l8192_id0_3_cond_3_2;
  reg _tmp_590;
  reg _ram_w4_l8192_id0_4_cond_2_1;
  reg _ram_w4_l8192_id0_4_cond_3_1;
  reg _ram_w4_l8192_id0_4_cond_3_2;
  reg _tmp_591;
  reg _ram_w4_l8192_id0_5_cond_2_1;
  reg _ram_w4_l8192_id0_5_cond_3_1;
  reg _ram_w4_l8192_id0_5_cond_3_2;
  reg _tmp_592;
  reg _ram_w4_l8192_id0_6_cond_2_1;
  reg _ram_w4_l8192_id0_6_cond_3_1;
  reg _ram_w4_l8192_id0_6_cond_3_2;
  reg _tmp_593;
  reg _ram_w4_l8192_id0_7_cond_2_1;
  reg _ram_w4_l8192_id0_7_cond_3_1;
  reg _ram_w4_l8192_id0_7_cond_3_2;
  wire signed [4-1:0] _tmp_594;
  wire _tmp_595;
  assign _tmp_594 = (__tmp_585_2 == 0)? ram_w4_l8192_id0_0_0_rdata : 
                    (__tmp_585_2 == 1)? ram_w4_l8192_id0_1_0_rdata : 
                    (__tmp_585_2 == 2)? ram_w4_l8192_id0_2_0_rdata : 
                    (__tmp_585_2 == 3)? ram_w4_l8192_id0_3_0_rdata : 
                    (__tmp_585_2 == 4)? ram_w4_l8192_id0_4_0_rdata : 
                    (__tmp_585_2 == 5)? ram_w4_l8192_id0_5_0_rdata : 
                    (__tmp_585_2 == 6)? ram_w4_l8192_id0_6_0_rdata : 
                    (__tmp_585_2 == 7)? ram_w4_l8192_id0_7_0_rdata : 0;
  assign _tmp_595 = _tmp_586;
  assign _stream_conv2d_16_source_28_source_ram_rdata = (_stream_conv2d_16_source_28_source_ram_sel == 12)? _tmp_594 : 0;
  localparam _tmp_596 = 1;
  wire [_tmp_596-1:0] _tmp_597;
  assign _tmp_597 = _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
  reg [_tmp_596-1:0] __tmp_597_1;
  reg [4-1:0] __variable_wdata_502;
  assign stream_conv2d_16_source_28_data = __variable_wdata_502;
  reg [32-1:0] _stream_conv2d_16_source_28_source_pat_fsm_11;
  localparam _stream_conv2d_16_source_28_source_pat_fsm_11_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_28_source_pat_all_offset;
  assign _stream_conv2d_16_source_28_source_pat_all_offset = _stream_conv2d_16_source_28_source_offset_buf + _source_stream_conv2d_16_source_28_pat_cur_offset_0 + _source_stream_conv2d_16_source_28_pat_cur_offset_1 + _source_stream_conv2d_16_source_28_pat_cur_offset_2 + _source_stream_conv2d_16_source_28_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_29_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_29_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_29_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_29_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_29_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_29_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_29_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_29_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_29_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_29_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_29_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_29_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_29_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_29_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_29_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_29_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_29_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_29_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_29_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_29_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_29_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_29_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_29_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_29_pat_stride_buf_3;
  reg _set_flag_598;
  wire [3-1:0] _tmp_599;
  assign _tmp_599 = _stream_conv2d_16_source_29_source_ram_raddr;
  reg [3-1:0] __tmp_599_1;
  reg [3-1:0] __tmp_599_2;
  reg _tmp_600;
  reg _ram_w4_l8192_id1_0_cond_1_1;
  reg _ram_w4_l8192_id1_0_cond_2_1;
  reg _ram_w4_l8192_id1_0_cond_2_2;
  reg _tmp_601;
  reg _ram_w4_l8192_id1_1_cond_1_1;
  reg _ram_w4_l8192_id1_1_cond_2_1;
  reg _ram_w4_l8192_id1_1_cond_2_2;
  reg _tmp_602;
  reg _ram_w4_l8192_id1_2_cond_1_1;
  reg _ram_w4_l8192_id1_2_cond_2_1;
  reg _ram_w4_l8192_id1_2_cond_2_2;
  reg _tmp_603;
  reg _ram_w4_l8192_id1_3_cond_1_1;
  reg _ram_w4_l8192_id1_3_cond_2_1;
  reg _ram_w4_l8192_id1_3_cond_2_2;
  reg _tmp_604;
  reg _ram_w4_l8192_id1_4_cond_1_1;
  reg _ram_w4_l8192_id1_4_cond_2_1;
  reg _ram_w4_l8192_id1_4_cond_2_2;
  reg _tmp_605;
  reg _ram_w4_l8192_id1_5_cond_1_1;
  reg _ram_w4_l8192_id1_5_cond_2_1;
  reg _ram_w4_l8192_id1_5_cond_2_2;
  reg _tmp_606;
  reg _ram_w4_l8192_id1_6_cond_1_1;
  reg _ram_w4_l8192_id1_6_cond_2_1;
  reg _ram_w4_l8192_id1_6_cond_2_2;
  reg _tmp_607;
  reg _ram_w4_l8192_id1_7_cond_1_1;
  reg _ram_w4_l8192_id1_7_cond_2_1;
  reg _ram_w4_l8192_id1_7_cond_2_2;
  wire signed [4-1:0] _tmp_608;
  wire _tmp_609;
  assign _tmp_608 = (__tmp_599_2 == 0)? ram_w4_l8192_id1_0_0_rdata : 
                    (__tmp_599_2 == 1)? ram_w4_l8192_id1_1_0_rdata : 
                    (__tmp_599_2 == 2)? ram_w4_l8192_id1_2_0_rdata : 
                    (__tmp_599_2 == 3)? ram_w4_l8192_id1_3_0_rdata : 
                    (__tmp_599_2 == 4)? ram_w4_l8192_id1_4_0_rdata : 
                    (__tmp_599_2 == 5)? ram_w4_l8192_id1_5_0_rdata : 
                    (__tmp_599_2 == 6)? ram_w4_l8192_id1_6_0_rdata : 
                    (__tmp_599_2 == 7)? ram_w4_l8192_id1_7_0_rdata : 0;
  assign _tmp_609 = _tmp_600;
  assign _stream_conv2d_16_source_29_source_ram_rdata = (_stream_conv2d_16_source_29_source_ram_sel == 13)? _tmp_608 : 0;
  localparam _tmp_610 = 1;
  wire [_tmp_610-1:0] _tmp_611;
  assign _tmp_611 = _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
  reg [_tmp_610-1:0] __tmp_611_1;
  reg [4-1:0] __variable_wdata_503;
  assign stream_conv2d_16_source_29_data = __variable_wdata_503;
  reg [32-1:0] _stream_conv2d_16_source_29_source_pat_fsm_12;
  localparam _stream_conv2d_16_source_29_source_pat_fsm_12_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_29_source_pat_all_offset;
  assign _stream_conv2d_16_source_29_source_pat_all_offset = _stream_conv2d_16_source_29_source_offset_buf + _source_stream_conv2d_16_source_29_pat_cur_offset_0 + _source_stream_conv2d_16_source_29_pat_cur_offset_1 + _source_stream_conv2d_16_source_29_pat_cur_offset_2 + _source_stream_conv2d_16_source_29_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_30_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_30_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_30_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_30_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_30_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_30_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_30_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_30_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_30_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_30_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_30_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_30_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_30_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_30_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_30_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_30_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_30_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_30_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_30_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_30_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_30_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_30_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_30_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_30_pat_stride_buf_3;
  reg _set_flag_612;
  wire [3-1:0] _tmp_613;
  assign _tmp_613 = _stream_conv2d_16_source_30_source_ram_raddr;
  reg [3-1:0] __tmp_613_1;
  reg [3-1:0] __tmp_613_2;
  reg _tmp_614;
  reg _ram_w4_l8192_id2_0_cond_1_1;
  reg _ram_w4_l8192_id2_0_cond_2_1;
  reg _ram_w4_l8192_id2_0_cond_2_2;
  reg _tmp_615;
  reg _ram_w4_l8192_id2_1_cond_1_1;
  reg _ram_w4_l8192_id2_1_cond_2_1;
  reg _ram_w4_l8192_id2_1_cond_2_2;
  reg _tmp_616;
  reg _ram_w4_l8192_id2_2_cond_1_1;
  reg _ram_w4_l8192_id2_2_cond_2_1;
  reg _ram_w4_l8192_id2_2_cond_2_2;
  reg _tmp_617;
  reg _ram_w4_l8192_id2_3_cond_1_1;
  reg _ram_w4_l8192_id2_3_cond_2_1;
  reg _ram_w4_l8192_id2_3_cond_2_2;
  reg _tmp_618;
  reg _ram_w4_l8192_id2_4_cond_1_1;
  reg _ram_w4_l8192_id2_4_cond_2_1;
  reg _ram_w4_l8192_id2_4_cond_2_2;
  reg _tmp_619;
  reg _ram_w4_l8192_id2_5_cond_1_1;
  reg _ram_w4_l8192_id2_5_cond_2_1;
  reg _ram_w4_l8192_id2_5_cond_2_2;
  reg _tmp_620;
  reg _ram_w4_l8192_id2_6_cond_1_1;
  reg _ram_w4_l8192_id2_6_cond_2_1;
  reg _ram_w4_l8192_id2_6_cond_2_2;
  reg _tmp_621;
  reg _ram_w4_l8192_id2_7_cond_1_1;
  reg _ram_w4_l8192_id2_7_cond_2_1;
  reg _ram_w4_l8192_id2_7_cond_2_2;
  wire signed [4-1:0] _tmp_622;
  wire _tmp_623;
  assign _tmp_622 = (__tmp_613_2 == 0)? ram_w4_l8192_id2_0_0_rdata : 
                    (__tmp_613_2 == 1)? ram_w4_l8192_id2_1_0_rdata : 
                    (__tmp_613_2 == 2)? ram_w4_l8192_id2_2_0_rdata : 
                    (__tmp_613_2 == 3)? ram_w4_l8192_id2_3_0_rdata : 
                    (__tmp_613_2 == 4)? ram_w4_l8192_id2_4_0_rdata : 
                    (__tmp_613_2 == 5)? ram_w4_l8192_id2_5_0_rdata : 
                    (__tmp_613_2 == 6)? ram_w4_l8192_id2_6_0_rdata : 
                    (__tmp_613_2 == 7)? ram_w4_l8192_id2_7_0_rdata : 0;
  assign _tmp_623 = _tmp_614;
  assign _stream_conv2d_16_source_30_source_ram_rdata = (_stream_conv2d_16_source_30_source_ram_sel == 14)? _tmp_622 : 0;
  localparam _tmp_624 = 1;
  wire [_tmp_624-1:0] _tmp_625;
  assign _tmp_625 = _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
  reg [_tmp_624-1:0] __tmp_625_1;
  reg [4-1:0] __variable_wdata_504;
  assign stream_conv2d_16_source_30_data = __variable_wdata_504;
  reg [32-1:0] _stream_conv2d_16_source_30_source_pat_fsm_13;
  localparam _stream_conv2d_16_source_30_source_pat_fsm_13_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_30_source_pat_all_offset;
  assign _stream_conv2d_16_source_30_source_pat_all_offset = _stream_conv2d_16_source_30_source_offset_buf + _source_stream_conv2d_16_source_30_pat_cur_offset_0 + _source_stream_conv2d_16_source_30_pat_cur_offset_1 + _source_stream_conv2d_16_source_30_pat_cur_offset_2 + _source_stream_conv2d_16_source_30_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_31_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_31_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_31_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_31_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_31_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_31_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_31_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_31_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_31_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_31_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_31_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_31_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_31_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_31_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_31_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_31_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_31_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_31_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_31_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_31_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_31_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_31_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_31_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_31_pat_stride_buf_3;
  reg _set_flag_626;
  wire [3-1:0] _tmp_627;
  assign _tmp_627 = _stream_conv2d_16_source_31_source_ram_raddr;
  reg [3-1:0] __tmp_627_1;
  reg [3-1:0] __tmp_627_2;
  reg _tmp_628;
  reg _ram_w4_l8192_id3_0_cond_1_1;
  reg _ram_w4_l8192_id3_0_cond_2_1;
  reg _ram_w4_l8192_id3_0_cond_2_2;
  reg _tmp_629;
  reg _ram_w4_l8192_id3_1_cond_1_1;
  reg _ram_w4_l8192_id3_1_cond_2_1;
  reg _ram_w4_l8192_id3_1_cond_2_2;
  reg _tmp_630;
  reg _ram_w4_l8192_id3_2_cond_1_1;
  reg _ram_w4_l8192_id3_2_cond_2_1;
  reg _ram_w4_l8192_id3_2_cond_2_2;
  reg _tmp_631;
  reg _ram_w4_l8192_id3_3_cond_1_1;
  reg _ram_w4_l8192_id3_3_cond_2_1;
  reg _ram_w4_l8192_id3_3_cond_2_2;
  reg _tmp_632;
  reg _ram_w4_l8192_id3_4_cond_1_1;
  reg _ram_w4_l8192_id3_4_cond_2_1;
  reg _ram_w4_l8192_id3_4_cond_2_2;
  reg _tmp_633;
  reg _ram_w4_l8192_id3_5_cond_1_1;
  reg _ram_w4_l8192_id3_5_cond_2_1;
  reg _ram_w4_l8192_id3_5_cond_2_2;
  reg _tmp_634;
  reg _ram_w4_l8192_id3_6_cond_1_1;
  reg _ram_w4_l8192_id3_6_cond_2_1;
  reg _ram_w4_l8192_id3_6_cond_2_2;
  reg _tmp_635;
  reg _ram_w4_l8192_id3_7_cond_1_1;
  reg _ram_w4_l8192_id3_7_cond_2_1;
  reg _ram_w4_l8192_id3_7_cond_2_2;
  wire signed [4-1:0] _tmp_636;
  wire _tmp_637;
  assign _tmp_636 = (__tmp_627_2 == 0)? ram_w4_l8192_id3_0_0_rdata : 
                    (__tmp_627_2 == 1)? ram_w4_l8192_id3_1_0_rdata : 
                    (__tmp_627_2 == 2)? ram_w4_l8192_id3_2_0_rdata : 
                    (__tmp_627_2 == 3)? ram_w4_l8192_id3_3_0_rdata : 
                    (__tmp_627_2 == 4)? ram_w4_l8192_id3_4_0_rdata : 
                    (__tmp_627_2 == 5)? ram_w4_l8192_id3_5_0_rdata : 
                    (__tmp_627_2 == 6)? ram_w4_l8192_id3_6_0_rdata : 
                    (__tmp_627_2 == 7)? ram_w4_l8192_id3_7_0_rdata : 0;
  assign _tmp_637 = _tmp_628;
  assign _stream_conv2d_16_source_31_source_ram_rdata = (_stream_conv2d_16_source_31_source_ram_sel == 15)? _tmp_636 : 0;
  localparam _tmp_638 = 1;
  wire [_tmp_638-1:0] _tmp_639;
  assign _tmp_639 = _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
  reg [_tmp_638-1:0] __tmp_639_1;
  reg [4-1:0] __variable_wdata_505;
  assign stream_conv2d_16_source_31_data = __variable_wdata_505;
  reg [32-1:0] _stream_conv2d_16_source_31_source_pat_fsm_14;
  localparam _stream_conv2d_16_source_31_source_pat_fsm_14_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_31_source_pat_all_offset;
  assign _stream_conv2d_16_source_31_source_pat_all_offset = _stream_conv2d_16_source_31_source_offset_buf + _source_stream_conv2d_16_source_31_pat_cur_offset_0 + _source_stream_conv2d_16_source_31_pat_cur_offset_1 + _source_stream_conv2d_16_source_31_pat_cur_offset_2 + _source_stream_conv2d_16_source_31_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_32_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_32_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_32_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_32_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_32_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_32_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_32_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_32_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_32_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_32_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_32_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_32_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_32_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_32_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_32_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_32_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_32_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_32_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_32_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_32_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_32_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_32_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_32_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_32_pat_stride_buf_3;
  reg _set_flag_640;
  wire [3-1:0] _tmp_641;
  assign _tmp_641 = _stream_conv2d_16_source_32_source_ram_raddr;
  reg [3-1:0] __tmp_641_1;
  reg [3-1:0] __tmp_641_2;
  reg _tmp_642;
  reg _ram_w4_l8192_id4_0_cond_1_1;
  reg _ram_w4_l8192_id4_0_cond_2_1;
  reg _ram_w4_l8192_id4_0_cond_2_2;
  reg _tmp_643;
  reg _ram_w4_l8192_id4_1_cond_1_1;
  reg _ram_w4_l8192_id4_1_cond_2_1;
  reg _ram_w4_l8192_id4_1_cond_2_2;
  reg _tmp_644;
  reg _ram_w4_l8192_id4_2_cond_1_1;
  reg _ram_w4_l8192_id4_2_cond_2_1;
  reg _ram_w4_l8192_id4_2_cond_2_2;
  reg _tmp_645;
  reg _ram_w4_l8192_id4_3_cond_1_1;
  reg _ram_w4_l8192_id4_3_cond_2_1;
  reg _ram_w4_l8192_id4_3_cond_2_2;
  reg _tmp_646;
  reg _ram_w4_l8192_id4_4_cond_1_1;
  reg _ram_w4_l8192_id4_4_cond_2_1;
  reg _ram_w4_l8192_id4_4_cond_2_2;
  reg _tmp_647;
  reg _ram_w4_l8192_id4_5_cond_1_1;
  reg _ram_w4_l8192_id4_5_cond_2_1;
  reg _ram_w4_l8192_id4_5_cond_2_2;
  reg _tmp_648;
  reg _ram_w4_l8192_id4_6_cond_1_1;
  reg _ram_w4_l8192_id4_6_cond_2_1;
  reg _ram_w4_l8192_id4_6_cond_2_2;
  reg _tmp_649;
  reg _ram_w4_l8192_id4_7_cond_1_1;
  reg _ram_w4_l8192_id4_7_cond_2_1;
  reg _ram_w4_l8192_id4_7_cond_2_2;
  wire signed [4-1:0] _tmp_650;
  wire _tmp_651;
  assign _tmp_650 = (__tmp_641_2 == 0)? ram_w4_l8192_id4_0_0_rdata : 
                    (__tmp_641_2 == 1)? ram_w4_l8192_id4_1_0_rdata : 
                    (__tmp_641_2 == 2)? ram_w4_l8192_id4_2_0_rdata : 
                    (__tmp_641_2 == 3)? ram_w4_l8192_id4_3_0_rdata : 
                    (__tmp_641_2 == 4)? ram_w4_l8192_id4_4_0_rdata : 
                    (__tmp_641_2 == 5)? ram_w4_l8192_id4_5_0_rdata : 
                    (__tmp_641_2 == 6)? ram_w4_l8192_id4_6_0_rdata : 
                    (__tmp_641_2 == 7)? ram_w4_l8192_id4_7_0_rdata : 0;
  assign _tmp_651 = _tmp_642;
  assign _stream_conv2d_16_source_32_source_ram_rdata = (_stream_conv2d_16_source_32_source_ram_sel == 16)? _tmp_650 : 0;
  localparam _tmp_652 = 1;
  wire [_tmp_652-1:0] _tmp_653;
  assign _tmp_653 = _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
  reg [_tmp_652-1:0] __tmp_653_1;
  reg [4-1:0] __variable_wdata_506;
  assign stream_conv2d_16_source_32_data = __variable_wdata_506;
  reg [32-1:0] _stream_conv2d_16_source_32_source_pat_fsm_15;
  localparam _stream_conv2d_16_source_32_source_pat_fsm_15_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_32_source_pat_all_offset;
  assign _stream_conv2d_16_source_32_source_pat_all_offset = _stream_conv2d_16_source_32_source_offset_buf + _source_stream_conv2d_16_source_32_pat_cur_offset_0 + _source_stream_conv2d_16_source_32_pat_cur_offset_1 + _source_stream_conv2d_16_source_32_pat_cur_offset_2 + _source_stream_conv2d_16_source_32_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_33_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_33_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_33_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_33_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_33_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_33_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_33_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_33_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_33_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_33_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_33_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_33_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_33_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_33_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_33_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_33_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_33_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_33_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_33_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_33_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_33_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_33_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_33_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_33_pat_stride_buf_3;
  reg _set_flag_654;
  wire [3-1:0] _tmp_655;
  assign _tmp_655 = _stream_conv2d_16_source_33_source_ram_raddr;
  reg [3-1:0] __tmp_655_1;
  reg [3-1:0] __tmp_655_2;
  reg _tmp_656;
  reg _ram_w4_l8192_id5_0_cond_1_1;
  reg _ram_w4_l8192_id5_0_cond_2_1;
  reg _ram_w4_l8192_id5_0_cond_2_2;
  reg _tmp_657;
  reg _ram_w4_l8192_id5_1_cond_1_1;
  reg _ram_w4_l8192_id5_1_cond_2_1;
  reg _ram_w4_l8192_id5_1_cond_2_2;
  reg _tmp_658;
  reg _ram_w4_l8192_id5_2_cond_1_1;
  reg _ram_w4_l8192_id5_2_cond_2_1;
  reg _ram_w4_l8192_id5_2_cond_2_2;
  reg _tmp_659;
  reg _ram_w4_l8192_id5_3_cond_1_1;
  reg _ram_w4_l8192_id5_3_cond_2_1;
  reg _ram_w4_l8192_id5_3_cond_2_2;
  reg _tmp_660;
  reg _ram_w4_l8192_id5_4_cond_1_1;
  reg _ram_w4_l8192_id5_4_cond_2_1;
  reg _ram_w4_l8192_id5_4_cond_2_2;
  reg _tmp_661;
  reg _ram_w4_l8192_id5_5_cond_1_1;
  reg _ram_w4_l8192_id5_5_cond_2_1;
  reg _ram_w4_l8192_id5_5_cond_2_2;
  reg _tmp_662;
  reg _ram_w4_l8192_id5_6_cond_1_1;
  reg _ram_w4_l8192_id5_6_cond_2_1;
  reg _ram_w4_l8192_id5_6_cond_2_2;
  reg _tmp_663;
  reg _ram_w4_l8192_id5_7_cond_1_1;
  reg _ram_w4_l8192_id5_7_cond_2_1;
  reg _ram_w4_l8192_id5_7_cond_2_2;
  wire signed [4-1:0] _tmp_664;
  wire _tmp_665;
  assign _tmp_664 = (__tmp_655_2 == 0)? ram_w4_l8192_id5_0_0_rdata : 
                    (__tmp_655_2 == 1)? ram_w4_l8192_id5_1_0_rdata : 
                    (__tmp_655_2 == 2)? ram_w4_l8192_id5_2_0_rdata : 
                    (__tmp_655_2 == 3)? ram_w4_l8192_id5_3_0_rdata : 
                    (__tmp_655_2 == 4)? ram_w4_l8192_id5_4_0_rdata : 
                    (__tmp_655_2 == 5)? ram_w4_l8192_id5_5_0_rdata : 
                    (__tmp_655_2 == 6)? ram_w4_l8192_id5_6_0_rdata : 
                    (__tmp_655_2 == 7)? ram_w4_l8192_id5_7_0_rdata : 0;
  assign _tmp_665 = _tmp_656;
  assign _stream_conv2d_16_source_33_source_ram_rdata = (_stream_conv2d_16_source_33_source_ram_sel == 17)? _tmp_664 : 0;
  localparam _tmp_666 = 1;
  wire [_tmp_666-1:0] _tmp_667;
  assign _tmp_667 = _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
  reg [_tmp_666-1:0] __tmp_667_1;
  reg [4-1:0] __variable_wdata_507;
  assign stream_conv2d_16_source_33_data = __variable_wdata_507;
  reg [32-1:0] _stream_conv2d_16_source_33_source_pat_fsm_16;
  localparam _stream_conv2d_16_source_33_source_pat_fsm_16_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_33_source_pat_all_offset;
  assign _stream_conv2d_16_source_33_source_pat_all_offset = _stream_conv2d_16_source_33_source_offset_buf + _source_stream_conv2d_16_source_33_pat_cur_offset_0 + _source_stream_conv2d_16_source_33_pat_cur_offset_1 + _source_stream_conv2d_16_source_33_pat_cur_offset_2 + _source_stream_conv2d_16_source_33_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_34_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_34_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_34_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_34_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_34_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_34_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_34_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_34_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_34_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_34_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_34_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_34_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_34_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_34_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_34_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_34_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_34_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_34_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_34_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_34_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_34_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_34_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_34_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_34_pat_stride_buf_3;
  reg _set_flag_668;
  wire [3-1:0] _tmp_669;
  assign _tmp_669 = _stream_conv2d_16_source_34_source_ram_raddr;
  reg [3-1:0] __tmp_669_1;
  reg [3-1:0] __tmp_669_2;
  reg _tmp_670;
  reg _ram_w4_l8192_id6_0_cond_1_1;
  reg _ram_w4_l8192_id6_0_cond_2_1;
  reg _ram_w4_l8192_id6_0_cond_2_2;
  reg _tmp_671;
  reg _ram_w4_l8192_id6_1_cond_1_1;
  reg _ram_w4_l8192_id6_1_cond_2_1;
  reg _ram_w4_l8192_id6_1_cond_2_2;
  reg _tmp_672;
  reg _ram_w4_l8192_id6_2_cond_1_1;
  reg _ram_w4_l8192_id6_2_cond_2_1;
  reg _ram_w4_l8192_id6_2_cond_2_2;
  reg _tmp_673;
  reg _ram_w4_l8192_id6_3_cond_1_1;
  reg _ram_w4_l8192_id6_3_cond_2_1;
  reg _ram_w4_l8192_id6_3_cond_2_2;
  reg _tmp_674;
  reg _ram_w4_l8192_id6_4_cond_1_1;
  reg _ram_w4_l8192_id6_4_cond_2_1;
  reg _ram_w4_l8192_id6_4_cond_2_2;
  reg _tmp_675;
  reg _ram_w4_l8192_id6_5_cond_1_1;
  reg _ram_w4_l8192_id6_5_cond_2_1;
  reg _ram_w4_l8192_id6_5_cond_2_2;
  reg _tmp_676;
  reg _ram_w4_l8192_id6_6_cond_1_1;
  reg _ram_w4_l8192_id6_6_cond_2_1;
  reg _ram_w4_l8192_id6_6_cond_2_2;
  reg _tmp_677;
  reg _ram_w4_l8192_id6_7_cond_1_1;
  reg _ram_w4_l8192_id6_7_cond_2_1;
  reg _ram_w4_l8192_id6_7_cond_2_2;
  wire signed [4-1:0] _tmp_678;
  wire _tmp_679;
  assign _tmp_678 = (__tmp_669_2 == 0)? ram_w4_l8192_id6_0_0_rdata : 
                    (__tmp_669_2 == 1)? ram_w4_l8192_id6_1_0_rdata : 
                    (__tmp_669_2 == 2)? ram_w4_l8192_id6_2_0_rdata : 
                    (__tmp_669_2 == 3)? ram_w4_l8192_id6_3_0_rdata : 
                    (__tmp_669_2 == 4)? ram_w4_l8192_id6_4_0_rdata : 
                    (__tmp_669_2 == 5)? ram_w4_l8192_id6_5_0_rdata : 
                    (__tmp_669_2 == 6)? ram_w4_l8192_id6_6_0_rdata : 
                    (__tmp_669_2 == 7)? ram_w4_l8192_id6_7_0_rdata : 0;
  assign _tmp_679 = _tmp_670;
  assign _stream_conv2d_16_source_34_source_ram_rdata = (_stream_conv2d_16_source_34_source_ram_sel == 18)? _tmp_678 : 0;
  localparam _tmp_680 = 1;
  wire [_tmp_680-1:0] _tmp_681;
  assign _tmp_681 = _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
  reg [_tmp_680-1:0] __tmp_681_1;
  reg [4-1:0] __variable_wdata_508;
  assign stream_conv2d_16_source_34_data = __variable_wdata_508;
  reg [32-1:0] _stream_conv2d_16_source_34_source_pat_fsm_17;
  localparam _stream_conv2d_16_source_34_source_pat_fsm_17_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_34_source_pat_all_offset;
  assign _stream_conv2d_16_source_34_source_pat_all_offset = _stream_conv2d_16_source_34_source_offset_buf + _source_stream_conv2d_16_source_34_pat_cur_offset_0 + _source_stream_conv2d_16_source_34_pat_cur_offset_1 + _source_stream_conv2d_16_source_34_pat_cur_offset_2 + _source_stream_conv2d_16_source_34_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_35_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_35_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_35_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_35_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_35_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_35_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_35_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_35_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_35_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_35_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_35_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_35_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_35_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_35_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_35_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_35_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_35_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_35_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_35_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_35_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_35_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_35_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_35_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_35_pat_stride_buf_3;
  reg _set_flag_682;
  wire [3-1:0] _tmp_683;
  assign _tmp_683 = _stream_conv2d_16_source_35_source_ram_raddr;
  reg [3-1:0] __tmp_683_1;
  reg [3-1:0] __tmp_683_2;
  reg _tmp_684;
  reg _ram_w4_l8192_id7_0_cond_1_1;
  reg _ram_w4_l8192_id7_0_cond_2_1;
  reg _ram_w4_l8192_id7_0_cond_2_2;
  reg _tmp_685;
  reg _ram_w4_l8192_id7_1_cond_1_1;
  reg _ram_w4_l8192_id7_1_cond_2_1;
  reg _ram_w4_l8192_id7_1_cond_2_2;
  reg _tmp_686;
  reg _ram_w4_l8192_id7_2_cond_1_1;
  reg _ram_w4_l8192_id7_2_cond_2_1;
  reg _ram_w4_l8192_id7_2_cond_2_2;
  reg _tmp_687;
  reg _ram_w4_l8192_id7_3_cond_1_1;
  reg _ram_w4_l8192_id7_3_cond_2_1;
  reg _ram_w4_l8192_id7_3_cond_2_2;
  reg _tmp_688;
  reg _ram_w4_l8192_id7_4_cond_1_1;
  reg _ram_w4_l8192_id7_4_cond_2_1;
  reg _ram_w4_l8192_id7_4_cond_2_2;
  reg _tmp_689;
  reg _ram_w4_l8192_id7_5_cond_1_1;
  reg _ram_w4_l8192_id7_5_cond_2_1;
  reg _ram_w4_l8192_id7_5_cond_2_2;
  reg _tmp_690;
  reg _ram_w4_l8192_id7_6_cond_1_1;
  reg _ram_w4_l8192_id7_6_cond_2_1;
  reg _ram_w4_l8192_id7_6_cond_2_2;
  reg _tmp_691;
  reg _ram_w4_l8192_id7_7_cond_1_1;
  reg _ram_w4_l8192_id7_7_cond_2_1;
  reg _ram_w4_l8192_id7_7_cond_2_2;
  wire signed [4-1:0] _tmp_692;
  wire _tmp_693;
  assign _tmp_692 = (__tmp_683_2 == 0)? ram_w4_l8192_id7_0_0_rdata : 
                    (__tmp_683_2 == 1)? ram_w4_l8192_id7_1_0_rdata : 
                    (__tmp_683_2 == 2)? ram_w4_l8192_id7_2_0_rdata : 
                    (__tmp_683_2 == 3)? ram_w4_l8192_id7_3_0_rdata : 
                    (__tmp_683_2 == 4)? ram_w4_l8192_id7_4_0_rdata : 
                    (__tmp_683_2 == 5)? ram_w4_l8192_id7_5_0_rdata : 
                    (__tmp_683_2 == 6)? ram_w4_l8192_id7_6_0_rdata : 
                    (__tmp_683_2 == 7)? ram_w4_l8192_id7_7_0_rdata : 0;
  assign _tmp_693 = _tmp_684;
  assign _stream_conv2d_16_source_35_source_ram_rdata = (_stream_conv2d_16_source_35_source_ram_sel == 19)? _tmp_692 : 0;
  localparam _tmp_694 = 1;
  wire [_tmp_694-1:0] _tmp_695;
  assign _tmp_695 = _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
  reg [_tmp_694-1:0] __tmp_695_1;
  reg [4-1:0] __variable_wdata_509;
  assign stream_conv2d_16_source_35_data = __variable_wdata_509;
  reg [32-1:0] _stream_conv2d_16_source_35_source_pat_fsm_18;
  localparam _stream_conv2d_16_source_35_source_pat_fsm_18_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_35_source_pat_all_offset;
  assign _stream_conv2d_16_source_35_source_pat_all_offset = _stream_conv2d_16_source_35_source_offset_buf + _source_stream_conv2d_16_source_35_pat_cur_offset_0 + _source_stream_conv2d_16_source_35_pat_cur_offset_1 + _source_stream_conv2d_16_source_35_pat_cur_offset_2 + _source_stream_conv2d_16_source_35_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_16_source_36_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_16_source_36_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_16_source_36_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_16_source_36_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_16_source_36_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_16_source_36_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_16_source_36_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_16_source_36_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_16_source_36_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_16_source_36_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_16_source_36_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_16_source_36_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_16_source_36_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_16_source_36_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_16_source_36_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_16_source_36_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_16_source_36_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_16_source_36_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_16_source_36_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_16_source_36_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_16_source_36_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_16_source_36_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_16_source_36_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_16_source_36_pat_stride_buf_3;
  reg _set_flag_696;
  wire [3-1:0] _tmp_697;
  assign _tmp_697 = _stream_conv2d_16_source_36_source_ram_raddr;
  reg [3-1:0] __tmp_697_1;
  reg [3-1:0] __tmp_697_2;
  reg _tmp_698;
  reg _ram_w4_l8192_id8_0_cond_1_1;
  reg _ram_w4_l8192_id8_0_cond_2_1;
  reg _ram_w4_l8192_id8_0_cond_2_2;
  reg _tmp_699;
  reg _ram_w4_l8192_id8_1_cond_1_1;
  reg _ram_w4_l8192_id8_1_cond_2_1;
  reg _ram_w4_l8192_id8_1_cond_2_2;
  reg _tmp_700;
  reg _ram_w4_l8192_id8_2_cond_1_1;
  reg _ram_w4_l8192_id8_2_cond_2_1;
  reg _ram_w4_l8192_id8_2_cond_2_2;
  reg _tmp_701;
  reg _ram_w4_l8192_id8_3_cond_1_1;
  reg _ram_w4_l8192_id8_3_cond_2_1;
  reg _ram_w4_l8192_id8_3_cond_2_2;
  reg _tmp_702;
  reg _ram_w4_l8192_id8_4_cond_1_1;
  reg _ram_w4_l8192_id8_4_cond_2_1;
  reg _ram_w4_l8192_id8_4_cond_2_2;
  reg _tmp_703;
  reg _ram_w4_l8192_id8_5_cond_1_1;
  reg _ram_w4_l8192_id8_5_cond_2_1;
  reg _ram_w4_l8192_id8_5_cond_2_2;
  reg _tmp_704;
  reg _ram_w4_l8192_id8_6_cond_1_1;
  reg _ram_w4_l8192_id8_6_cond_2_1;
  reg _ram_w4_l8192_id8_6_cond_2_2;
  reg _tmp_705;
  reg _ram_w4_l8192_id8_7_cond_1_1;
  reg _ram_w4_l8192_id8_7_cond_2_1;
  reg _ram_w4_l8192_id8_7_cond_2_2;
  wire signed [4-1:0] _tmp_706;
  wire _tmp_707;
  assign _tmp_706 = (__tmp_697_2 == 0)? ram_w4_l8192_id8_0_0_rdata : 
                    (__tmp_697_2 == 1)? ram_w4_l8192_id8_1_0_rdata : 
                    (__tmp_697_2 == 2)? ram_w4_l8192_id8_2_0_rdata : 
                    (__tmp_697_2 == 3)? ram_w4_l8192_id8_3_0_rdata : 
                    (__tmp_697_2 == 4)? ram_w4_l8192_id8_4_0_rdata : 
                    (__tmp_697_2 == 5)? ram_w4_l8192_id8_5_0_rdata : 
                    (__tmp_697_2 == 6)? ram_w4_l8192_id8_6_0_rdata : 
                    (__tmp_697_2 == 7)? ram_w4_l8192_id8_7_0_rdata : 0;
  assign _tmp_707 = _tmp_698;
  assign _stream_conv2d_16_source_36_source_ram_rdata = (_stream_conv2d_16_source_36_source_ram_sel == 20)? _tmp_706 : 0;
  localparam _tmp_708 = 1;
  wire [_tmp_708-1:0] _tmp_709;
  assign _tmp_709 = _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
  reg [_tmp_708-1:0] __tmp_709_1;
  reg [4-1:0] __variable_wdata_510;
  assign stream_conv2d_16_source_36_data = __variable_wdata_510;
  reg [32-1:0] _stream_conv2d_16_source_36_source_pat_fsm_19;
  localparam _stream_conv2d_16_source_36_source_pat_fsm_19_init = 0;
  wire [32-1:0] _stream_conv2d_16_source_36_source_pat_all_offset;
  assign _stream_conv2d_16_source_36_source_pat_all_offset = _stream_conv2d_16_source_36_source_offset_buf + _source_stream_conv2d_16_source_36_pat_cur_offset_0 + _source_stream_conv2d_16_source_36_pat_cur_offset_1 + _source_stream_conv2d_16_source_36_pat_cur_offset_2 + _source_stream_conv2d_16_source_36_pat_cur_offset_3;
  reg _set_flag_710;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_1;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_2;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_3;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_4;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_5;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_6;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_7;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_8;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_9;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_10;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_11;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_12;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_13;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_14;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_15;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_16;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_17;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_18;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_19;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_20;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_21;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_22;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_23;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_24;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_25;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_26;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_27;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_28;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_29;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_30;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_31;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_32;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_33;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_34;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_35;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_36;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_37;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_38;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_39;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_40;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_41;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_42;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_43;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_44;
  reg [32-1:0] __stream_conv2d_16_sink_37_sink_offset_0_45;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_1;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_2;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_3;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_4;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_5;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_6;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_7;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_8;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_9;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_10;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_11;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_12;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_13;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_14;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_15;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_16;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_17;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_18;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_19;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_20;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_21;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_22;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_23;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_24;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_25;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_26;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_27;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_28;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_29;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_30;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_31;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_32;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_33;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_34;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_35;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_36;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_37;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_38;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_39;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_40;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_41;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_42;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_43;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_44;
  reg [33-1:0] __stream_conv2d_16_sink_37_sink_size_1_45;
  reg __stream_seq_14_cond_2_1;
  reg __stream_seq_14_cond_2_2;
  reg __stream_seq_14_cond_2_3;
  reg __stream_seq_14_cond_2_4;
  reg __stream_seq_14_cond_2_5;
  reg __stream_seq_14_cond_2_6;
  reg __stream_seq_14_cond_2_7;
  reg __stream_seq_14_cond_2_8;
  reg __stream_seq_14_cond_2_9;
  reg __stream_seq_14_cond_2_10;
  reg __stream_seq_14_cond_2_11;
  reg __stream_seq_14_cond_2_12;
  reg __stream_seq_14_cond_2_13;
  reg __stream_seq_14_cond_2_14;
  reg __stream_seq_14_cond_2_15;
  reg __stream_seq_14_cond_2_16;
  reg __stream_seq_14_cond_2_17;
  reg __stream_seq_14_cond_2_18;
  reg __stream_seq_14_cond_2_19;
  reg __stream_seq_14_cond_2_20;
  reg __stream_seq_14_cond_2_21;
  reg __stream_seq_14_cond_2_22;
  reg __stream_seq_14_cond_2_23;
  reg __stream_seq_14_cond_2_24;
  reg __stream_seq_14_cond_2_25;
  reg __stream_seq_14_cond_2_26;
  reg __stream_seq_14_cond_2_27;
  reg __stream_seq_14_cond_2_28;
  reg __stream_seq_14_cond_2_29;
  reg __stream_seq_14_cond_2_30;
  reg __stream_seq_14_cond_2_31;
  reg __stream_seq_14_cond_2_32;
  reg __stream_seq_14_cond_2_33;
  reg __stream_seq_14_cond_2_34;
  reg __stream_seq_14_cond_2_35;
  reg __stream_seq_14_cond_2_36;
  reg __stream_seq_14_cond_2_37;
  reg __stream_seq_14_cond_2_38;
  reg __stream_seq_14_cond_2_39;
  reg __stream_seq_14_cond_2_40;
  reg __stream_seq_14_cond_2_41;
  reg __stream_seq_14_cond_2_42;
  reg __stream_seq_14_cond_2_43;
  reg __stream_seq_14_cond_2_44;
  reg __stream_seq_14_cond_2_45;
  reg __set_flag_710_1;
  reg __set_flag_710_2;
  reg __set_flag_710_3;
  reg __set_flag_710_4;
  reg __set_flag_710_5;
  reg __set_flag_710_6;
  reg __set_flag_710_7;
  reg __set_flag_710_8;
  reg __set_flag_710_9;
  reg __set_flag_710_10;
  reg __set_flag_710_11;
  reg __set_flag_710_12;
  reg __set_flag_710_13;
  reg __set_flag_710_14;
  reg __set_flag_710_15;
  reg __set_flag_710_16;
  reg __set_flag_710_17;
  reg __set_flag_710_18;
  reg __set_flag_710_19;
  reg __set_flag_710_20;
  reg __set_flag_710_21;
  reg __set_flag_710_22;
  reg __set_flag_710_23;
  reg __set_flag_710_24;
  reg __set_flag_710_25;
  reg __set_flag_710_26;
  reg __set_flag_710_27;
  reg __set_flag_710_28;
  reg __set_flag_710_29;
  reg __set_flag_710_30;
  reg __set_flag_710_31;
  reg __set_flag_710_32;
  reg __set_flag_710_33;
  reg __set_flag_710_34;
  reg __set_flag_710_35;
  reg __set_flag_710_36;
  reg __set_flag_710_37;
  reg __set_flag_710_38;
  reg __set_flag_710_39;
  reg __set_flag_710_40;
  reg __set_flag_710_41;
  reg __set_flag_710_42;
  reg __set_flag_710_43;
  reg __set_flag_710_44;
  reg __set_flag_710_45;
  wire [2-1:0] _tmp_711;
  assign _tmp_711 = _stream_conv2d_16_sink_37_sink_waddr;
  reg _ram_w8_l2048_id11_0_cond_0_1;
  reg _ram_w8_l2048_id11_1_cond_0_1;
  reg _ram_w8_l2048_id11_2_cond_0_1;
  reg _ram_w8_l2048_id11_3_cond_0_1;
  reg __stream_conv2d_16_start_1;
  reg __stream_conv2d_16_start_2;
  reg __stream_conv2d_16_start_3;
  reg __stream_conv2d_16_start_4;
  reg __stream_conv2d_16_start_5;
  reg __stream_conv2d_16_start_6;
  reg __stream_conv2d_16_start_7;
  reg __stream_conv2d_16_start_8;
  reg __stream_conv2d_16_start_9;
  reg __stream_conv2d_16_start_10;
  reg __stream_conv2d_16_start_11;
  reg __stream_conv2d_16_start_12;
  reg __stream_conv2d_16_start_13;
  reg __stream_conv2d_16_start_14;
  reg __stream_conv2d_16_start_15;
  reg __stream_conv2d_16_start_16;
  reg __stream_conv2d_16_start_17;
  reg __stream_conv2d_16_start_18;
  reg __stream_conv2d_16_start_19;
  reg __stream_conv2d_16_start_20;
  reg __stream_conv2d_16_start_21;
  reg __stream_conv2d_16_start_22;
  reg __stream_conv2d_16_start_23;
  reg __stream_conv2d_16_start_24;
  reg __stream_conv2d_16_start_25;
  reg __stream_conv2d_16_start_26;
  reg __stream_conv2d_16_start_27;
  reg __stream_conv2d_16_start_28;
  reg __stream_conv2d_16_start_29;
  reg __stream_conv2d_16_start_30;
  reg __stream_conv2d_16_start_31;
  reg __stream_conv2d_16_start_32;
  reg __stream_conv2d_16_start_33;
  reg __stream_conv2d_16_start_34;
  reg __stream_conv2d_16_start_35;
  reg __stream_conv2d_16_start_36;
  reg __stream_conv2d_16_start_37;
  reg __stream_conv2d_16_start_38;
  reg __stream_conv2d_16_start_39;
  reg __stream_conv2d_16_start_40;
  reg __stream_conv2d_16_start_41;
  reg __stream_conv2d_16_start_42;
  reg __stream_conv2d_16_start_43;
  reg __stream_conv2d_16_start_44;
  reg __stream_conv2d_16_start_45;
  reg __stream_conv2d_16_start_46;
  reg [32-1:0] _stream_conv2d_16_sink_37_sink_fsm_20;
  localparam _stream_conv2d_16_sink_37_sink_fsm_20_init = 0;
  assign _stream_conv2d_16_start_flag = ((conv2d_16_comp_fsm == 4) && !_stream_conv2d_16_source_busy)? 1 : 0;
  localparam _tmp_712 = 1;
  wire [_tmp_712-1:0] _tmp_713;
  assign _tmp_713 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_712-1:0] __tmp_713_1;
  reg [_tmp_712-1:0] __tmp_713_2;
  reg [_tmp_712-1:0] __tmp_713_3;
  reg [_tmp_712-1:0] __tmp_713_4;
  reg [_tmp_712-1:0] __tmp_713_5;
  localparam _tmp_714 = 1;
  wire [_tmp_714-1:0] _tmp_715;
  assign _tmp_715 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_714-1:0] __tmp_715_1;
  reg [_tmp_714-1:0] __tmp_715_2;
  reg [_tmp_714-1:0] __tmp_715_3;
  reg [_tmp_714-1:0] __tmp_715_4;
  reg [_tmp_714-1:0] __tmp_715_5;
  reg [_tmp_714-1:0] __tmp_715_6;
  reg [_tmp_714-1:0] __tmp_715_7;
  reg [_tmp_714-1:0] __tmp_715_8;
  reg [_tmp_714-1:0] __tmp_715_9;
  reg [_tmp_714-1:0] __tmp_715_10;
  reg [_tmp_714-1:0] __tmp_715_11;
  reg [_tmp_714-1:0] __tmp_715_12;
  localparam _tmp_716 = 1;
  wire [_tmp_716-1:0] _tmp_717;
  assign _tmp_717 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_716-1:0] __tmp_717_1;
  reg [_tmp_716-1:0] __tmp_717_2;
  reg [_tmp_716-1:0] __tmp_717_3;
  reg [_tmp_716-1:0] __tmp_717_4;
  reg [_tmp_716-1:0] __tmp_717_5;
  reg [_tmp_716-1:0] __tmp_717_6;
  reg [_tmp_716-1:0] __tmp_717_7;
  reg [_tmp_716-1:0] __tmp_717_8;
  reg [_tmp_716-1:0] __tmp_717_9;
  reg [_tmp_716-1:0] __tmp_717_10;
  reg [_tmp_716-1:0] __tmp_717_11;
  reg [_tmp_716-1:0] __tmp_717_12;
  localparam _tmp_718 = 1;
  wire [_tmp_718-1:0] _tmp_719;
  assign _tmp_719 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_718-1:0] __tmp_719_1;
  reg [_tmp_718-1:0] __tmp_719_2;
  reg [_tmp_718-1:0] __tmp_719_3;
  reg [_tmp_718-1:0] __tmp_719_4;
  reg [_tmp_718-1:0] __tmp_719_5;
  reg [_tmp_718-1:0] __tmp_719_6;
  reg [_tmp_718-1:0] __tmp_719_7;
  reg [_tmp_718-1:0] __tmp_719_8;
  reg [_tmp_718-1:0] __tmp_719_9;
  reg [_tmp_718-1:0] __tmp_719_10;
  reg [_tmp_718-1:0] __tmp_719_11;
  reg [_tmp_718-1:0] __tmp_719_12;
  localparam _tmp_720 = 1;
  wire [_tmp_720-1:0] _tmp_721;
  assign _tmp_721 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_720-1:0] __tmp_721_1;
  reg [_tmp_720-1:0] __tmp_721_2;
  reg [_tmp_720-1:0] __tmp_721_3;
  reg [_tmp_720-1:0] __tmp_721_4;
  reg [_tmp_720-1:0] __tmp_721_5;
  reg [_tmp_720-1:0] __tmp_721_6;
  reg [_tmp_720-1:0] __tmp_721_7;
  reg [_tmp_720-1:0] __tmp_721_8;
  reg [_tmp_720-1:0] __tmp_721_9;
  reg [_tmp_720-1:0] __tmp_721_10;
  reg [_tmp_720-1:0] __tmp_721_11;
  reg [_tmp_720-1:0] __tmp_721_12;
  localparam _tmp_722 = 1;
  wire [_tmp_722-1:0] _tmp_723;
  assign _tmp_723 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_722-1:0] __tmp_723_1;
  reg [_tmp_722-1:0] __tmp_723_2;
  reg [_tmp_722-1:0] __tmp_723_3;
  reg [_tmp_722-1:0] __tmp_723_4;
  reg [_tmp_722-1:0] __tmp_723_5;
  reg [_tmp_722-1:0] __tmp_723_6;
  reg [_tmp_722-1:0] __tmp_723_7;
  reg [_tmp_722-1:0] __tmp_723_8;
  reg [_tmp_722-1:0] __tmp_723_9;
  reg [_tmp_722-1:0] __tmp_723_10;
  reg [_tmp_722-1:0] __tmp_723_11;
  reg [_tmp_722-1:0] __tmp_723_12;
  localparam _tmp_724 = 1;
  wire [_tmp_724-1:0] _tmp_725;
  assign _tmp_725 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_724-1:0] __tmp_725_1;
  reg [_tmp_724-1:0] __tmp_725_2;
  reg [_tmp_724-1:0] __tmp_725_3;
  reg [_tmp_724-1:0] __tmp_725_4;
  reg [_tmp_724-1:0] __tmp_725_5;
  reg [_tmp_724-1:0] __tmp_725_6;
  reg [_tmp_724-1:0] __tmp_725_7;
  reg [_tmp_724-1:0] __tmp_725_8;
  reg [_tmp_724-1:0] __tmp_725_9;
  reg [_tmp_724-1:0] __tmp_725_10;
  reg [_tmp_724-1:0] __tmp_725_11;
  reg [_tmp_724-1:0] __tmp_725_12;
  localparam _tmp_726 = 1;
  wire [_tmp_726-1:0] _tmp_727;
  assign _tmp_727 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_726-1:0] __tmp_727_1;
  reg [_tmp_726-1:0] __tmp_727_2;
  reg [_tmp_726-1:0] __tmp_727_3;
  reg [_tmp_726-1:0] __tmp_727_4;
  reg [_tmp_726-1:0] __tmp_727_5;
  reg [_tmp_726-1:0] __tmp_727_6;
  reg [_tmp_726-1:0] __tmp_727_7;
  reg [_tmp_726-1:0] __tmp_727_8;
  reg [_tmp_726-1:0] __tmp_727_9;
  reg [_tmp_726-1:0] __tmp_727_10;
  reg [_tmp_726-1:0] __tmp_727_11;
  reg [_tmp_726-1:0] __tmp_727_12;
  localparam _tmp_728 = 1;
  wire [_tmp_728-1:0] _tmp_729;
  assign _tmp_729 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_728-1:0] __tmp_729_1;
  reg [_tmp_728-1:0] __tmp_729_2;
  reg [_tmp_728-1:0] __tmp_729_3;
  reg [_tmp_728-1:0] __tmp_729_4;
  reg [_tmp_728-1:0] __tmp_729_5;
  reg [_tmp_728-1:0] __tmp_729_6;
  reg [_tmp_728-1:0] __tmp_729_7;
  reg [_tmp_728-1:0] __tmp_729_8;
  reg [_tmp_728-1:0] __tmp_729_9;
  reg [_tmp_728-1:0] __tmp_729_10;
  reg [_tmp_728-1:0] __tmp_729_11;
  reg [_tmp_728-1:0] __tmp_729_12;
  localparam _tmp_730 = 1;
  wire [_tmp_730-1:0] _tmp_731;
  assign _tmp_731 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_730-1:0] __tmp_731_1;
  reg [_tmp_730-1:0] __tmp_731_2;
  reg [_tmp_730-1:0] __tmp_731_3;
  reg [_tmp_730-1:0] __tmp_731_4;
  reg [_tmp_730-1:0] __tmp_731_5;
  reg [_tmp_730-1:0] __tmp_731_6;
  reg [_tmp_730-1:0] __tmp_731_7;
  reg [_tmp_730-1:0] __tmp_731_8;
  reg [_tmp_730-1:0] __tmp_731_9;
  reg [_tmp_730-1:0] __tmp_731_10;
  reg [_tmp_730-1:0] __tmp_731_11;
  reg [_tmp_730-1:0] __tmp_731_12;
  localparam _tmp_732 = 1;
  wire [_tmp_732-1:0] _tmp_733;
  assign _tmp_733 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_732-1:0] __tmp_733_1;
  reg [_tmp_732-1:0] __tmp_733_2;
  reg [_tmp_732-1:0] __tmp_733_3;
  reg [_tmp_732-1:0] __tmp_733_4;
  reg [_tmp_732-1:0] __tmp_733_5;
  reg [_tmp_732-1:0] __tmp_733_6;
  reg [_tmp_732-1:0] __tmp_733_7;
  reg [_tmp_732-1:0] __tmp_733_8;
  reg [_tmp_732-1:0] __tmp_733_9;
  reg [_tmp_732-1:0] __tmp_733_10;
  reg [_tmp_732-1:0] __tmp_733_11;
  reg [_tmp_732-1:0] __tmp_733_12;
  localparam _tmp_734 = 1;
  wire [_tmp_734-1:0] _tmp_735;
  assign _tmp_735 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_734-1:0] __tmp_735_1;
  reg [_tmp_734-1:0] __tmp_735_2;
  reg [_tmp_734-1:0] __tmp_735_3;
  reg [_tmp_734-1:0] __tmp_735_4;
  reg [_tmp_734-1:0] __tmp_735_5;
  reg [_tmp_734-1:0] __tmp_735_6;
  reg [_tmp_734-1:0] __tmp_735_7;
  reg [_tmp_734-1:0] __tmp_735_8;
  reg [_tmp_734-1:0] __tmp_735_9;
  reg [_tmp_734-1:0] __tmp_735_10;
  reg [_tmp_734-1:0] __tmp_735_11;
  reg [_tmp_734-1:0] __tmp_735_12;
  localparam _tmp_736 = 1;
  wire [_tmp_736-1:0] _tmp_737;
  assign _tmp_737 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_736-1:0] __tmp_737_1;
  reg [_tmp_736-1:0] __tmp_737_2;
  reg [_tmp_736-1:0] __tmp_737_3;
  reg [_tmp_736-1:0] __tmp_737_4;
  reg [_tmp_736-1:0] __tmp_737_5;
  reg [_tmp_736-1:0] __tmp_737_6;
  reg [_tmp_736-1:0] __tmp_737_7;
  reg [_tmp_736-1:0] __tmp_737_8;
  reg [_tmp_736-1:0] __tmp_737_9;
  reg [_tmp_736-1:0] __tmp_737_10;
  reg [_tmp_736-1:0] __tmp_737_11;
  reg [_tmp_736-1:0] __tmp_737_12;
  localparam _tmp_738 = 1;
  wire [_tmp_738-1:0] _tmp_739;
  assign _tmp_739 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_738-1:0] __tmp_739_1;
  reg [_tmp_738-1:0] __tmp_739_2;
  reg [_tmp_738-1:0] __tmp_739_3;
  reg [_tmp_738-1:0] __tmp_739_4;
  reg [_tmp_738-1:0] __tmp_739_5;
  reg [_tmp_738-1:0] __tmp_739_6;
  reg [_tmp_738-1:0] __tmp_739_7;
  reg [_tmp_738-1:0] __tmp_739_8;
  reg [_tmp_738-1:0] __tmp_739_9;
  reg [_tmp_738-1:0] __tmp_739_10;
  reg [_tmp_738-1:0] __tmp_739_11;
  reg [_tmp_738-1:0] __tmp_739_12;
  localparam _tmp_740 = 1;
  wire [_tmp_740-1:0] _tmp_741;
  assign _tmp_741 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_740-1:0] __tmp_741_1;
  reg [_tmp_740-1:0] __tmp_741_2;
  reg [_tmp_740-1:0] __tmp_741_3;
  reg [_tmp_740-1:0] __tmp_741_4;
  reg [_tmp_740-1:0] __tmp_741_5;
  reg [_tmp_740-1:0] __tmp_741_6;
  reg [_tmp_740-1:0] __tmp_741_7;
  reg [_tmp_740-1:0] __tmp_741_8;
  reg [_tmp_740-1:0] __tmp_741_9;
  reg [_tmp_740-1:0] __tmp_741_10;
  reg [_tmp_740-1:0] __tmp_741_11;
  reg [_tmp_740-1:0] __tmp_741_12;
  localparam _tmp_742 = 1;
  wire [_tmp_742-1:0] _tmp_743;
  assign _tmp_743 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_742-1:0] __tmp_743_1;
  reg [_tmp_742-1:0] __tmp_743_2;
  reg [_tmp_742-1:0] __tmp_743_3;
  reg [_tmp_742-1:0] __tmp_743_4;
  reg [_tmp_742-1:0] __tmp_743_5;
  reg [_tmp_742-1:0] __tmp_743_6;
  reg [_tmp_742-1:0] __tmp_743_7;
  reg [_tmp_742-1:0] __tmp_743_8;
  reg [_tmp_742-1:0] __tmp_743_9;
  reg [_tmp_742-1:0] __tmp_743_10;
  reg [_tmp_742-1:0] __tmp_743_11;
  reg [_tmp_742-1:0] __tmp_743_12;
  localparam _tmp_744 = 1;
  wire [_tmp_744-1:0] _tmp_745;
  assign _tmp_745 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_744-1:0] __tmp_745_1;
  reg [_tmp_744-1:0] __tmp_745_2;
  reg [_tmp_744-1:0] __tmp_745_3;
  reg [_tmp_744-1:0] __tmp_745_4;
  reg [_tmp_744-1:0] __tmp_745_5;
  reg [_tmp_744-1:0] __tmp_745_6;
  reg [_tmp_744-1:0] __tmp_745_7;
  reg [_tmp_744-1:0] __tmp_745_8;
  reg [_tmp_744-1:0] __tmp_745_9;
  reg [_tmp_744-1:0] __tmp_745_10;
  reg [_tmp_744-1:0] __tmp_745_11;
  reg [_tmp_744-1:0] __tmp_745_12;
  localparam _tmp_746 = 1;
  wire [_tmp_746-1:0] _tmp_747;
  assign _tmp_747 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_746-1:0] __tmp_747_1;
  reg [_tmp_746-1:0] __tmp_747_2;
  reg [_tmp_746-1:0] __tmp_747_3;
  reg [_tmp_746-1:0] __tmp_747_4;
  reg [_tmp_746-1:0] __tmp_747_5;
  reg [_tmp_746-1:0] __tmp_747_6;
  reg [_tmp_746-1:0] __tmp_747_7;
  reg [_tmp_746-1:0] __tmp_747_8;
  reg [_tmp_746-1:0] __tmp_747_9;
  reg [_tmp_746-1:0] __tmp_747_10;
  reg [_tmp_746-1:0] __tmp_747_11;
  reg [_tmp_746-1:0] __tmp_747_12;
  localparam _tmp_748 = 1;
  wire [_tmp_748-1:0] _tmp_749;
  assign _tmp_749 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_748-1:0] __tmp_749_1;
  reg [_tmp_748-1:0] __tmp_749_2;
  reg [_tmp_748-1:0] __tmp_749_3;
  reg [_tmp_748-1:0] __tmp_749_4;
  reg [_tmp_748-1:0] __tmp_749_5;
  reg [_tmp_748-1:0] __tmp_749_6;
  reg [_tmp_748-1:0] __tmp_749_7;
  reg [_tmp_748-1:0] __tmp_749_8;
  reg [_tmp_748-1:0] __tmp_749_9;
  reg [_tmp_748-1:0] __tmp_749_10;
  reg [_tmp_748-1:0] __tmp_749_11;
  reg [_tmp_748-1:0] __tmp_749_12;
  localparam _tmp_750 = 1;
  wire [_tmp_750-1:0] _tmp_751;
  assign _tmp_751 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_750-1:0] __tmp_751_1;
  reg [_tmp_750-1:0] __tmp_751_2;
  reg [_tmp_750-1:0] __tmp_751_3;
  reg [_tmp_750-1:0] __tmp_751_4;
  reg [_tmp_750-1:0] __tmp_751_5;
  reg [_tmp_750-1:0] __tmp_751_6;
  reg [_tmp_750-1:0] __tmp_751_7;
  reg [_tmp_750-1:0] __tmp_751_8;
  reg [_tmp_750-1:0] __tmp_751_9;
  reg [_tmp_750-1:0] __tmp_751_10;
  reg [_tmp_750-1:0] __tmp_751_11;
  reg [_tmp_750-1:0] __tmp_751_12;
  localparam _tmp_752 = 1;
  wire [_tmp_752-1:0] _tmp_753;
  assign _tmp_753 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_752-1:0] __tmp_753_1;
  reg [_tmp_752-1:0] __tmp_753_2;
  reg [_tmp_752-1:0] __tmp_753_3;
  reg [_tmp_752-1:0] __tmp_753_4;
  reg [_tmp_752-1:0] __tmp_753_5;
  reg [_tmp_752-1:0] __tmp_753_6;
  reg [_tmp_752-1:0] __tmp_753_7;
  reg [_tmp_752-1:0] __tmp_753_8;
  reg [_tmp_752-1:0] __tmp_753_9;
  reg [_tmp_752-1:0] __tmp_753_10;
  reg [_tmp_752-1:0] __tmp_753_11;
  reg [_tmp_752-1:0] __tmp_753_12;
  localparam _tmp_754 = 1;
  wire [_tmp_754-1:0] _tmp_755;
  assign _tmp_755 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_754-1:0] __tmp_755_1;
  reg [_tmp_754-1:0] __tmp_755_2;
  reg [_tmp_754-1:0] __tmp_755_3;
  reg [_tmp_754-1:0] __tmp_755_4;
  reg [_tmp_754-1:0] __tmp_755_5;
  reg [_tmp_754-1:0] __tmp_755_6;
  reg [_tmp_754-1:0] __tmp_755_7;
  reg [_tmp_754-1:0] __tmp_755_8;
  reg [_tmp_754-1:0] __tmp_755_9;
  reg [_tmp_754-1:0] __tmp_755_10;
  reg [_tmp_754-1:0] __tmp_755_11;
  reg [_tmp_754-1:0] __tmp_755_12;
  localparam _tmp_756 = 1;
  wire [_tmp_756-1:0] _tmp_757;
  assign _tmp_757 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_756-1:0] __tmp_757_1;
  reg [_tmp_756-1:0] __tmp_757_2;
  reg [_tmp_756-1:0] __tmp_757_3;
  reg [_tmp_756-1:0] __tmp_757_4;
  reg [_tmp_756-1:0] __tmp_757_5;
  reg [_tmp_756-1:0] __tmp_757_6;
  reg [_tmp_756-1:0] __tmp_757_7;
  reg [_tmp_756-1:0] __tmp_757_8;
  reg [_tmp_756-1:0] __tmp_757_9;
  reg [_tmp_756-1:0] __tmp_757_10;
  reg [_tmp_756-1:0] __tmp_757_11;
  reg [_tmp_756-1:0] __tmp_757_12;
  localparam _tmp_758 = 1;
  wire [_tmp_758-1:0] _tmp_759;
  assign _tmp_759 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_758-1:0] __tmp_759_1;
  reg [_tmp_758-1:0] __tmp_759_2;
  reg [_tmp_758-1:0] __tmp_759_3;
  reg [_tmp_758-1:0] __tmp_759_4;
  reg [_tmp_758-1:0] __tmp_759_5;
  reg [_tmp_758-1:0] __tmp_759_6;
  reg [_tmp_758-1:0] __tmp_759_7;
  reg [_tmp_758-1:0] __tmp_759_8;
  reg [_tmp_758-1:0] __tmp_759_9;
  reg [_tmp_758-1:0] __tmp_759_10;
  reg [_tmp_758-1:0] __tmp_759_11;
  reg [_tmp_758-1:0] __tmp_759_12;
  localparam _tmp_760 = 1;
  wire [_tmp_760-1:0] _tmp_761;
  assign _tmp_761 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_760-1:0] __tmp_761_1;
  reg [_tmp_760-1:0] __tmp_761_2;
  reg [_tmp_760-1:0] __tmp_761_3;
  reg [_tmp_760-1:0] __tmp_761_4;
  reg [_tmp_760-1:0] __tmp_761_5;
  reg [_tmp_760-1:0] __tmp_761_6;
  reg [_tmp_760-1:0] __tmp_761_7;
  reg [_tmp_760-1:0] __tmp_761_8;
  reg [_tmp_760-1:0] __tmp_761_9;
  reg [_tmp_760-1:0] __tmp_761_10;
  reg [_tmp_760-1:0] __tmp_761_11;
  reg [_tmp_760-1:0] __tmp_761_12;
  localparam _tmp_762 = 1;
  wire [_tmp_762-1:0] _tmp_763;
  assign _tmp_763 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_762-1:0] __tmp_763_1;
  reg [_tmp_762-1:0] __tmp_763_2;
  reg [_tmp_762-1:0] __tmp_763_3;
  reg [_tmp_762-1:0] __tmp_763_4;
  reg [_tmp_762-1:0] __tmp_763_5;
  reg [_tmp_762-1:0] __tmp_763_6;
  reg [_tmp_762-1:0] __tmp_763_7;
  reg [_tmp_762-1:0] __tmp_763_8;
  reg [_tmp_762-1:0] __tmp_763_9;
  reg [_tmp_762-1:0] __tmp_763_10;
  reg [_tmp_762-1:0] __tmp_763_11;
  reg [_tmp_762-1:0] __tmp_763_12;
  localparam _tmp_764 = 1;
  wire [_tmp_764-1:0] _tmp_765;
  assign _tmp_765 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_764-1:0] __tmp_765_1;
  reg [_tmp_764-1:0] __tmp_765_2;
  reg [_tmp_764-1:0] __tmp_765_3;
  reg [_tmp_764-1:0] __tmp_765_4;
  reg [_tmp_764-1:0] __tmp_765_5;
  reg [_tmp_764-1:0] __tmp_765_6;
  reg [_tmp_764-1:0] __tmp_765_7;
  reg [_tmp_764-1:0] __tmp_765_8;
  reg [_tmp_764-1:0] __tmp_765_9;
  reg [_tmp_764-1:0] __tmp_765_10;
  reg [_tmp_764-1:0] __tmp_765_11;
  reg [_tmp_764-1:0] __tmp_765_12;
  localparam _tmp_766 = 1;
  wire [_tmp_766-1:0] _tmp_767;
  assign _tmp_767 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_766-1:0] __tmp_767_1;
  reg [_tmp_766-1:0] __tmp_767_2;
  reg [_tmp_766-1:0] __tmp_767_3;
  reg [_tmp_766-1:0] __tmp_767_4;
  reg [_tmp_766-1:0] __tmp_767_5;
  reg [_tmp_766-1:0] __tmp_767_6;
  reg [_tmp_766-1:0] __tmp_767_7;
  reg [_tmp_766-1:0] __tmp_767_8;
  reg [_tmp_766-1:0] __tmp_767_9;
  reg [_tmp_766-1:0] __tmp_767_10;
  reg [_tmp_766-1:0] __tmp_767_11;
  reg [_tmp_766-1:0] __tmp_767_12;
  localparam _tmp_768 = 1;
  wire [_tmp_768-1:0] _tmp_769;
  assign _tmp_769 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_768-1:0] __tmp_769_1;
  reg [_tmp_768-1:0] __tmp_769_2;
  reg [_tmp_768-1:0] __tmp_769_3;
  reg [_tmp_768-1:0] __tmp_769_4;
  reg [_tmp_768-1:0] __tmp_769_5;
  reg [_tmp_768-1:0] __tmp_769_6;
  reg [_tmp_768-1:0] __tmp_769_7;
  reg [_tmp_768-1:0] __tmp_769_8;
  reg [_tmp_768-1:0] __tmp_769_9;
  reg [_tmp_768-1:0] __tmp_769_10;
  reg [_tmp_768-1:0] __tmp_769_11;
  reg [_tmp_768-1:0] __tmp_769_12;
  reg [_tmp_768-1:0] __tmp_769_13;
  reg [_tmp_768-1:0] __tmp_769_14;
  reg [_tmp_768-1:0] __tmp_769_15;
  reg [_tmp_768-1:0] __tmp_769_16;
  reg [_tmp_768-1:0] __tmp_769_17;
  reg [_tmp_768-1:0] __tmp_769_18;
  reg [_tmp_768-1:0] __tmp_769_19;
  reg [_tmp_768-1:0] __tmp_769_20;
  reg [_tmp_768-1:0] __tmp_769_21;
  reg [_tmp_768-1:0] __tmp_769_22;
  localparam _tmp_770 = 1;
  wire [_tmp_770-1:0] _tmp_771;
  assign _tmp_771 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_770-1:0] __tmp_771_1;
  reg [_tmp_770-1:0] __tmp_771_2;
  reg [_tmp_770-1:0] __tmp_771_3;
  reg [_tmp_770-1:0] __tmp_771_4;
  reg [_tmp_770-1:0] __tmp_771_5;
  reg [_tmp_770-1:0] __tmp_771_6;
  reg [_tmp_770-1:0] __tmp_771_7;
  reg [_tmp_770-1:0] __tmp_771_8;
  reg [_tmp_770-1:0] __tmp_771_9;
  reg [_tmp_770-1:0] __tmp_771_10;
  reg [_tmp_770-1:0] __tmp_771_11;
  reg [_tmp_770-1:0] __tmp_771_12;
  reg [_tmp_770-1:0] __tmp_771_13;
  reg [_tmp_770-1:0] __tmp_771_14;
  reg [_tmp_770-1:0] __tmp_771_15;
  reg [_tmp_770-1:0] __tmp_771_16;
  reg [_tmp_770-1:0] __tmp_771_17;
  reg [_tmp_770-1:0] __tmp_771_18;
  reg [_tmp_770-1:0] __tmp_771_19;
  reg [_tmp_770-1:0] __tmp_771_20;
  reg [_tmp_770-1:0] __tmp_771_21;
  reg [_tmp_770-1:0] __tmp_771_22;
  localparam _tmp_772 = 1;
  wire [_tmp_772-1:0] _tmp_773;
  assign _tmp_773 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_772-1:0] __tmp_773_1;
  reg [_tmp_772-1:0] __tmp_773_2;
  reg [_tmp_772-1:0] __tmp_773_3;
  reg [_tmp_772-1:0] __tmp_773_4;
  reg [_tmp_772-1:0] __tmp_773_5;
  reg [_tmp_772-1:0] __tmp_773_6;
  reg [_tmp_772-1:0] __tmp_773_7;
  reg [_tmp_772-1:0] __tmp_773_8;
  reg [_tmp_772-1:0] __tmp_773_9;
  reg [_tmp_772-1:0] __tmp_773_10;
  reg [_tmp_772-1:0] __tmp_773_11;
  reg [_tmp_772-1:0] __tmp_773_12;
  reg [_tmp_772-1:0] __tmp_773_13;
  reg [_tmp_772-1:0] __tmp_773_14;
  reg [_tmp_772-1:0] __tmp_773_15;
  reg [_tmp_772-1:0] __tmp_773_16;
  reg [_tmp_772-1:0] __tmp_773_17;
  reg [_tmp_772-1:0] __tmp_773_18;
  reg [_tmp_772-1:0] __tmp_773_19;
  reg [_tmp_772-1:0] __tmp_773_20;
  reg [_tmp_772-1:0] __tmp_773_21;
  reg [_tmp_772-1:0] __tmp_773_22;
  localparam _tmp_774 = 1;
  wire [_tmp_774-1:0] _tmp_775;
  assign _tmp_775 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_774-1:0] __tmp_775_1;
  reg [_tmp_774-1:0] __tmp_775_2;
  reg [_tmp_774-1:0] __tmp_775_3;
  reg [_tmp_774-1:0] __tmp_775_4;
  reg [_tmp_774-1:0] __tmp_775_5;
  reg [_tmp_774-1:0] __tmp_775_6;
  reg [_tmp_774-1:0] __tmp_775_7;
  reg [_tmp_774-1:0] __tmp_775_8;
  reg [_tmp_774-1:0] __tmp_775_9;
  reg [_tmp_774-1:0] __tmp_775_10;
  reg [_tmp_774-1:0] __tmp_775_11;
  reg [_tmp_774-1:0] __tmp_775_12;
  reg [_tmp_774-1:0] __tmp_775_13;
  reg [_tmp_774-1:0] __tmp_775_14;
  reg [_tmp_774-1:0] __tmp_775_15;
  reg [_tmp_774-1:0] __tmp_775_16;
  reg [_tmp_774-1:0] __tmp_775_17;
  reg [_tmp_774-1:0] __tmp_775_18;
  reg [_tmp_774-1:0] __tmp_775_19;
  reg [_tmp_774-1:0] __tmp_775_20;
  reg [_tmp_774-1:0] __tmp_775_21;
  reg [_tmp_774-1:0] __tmp_775_22;
  localparam _tmp_776 = 1;
  wire [_tmp_776-1:0] _tmp_777;
  assign _tmp_777 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_776-1:0] __tmp_777_1;
  reg [_tmp_776-1:0] __tmp_777_2;
  reg [_tmp_776-1:0] __tmp_777_3;
  reg [_tmp_776-1:0] __tmp_777_4;
  reg [_tmp_776-1:0] __tmp_777_5;
  reg [_tmp_776-1:0] __tmp_777_6;
  reg [_tmp_776-1:0] __tmp_777_7;
  reg [_tmp_776-1:0] __tmp_777_8;
  reg [_tmp_776-1:0] __tmp_777_9;
  reg [_tmp_776-1:0] __tmp_777_10;
  reg [_tmp_776-1:0] __tmp_777_11;
  reg [_tmp_776-1:0] __tmp_777_12;
  reg [_tmp_776-1:0] __tmp_777_13;
  reg [_tmp_776-1:0] __tmp_777_14;
  reg [_tmp_776-1:0] __tmp_777_15;
  reg [_tmp_776-1:0] __tmp_777_16;
  reg [_tmp_776-1:0] __tmp_777_17;
  reg [_tmp_776-1:0] __tmp_777_18;
  reg [_tmp_776-1:0] __tmp_777_19;
  reg [_tmp_776-1:0] __tmp_777_20;
  reg [_tmp_776-1:0] __tmp_777_21;
  reg [_tmp_776-1:0] __tmp_777_22;
  localparam _tmp_778 = 1;
  wire [_tmp_778-1:0] _tmp_779;
  assign _tmp_779 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_778-1:0] __tmp_779_1;
  reg [_tmp_778-1:0] __tmp_779_2;
  reg [_tmp_778-1:0] __tmp_779_3;
  reg [_tmp_778-1:0] __tmp_779_4;
  reg [_tmp_778-1:0] __tmp_779_5;
  reg [_tmp_778-1:0] __tmp_779_6;
  reg [_tmp_778-1:0] __tmp_779_7;
  reg [_tmp_778-1:0] __tmp_779_8;
  reg [_tmp_778-1:0] __tmp_779_9;
  reg [_tmp_778-1:0] __tmp_779_10;
  reg [_tmp_778-1:0] __tmp_779_11;
  reg [_tmp_778-1:0] __tmp_779_12;
  reg [_tmp_778-1:0] __tmp_779_13;
  reg [_tmp_778-1:0] __tmp_779_14;
  reg [_tmp_778-1:0] __tmp_779_15;
  reg [_tmp_778-1:0] __tmp_779_16;
  reg [_tmp_778-1:0] __tmp_779_17;
  reg [_tmp_778-1:0] __tmp_779_18;
  reg [_tmp_778-1:0] __tmp_779_19;
  reg [_tmp_778-1:0] __tmp_779_20;
  reg [_tmp_778-1:0] __tmp_779_21;
  reg [_tmp_778-1:0] __tmp_779_22;
  localparam _tmp_780 = 1;
  wire [_tmp_780-1:0] _tmp_781;
  assign _tmp_781 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_780-1:0] __tmp_781_1;
  reg [_tmp_780-1:0] __tmp_781_2;
  reg [_tmp_780-1:0] __tmp_781_3;
  reg [_tmp_780-1:0] __tmp_781_4;
  reg [_tmp_780-1:0] __tmp_781_5;
  reg [_tmp_780-1:0] __tmp_781_6;
  reg [_tmp_780-1:0] __tmp_781_7;
  reg [_tmp_780-1:0] __tmp_781_8;
  reg [_tmp_780-1:0] __tmp_781_9;
  reg [_tmp_780-1:0] __tmp_781_10;
  reg [_tmp_780-1:0] __tmp_781_11;
  reg [_tmp_780-1:0] __tmp_781_12;
  reg [_tmp_780-1:0] __tmp_781_13;
  reg [_tmp_780-1:0] __tmp_781_14;
  reg [_tmp_780-1:0] __tmp_781_15;
  reg [_tmp_780-1:0] __tmp_781_16;
  reg [_tmp_780-1:0] __tmp_781_17;
  reg [_tmp_780-1:0] __tmp_781_18;
  reg [_tmp_780-1:0] __tmp_781_19;
  reg [_tmp_780-1:0] __tmp_781_20;
  reg [_tmp_780-1:0] __tmp_781_21;
  reg [_tmp_780-1:0] __tmp_781_22;
  localparam _tmp_782 = 1;
  wire [_tmp_782-1:0] _tmp_783;
  assign _tmp_783 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_782-1:0] __tmp_783_1;
  reg [_tmp_782-1:0] __tmp_783_2;
  reg [_tmp_782-1:0] __tmp_783_3;
  reg [_tmp_782-1:0] __tmp_783_4;
  reg [_tmp_782-1:0] __tmp_783_5;
  reg [_tmp_782-1:0] __tmp_783_6;
  reg [_tmp_782-1:0] __tmp_783_7;
  reg [_tmp_782-1:0] __tmp_783_8;
  reg [_tmp_782-1:0] __tmp_783_9;
  reg [_tmp_782-1:0] __tmp_783_10;
  reg [_tmp_782-1:0] __tmp_783_11;
  reg [_tmp_782-1:0] __tmp_783_12;
  reg [_tmp_782-1:0] __tmp_783_13;
  reg [_tmp_782-1:0] __tmp_783_14;
  reg [_tmp_782-1:0] __tmp_783_15;
  reg [_tmp_782-1:0] __tmp_783_16;
  reg [_tmp_782-1:0] __tmp_783_17;
  reg [_tmp_782-1:0] __tmp_783_18;
  reg [_tmp_782-1:0] __tmp_783_19;
  reg [_tmp_782-1:0] __tmp_783_20;
  reg [_tmp_782-1:0] __tmp_783_21;
  reg [_tmp_782-1:0] __tmp_783_22;
  localparam _tmp_784 = 1;
  wire [_tmp_784-1:0] _tmp_785;
  assign _tmp_785 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_784-1:0] __tmp_785_1;
  reg [_tmp_784-1:0] __tmp_785_2;
  reg [_tmp_784-1:0] __tmp_785_3;
  reg [_tmp_784-1:0] __tmp_785_4;
  reg [_tmp_784-1:0] __tmp_785_5;
  reg [_tmp_784-1:0] __tmp_785_6;
  reg [_tmp_784-1:0] __tmp_785_7;
  reg [_tmp_784-1:0] __tmp_785_8;
  reg [_tmp_784-1:0] __tmp_785_9;
  reg [_tmp_784-1:0] __tmp_785_10;
  reg [_tmp_784-1:0] __tmp_785_11;
  reg [_tmp_784-1:0] __tmp_785_12;
  reg [_tmp_784-1:0] __tmp_785_13;
  reg [_tmp_784-1:0] __tmp_785_14;
  reg [_tmp_784-1:0] __tmp_785_15;
  reg [_tmp_784-1:0] __tmp_785_16;
  reg [_tmp_784-1:0] __tmp_785_17;
  reg [_tmp_784-1:0] __tmp_785_18;
  reg [_tmp_784-1:0] __tmp_785_19;
  reg [_tmp_784-1:0] __tmp_785_20;
  reg [_tmp_784-1:0] __tmp_785_21;
  reg [_tmp_784-1:0] __tmp_785_22;
  localparam _tmp_786 = 1;
  wire [_tmp_786-1:0] _tmp_787;
  assign _tmp_787 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_786-1:0] __tmp_787_1;
  reg [_tmp_786-1:0] __tmp_787_2;
  reg [_tmp_786-1:0] __tmp_787_3;
  reg [_tmp_786-1:0] __tmp_787_4;
  reg [_tmp_786-1:0] __tmp_787_5;
  reg [_tmp_786-1:0] __tmp_787_6;
  reg [_tmp_786-1:0] __tmp_787_7;
  reg [_tmp_786-1:0] __tmp_787_8;
  reg [_tmp_786-1:0] __tmp_787_9;
  reg [_tmp_786-1:0] __tmp_787_10;
  reg [_tmp_786-1:0] __tmp_787_11;
  reg [_tmp_786-1:0] __tmp_787_12;
  reg [_tmp_786-1:0] __tmp_787_13;
  reg [_tmp_786-1:0] __tmp_787_14;
  reg [_tmp_786-1:0] __tmp_787_15;
  reg [_tmp_786-1:0] __tmp_787_16;
  reg [_tmp_786-1:0] __tmp_787_17;
  reg [_tmp_786-1:0] __tmp_787_18;
  reg [_tmp_786-1:0] __tmp_787_19;
  reg [_tmp_786-1:0] __tmp_787_20;
  reg [_tmp_786-1:0] __tmp_787_21;
  reg [_tmp_786-1:0] __tmp_787_22;
  reg [_tmp_786-1:0] __tmp_787_23;
  reg [_tmp_786-1:0] __tmp_787_24;
  reg [_tmp_786-1:0] __tmp_787_25;
  reg [_tmp_786-1:0] __tmp_787_26;
  reg [_tmp_786-1:0] __tmp_787_27;
  reg [_tmp_786-1:0] __tmp_787_28;
  localparam _tmp_788 = 1;
  wire [_tmp_788-1:0] _tmp_789;
  assign _tmp_789 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_788-1:0] __tmp_789_1;
  reg [_tmp_788-1:0] __tmp_789_2;
  reg [_tmp_788-1:0] __tmp_789_3;
  reg [_tmp_788-1:0] __tmp_789_4;
  reg [_tmp_788-1:0] __tmp_789_5;
  reg [_tmp_788-1:0] __tmp_789_6;
  reg [_tmp_788-1:0] __tmp_789_7;
  reg [_tmp_788-1:0] __tmp_789_8;
  reg [_tmp_788-1:0] __tmp_789_9;
  reg [_tmp_788-1:0] __tmp_789_10;
  reg [_tmp_788-1:0] __tmp_789_11;
  reg [_tmp_788-1:0] __tmp_789_12;
  reg [_tmp_788-1:0] __tmp_789_13;
  reg [_tmp_788-1:0] __tmp_789_14;
  reg [_tmp_788-1:0] __tmp_789_15;
  reg [_tmp_788-1:0] __tmp_789_16;
  reg [_tmp_788-1:0] __tmp_789_17;
  reg [_tmp_788-1:0] __tmp_789_18;
  reg [_tmp_788-1:0] __tmp_789_19;
  reg [_tmp_788-1:0] __tmp_789_20;
  reg [_tmp_788-1:0] __tmp_789_21;
  reg [_tmp_788-1:0] __tmp_789_22;
  reg [_tmp_788-1:0] __tmp_789_23;
  reg [_tmp_788-1:0] __tmp_789_24;
  reg [_tmp_788-1:0] __tmp_789_25;
  reg [_tmp_788-1:0] __tmp_789_26;
  localparam _tmp_790 = 1;
  wire [_tmp_790-1:0] _tmp_791;
  assign _tmp_791 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_790-1:0] __tmp_791_1;
  reg [_tmp_790-1:0] __tmp_791_2;
  reg [_tmp_790-1:0] __tmp_791_3;
  reg [_tmp_790-1:0] __tmp_791_4;
  reg [_tmp_790-1:0] __tmp_791_5;
  reg [_tmp_790-1:0] __tmp_791_6;
  reg [_tmp_790-1:0] __tmp_791_7;
  reg [_tmp_790-1:0] __tmp_791_8;
  reg [_tmp_790-1:0] __tmp_791_9;
  reg [_tmp_790-1:0] __tmp_791_10;
  reg [_tmp_790-1:0] __tmp_791_11;
  reg [_tmp_790-1:0] __tmp_791_12;
  reg [_tmp_790-1:0] __tmp_791_13;
  reg [_tmp_790-1:0] __tmp_791_14;
  reg [_tmp_790-1:0] __tmp_791_15;
  reg [_tmp_790-1:0] __tmp_791_16;
  reg [_tmp_790-1:0] __tmp_791_17;
  reg [_tmp_790-1:0] __tmp_791_18;
  reg [_tmp_790-1:0] __tmp_791_19;
  reg [_tmp_790-1:0] __tmp_791_20;
  reg [_tmp_790-1:0] __tmp_791_21;
  reg [_tmp_790-1:0] __tmp_791_22;
  reg [_tmp_790-1:0] __tmp_791_23;
  reg [_tmp_790-1:0] __tmp_791_24;
  reg [_tmp_790-1:0] __tmp_791_25;
  reg [_tmp_790-1:0] __tmp_791_26;
  localparam _tmp_792 = 1;
  wire [_tmp_792-1:0] _tmp_793;
  assign _tmp_793 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_792-1:0] __tmp_793_1;
  reg [_tmp_792-1:0] __tmp_793_2;
  reg [_tmp_792-1:0] __tmp_793_3;
  reg [_tmp_792-1:0] __tmp_793_4;
  reg [_tmp_792-1:0] __tmp_793_5;
  reg [_tmp_792-1:0] __tmp_793_6;
  reg [_tmp_792-1:0] __tmp_793_7;
  reg [_tmp_792-1:0] __tmp_793_8;
  reg [_tmp_792-1:0] __tmp_793_9;
  reg [_tmp_792-1:0] __tmp_793_10;
  reg [_tmp_792-1:0] __tmp_793_11;
  reg [_tmp_792-1:0] __tmp_793_12;
  reg [_tmp_792-1:0] __tmp_793_13;
  reg [_tmp_792-1:0] __tmp_793_14;
  reg [_tmp_792-1:0] __tmp_793_15;
  reg [_tmp_792-1:0] __tmp_793_16;
  reg [_tmp_792-1:0] __tmp_793_17;
  reg [_tmp_792-1:0] __tmp_793_18;
  reg [_tmp_792-1:0] __tmp_793_19;
  reg [_tmp_792-1:0] __tmp_793_20;
  reg [_tmp_792-1:0] __tmp_793_21;
  reg [_tmp_792-1:0] __tmp_793_22;
  reg [_tmp_792-1:0] __tmp_793_23;
  reg [_tmp_792-1:0] __tmp_793_24;
  reg [_tmp_792-1:0] __tmp_793_25;
  reg [_tmp_792-1:0] __tmp_793_26;
  localparam _tmp_794 = 1;
  wire [_tmp_794-1:0] _tmp_795;
  assign _tmp_795 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_794-1:0] __tmp_795_1;
  reg [_tmp_794-1:0] __tmp_795_2;
  reg [_tmp_794-1:0] __tmp_795_3;
  reg [_tmp_794-1:0] __tmp_795_4;
  reg [_tmp_794-1:0] __tmp_795_5;
  reg [_tmp_794-1:0] __tmp_795_6;
  reg [_tmp_794-1:0] __tmp_795_7;
  reg [_tmp_794-1:0] __tmp_795_8;
  reg [_tmp_794-1:0] __tmp_795_9;
  reg [_tmp_794-1:0] __tmp_795_10;
  reg [_tmp_794-1:0] __tmp_795_11;
  reg [_tmp_794-1:0] __tmp_795_12;
  reg [_tmp_794-1:0] __tmp_795_13;
  reg [_tmp_794-1:0] __tmp_795_14;
  reg [_tmp_794-1:0] __tmp_795_15;
  reg [_tmp_794-1:0] __tmp_795_16;
  reg [_tmp_794-1:0] __tmp_795_17;
  reg [_tmp_794-1:0] __tmp_795_18;
  reg [_tmp_794-1:0] __tmp_795_19;
  reg [_tmp_794-1:0] __tmp_795_20;
  reg [_tmp_794-1:0] __tmp_795_21;
  reg [_tmp_794-1:0] __tmp_795_22;
  reg [_tmp_794-1:0] __tmp_795_23;
  reg [_tmp_794-1:0] __tmp_795_24;
  reg [_tmp_794-1:0] __tmp_795_25;
  reg [_tmp_794-1:0] __tmp_795_26;
  reg [_tmp_794-1:0] __tmp_795_27;
  reg [_tmp_794-1:0] __tmp_795_28;
  reg [_tmp_794-1:0] __tmp_795_29;
  reg [_tmp_794-1:0] __tmp_795_30;
  reg [_tmp_794-1:0] __tmp_795_31;
  reg [_tmp_794-1:0] __tmp_795_32;
  reg [_tmp_794-1:0] __tmp_795_33;
  reg [_tmp_794-1:0] __tmp_795_34;
  localparam _tmp_796 = 1;
  wire [_tmp_796-1:0] _tmp_797;
  assign _tmp_797 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_796-1:0] __tmp_797_1;
  reg [_tmp_796-1:0] __tmp_797_2;
  reg [_tmp_796-1:0] __tmp_797_3;
  reg [_tmp_796-1:0] __tmp_797_4;
  reg [_tmp_796-1:0] __tmp_797_5;
  reg [_tmp_796-1:0] __tmp_797_6;
  reg [_tmp_796-1:0] __tmp_797_7;
  reg [_tmp_796-1:0] __tmp_797_8;
  reg [_tmp_796-1:0] __tmp_797_9;
  reg [_tmp_796-1:0] __tmp_797_10;
  reg [_tmp_796-1:0] __tmp_797_11;
  reg [_tmp_796-1:0] __tmp_797_12;
  reg [_tmp_796-1:0] __tmp_797_13;
  reg [_tmp_796-1:0] __tmp_797_14;
  reg [_tmp_796-1:0] __tmp_797_15;
  reg [_tmp_796-1:0] __tmp_797_16;
  reg [_tmp_796-1:0] __tmp_797_17;
  reg [_tmp_796-1:0] __tmp_797_18;
  reg [_tmp_796-1:0] __tmp_797_19;
  reg [_tmp_796-1:0] __tmp_797_20;
  reg [_tmp_796-1:0] __tmp_797_21;
  reg [_tmp_796-1:0] __tmp_797_22;
  reg [_tmp_796-1:0] __tmp_797_23;
  reg [_tmp_796-1:0] __tmp_797_24;
  reg [_tmp_796-1:0] __tmp_797_25;
  reg [_tmp_796-1:0] __tmp_797_26;
  reg [_tmp_796-1:0] __tmp_797_27;
  reg [_tmp_796-1:0] __tmp_797_28;
  reg [_tmp_796-1:0] __tmp_797_29;
  reg [_tmp_796-1:0] __tmp_797_30;
  reg [_tmp_796-1:0] __tmp_797_31;
  reg [_tmp_796-1:0] __tmp_797_32;
  reg [_tmp_796-1:0] __tmp_797_33;
  reg [_tmp_796-1:0] __tmp_797_34;
  localparam _tmp_798 = 1;
  wire [_tmp_798-1:0] _tmp_799;
  assign _tmp_799 = (_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag;
  reg [_tmp_798-1:0] __tmp_799_1;
  reg [_tmp_798-1:0] __tmp_799_2;
  reg [_tmp_798-1:0] __tmp_799_3;
  reg [_tmp_798-1:0] __tmp_799_4;
  reg [_tmp_798-1:0] __tmp_799_5;
  reg [_tmp_798-1:0] __tmp_799_6;
  reg [_tmp_798-1:0] __tmp_799_7;
  reg [_tmp_798-1:0] __tmp_799_8;
  reg [_tmp_798-1:0] __tmp_799_9;
  reg [_tmp_798-1:0] __tmp_799_10;
  reg [_tmp_798-1:0] __tmp_799_11;
  reg [_tmp_798-1:0] __tmp_799_12;
  reg [_tmp_798-1:0] __tmp_799_13;
  reg [_tmp_798-1:0] __tmp_799_14;
  reg [_tmp_798-1:0] __tmp_799_15;
  reg [_tmp_798-1:0] __tmp_799_16;
  reg [_tmp_798-1:0] __tmp_799_17;
  reg [_tmp_798-1:0] __tmp_799_18;
  reg [_tmp_798-1:0] __tmp_799_19;
  reg [_tmp_798-1:0] __tmp_799_20;
  reg [_tmp_798-1:0] __tmp_799_21;
  reg [_tmp_798-1:0] __tmp_799_22;
  reg [_tmp_798-1:0] __tmp_799_23;
  reg [_tmp_798-1:0] __tmp_799_24;
  reg [_tmp_798-1:0] __tmp_799_25;
  reg [_tmp_798-1:0] __tmp_799_26;
  reg [_tmp_798-1:0] __tmp_799_27;
  reg [_tmp_798-1:0] __tmp_799_28;
  reg [_tmp_798-1:0] __tmp_799_29;
  reg [_tmp_798-1:0] __tmp_799_30;
  reg [_tmp_798-1:0] __tmp_799_31;
  reg [_tmp_798-1:0] __tmp_799_32;
  reg [_tmp_798-1:0] __tmp_799_33;
  reg [_tmp_798-1:0] __tmp_799_34;
  wire _stream_conv2d_16_done;
  assign _stream_conv2d_16_done = _stream_conv2d_16_source_10_idle && _stream_conv2d_16_source_12_idle && _stream_conv2d_16_source_14_idle && _stream_conv2d_16_source_19_idle && _stream_conv2d_16_source_20_idle && _stream_conv2d_16_source_21_idle && _stream_conv2d_16_source_22_idle && _stream_conv2d_16_source_23_idle && _stream_conv2d_16_source_24_idle && _stream_conv2d_16_source_25_idle && _stream_conv2d_16_source_26_idle && _stream_conv2d_16_source_27_idle && _stream_conv2d_16_source_28_idle && _stream_conv2d_16_source_29_idle && _stream_conv2d_16_source_30_idle && _stream_conv2d_16_source_31_idle && _stream_conv2d_16_source_32_idle && _stream_conv2d_16_source_33_idle && _stream_conv2d_16_source_34_idle && _stream_conv2d_16_source_35_idle && _stream_conv2d_16_source_36_idle && _stream_conv2d_16_source_6_idle && _stream_conv2d_16_source_8_idle;
  localparam _tmp_800 = 1;
  wire [_tmp_800-1:0] _tmp_801;
  assign _tmp_801 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_800-1:0] __tmp_801_1;
  localparam _tmp_802 = 1;
  wire [_tmp_802-1:0] _tmp_803;
  assign _tmp_803 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_802-1:0] __tmp_803_1;
  reg [_tmp_802-1:0] __tmp_803_2;
  reg [_tmp_802-1:0] __tmp_803_3;
  reg [_tmp_802-1:0] __tmp_803_4;
  reg [_tmp_802-1:0] __tmp_803_5;
  reg [_tmp_802-1:0] __tmp_803_6;
  reg [_tmp_802-1:0] __tmp_803_7;
  reg [_tmp_802-1:0] __tmp_803_8;
  reg [_tmp_802-1:0] __tmp_803_9;
  localparam _tmp_804 = 1;
  wire [_tmp_804-1:0] _tmp_805;
  assign _tmp_805 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_804-1:0] __tmp_805_1;
  reg [_tmp_804-1:0] __tmp_805_2;
  reg [_tmp_804-1:0] __tmp_805_3;
  reg [_tmp_804-1:0] __tmp_805_4;
  reg [_tmp_804-1:0] __tmp_805_5;
  reg [_tmp_804-1:0] __tmp_805_6;
  reg [_tmp_804-1:0] __tmp_805_7;
  reg [_tmp_804-1:0] __tmp_805_8;
  reg [_tmp_804-1:0] __tmp_805_9;
  localparam _tmp_806 = 1;
  wire [_tmp_806-1:0] _tmp_807;
  assign _tmp_807 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_806-1:0] __tmp_807_1;
  reg [_tmp_806-1:0] __tmp_807_2;
  reg [_tmp_806-1:0] __tmp_807_3;
  reg [_tmp_806-1:0] __tmp_807_4;
  reg [_tmp_806-1:0] __tmp_807_5;
  reg [_tmp_806-1:0] __tmp_807_6;
  reg [_tmp_806-1:0] __tmp_807_7;
  reg [_tmp_806-1:0] __tmp_807_8;
  reg [_tmp_806-1:0] __tmp_807_9;
  reg [4-1:0] _mul_4_sink_wait_count;
  localparam _tmp_808 = 1;
  wire [_tmp_808-1:0] _tmp_809;
  assign _tmp_809 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_808-1:0] __tmp_809_1;
  reg [_tmp_808-1:0] __tmp_809_2;
  reg [_tmp_808-1:0] __tmp_809_3;
  reg [_tmp_808-1:0] __tmp_809_4;
  reg [_tmp_808-1:0] __tmp_809_5;
  reg [_tmp_808-1:0] __tmp_809_6;
  reg [_tmp_808-1:0] __tmp_809_7;
  reg [_tmp_808-1:0] __tmp_809_8;
  reg [_tmp_808-1:0] __tmp_809_9;
  reg [_tmp_808-1:0] __tmp_809_10;
  reg [_tmp_808-1:0] __tmp_809_11;
  reg [_tmp_808-1:0] __tmp_809_12;
  localparam _tmp_810 = 1;
  wire [_tmp_810-1:0] _tmp_811;
  assign _tmp_811 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_810-1:0] __tmp_811_1;
  reg [_tmp_810-1:0] __tmp_811_2;
  reg [_tmp_810-1:0] __tmp_811_3;
  reg [_tmp_810-1:0] __tmp_811_4;
  reg [_tmp_810-1:0] __tmp_811_5;
  reg [_tmp_810-1:0] __tmp_811_6;
  reg [_tmp_810-1:0] __tmp_811_7;
  reg [_tmp_810-1:0] __tmp_811_8;
  reg [_tmp_810-1:0] __tmp_811_9;
  reg [_tmp_810-1:0] __tmp_811_10;
  reg [_tmp_810-1:0] __tmp_811_11;
  reg [_tmp_810-1:0] __tmp_811_12;
  localparam _tmp_812 = 1;
  wire [_tmp_812-1:0] _tmp_813;
  assign _tmp_813 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_812-1:0] __tmp_813_1;
  reg [_tmp_812-1:0] __tmp_813_2;
  reg [_tmp_812-1:0] __tmp_813_3;
  reg [_tmp_812-1:0] __tmp_813_4;
  reg [_tmp_812-1:0] __tmp_813_5;
  reg [_tmp_812-1:0] __tmp_813_6;
  reg [_tmp_812-1:0] __tmp_813_7;
  reg [_tmp_812-1:0] __tmp_813_8;
  reg [_tmp_812-1:0] __tmp_813_9;
  reg [_tmp_812-1:0] __tmp_813_10;
  reg [_tmp_812-1:0] __tmp_813_11;
  reg [_tmp_812-1:0] __tmp_813_12;
  localparam _tmp_814 = 1;
  wire [_tmp_814-1:0] _tmp_815;
  assign _tmp_815 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_814-1:0] __tmp_815_1;
  reg [_tmp_814-1:0] __tmp_815_2;
  reg [_tmp_814-1:0] __tmp_815_3;
  reg [_tmp_814-1:0] __tmp_815_4;
  reg [_tmp_814-1:0] __tmp_815_5;
  reg [_tmp_814-1:0] __tmp_815_6;
  reg [_tmp_814-1:0] __tmp_815_7;
  reg [_tmp_814-1:0] __tmp_815_8;
  reg [_tmp_814-1:0] __tmp_815_9;
  localparam _tmp_816 = 1;
  wire [_tmp_816-1:0] _tmp_817;
  assign _tmp_817 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_816-1:0] __tmp_817_1;
  reg [_tmp_816-1:0] __tmp_817_2;
  reg [_tmp_816-1:0] __tmp_817_3;
  reg [_tmp_816-1:0] __tmp_817_4;
  reg [_tmp_816-1:0] __tmp_817_5;
  reg [_tmp_816-1:0] __tmp_817_6;
  reg [_tmp_816-1:0] __tmp_817_7;
  reg [_tmp_816-1:0] __tmp_817_8;
  reg [_tmp_816-1:0] __tmp_817_9;
  localparam _tmp_818 = 1;
  wire [_tmp_818-1:0] _tmp_819;
  assign _tmp_819 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_818-1:0] __tmp_819_1;
  reg [_tmp_818-1:0] __tmp_819_2;
  reg [_tmp_818-1:0] __tmp_819_3;
  reg [_tmp_818-1:0] __tmp_819_4;
  reg [_tmp_818-1:0] __tmp_819_5;
  reg [_tmp_818-1:0] __tmp_819_6;
  reg [_tmp_818-1:0] __tmp_819_7;
  reg [_tmp_818-1:0] __tmp_819_8;
  reg [_tmp_818-1:0] __tmp_819_9;
  reg [4-1:0] _mul_5_sink_wait_count;
  localparam _tmp_820 = 1;
  wire [_tmp_820-1:0] _tmp_821;
  assign _tmp_821 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_820-1:0] __tmp_821_1;
  reg [_tmp_820-1:0] __tmp_821_2;
  reg [_tmp_820-1:0] __tmp_821_3;
  reg [_tmp_820-1:0] __tmp_821_4;
  reg [_tmp_820-1:0] __tmp_821_5;
  reg [_tmp_820-1:0] __tmp_821_6;
  reg [_tmp_820-1:0] __tmp_821_7;
  reg [_tmp_820-1:0] __tmp_821_8;
  reg [_tmp_820-1:0] __tmp_821_9;
  reg [_tmp_820-1:0] __tmp_821_10;
  reg [_tmp_820-1:0] __tmp_821_11;
  reg [_tmp_820-1:0] __tmp_821_12;
  localparam _tmp_822 = 1;
  wire [_tmp_822-1:0] _tmp_823;
  assign _tmp_823 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_822-1:0] __tmp_823_1;
  reg [_tmp_822-1:0] __tmp_823_2;
  reg [_tmp_822-1:0] __tmp_823_3;
  reg [_tmp_822-1:0] __tmp_823_4;
  reg [_tmp_822-1:0] __tmp_823_5;
  reg [_tmp_822-1:0] __tmp_823_6;
  reg [_tmp_822-1:0] __tmp_823_7;
  reg [_tmp_822-1:0] __tmp_823_8;
  reg [_tmp_822-1:0] __tmp_823_9;
  reg [_tmp_822-1:0] __tmp_823_10;
  reg [_tmp_822-1:0] __tmp_823_11;
  reg [_tmp_822-1:0] __tmp_823_12;
  localparam _tmp_824 = 1;
  wire [_tmp_824-1:0] _tmp_825;
  assign _tmp_825 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_824-1:0] __tmp_825_1;
  reg [_tmp_824-1:0] __tmp_825_2;
  reg [_tmp_824-1:0] __tmp_825_3;
  reg [_tmp_824-1:0] __tmp_825_4;
  reg [_tmp_824-1:0] __tmp_825_5;
  reg [_tmp_824-1:0] __tmp_825_6;
  reg [_tmp_824-1:0] __tmp_825_7;
  reg [_tmp_824-1:0] __tmp_825_8;
  reg [_tmp_824-1:0] __tmp_825_9;
  reg [_tmp_824-1:0] __tmp_825_10;
  reg [_tmp_824-1:0] __tmp_825_11;
  reg [_tmp_824-1:0] __tmp_825_12;
  localparam _tmp_826 = 1;
  wire [_tmp_826-1:0] _tmp_827;
  assign _tmp_827 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_826-1:0] __tmp_827_1;
  reg [_tmp_826-1:0] __tmp_827_2;
  reg [_tmp_826-1:0] __tmp_827_3;
  reg [_tmp_826-1:0] __tmp_827_4;
  reg [_tmp_826-1:0] __tmp_827_5;
  reg [_tmp_826-1:0] __tmp_827_6;
  reg [_tmp_826-1:0] __tmp_827_7;
  reg [_tmp_826-1:0] __tmp_827_8;
  reg [_tmp_826-1:0] __tmp_827_9;
  localparam _tmp_828 = 1;
  wire [_tmp_828-1:0] _tmp_829;
  assign _tmp_829 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_828-1:0] __tmp_829_1;
  reg [_tmp_828-1:0] __tmp_829_2;
  reg [_tmp_828-1:0] __tmp_829_3;
  reg [_tmp_828-1:0] __tmp_829_4;
  reg [_tmp_828-1:0] __tmp_829_5;
  reg [_tmp_828-1:0] __tmp_829_6;
  reg [_tmp_828-1:0] __tmp_829_7;
  reg [_tmp_828-1:0] __tmp_829_8;
  reg [_tmp_828-1:0] __tmp_829_9;
  localparam _tmp_830 = 1;
  wire [_tmp_830-1:0] _tmp_831;
  assign _tmp_831 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_830-1:0] __tmp_831_1;
  reg [_tmp_830-1:0] __tmp_831_2;
  reg [_tmp_830-1:0] __tmp_831_3;
  reg [_tmp_830-1:0] __tmp_831_4;
  reg [_tmp_830-1:0] __tmp_831_5;
  reg [_tmp_830-1:0] __tmp_831_6;
  reg [_tmp_830-1:0] __tmp_831_7;
  reg [_tmp_830-1:0] __tmp_831_8;
  reg [_tmp_830-1:0] __tmp_831_9;
  reg [4-1:0] _mul_6_sink_wait_count;
  localparam _tmp_832 = 1;
  wire [_tmp_832-1:0] _tmp_833;
  assign _tmp_833 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_832-1:0] __tmp_833_1;
  reg [_tmp_832-1:0] __tmp_833_2;
  reg [_tmp_832-1:0] __tmp_833_3;
  reg [_tmp_832-1:0] __tmp_833_4;
  reg [_tmp_832-1:0] __tmp_833_5;
  reg [_tmp_832-1:0] __tmp_833_6;
  reg [_tmp_832-1:0] __tmp_833_7;
  reg [_tmp_832-1:0] __tmp_833_8;
  reg [_tmp_832-1:0] __tmp_833_9;
  reg [_tmp_832-1:0] __tmp_833_10;
  reg [_tmp_832-1:0] __tmp_833_11;
  reg [_tmp_832-1:0] __tmp_833_12;
  localparam _tmp_834 = 1;
  wire [_tmp_834-1:0] _tmp_835;
  assign _tmp_835 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_834-1:0] __tmp_835_1;
  reg [_tmp_834-1:0] __tmp_835_2;
  reg [_tmp_834-1:0] __tmp_835_3;
  reg [_tmp_834-1:0] __tmp_835_4;
  reg [_tmp_834-1:0] __tmp_835_5;
  reg [_tmp_834-1:0] __tmp_835_6;
  reg [_tmp_834-1:0] __tmp_835_7;
  reg [_tmp_834-1:0] __tmp_835_8;
  reg [_tmp_834-1:0] __tmp_835_9;
  reg [_tmp_834-1:0] __tmp_835_10;
  reg [_tmp_834-1:0] __tmp_835_11;
  reg [_tmp_834-1:0] __tmp_835_12;
  localparam _tmp_836 = 1;
  wire [_tmp_836-1:0] _tmp_837;
  assign _tmp_837 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_836-1:0] __tmp_837_1;
  reg [_tmp_836-1:0] __tmp_837_2;
  reg [_tmp_836-1:0] __tmp_837_3;
  reg [_tmp_836-1:0] __tmp_837_4;
  reg [_tmp_836-1:0] __tmp_837_5;
  reg [_tmp_836-1:0] __tmp_837_6;
  reg [_tmp_836-1:0] __tmp_837_7;
  reg [_tmp_836-1:0] __tmp_837_8;
  reg [_tmp_836-1:0] __tmp_837_9;
  reg [_tmp_836-1:0] __tmp_837_10;
  reg [_tmp_836-1:0] __tmp_837_11;
  reg [_tmp_836-1:0] __tmp_837_12;
  localparam _tmp_838 = 1;
  wire [_tmp_838-1:0] _tmp_839;
  assign _tmp_839 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_838-1:0] __tmp_839_1;
  reg [_tmp_838-1:0] __tmp_839_2;
  reg [_tmp_838-1:0] __tmp_839_3;
  reg [_tmp_838-1:0] __tmp_839_4;
  reg [_tmp_838-1:0] __tmp_839_5;
  reg [_tmp_838-1:0] __tmp_839_6;
  reg [_tmp_838-1:0] __tmp_839_7;
  reg [_tmp_838-1:0] __tmp_839_8;
  reg [_tmp_838-1:0] __tmp_839_9;
  localparam _tmp_840 = 1;
  wire [_tmp_840-1:0] _tmp_841;
  assign _tmp_841 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_840-1:0] __tmp_841_1;
  reg [_tmp_840-1:0] __tmp_841_2;
  reg [_tmp_840-1:0] __tmp_841_3;
  reg [_tmp_840-1:0] __tmp_841_4;
  reg [_tmp_840-1:0] __tmp_841_5;
  reg [_tmp_840-1:0] __tmp_841_6;
  reg [_tmp_840-1:0] __tmp_841_7;
  reg [_tmp_840-1:0] __tmp_841_8;
  reg [_tmp_840-1:0] __tmp_841_9;
  localparam _tmp_842 = 1;
  wire [_tmp_842-1:0] _tmp_843;
  assign _tmp_843 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_842-1:0] __tmp_843_1;
  reg [_tmp_842-1:0] __tmp_843_2;
  reg [_tmp_842-1:0] __tmp_843_3;
  reg [_tmp_842-1:0] __tmp_843_4;
  reg [_tmp_842-1:0] __tmp_843_5;
  reg [_tmp_842-1:0] __tmp_843_6;
  reg [_tmp_842-1:0] __tmp_843_7;
  reg [_tmp_842-1:0] __tmp_843_8;
  reg [_tmp_842-1:0] __tmp_843_9;
  reg [4-1:0] _mul_7_sink_wait_count;
  localparam _tmp_844 = 1;
  wire [_tmp_844-1:0] _tmp_845;
  assign _tmp_845 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_844-1:0] __tmp_845_1;
  reg [_tmp_844-1:0] __tmp_845_2;
  reg [_tmp_844-1:0] __tmp_845_3;
  reg [_tmp_844-1:0] __tmp_845_4;
  reg [_tmp_844-1:0] __tmp_845_5;
  reg [_tmp_844-1:0] __tmp_845_6;
  reg [_tmp_844-1:0] __tmp_845_7;
  reg [_tmp_844-1:0] __tmp_845_8;
  reg [_tmp_844-1:0] __tmp_845_9;
  reg [_tmp_844-1:0] __tmp_845_10;
  reg [_tmp_844-1:0] __tmp_845_11;
  reg [_tmp_844-1:0] __tmp_845_12;
  localparam _tmp_846 = 1;
  wire [_tmp_846-1:0] _tmp_847;
  assign _tmp_847 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_846-1:0] __tmp_847_1;
  reg [_tmp_846-1:0] __tmp_847_2;
  reg [_tmp_846-1:0] __tmp_847_3;
  reg [_tmp_846-1:0] __tmp_847_4;
  reg [_tmp_846-1:0] __tmp_847_5;
  reg [_tmp_846-1:0] __tmp_847_6;
  reg [_tmp_846-1:0] __tmp_847_7;
  reg [_tmp_846-1:0] __tmp_847_8;
  reg [_tmp_846-1:0] __tmp_847_9;
  reg [_tmp_846-1:0] __tmp_847_10;
  reg [_tmp_846-1:0] __tmp_847_11;
  reg [_tmp_846-1:0] __tmp_847_12;
  localparam _tmp_848 = 1;
  wire [_tmp_848-1:0] _tmp_849;
  assign _tmp_849 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_848-1:0] __tmp_849_1;
  reg [_tmp_848-1:0] __tmp_849_2;
  reg [_tmp_848-1:0] __tmp_849_3;
  reg [_tmp_848-1:0] __tmp_849_4;
  reg [_tmp_848-1:0] __tmp_849_5;
  reg [_tmp_848-1:0] __tmp_849_6;
  reg [_tmp_848-1:0] __tmp_849_7;
  reg [_tmp_848-1:0] __tmp_849_8;
  reg [_tmp_848-1:0] __tmp_849_9;
  reg [_tmp_848-1:0] __tmp_849_10;
  reg [_tmp_848-1:0] __tmp_849_11;
  reg [_tmp_848-1:0] __tmp_849_12;
  localparam _tmp_850 = 1;
  wire [_tmp_850-1:0] _tmp_851;
  assign _tmp_851 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_850-1:0] __tmp_851_1;
  reg [_tmp_850-1:0] __tmp_851_2;
  reg [_tmp_850-1:0] __tmp_851_3;
  reg [_tmp_850-1:0] __tmp_851_4;
  reg [_tmp_850-1:0] __tmp_851_5;
  reg [_tmp_850-1:0] __tmp_851_6;
  reg [_tmp_850-1:0] __tmp_851_7;
  reg [_tmp_850-1:0] __tmp_851_8;
  reg [_tmp_850-1:0] __tmp_851_9;
  localparam _tmp_852 = 1;
  wire [_tmp_852-1:0] _tmp_853;
  assign _tmp_853 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_852-1:0] __tmp_853_1;
  reg [_tmp_852-1:0] __tmp_853_2;
  reg [_tmp_852-1:0] __tmp_853_3;
  reg [_tmp_852-1:0] __tmp_853_4;
  reg [_tmp_852-1:0] __tmp_853_5;
  reg [_tmp_852-1:0] __tmp_853_6;
  reg [_tmp_852-1:0] __tmp_853_7;
  reg [_tmp_852-1:0] __tmp_853_8;
  reg [_tmp_852-1:0] __tmp_853_9;
  localparam _tmp_854 = 1;
  wire [_tmp_854-1:0] _tmp_855;
  assign _tmp_855 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_854-1:0] __tmp_855_1;
  reg [_tmp_854-1:0] __tmp_855_2;
  reg [_tmp_854-1:0] __tmp_855_3;
  reg [_tmp_854-1:0] __tmp_855_4;
  reg [_tmp_854-1:0] __tmp_855_5;
  reg [_tmp_854-1:0] __tmp_855_6;
  reg [_tmp_854-1:0] __tmp_855_7;
  reg [_tmp_854-1:0] __tmp_855_8;
  reg [_tmp_854-1:0] __tmp_855_9;
  reg [4-1:0] _mul_8_sink_wait_count;
  localparam _tmp_856 = 1;
  wire [_tmp_856-1:0] _tmp_857;
  assign _tmp_857 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_856-1:0] __tmp_857_1;
  reg [_tmp_856-1:0] __tmp_857_2;
  reg [_tmp_856-1:0] __tmp_857_3;
  reg [_tmp_856-1:0] __tmp_857_4;
  reg [_tmp_856-1:0] __tmp_857_5;
  reg [_tmp_856-1:0] __tmp_857_6;
  reg [_tmp_856-1:0] __tmp_857_7;
  reg [_tmp_856-1:0] __tmp_857_8;
  reg [_tmp_856-1:0] __tmp_857_9;
  reg [_tmp_856-1:0] __tmp_857_10;
  reg [_tmp_856-1:0] __tmp_857_11;
  reg [_tmp_856-1:0] __tmp_857_12;
  localparam _tmp_858 = 1;
  wire [_tmp_858-1:0] _tmp_859;
  assign _tmp_859 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_858-1:0] __tmp_859_1;
  reg [_tmp_858-1:0] __tmp_859_2;
  reg [_tmp_858-1:0] __tmp_859_3;
  reg [_tmp_858-1:0] __tmp_859_4;
  reg [_tmp_858-1:0] __tmp_859_5;
  reg [_tmp_858-1:0] __tmp_859_6;
  reg [_tmp_858-1:0] __tmp_859_7;
  reg [_tmp_858-1:0] __tmp_859_8;
  reg [_tmp_858-1:0] __tmp_859_9;
  reg [_tmp_858-1:0] __tmp_859_10;
  reg [_tmp_858-1:0] __tmp_859_11;
  reg [_tmp_858-1:0] __tmp_859_12;
  localparam _tmp_860 = 1;
  wire [_tmp_860-1:0] _tmp_861;
  assign _tmp_861 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_860-1:0] __tmp_861_1;
  reg [_tmp_860-1:0] __tmp_861_2;
  reg [_tmp_860-1:0] __tmp_861_3;
  reg [_tmp_860-1:0] __tmp_861_4;
  reg [_tmp_860-1:0] __tmp_861_5;
  reg [_tmp_860-1:0] __tmp_861_6;
  reg [_tmp_860-1:0] __tmp_861_7;
  reg [_tmp_860-1:0] __tmp_861_8;
  reg [_tmp_860-1:0] __tmp_861_9;
  reg [_tmp_860-1:0] __tmp_861_10;
  reg [_tmp_860-1:0] __tmp_861_11;
  reg [_tmp_860-1:0] __tmp_861_12;
  localparam _tmp_862 = 1;
  wire [_tmp_862-1:0] _tmp_863;
  assign _tmp_863 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_862-1:0] __tmp_863_1;
  reg [_tmp_862-1:0] __tmp_863_2;
  reg [_tmp_862-1:0] __tmp_863_3;
  reg [_tmp_862-1:0] __tmp_863_4;
  reg [_tmp_862-1:0] __tmp_863_5;
  reg [_tmp_862-1:0] __tmp_863_6;
  reg [_tmp_862-1:0] __tmp_863_7;
  reg [_tmp_862-1:0] __tmp_863_8;
  reg [_tmp_862-1:0] __tmp_863_9;
  localparam _tmp_864 = 1;
  wire [_tmp_864-1:0] _tmp_865;
  assign _tmp_865 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_864-1:0] __tmp_865_1;
  reg [_tmp_864-1:0] __tmp_865_2;
  reg [_tmp_864-1:0] __tmp_865_3;
  reg [_tmp_864-1:0] __tmp_865_4;
  reg [_tmp_864-1:0] __tmp_865_5;
  reg [_tmp_864-1:0] __tmp_865_6;
  reg [_tmp_864-1:0] __tmp_865_7;
  reg [_tmp_864-1:0] __tmp_865_8;
  reg [_tmp_864-1:0] __tmp_865_9;
  localparam _tmp_866 = 1;
  wire [_tmp_866-1:0] _tmp_867;
  assign _tmp_867 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_866-1:0] __tmp_867_1;
  reg [_tmp_866-1:0] __tmp_867_2;
  reg [_tmp_866-1:0] __tmp_867_3;
  reg [_tmp_866-1:0] __tmp_867_4;
  reg [_tmp_866-1:0] __tmp_867_5;
  reg [_tmp_866-1:0] __tmp_867_6;
  reg [_tmp_866-1:0] __tmp_867_7;
  reg [_tmp_866-1:0] __tmp_867_8;
  reg [_tmp_866-1:0] __tmp_867_9;
  reg [4-1:0] _mul_9_sink_wait_count;
  localparam _tmp_868 = 1;
  wire [_tmp_868-1:0] _tmp_869;
  assign _tmp_869 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_868-1:0] __tmp_869_1;
  reg [_tmp_868-1:0] __tmp_869_2;
  reg [_tmp_868-1:0] __tmp_869_3;
  reg [_tmp_868-1:0] __tmp_869_4;
  reg [_tmp_868-1:0] __tmp_869_5;
  reg [_tmp_868-1:0] __tmp_869_6;
  reg [_tmp_868-1:0] __tmp_869_7;
  reg [_tmp_868-1:0] __tmp_869_8;
  reg [_tmp_868-1:0] __tmp_869_9;
  reg [_tmp_868-1:0] __tmp_869_10;
  reg [_tmp_868-1:0] __tmp_869_11;
  reg [_tmp_868-1:0] __tmp_869_12;
  localparam _tmp_870 = 1;
  wire [_tmp_870-1:0] _tmp_871;
  assign _tmp_871 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_870-1:0] __tmp_871_1;
  reg [_tmp_870-1:0] __tmp_871_2;
  reg [_tmp_870-1:0] __tmp_871_3;
  reg [_tmp_870-1:0] __tmp_871_4;
  reg [_tmp_870-1:0] __tmp_871_5;
  reg [_tmp_870-1:0] __tmp_871_6;
  reg [_tmp_870-1:0] __tmp_871_7;
  reg [_tmp_870-1:0] __tmp_871_8;
  reg [_tmp_870-1:0] __tmp_871_9;
  reg [_tmp_870-1:0] __tmp_871_10;
  reg [_tmp_870-1:0] __tmp_871_11;
  reg [_tmp_870-1:0] __tmp_871_12;
  localparam _tmp_872 = 1;
  wire [_tmp_872-1:0] _tmp_873;
  assign _tmp_873 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_872-1:0] __tmp_873_1;
  reg [_tmp_872-1:0] __tmp_873_2;
  reg [_tmp_872-1:0] __tmp_873_3;
  reg [_tmp_872-1:0] __tmp_873_4;
  reg [_tmp_872-1:0] __tmp_873_5;
  reg [_tmp_872-1:0] __tmp_873_6;
  reg [_tmp_872-1:0] __tmp_873_7;
  reg [_tmp_872-1:0] __tmp_873_8;
  reg [_tmp_872-1:0] __tmp_873_9;
  reg [_tmp_872-1:0] __tmp_873_10;
  reg [_tmp_872-1:0] __tmp_873_11;
  reg [_tmp_872-1:0] __tmp_873_12;
  localparam _tmp_874 = 1;
  wire [_tmp_874-1:0] _tmp_875;
  assign _tmp_875 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_874-1:0] __tmp_875_1;
  reg [_tmp_874-1:0] __tmp_875_2;
  reg [_tmp_874-1:0] __tmp_875_3;
  reg [_tmp_874-1:0] __tmp_875_4;
  reg [_tmp_874-1:0] __tmp_875_5;
  reg [_tmp_874-1:0] __tmp_875_6;
  reg [_tmp_874-1:0] __tmp_875_7;
  reg [_tmp_874-1:0] __tmp_875_8;
  reg [_tmp_874-1:0] __tmp_875_9;
  localparam _tmp_876 = 1;
  wire [_tmp_876-1:0] _tmp_877;
  assign _tmp_877 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_876-1:0] __tmp_877_1;
  reg [_tmp_876-1:0] __tmp_877_2;
  reg [_tmp_876-1:0] __tmp_877_3;
  reg [_tmp_876-1:0] __tmp_877_4;
  reg [_tmp_876-1:0] __tmp_877_5;
  reg [_tmp_876-1:0] __tmp_877_6;
  reg [_tmp_876-1:0] __tmp_877_7;
  reg [_tmp_876-1:0] __tmp_877_8;
  reg [_tmp_876-1:0] __tmp_877_9;
  localparam _tmp_878 = 1;
  wire [_tmp_878-1:0] _tmp_879;
  assign _tmp_879 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_878-1:0] __tmp_879_1;
  reg [_tmp_878-1:0] __tmp_879_2;
  reg [_tmp_878-1:0] __tmp_879_3;
  reg [_tmp_878-1:0] __tmp_879_4;
  reg [_tmp_878-1:0] __tmp_879_5;
  reg [_tmp_878-1:0] __tmp_879_6;
  reg [_tmp_878-1:0] __tmp_879_7;
  reg [_tmp_878-1:0] __tmp_879_8;
  reg [_tmp_878-1:0] __tmp_879_9;
  reg [4-1:0] _mul_10_sink_wait_count;
  localparam _tmp_880 = 1;
  wire [_tmp_880-1:0] _tmp_881;
  assign _tmp_881 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_880-1:0] __tmp_881_1;
  reg [_tmp_880-1:0] __tmp_881_2;
  reg [_tmp_880-1:0] __tmp_881_3;
  reg [_tmp_880-1:0] __tmp_881_4;
  reg [_tmp_880-1:0] __tmp_881_5;
  reg [_tmp_880-1:0] __tmp_881_6;
  reg [_tmp_880-1:0] __tmp_881_7;
  reg [_tmp_880-1:0] __tmp_881_8;
  reg [_tmp_880-1:0] __tmp_881_9;
  reg [_tmp_880-1:0] __tmp_881_10;
  reg [_tmp_880-1:0] __tmp_881_11;
  reg [_tmp_880-1:0] __tmp_881_12;
  localparam _tmp_882 = 1;
  wire [_tmp_882-1:0] _tmp_883;
  assign _tmp_883 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_882-1:0] __tmp_883_1;
  reg [_tmp_882-1:0] __tmp_883_2;
  reg [_tmp_882-1:0] __tmp_883_3;
  reg [_tmp_882-1:0] __tmp_883_4;
  reg [_tmp_882-1:0] __tmp_883_5;
  reg [_tmp_882-1:0] __tmp_883_6;
  reg [_tmp_882-1:0] __tmp_883_7;
  reg [_tmp_882-1:0] __tmp_883_8;
  reg [_tmp_882-1:0] __tmp_883_9;
  reg [_tmp_882-1:0] __tmp_883_10;
  reg [_tmp_882-1:0] __tmp_883_11;
  reg [_tmp_882-1:0] __tmp_883_12;
  localparam _tmp_884 = 1;
  wire [_tmp_884-1:0] _tmp_885;
  assign _tmp_885 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_884-1:0] __tmp_885_1;
  reg [_tmp_884-1:0] __tmp_885_2;
  reg [_tmp_884-1:0] __tmp_885_3;
  reg [_tmp_884-1:0] __tmp_885_4;
  reg [_tmp_884-1:0] __tmp_885_5;
  reg [_tmp_884-1:0] __tmp_885_6;
  reg [_tmp_884-1:0] __tmp_885_7;
  reg [_tmp_884-1:0] __tmp_885_8;
  reg [_tmp_884-1:0] __tmp_885_9;
  reg [_tmp_884-1:0] __tmp_885_10;
  reg [_tmp_884-1:0] __tmp_885_11;
  reg [_tmp_884-1:0] __tmp_885_12;
  localparam _tmp_886 = 1;
  wire [_tmp_886-1:0] _tmp_887;
  assign _tmp_887 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_886-1:0] __tmp_887_1;
  reg [_tmp_886-1:0] __tmp_887_2;
  reg [_tmp_886-1:0] __tmp_887_3;
  reg [_tmp_886-1:0] __tmp_887_4;
  reg [_tmp_886-1:0] __tmp_887_5;
  reg [_tmp_886-1:0] __tmp_887_6;
  reg [_tmp_886-1:0] __tmp_887_7;
  reg [_tmp_886-1:0] __tmp_887_8;
  reg [_tmp_886-1:0] __tmp_887_9;
  localparam _tmp_888 = 1;
  wire [_tmp_888-1:0] _tmp_889;
  assign _tmp_889 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_888-1:0] __tmp_889_1;
  reg [_tmp_888-1:0] __tmp_889_2;
  reg [_tmp_888-1:0] __tmp_889_3;
  reg [_tmp_888-1:0] __tmp_889_4;
  reg [_tmp_888-1:0] __tmp_889_5;
  reg [_tmp_888-1:0] __tmp_889_6;
  reg [_tmp_888-1:0] __tmp_889_7;
  reg [_tmp_888-1:0] __tmp_889_8;
  reg [_tmp_888-1:0] __tmp_889_9;
  localparam _tmp_890 = 1;
  wire [_tmp_890-1:0] _tmp_891;
  assign _tmp_891 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_890-1:0] __tmp_891_1;
  reg [_tmp_890-1:0] __tmp_891_2;
  reg [_tmp_890-1:0] __tmp_891_3;
  reg [_tmp_890-1:0] __tmp_891_4;
  reg [_tmp_890-1:0] __tmp_891_5;
  reg [_tmp_890-1:0] __tmp_891_6;
  reg [_tmp_890-1:0] __tmp_891_7;
  reg [_tmp_890-1:0] __tmp_891_8;
  reg [_tmp_890-1:0] __tmp_891_9;
  reg [4-1:0] _mul_11_sink_wait_count;
  localparam _tmp_892 = 1;
  wire [_tmp_892-1:0] _tmp_893;
  assign _tmp_893 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_892-1:0] __tmp_893_1;
  reg [_tmp_892-1:0] __tmp_893_2;
  reg [_tmp_892-1:0] __tmp_893_3;
  reg [_tmp_892-1:0] __tmp_893_4;
  reg [_tmp_892-1:0] __tmp_893_5;
  reg [_tmp_892-1:0] __tmp_893_6;
  reg [_tmp_892-1:0] __tmp_893_7;
  reg [_tmp_892-1:0] __tmp_893_8;
  reg [_tmp_892-1:0] __tmp_893_9;
  reg [_tmp_892-1:0] __tmp_893_10;
  reg [_tmp_892-1:0] __tmp_893_11;
  reg [_tmp_892-1:0] __tmp_893_12;
  localparam _tmp_894 = 1;
  wire [_tmp_894-1:0] _tmp_895;
  assign _tmp_895 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_894-1:0] __tmp_895_1;
  reg [_tmp_894-1:0] __tmp_895_2;
  reg [_tmp_894-1:0] __tmp_895_3;
  reg [_tmp_894-1:0] __tmp_895_4;
  reg [_tmp_894-1:0] __tmp_895_5;
  reg [_tmp_894-1:0] __tmp_895_6;
  reg [_tmp_894-1:0] __tmp_895_7;
  reg [_tmp_894-1:0] __tmp_895_8;
  reg [_tmp_894-1:0] __tmp_895_9;
  reg [_tmp_894-1:0] __tmp_895_10;
  reg [_tmp_894-1:0] __tmp_895_11;
  reg [_tmp_894-1:0] __tmp_895_12;
  localparam _tmp_896 = 1;
  wire [_tmp_896-1:0] _tmp_897;
  assign _tmp_897 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_896-1:0] __tmp_897_1;
  reg [_tmp_896-1:0] __tmp_897_2;
  reg [_tmp_896-1:0] __tmp_897_3;
  reg [_tmp_896-1:0] __tmp_897_4;
  reg [_tmp_896-1:0] __tmp_897_5;
  reg [_tmp_896-1:0] __tmp_897_6;
  reg [_tmp_896-1:0] __tmp_897_7;
  reg [_tmp_896-1:0] __tmp_897_8;
  reg [_tmp_896-1:0] __tmp_897_9;
  reg [_tmp_896-1:0] __tmp_897_10;
  reg [_tmp_896-1:0] __tmp_897_11;
  reg [_tmp_896-1:0] __tmp_897_12;
  localparam _tmp_898 = 1;
  wire [_tmp_898-1:0] _tmp_899;
  assign _tmp_899 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_898-1:0] __tmp_899_1;
  reg [_tmp_898-1:0] __tmp_899_2;
  reg [_tmp_898-1:0] __tmp_899_3;
  reg [_tmp_898-1:0] __tmp_899_4;
  reg [_tmp_898-1:0] __tmp_899_5;
  reg [_tmp_898-1:0] __tmp_899_6;
  reg [_tmp_898-1:0] __tmp_899_7;
  reg [_tmp_898-1:0] __tmp_899_8;
  reg [_tmp_898-1:0] __tmp_899_9;
  localparam _tmp_900 = 1;
  wire [_tmp_900-1:0] _tmp_901;
  assign _tmp_901 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_900-1:0] __tmp_901_1;
  reg [_tmp_900-1:0] __tmp_901_2;
  reg [_tmp_900-1:0] __tmp_901_3;
  reg [_tmp_900-1:0] __tmp_901_4;
  reg [_tmp_900-1:0] __tmp_901_5;
  reg [_tmp_900-1:0] __tmp_901_6;
  reg [_tmp_900-1:0] __tmp_901_7;
  reg [_tmp_900-1:0] __tmp_901_8;
  reg [_tmp_900-1:0] __tmp_901_9;
  localparam _tmp_902 = 1;
  wire [_tmp_902-1:0] _tmp_903;
  assign _tmp_903 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_902-1:0] __tmp_903_1;
  reg [_tmp_902-1:0] __tmp_903_2;
  reg [_tmp_902-1:0] __tmp_903_3;
  reg [_tmp_902-1:0] __tmp_903_4;
  reg [_tmp_902-1:0] __tmp_903_5;
  reg [_tmp_902-1:0] __tmp_903_6;
  reg [_tmp_902-1:0] __tmp_903_7;
  reg [_tmp_902-1:0] __tmp_903_8;
  reg [_tmp_902-1:0] __tmp_903_9;
  reg [4-1:0] _mul_12_sink_wait_count;
  localparam _tmp_904 = 1;
  wire [_tmp_904-1:0] _tmp_905;
  assign _tmp_905 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_904-1:0] __tmp_905_1;
  reg [_tmp_904-1:0] __tmp_905_2;
  reg [_tmp_904-1:0] __tmp_905_3;
  reg [_tmp_904-1:0] __tmp_905_4;
  reg [_tmp_904-1:0] __tmp_905_5;
  reg [_tmp_904-1:0] __tmp_905_6;
  reg [_tmp_904-1:0] __tmp_905_7;
  reg [_tmp_904-1:0] __tmp_905_8;
  reg [_tmp_904-1:0] __tmp_905_9;
  reg [_tmp_904-1:0] __tmp_905_10;
  reg [_tmp_904-1:0] __tmp_905_11;
  reg [_tmp_904-1:0] __tmp_905_12;
  localparam _tmp_906 = 1;
  wire [_tmp_906-1:0] _tmp_907;
  assign _tmp_907 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_906-1:0] __tmp_907_1;
  reg [_tmp_906-1:0] __tmp_907_2;
  reg [_tmp_906-1:0] __tmp_907_3;
  reg [_tmp_906-1:0] __tmp_907_4;
  reg [_tmp_906-1:0] __tmp_907_5;
  reg [_tmp_906-1:0] __tmp_907_6;
  reg [_tmp_906-1:0] __tmp_907_7;
  reg [_tmp_906-1:0] __tmp_907_8;
  reg [_tmp_906-1:0] __tmp_907_9;
  reg [_tmp_906-1:0] __tmp_907_10;
  reg [_tmp_906-1:0] __tmp_907_11;
  reg [_tmp_906-1:0] __tmp_907_12;
  localparam _tmp_908 = 1;
  wire [_tmp_908-1:0] _tmp_909;
  assign _tmp_909 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_908-1:0] __tmp_909_1;
  reg [_tmp_908-1:0] __tmp_909_2;
  reg [_tmp_908-1:0] __tmp_909_3;
  reg [_tmp_908-1:0] __tmp_909_4;
  reg [_tmp_908-1:0] __tmp_909_5;
  reg [_tmp_908-1:0] __tmp_909_6;
  reg [_tmp_908-1:0] __tmp_909_7;
  reg [_tmp_908-1:0] __tmp_909_8;
  reg [_tmp_908-1:0] __tmp_909_9;
  reg [_tmp_908-1:0] __tmp_909_10;
  reg [_tmp_908-1:0] __tmp_909_11;
  reg [_tmp_908-1:0] __tmp_909_12;
  localparam _tmp_910 = 1;
  wire [_tmp_910-1:0] _tmp_911;
  assign _tmp_911 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_910-1:0] __tmp_911_1;
  reg [_tmp_910-1:0] __tmp_911_2;
  reg [_tmp_910-1:0] __tmp_911_3;
  reg [_tmp_910-1:0] __tmp_911_4;
  reg [_tmp_910-1:0] __tmp_911_5;
  reg [_tmp_910-1:0] __tmp_911_6;
  reg [_tmp_910-1:0] __tmp_911_7;
  reg [_tmp_910-1:0] __tmp_911_8;
  reg [_tmp_910-1:0] __tmp_911_9;
  reg [_tmp_910-1:0] __tmp_911_10;
  reg [_tmp_910-1:0] __tmp_911_11;
  reg [_tmp_910-1:0] __tmp_911_12;
  reg [_tmp_910-1:0] __tmp_911_13;
  reg [_tmp_910-1:0] __tmp_911_14;
  reg [_tmp_910-1:0] __tmp_911_15;
  reg [_tmp_910-1:0] __tmp_911_16;
  reg [_tmp_910-1:0] __tmp_911_17;
  reg [_tmp_910-1:0] __tmp_911_18;
  reg [_tmp_910-1:0] __tmp_911_19;
  localparam _tmp_912 = 1;
  wire [_tmp_912-1:0] _tmp_913;
  assign _tmp_913 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_912-1:0] __tmp_913_1;
  reg [_tmp_912-1:0] __tmp_913_2;
  reg [_tmp_912-1:0] __tmp_913_3;
  reg [_tmp_912-1:0] __tmp_913_4;
  reg [_tmp_912-1:0] __tmp_913_5;
  reg [_tmp_912-1:0] __tmp_913_6;
  reg [_tmp_912-1:0] __tmp_913_7;
  reg [_tmp_912-1:0] __tmp_913_8;
  reg [_tmp_912-1:0] __tmp_913_9;
  reg [_tmp_912-1:0] __tmp_913_10;
  reg [_tmp_912-1:0] __tmp_913_11;
  reg [_tmp_912-1:0] __tmp_913_12;
  reg [_tmp_912-1:0] __tmp_913_13;
  reg [_tmp_912-1:0] __tmp_913_14;
  reg [_tmp_912-1:0] __tmp_913_15;
  reg [_tmp_912-1:0] __tmp_913_16;
  reg [_tmp_912-1:0] __tmp_913_17;
  reg [_tmp_912-1:0] __tmp_913_18;
  reg [_tmp_912-1:0] __tmp_913_19;
  localparam _tmp_914 = 1;
  wire [_tmp_914-1:0] _tmp_915;
  assign _tmp_915 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_914-1:0] __tmp_915_1;
  reg [_tmp_914-1:0] __tmp_915_2;
  reg [_tmp_914-1:0] __tmp_915_3;
  reg [_tmp_914-1:0] __tmp_915_4;
  reg [_tmp_914-1:0] __tmp_915_5;
  reg [_tmp_914-1:0] __tmp_915_6;
  reg [_tmp_914-1:0] __tmp_915_7;
  reg [_tmp_914-1:0] __tmp_915_8;
  reg [_tmp_914-1:0] __tmp_915_9;
  reg [_tmp_914-1:0] __tmp_915_10;
  reg [_tmp_914-1:0] __tmp_915_11;
  reg [_tmp_914-1:0] __tmp_915_12;
  reg [_tmp_914-1:0] __tmp_915_13;
  reg [_tmp_914-1:0] __tmp_915_14;
  reg [_tmp_914-1:0] __tmp_915_15;
  reg [_tmp_914-1:0] __tmp_915_16;
  reg [_tmp_914-1:0] __tmp_915_17;
  reg [_tmp_914-1:0] __tmp_915_18;
  reg [_tmp_914-1:0] __tmp_915_19;
  localparam _tmp_916 = 1;
  wire [_tmp_916-1:0] _tmp_917;
  assign _tmp_917 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_916-1:0] __tmp_917_1;
  reg [_tmp_916-1:0] __tmp_917_2;
  reg [_tmp_916-1:0] __tmp_917_3;
  reg [_tmp_916-1:0] __tmp_917_4;
  reg [_tmp_916-1:0] __tmp_917_5;
  reg [_tmp_916-1:0] __tmp_917_6;
  reg [_tmp_916-1:0] __tmp_917_7;
  reg [_tmp_916-1:0] __tmp_917_8;
  reg [_tmp_916-1:0] __tmp_917_9;
  reg [_tmp_916-1:0] __tmp_917_10;
  reg [_tmp_916-1:0] __tmp_917_11;
  reg [_tmp_916-1:0] __tmp_917_12;
  reg [_tmp_916-1:0] __tmp_917_13;
  reg [_tmp_916-1:0] __tmp_917_14;
  reg [_tmp_916-1:0] __tmp_917_15;
  reg [_tmp_916-1:0] __tmp_917_16;
  reg [_tmp_916-1:0] __tmp_917_17;
  reg [_tmp_916-1:0] __tmp_917_18;
  reg [_tmp_916-1:0] __tmp_917_19;
  localparam _tmp_918 = 1;
  wire [_tmp_918-1:0] _tmp_919;
  assign _tmp_919 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_918-1:0] __tmp_919_1;
  reg [_tmp_918-1:0] __tmp_919_2;
  reg [_tmp_918-1:0] __tmp_919_3;
  reg [_tmp_918-1:0] __tmp_919_4;
  reg [_tmp_918-1:0] __tmp_919_5;
  reg [_tmp_918-1:0] __tmp_919_6;
  reg [_tmp_918-1:0] __tmp_919_7;
  reg [_tmp_918-1:0] __tmp_919_8;
  reg [_tmp_918-1:0] __tmp_919_9;
  reg [_tmp_918-1:0] __tmp_919_10;
  reg [_tmp_918-1:0] __tmp_919_11;
  reg [_tmp_918-1:0] __tmp_919_12;
  reg [_tmp_918-1:0] __tmp_919_13;
  reg [_tmp_918-1:0] __tmp_919_14;
  reg [_tmp_918-1:0] __tmp_919_15;
  reg [_tmp_918-1:0] __tmp_919_16;
  reg [_tmp_918-1:0] __tmp_919_17;
  reg [_tmp_918-1:0] __tmp_919_18;
  reg [_tmp_918-1:0] __tmp_919_19;
  localparam _tmp_920 = 1;
  wire [_tmp_920-1:0] _tmp_921;
  assign _tmp_921 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_920-1:0] __tmp_921_1;
  reg [_tmp_920-1:0] __tmp_921_2;
  reg [_tmp_920-1:0] __tmp_921_3;
  reg [_tmp_920-1:0] __tmp_921_4;
  reg [_tmp_920-1:0] __tmp_921_5;
  reg [_tmp_920-1:0] __tmp_921_6;
  reg [_tmp_920-1:0] __tmp_921_7;
  reg [_tmp_920-1:0] __tmp_921_8;
  reg [_tmp_920-1:0] __tmp_921_9;
  reg [_tmp_920-1:0] __tmp_921_10;
  reg [_tmp_920-1:0] __tmp_921_11;
  reg [_tmp_920-1:0] __tmp_921_12;
  reg [_tmp_920-1:0] __tmp_921_13;
  reg [_tmp_920-1:0] __tmp_921_14;
  reg [_tmp_920-1:0] __tmp_921_15;
  reg [_tmp_920-1:0] __tmp_921_16;
  reg [_tmp_920-1:0] __tmp_921_17;
  reg [_tmp_920-1:0] __tmp_921_18;
  reg [_tmp_920-1:0] __tmp_921_19;
  localparam _tmp_922 = 1;
  wire [_tmp_922-1:0] _tmp_923;
  assign _tmp_923 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_922-1:0] __tmp_923_1;
  reg [_tmp_922-1:0] __tmp_923_2;
  reg [_tmp_922-1:0] __tmp_923_3;
  reg [_tmp_922-1:0] __tmp_923_4;
  reg [_tmp_922-1:0] __tmp_923_5;
  reg [_tmp_922-1:0] __tmp_923_6;
  reg [_tmp_922-1:0] __tmp_923_7;
  reg [_tmp_922-1:0] __tmp_923_8;
  reg [_tmp_922-1:0] __tmp_923_9;
  reg [_tmp_922-1:0] __tmp_923_10;
  reg [_tmp_922-1:0] __tmp_923_11;
  reg [_tmp_922-1:0] __tmp_923_12;
  reg [_tmp_922-1:0] __tmp_923_13;
  reg [_tmp_922-1:0] __tmp_923_14;
  reg [_tmp_922-1:0] __tmp_923_15;
  reg [_tmp_922-1:0] __tmp_923_16;
  reg [_tmp_922-1:0] __tmp_923_17;
  reg [_tmp_922-1:0] __tmp_923_18;
  reg [_tmp_922-1:0] __tmp_923_19;
  localparam _tmp_924 = 1;
  wire [_tmp_924-1:0] _tmp_925;
  assign _tmp_925 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_924-1:0] __tmp_925_1;
  reg [_tmp_924-1:0] __tmp_925_2;
  reg [_tmp_924-1:0] __tmp_925_3;
  reg [_tmp_924-1:0] __tmp_925_4;
  reg [_tmp_924-1:0] __tmp_925_5;
  reg [_tmp_924-1:0] __tmp_925_6;
  reg [_tmp_924-1:0] __tmp_925_7;
  reg [_tmp_924-1:0] __tmp_925_8;
  reg [_tmp_924-1:0] __tmp_925_9;
  reg [_tmp_924-1:0] __tmp_925_10;
  reg [_tmp_924-1:0] __tmp_925_11;
  reg [_tmp_924-1:0] __tmp_925_12;
  reg [_tmp_924-1:0] __tmp_925_13;
  reg [_tmp_924-1:0] __tmp_925_14;
  reg [_tmp_924-1:0] __tmp_925_15;
  reg [_tmp_924-1:0] __tmp_925_16;
  reg [_tmp_924-1:0] __tmp_925_17;
  reg [_tmp_924-1:0] __tmp_925_18;
  reg [_tmp_924-1:0] __tmp_925_19;
  localparam _tmp_926 = 1;
  wire [_tmp_926-1:0] _tmp_927;
  assign _tmp_927 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_926-1:0] __tmp_927_1;
  reg [_tmp_926-1:0] __tmp_927_2;
  reg [_tmp_926-1:0] __tmp_927_3;
  reg [_tmp_926-1:0] __tmp_927_4;
  reg [_tmp_926-1:0] __tmp_927_5;
  reg [_tmp_926-1:0] __tmp_927_6;
  reg [_tmp_926-1:0] __tmp_927_7;
  reg [_tmp_926-1:0] __tmp_927_8;
  reg [_tmp_926-1:0] __tmp_927_9;
  reg [_tmp_926-1:0] __tmp_927_10;
  reg [_tmp_926-1:0] __tmp_927_11;
  reg [_tmp_926-1:0] __tmp_927_12;
  reg [_tmp_926-1:0] __tmp_927_13;
  reg [_tmp_926-1:0] __tmp_927_14;
  reg [_tmp_926-1:0] __tmp_927_15;
  reg [_tmp_926-1:0] __tmp_927_16;
  reg [_tmp_926-1:0] __tmp_927_17;
  reg [_tmp_926-1:0] __tmp_927_18;
  reg [_tmp_926-1:0] __tmp_927_19;
  reg [3-1:0] _add_tree_2_sink_wait_count;
  localparam _tmp_928 = 1;
  wire [_tmp_928-1:0] _tmp_929;
  assign _tmp_929 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_928-1:0] __tmp_929_1;
  reg [_tmp_928-1:0] __tmp_929_2;
  reg [_tmp_928-1:0] __tmp_929_3;
  reg [_tmp_928-1:0] __tmp_929_4;
  reg [_tmp_928-1:0] __tmp_929_5;
  reg [_tmp_928-1:0] __tmp_929_6;
  localparam _tmp_930 = 1;
  wire [_tmp_930-1:0] _tmp_931;
  assign _tmp_931 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_930-1:0] __tmp_931_1;
  reg [_tmp_930-1:0] __tmp_931_2;
  reg [_tmp_930-1:0] __tmp_931_3;
  reg [_tmp_930-1:0] __tmp_931_4;
  reg [_tmp_930-1:0] __tmp_931_5;
  reg [_tmp_930-1:0] __tmp_931_6;
  localparam _tmp_932 = 1;
  wire [_tmp_932-1:0] _tmp_933;
  assign _tmp_933 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_932-1:0] __tmp_933_1;
  reg [_tmp_932-1:0] __tmp_933_2;
  reg [_tmp_932-1:0] __tmp_933_3;
  reg [_tmp_932-1:0] __tmp_933_4;
  reg [_tmp_932-1:0] __tmp_933_5;
  reg [_tmp_932-1:0] __tmp_933_6;
  localparam _tmp_934 = 1;
  wire [_tmp_934-1:0] _tmp_935;
  assign _tmp_935 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_934-1:0] __tmp_935_1;
  reg [_tmp_934-1:0] __tmp_935_2;
  reg [_tmp_934-1:0] __tmp_935_3;
  reg [_tmp_934-1:0] __tmp_935_4;
  reg [_tmp_934-1:0] __tmp_935_5;
  reg [_tmp_934-1:0] __tmp_935_6;
  reg [_tmp_934-1:0] __tmp_935_7;
  reg [_tmp_934-1:0] __tmp_935_8;
  reg [_tmp_934-1:0] __tmp_935_9;
  reg [_tmp_934-1:0] __tmp_935_10;
  reg [_tmp_934-1:0] __tmp_935_11;
  reg [_tmp_934-1:0] __tmp_935_12;
  reg [_tmp_934-1:0] __tmp_935_13;
  reg [_tmp_934-1:0] __tmp_935_14;
  reg [_tmp_934-1:0] __tmp_935_15;
  reg [_tmp_934-1:0] __tmp_935_16;
  reg [_tmp_934-1:0] __tmp_935_17;
  reg [_tmp_934-1:0] __tmp_935_18;
  reg [_tmp_934-1:0] __tmp_935_19;
  reg [_tmp_934-1:0] __tmp_935_20;
  reg [_tmp_934-1:0] __tmp_935_21;
  reg [_tmp_934-1:0] __tmp_935_22;
  reg [_tmp_934-1:0] __tmp_935_23;
  reg [_tmp_934-1:0] __tmp_935_24;
  localparam _tmp_936 = 1;
  wire [_tmp_936-1:0] _tmp_937;
  assign _tmp_937 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_936-1:0] __tmp_937_1;
  reg [_tmp_936-1:0] __tmp_937_2;
  reg [_tmp_936-1:0] __tmp_937_3;
  reg [_tmp_936-1:0] __tmp_937_4;
  reg [_tmp_936-1:0] __tmp_937_5;
  reg [_tmp_936-1:0] __tmp_937_6;
  reg [_tmp_936-1:0] __tmp_937_7;
  reg [_tmp_936-1:0] __tmp_937_8;
  reg [_tmp_936-1:0] __tmp_937_9;
  reg [_tmp_936-1:0] __tmp_937_10;
  reg [_tmp_936-1:0] __tmp_937_11;
  reg [_tmp_936-1:0] __tmp_937_12;
  reg [_tmp_936-1:0] __tmp_937_13;
  reg [_tmp_936-1:0] __tmp_937_14;
  reg [_tmp_936-1:0] __tmp_937_15;
  reg [_tmp_936-1:0] __tmp_937_16;
  reg [_tmp_936-1:0] __tmp_937_17;
  reg [_tmp_936-1:0] __tmp_937_18;
  reg [_tmp_936-1:0] __tmp_937_19;
  reg [_tmp_936-1:0] __tmp_937_20;
  reg [_tmp_936-1:0] __tmp_937_21;
  reg [_tmp_936-1:0] __tmp_937_22;
  reg [_tmp_936-1:0] __tmp_937_23;
  localparam _tmp_938 = 1;
  wire [_tmp_938-1:0] _tmp_939;
  assign _tmp_939 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_938-1:0] __tmp_939_1;
  reg [_tmp_938-1:0] __tmp_939_2;
  reg [_tmp_938-1:0] __tmp_939_3;
  reg [_tmp_938-1:0] __tmp_939_4;
  reg [_tmp_938-1:0] __tmp_939_5;
  reg [_tmp_938-1:0] __tmp_939_6;
  reg [_tmp_938-1:0] __tmp_939_7;
  reg [_tmp_938-1:0] __tmp_939_8;
  reg [_tmp_938-1:0] __tmp_939_9;
  reg [_tmp_938-1:0] __tmp_939_10;
  reg [_tmp_938-1:0] __tmp_939_11;
  reg [_tmp_938-1:0] __tmp_939_12;
  reg [_tmp_938-1:0] __tmp_939_13;
  reg [_tmp_938-1:0] __tmp_939_14;
  reg [_tmp_938-1:0] __tmp_939_15;
  reg [_tmp_938-1:0] __tmp_939_16;
  reg [_tmp_938-1:0] __tmp_939_17;
  reg [_tmp_938-1:0] __tmp_939_18;
  reg [_tmp_938-1:0] __tmp_939_19;
  reg [_tmp_938-1:0] __tmp_939_20;
  reg [_tmp_938-1:0] __tmp_939_21;
  reg [_tmp_938-1:0] __tmp_939_22;
  reg [_tmp_938-1:0] __tmp_939_23;
  localparam _tmp_940 = 1;
  wire [_tmp_940-1:0] _tmp_941;
  assign _tmp_941 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_940-1:0] __tmp_941_1;
  reg [_tmp_940-1:0] __tmp_941_2;
  reg [_tmp_940-1:0] __tmp_941_3;
  reg [_tmp_940-1:0] __tmp_941_4;
  reg [_tmp_940-1:0] __tmp_941_5;
  reg [_tmp_940-1:0] __tmp_941_6;
  reg [_tmp_940-1:0] __tmp_941_7;
  reg [_tmp_940-1:0] __tmp_941_8;
  reg [_tmp_940-1:0] __tmp_941_9;
  reg [_tmp_940-1:0] __tmp_941_10;
  reg [_tmp_940-1:0] __tmp_941_11;
  reg [_tmp_940-1:0] __tmp_941_12;
  reg [_tmp_940-1:0] __tmp_941_13;
  reg [_tmp_940-1:0] __tmp_941_14;
  reg [_tmp_940-1:0] __tmp_941_15;
  reg [_tmp_940-1:0] __tmp_941_16;
  reg [_tmp_940-1:0] __tmp_941_17;
  reg [_tmp_940-1:0] __tmp_941_18;
  reg [_tmp_940-1:0] __tmp_941_19;
  reg [_tmp_940-1:0] __tmp_941_20;
  reg [_tmp_940-1:0] __tmp_941_21;
  reg [_tmp_940-1:0] __tmp_941_22;
  reg [_tmp_940-1:0] __tmp_941_23;
  reg [4-1:0] _acc_0_sink_wait_count;
  localparam _tmp_942 = 1;
  wire [_tmp_942-1:0] _tmp_943;
  assign _tmp_943 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_942-1:0] __tmp_943_1;
  reg [_tmp_942-1:0] __tmp_943_2;
  reg [_tmp_942-1:0] __tmp_943_3;
  reg [_tmp_942-1:0] __tmp_943_4;
  reg [_tmp_942-1:0] __tmp_943_5;
  reg [_tmp_942-1:0] __tmp_943_6;
  reg [_tmp_942-1:0] __tmp_943_7;
  reg [_tmp_942-1:0] __tmp_943_8;
  reg [_tmp_942-1:0] __tmp_943_9;
  localparam _tmp_944 = 1;
  wire [_tmp_944-1:0] _tmp_945;
  assign _tmp_945 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_944-1:0] __tmp_945_1;
  reg [_tmp_944-1:0] __tmp_945_2;
  reg [_tmp_944-1:0] __tmp_945_3;
  reg [_tmp_944-1:0] __tmp_945_4;
  reg [_tmp_944-1:0] __tmp_945_5;
  reg [_tmp_944-1:0] __tmp_945_6;
  reg [_tmp_944-1:0] __tmp_945_7;
  reg [_tmp_944-1:0] __tmp_945_8;
  reg [_tmp_944-1:0] __tmp_945_9;
  localparam _tmp_946 = 1;
  wire [_tmp_946-1:0] _tmp_947;
  assign _tmp_947 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_946-1:0] __tmp_947_1;
  reg [_tmp_946-1:0] __tmp_947_2;
  reg [_tmp_946-1:0] __tmp_947_3;
  reg [_tmp_946-1:0] __tmp_947_4;
  reg [_tmp_946-1:0] __tmp_947_5;
  reg [_tmp_946-1:0] __tmp_947_6;
  reg [_tmp_946-1:0] __tmp_947_7;
  reg [_tmp_946-1:0] __tmp_947_8;
  reg [_tmp_946-1:0] __tmp_947_9;
  localparam _tmp_948 = 1;
  wire [_tmp_948-1:0] _tmp_949;
  assign _tmp_949 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_948-1:0] __tmp_949_1;
  reg [_tmp_948-1:0] __tmp_949_2;
  reg [_tmp_948-1:0] __tmp_949_3;
  reg [_tmp_948-1:0] __tmp_949_4;
  reg [_tmp_948-1:0] __tmp_949_5;
  reg [_tmp_948-1:0] __tmp_949_6;
  reg [_tmp_948-1:0] __tmp_949_7;
  reg [_tmp_948-1:0] __tmp_949_8;
  reg [_tmp_948-1:0] __tmp_949_9;
  reg [_tmp_948-1:0] __tmp_949_10;
  reg [_tmp_948-1:0] __tmp_949_11;
  reg [_tmp_948-1:0] __tmp_949_12;
  reg [_tmp_948-1:0] __tmp_949_13;
  reg [_tmp_948-1:0] __tmp_949_14;
  reg [_tmp_948-1:0] __tmp_949_15;
  reg [_tmp_948-1:0] __tmp_949_16;
  reg [_tmp_948-1:0] __tmp_949_17;
  reg [_tmp_948-1:0] __tmp_949_18;
  reg [_tmp_948-1:0] __tmp_949_19;
  reg [_tmp_948-1:0] __tmp_949_20;
  reg [_tmp_948-1:0] __tmp_949_21;
  reg [_tmp_948-1:0] __tmp_949_22;
  reg [_tmp_948-1:0] __tmp_949_23;
  reg [_tmp_948-1:0] __tmp_949_24;
  reg [_tmp_948-1:0] __tmp_949_25;
  reg [_tmp_948-1:0] __tmp_949_26;
  reg [_tmp_948-1:0] __tmp_949_27;
  reg [_tmp_948-1:0] __tmp_949_28;
  reg [_tmp_948-1:0] __tmp_949_29;
  reg [_tmp_948-1:0] __tmp_949_30;
  reg [_tmp_948-1:0] __tmp_949_31;
  localparam _tmp_950 = 1;
  wire [_tmp_950-1:0] _tmp_951;
  assign _tmp_951 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_950-1:0] __tmp_951_1;
  reg [_tmp_950-1:0] __tmp_951_2;
  reg [_tmp_950-1:0] __tmp_951_3;
  reg [_tmp_950-1:0] __tmp_951_4;
  reg [_tmp_950-1:0] __tmp_951_5;
  reg [_tmp_950-1:0] __tmp_951_6;
  reg [_tmp_950-1:0] __tmp_951_7;
  reg [_tmp_950-1:0] __tmp_951_8;
  reg [_tmp_950-1:0] __tmp_951_9;
  reg [_tmp_950-1:0] __tmp_951_10;
  reg [_tmp_950-1:0] __tmp_951_11;
  reg [_tmp_950-1:0] __tmp_951_12;
  reg [_tmp_950-1:0] __tmp_951_13;
  reg [_tmp_950-1:0] __tmp_951_14;
  reg [_tmp_950-1:0] __tmp_951_15;
  reg [_tmp_950-1:0] __tmp_951_16;
  reg [_tmp_950-1:0] __tmp_951_17;
  reg [_tmp_950-1:0] __tmp_951_18;
  reg [_tmp_950-1:0] __tmp_951_19;
  reg [_tmp_950-1:0] __tmp_951_20;
  reg [_tmp_950-1:0] __tmp_951_21;
  reg [_tmp_950-1:0] __tmp_951_22;
  reg [_tmp_950-1:0] __tmp_951_23;
  reg [_tmp_950-1:0] __tmp_951_24;
  reg [_tmp_950-1:0] __tmp_951_25;
  reg [_tmp_950-1:0] __tmp_951_26;
  reg [_tmp_950-1:0] __tmp_951_27;
  reg [_tmp_950-1:0] __tmp_951_28;
  reg [_tmp_950-1:0] __tmp_951_29;
  reg [_tmp_950-1:0] __tmp_951_30;
  reg [_tmp_950-1:0] __tmp_951_31;
  localparam _tmp_952 = 1;
  wire [_tmp_952-1:0] _tmp_953;
  assign _tmp_953 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_952-1:0] __tmp_953_1;
  reg [_tmp_952-1:0] __tmp_953_2;
  reg [_tmp_952-1:0] __tmp_953_3;
  reg [_tmp_952-1:0] __tmp_953_4;
  reg [_tmp_952-1:0] __tmp_953_5;
  reg [_tmp_952-1:0] __tmp_953_6;
  reg [_tmp_952-1:0] __tmp_953_7;
  reg [_tmp_952-1:0] __tmp_953_8;
  reg [_tmp_952-1:0] __tmp_953_9;
  reg [_tmp_952-1:0] __tmp_953_10;
  reg [_tmp_952-1:0] __tmp_953_11;
  reg [_tmp_952-1:0] __tmp_953_12;
  reg [_tmp_952-1:0] __tmp_953_13;
  reg [_tmp_952-1:0] __tmp_953_14;
  reg [_tmp_952-1:0] __tmp_953_15;
  reg [_tmp_952-1:0] __tmp_953_16;
  reg [_tmp_952-1:0] __tmp_953_17;
  reg [_tmp_952-1:0] __tmp_953_18;
  reg [_tmp_952-1:0] __tmp_953_19;
  reg [_tmp_952-1:0] __tmp_953_20;
  reg [_tmp_952-1:0] __tmp_953_21;
  reg [_tmp_952-1:0] __tmp_953_22;
  reg [_tmp_952-1:0] __tmp_953_23;
  reg [_tmp_952-1:0] __tmp_953_24;
  reg [_tmp_952-1:0] __tmp_953_25;
  reg [_tmp_952-1:0] __tmp_953_26;
  reg [_tmp_952-1:0] __tmp_953_27;
  reg [_tmp_952-1:0] __tmp_953_28;
  reg [_tmp_952-1:0] __tmp_953_29;
  reg [_tmp_952-1:0] __tmp_953_30;
  reg [_tmp_952-1:0] __tmp_953_31;
  reg [4-1:0] _mul_rshift_clip_3_sink_wait_count;
  localparam _tmp_954 = 1;
  wire [_tmp_954-1:0] _tmp_955;
  assign _tmp_955 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_954-1:0] __tmp_955_1;
  reg [_tmp_954-1:0] __tmp_955_2;
  reg [_tmp_954-1:0] __tmp_955_3;
  reg [_tmp_954-1:0] __tmp_955_4;
  reg [_tmp_954-1:0] __tmp_955_5;
  reg [_tmp_954-1:0] __tmp_955_6;
  reg [_tmp_954-1:0] __tmp_955_7;
  reg [_tmp_954-1:0] __tmp_955_8;
  reg [_tmp_954-1:0] __tmp_955_9;
  reg [_tmp_954-1:0] __tmp_955_10;
  reg [_tmp_954-1:0] __tmp_955_11;
  reg [_tmp_954-1:0] __tmp_955_12;
  localparam _tmp_956 = 1;
  wire [_tmp_956-1:0] _tmp_957;
  assign _tmp_957 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_956-1:0] __tmp_957_1;
  reg [_tmp_956-1:0] __tmp_957_2;
  reg [_tmp_956-1:0] __tmp_957_3;
  reg [_tmp_956-1:0] __tmp_957_4;
  reg [_tmp_956-1:0] __tmp_957_5;
  reg [_tmp_956-1:0] __tmp_957_6;
  reg [_tmp_956-1:0] __tmp_957_7;
  reg [_tmp_956-1:0] __tmp_957_8;
  reg [_tmp_956-1:0] __tmp_957_9;
  reg [_tmp_956-1:0] __tmp_957_10;
  reg [_tmp_956-1:0] __tmp_957_11;
  reg [_tmp_956-1:0] __tmp_957_12;
  localparam _tmp_958 = 1;
  wire [_tmp_958-1:0] _tmp_959;
  assign _tmp_959 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_958-1:0] __tmp_959_1;
  reg [_tmp_958-1:0] __tmp_959_2;
  reg [_tmp_958-1:0] __tmp_959_3;
  reg [_tmp_958-1:0] __tmp_959_4;
  reg [_tmp_958-1:0] __tmp_959_5;
  reg [_tmp_958-1:0] __tmp_959_6;
  reg [_tmp_958-1:0] __tmp_959_7;
  reg [_tmp_958-1:0] __tmp_959_8;
  reg [_tmp_958-1:0] __tmp_959_9;
  reg [_tmp_958-1:0] __tmp_959_10;
  reg [_tmp_958-1:0] __tmp_959_11;
  reg [_tmp_958-1:0] __tmp_959_12;
  reg [6-1:0] _stream_conv2d_16_sink_wait_count;
  localparam _tmp_960 = 1;
  wire [_tmp_960-1:0] _tmp_961;
  assign _tmp_961 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_960-1:0] __tmp_961_1;
  reg [_tmp_960-1:0] __tmp_961_2;
  reg [_tmp_960-1:0] __tmp_961_3;
  reg [_tmp_960-1:0] __tmp_961_4;
  reg [_tmp_960-1:0] __tmp_961_5;
  reg [_tmp_960-1:0] __tmp_961_6;
  reg [_tmp_960-1:0] __tmp_961_7;
  reg [_tmp_960-1:0] __tmp_961_8;
  reg [_tmp_960-1:0] __tmp_961_9;
  reg [_tmp_960-1:0] __tmp_961_10;
  reg [_tmp_960-1:0] __tmp_961_11;
  reg [_tmp_960-1:0] __tmp_961_12;
  reg [_tmp_960-1:0] __tmp_961_13;
  reg [_tmp_960-1:0] __tmp_961_14;
  reg [_tmp_960-1:0] __tmp_961_15;
  reg [_tmp_960-1:0] __tmp_961_16;
  reg [_tmp_960-1:0] __tmp_961_17;
  reg [_tmp_960-1:0] __tmp_961_18;
  reg [_tmp_960-1:0] __tmp_961_19;
  reg [_tmp_960-1:0] __tmp_961_20;
  reg [_tmp_960-1:0] __tmp_961_21;
  reg [_tmp_960-1:0] __tmp_961_22;
  reg [_tmp_960-1:0] __tmp_961_23;
  reg [_tmp_960-1:0] __tmp_961_24;
  reg [_tmp_960-1:0] __tmp_961_25;
  reg [_tmp_960-1:0] __tmp_961_26;
  reg [_tmp_960-1:0] __tmp_961_27;
  reg [_tmp_960-1:0] __tmp_961_28;
  reg [_tmp_960-1:0] __tmp_961_29;
  reg [_tmp_960-1:0] __tmp_961_30;
  reg [_tmp_960-1:0] __tmp_961_31;
  reg [_tmp_960-1:0] __tmp_961_32;
  reg [_tmp_960-1:0] __tmp_961_33;
  reg [_tmp_960-1:0] __tmp_961_34;
  reg [_tmp_960-1:0] __tmp_961_35;
  reg [_tmp_960-1:0] __tmp_961_36;
  reg [_tmp_960-1:0] __tmp_961_37;
  reg [_tmp_960-1:0] __tmp_961_38;
  reg [_tmp_960-1:0] __tmp_961_39;
  reg [_tmp_960-1:0] __tmp_961_40;
  reg [_tmp_960-1:0] __tmp_961_41;
  reg [_tmp_960-1:0] __tmp_961_42;
  reg [_tmp_960-1:0] __tmp_961_43;
  reg [_tmp_960-1:0] __tmp_961_44;
  reg [_tmp_960-1:0] __tmp_961_45;
  reg [_tmp_960-1:0] __tmp_961_46;
  localparam _tmp_962 = 1;
  wire [_tmp_962-1:0] _tmp_963;
  assign _tmp_963 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_962-1:0] __tmp_963_1;
  reg [_tmp_962-1:0] __tmp_963_2;
  reg [_tmp_962-1:0] __tmp_963_3;
  reg [_tmp_962-1:0] __tmp_963_4;
  reg [_tmp_962-1:0] __tmp_963_5;
  reg [_tmp_962-1:0] __tmp_963_6;
  reg [_tmp_962-1:0] __tmp_963_7;
  reg [_tmp_962-1:0] __tmp_963_8;
  reg [_tmp_962-1:0] __tmp_963_9;
  reg [_tmp_962-1:0] __tmp_963_10;
  reg [_tmp_962-1:0] __tmp_963_11;
  reg [_tmp_962-1:0] __tmp_963_12;
  reg [_tmp_962-1:0] __tmp_963_13;
  reg [_tmp_962-1:0] __tmp_963_14;
  reg [_tmp_962-1:0] __tmp_963_15;
  reg [_tmp_962-1:0] __tmp_963_16;
  reg [_tmp_962-1:0] __tmp_963_17;
  reg [_tmp_962-1:0] __tmp_963_18;
  reg [_tmp_962-1:0] __tmp_963_19;
  reg [_tmp_962-1:0] __tmp_963_20;
  reg [_tmp_962-1:0] __tmp_963_21;
  reg [_tmp_962-1:0] __tmp_963_22;
  reg [_tmp_962-1:0] __tmp_963_23;
  reg [_tmp_962-1:0] __tmp_963_24;
  reg [_tmp_962-1:0] __tmp_963_25;
  reg [_tmp_962-1:0] __tmp_963_26;
  reg [_tmp_962-1:0] __tmp_963_27;
  reg [_tmp_962-1:0] __tmp_963_28;
  reg [_tmp_962-1:0] __tmp_963_29;
  reg [_tmp_962-1:0] __tmp_963_30;
  reg [_tmp_962-1:0] __tmp_963_31;
  reg [_tmp_962-1:0] __tmp_963_32;
  reg [_tmp_962-1:0] __tmp_963_33;
  reg [_tmp_962-1:0] __tmp_963_34;
  reg [_tmp_962-1:0] __tmp_963_35;
  reg [_tmp_962-1:0] __tmp_963_36;
  reg [_tmp_962-1:0] __tmp_963_37;
  reg [_tmp_962-1:0] __tmp_963_38;
  reg [_tmp_962-1:0] __tmp_963_39;
  reg [_tmp_962-1:0] __tmp_963_40;
  reg [_tmp_962-1:0] __tmp_963_41;
  reg [_tmp_962-1:0] __tmp_963_42;
  reg [_tmp_962-1:0] __tmp_963_43;
  reg [_tmp_962-1:0] __tmp_963_44;
  reg [_tmp_962-1:0] __tmp_963_45;
  reg [_tmp_962-1:0] __tmp_963_46;
  localparam _tmp_964 = 1;
  wire [_tmp_964-1:0] _tmp_965;
  assign _tmp_965 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_964-1:0] __tmp_965_1;
  reg [_tmp_964-1:0] __tmp_965_2;
  reg [_tmp_964-1:0] __tmp_965_3;
  reg [_tmp_964-1:0] __tmp_965_4;
  reg [_tmp_964-1:0] __tmp_965_5;
  reg [_tmp_964-1:0] __tmp_965_6;
  reg [_tmp_964-1:0] __tmp_965_7;
  reg [_tmp_964-1:0] __tmp_965_8;
  reg [_tmp_964-1:0] __tmp_965_9;
  reg [_tmp_964-1:0] __tmp_965_10;
  reg [_tmp_964-1:0] __tmp_965_11;
  reg [_tmp_964-1:0] __tmp_965_12;
  reg [_tmp_964-1:0] __tmp_965_13;
  reg [_tmp_964-1:0] __tmp_965_14;
  reg [_tmp_964-1:0] __tmp_965_15;
  reg [_tmp_964-1:0] __tmp_965_16;
  reg [_tmp_964-1:0] __tmp_965_17;
  reg [_tmp_964-1:0] __tmp_965_18;
  reg [_tmp_964-1:0] __tmp_965_19;
  reg [_tmp_964-1:0] __tmp_965_20;
  reg [_tmp_964-1:0] __tmp_965_21;
  reg [_tmp_964-1:0] __tmp_965_22;
  reg [_tmp_964-1:0] __tmp_965_23;
  reg [_tmp_964-1:0] __tmp_965_24;
  reg [_tmp_964-1:0] __tmp_965_25;
  reg [_tmp_964-1:0] __tmp_965_26;
  reg [_tmp_964-1:0] __tmp_965_27;
  reg [_tmp_964-1:0] __tmp_965_28;
  reg [_tmp_964-1:0] __tmp_965_29;
  reg [_tmp_964-1:0] __tmp_965_30;
  reg [_tmp_964-1:0] __tmp_965_31;
  reg [_tmp_964-1:0] __tmp_965_32;
  reg [_tmp_964-1:0] __tmp_965_33;
  reg [_tmp_964-1:0] __tmp_965_34;
  reg [_tmp_964-1:0] __tmp_965_35;
  reg [_tmp_964-1:0] __tmp_965_36;
  reg [_tmp_964-1:0] __tmp_965_37;
  reg [_tmp_964-1:0] __tmp_965_38;
  reg [_tmp_964-1:0] __tmp_965_39;
  reg [_tmp_964-1:0] __tmp_965_40;
  reg [_tmp_964-1:0] __tmp_965_41;
  reg [_tmp_964-1:0] __tmp_965_42;
  reg [_tmp_964-1:0] __tmp_965_43;
  reg [_tmp_964-1:0] __tmp_965_44;
  reg [_tmp_964-1:0] __tmp_965_45;
  reg [_tmp_964-1:0] __tmp_965_46;
  localparam _tmp_966 = 1;
  wire [_tmp_966-1:0] _tmp_967;
  assign _tmp_967 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_966-1:0] __tmp_967_1;
  reg [_tmp_966-1:0] __tmp_967_2;
  reg [_tmp_966-1:0] __tmp_967_3;
  reg [_tmp_966-1:0] __tmp_967_4;
  reg [_tmp_966-1:0] __tmp_967_5;
  reg [_tmp_966-1:0] __tmp_967_6;
  reg [_tmp_966-1:0] __tmp_967_7;
  reg [_tmp_966-1:0] __tmp_967_8;
  reg [_tmp_966-1:0] __tmp_967_9;
  reg [_tmp_966-1:0] __tmp_967_10;
  reg [_tmp_966-1:0] __tmp_967_11;
  reg [_tmp_966-1:0] __tmp_967_12;
  reg [_tmp_966-1:0] __tmp_967_13;
  reg [_tmp_966-1:0] __tmp_967_14;
  reg [_tmp_966-1:0] __tmp_967_15;
  reg [_tmp_966-1:0] __tmp_967_16;
  reg [_tmp_966-1:0] __tmp_967_17;
  reg [_tmp_966-1:0] __tmp_967_18;
  reg [_tmp_966-1:0] __tmp_967_19;
  reg [_tmp_966-1:0] __tmp_967_20;
  reg [_tmp_966-1:0] __tmp_967_21;
  reg [_tmp_966-1:0] __tmp_967_22;
  reg [_tmp_966-1:0] __tmp_967_23;
  reg [_tmp_966-1:0] __tmp_967_24;
  reg [_tmp_966-1:0] __tmp_967_25;
  reg [_tmp_966-1:0] __tmp_967_26;
  reg [_tmp_966-1:0] __tmp_967_27;
  reg [_tmp_966-1:0] __tmp_967_28;
  reg [_tmp_966-1:0] __tmp_967_29;
  reg [_tmp_966-1:0] __tmp_967_30;
  reg [_tmp_966-1:0] __tmp_967_31;
  reg [_tmp_966-1:0] __tmp_967_32;
  reg [_tmp_966-1:0] __tmp_967_33;
  reg [_tmp_966-1:0] __tmp_967_34;
  reg [_tmp_966-1:0] __tmp_967_35;
  reg [_tmp_966-1:0] __tmp_967_36;
  reg [_tmp_966-1:0] __tmp_967_37;
  reg [_tmp_966-1:0] __tmp_967_38;
  reg [_tmp_966-1:0] __tmp_967_39;
  reg [_tmp_966-1:0] __tmp_967_40;
  reg [_tmp_966-1:0] __tmp_967_41;
  reg [_tmp_966-1:0] __tmp_967_42;
  reg [_tmp_966-1:0] __tmp_967_43;
  reg [_tmp_966-1:0] __tmp_967_44;
  reg [_tmp_966-1:0] __tmp_967_45;
  reg [_tmp_966-1:0] __tmp_967_46;
  localparam _tmp_968 = 1;
  wire [_tmp_968-1:0] _tmp_969;
  assign _tmp_969 = _stream_conv2d_16_fsm == 3;
  reg [_tmp_968-1:0] __tmp_969_1;
  reg [_tmp_968-1:0] __tmp_969_2;
  reg [_tmp_968-1:0] __tmp_969_3;
  reg [_tmp_968-1:0] __tmp_969_4;
  reg [_tmp_968-1:0] __tmp_969_5;
  reg [_tmp_968-1:0] __tmp_969_6;
  reg [_tmp_968-1:0] __tmp_969_7;
  reg [_tmp_968-1:0] __tmp_969_8;
  reg [_tmp_968-1:0] __tmp_969_9;
  reg [_tmp_968-1:0] __tmp_969_10;
  reg [_tmp_968-1:0] __tmp_969_11;
  reg [_tmp_968-1:0] __tmp_969_12;
  reg [_tmp_968-1:0] __tmp_969_13;
  reg [_tmp_968-1:0] __tmp_969_14;
  reg [_tmp_968-1:0] __tmp_969_15;
  reg [_tmp_968-1:0] __tmp_969_16;
  reg [_tmp_968-1:0] __tmp_969_17;
  reg [_tmp_968-1:0] __tmp_969_18;
  reg [_tmp_968-1:0] __tmp_969_19;
  reg [_tmp_968-1:0] __tmp_969_20;
  reg [_tmp_968-1:0] __tmp_969_21;
  reg [_tmp_968-1:0] __tmp_969_22;
  reg [_tmp_968-1:0] __tmp_969_23;
  reg [_tmp_968-1:0] __tmp_969_24;
  reg [_tmp_968-1:0] __tmp_969_25;
  reg [_tmp_968-1:0] __tmp_969_26;
  reg [_tmp_968-1:0] __tmp_969_27;
  reg [_tmp_968-1:0] __tmp_969_28;
  reg [_tmp_968-1:0] __tmp_969_29;
  reg [_tmp_968-1:0] __tmp_969_30;
  reg [_tmp_968-1:0] __tmp_969_31;
  reg [_tmp_968-1:0] __tmp_969_32;
  reg [_tmp_968-1:0] __tmp_969_33;
  reg [_tmp_968-1:0] __tmp_969_34;
  reg [_tmp_968-1:0] __tmp_969_35;
  reg [_tmp_968-1:0] __tmp_969_36;
  reg [_tmp_968-1:0] __tmp_969_37;
  reg [_tmp_968-1:0] __tmp_969_38;
  reg [_tmp_968-1:0] __tmp_969_39;
  reg [_tmp_968-1:0] __tmp_969_40;
  reg [_tmp_968-1:0] __tmp_969_41;
  reg [_tmp_968-1:0] __tmp_969_42;
  wire conv2d_16_dma_out_mask_0;
  assign conv2d_16_dma_out_mask_0 = conv2d_16_out_row_count + 0 >= cparam_conv2d_16_out_num_row;
  reg axim_flag_970;
  reg _control_conv2d_16_cond_48_10_1;
  reg _maxi_ram_w8_l2048_id11_1_write_start;
  reg [8-1:0] _maxi_ram_w8_l2048_id11_1_write_op_sel;
  reg [32-1:0] _maxi_ram_w8_l2048_id11_1_write_local_addr;
  reg [32-1:0] _maxi_ram_w8_l2048_id11_1_write_global_addr;
  reg [33-1:0] _maxi_ram_w8_l2048_id11_1_write_size;
  reg [32-1:0] _maxi_ram_w8_l2048_id11_1_write_local_stride;
  reg [32-1:0] _maxi_write_fsm;
  localparam _maxi_write_fsm_init = 0;
  reg [32-1:0] _maxi_write_cur_global_addr;
  reg [33-1:0] _maxi_write_cur_size;
  reg [33-1:0] _maxi_write_rest_size;
  reg _tmp_971;
  reg _tmp_972;
  wire _tmp_973;
  wire _tmp_974;
  assign _tmp_974 = 1;
  localparam _tmp_975 = 1;
  wire [_tmp_975-1:0] _tmp_976;
  assign _tmp_976 = (_tmp_973 || !_tmp_971) && (_tmp_974 || !_tmp_972);
  reg [_tmp_975-1:0] __tmp_976_1;
  wire signed [8-1:0] _tmp_977;
  reg signed [8-1:0] __tmp_977_1;
  assign _tmp_977 = (__tmp_976_1)? ram_w8_l2048_id11_0_1_rdata : __tmp_977_1;
  reg _tmp_978;
  reg _tmp_979;
  reg _tmp_980;
  reg _tmp_981;
  reg [34-1:0] _tmp_982;
  reg _tmp_983;
  reg _tmp_984;
  wire _tmp_985;
  wire _tmp_986;
  assign _tmp_986 = 1;
  localparam _tmp_987 = 1;
  wire [_tmp_987-1:0] _tmp_988;
  assign _tmp_988 = (_tmp_985 || !_tmp_983) && (_tmp_986 || !_tmp_984);
  reg [_tmp_987-1:0] __tmp_988_1;
  wire signed [8-1:0] _tmp_989;
  reg signed [8-1:0] __tmp_989_1;
  assign _tmp_989 = (__tmp_988_1)? ram_w8_l2048_id11_1_1_rdata : __tmp_989_1;
  reg _tmp_990;
  reg _tmp_991;
  reg _tmp_992;
  reg _tmp_993;
  reg [34-1:0] _tmp_994;
  reg _tmp_995;
  reg _tmp_996;
  wire _tmp_997;
  wire _tmp_998;
  assign _tmp_998 = 1;
  localparam _tmp_999 = 1;
  wire [_tmp_999-1:0] _tmp_1000;
  assign _tmp_1000 = (_tmp_997 || !_tmp_995) && (_tmp_998 || !_tmp_996);
  reg [_tmp_999-1:0] __tmp_1000_1;
  wire signed [8-1:0] _tmp_1001;
  reg signed [8-1:0] __tmp_1001_1;
  assign _tmp_1001 = (__tmp_1000_1)? ram_w8_l2048_id11_2_1_rdata : __tmp_1001_1;
  reg _tmp_1002;
  reg _tmp_1003;
  reg _tmp_1004;
  reg _tmp_1005;
  reg [34-1:0] _tmp_1006;
  reg _tmp_1007;
  reg _tmp_1008;
  wire _tmp_1009;
  wire _tmp_1010;
  assign _tmp_1010 = 1;
  localparam _tmp_1011 = 1;
  wire [_tmp_1011-1:0] _tmp_1012;
  assign _tmp_1012 = (_tmp_1009 || !_tmp_1007) && (_tmp_1010 || !_tmp_1008);
  reg [_tmp_1011-1:0] __tmp_1012_1;
  wire signed [8-1:0] _tmp_1013;
  reg signed [8-1:0] __tmp_1013_1;
  assign _tmp_1013 = (__tmp_1012_1)? ram_w8_l2048_id11_3_1_rdata : __tmp_1013_1;
  reg _tmp_1014;
  reg _tmp_1015;
  reg _tmp_1016;
  reg _tmp_1017;
  reg [34-1:0] _tmp_1018;
  reg [9-1:0] _tmp_1019;
  reg _maxi_cond_1_1;
  reg _tmp_1020;
  wire [32-1:0] _dataflow_cat_odata_98;
  wire _dataflow_cat_ovalid_98;
  wire _dataflow_cat_oready_98;
  assign _dataflow_cat_oready_98 = (_maxi_write_fsm == 3) && (_maxi_write_op_sel == 1) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid));
  reg _maxi_cond_2_1;
  reg axim_flag_1021;
  reg [32-1:0] _d1__maxi_write_fsm;
  reg __maxi_write_fsm_cond_4_0_1;
  wire conv2d_16_update_filter;
  assign conv2d_16_update_filter = (cparam_conv2d_16_data_stationary == 0) && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_bat_count >= cparam_conv2d_16_max_bat_count) || (cparam_conv2d_16_data_stationary == 1) && !cparam_conv2d_16_keep_filter;
  wire conv2d_16_update_act;
  assign conv2d_16_update_act = (cparam_conv2d_16_data_stationary == 1) && (conv2d_16_och_count >= cparam_conv2d_16_max_och_count) || (cparam_conv2d_16_data_stationary == 0);
  wire conv2d_16_mux_next_dma_flag_0;
  assign conv2d_16_mux_next_dma_flag_0 = (conv2d_16_row_select == 0)? (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)? 1 : cparam_conv2d_16_dma_flag_conds_0 : 
                                         (conv2d_16_row_select == 1)? (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)? 1 : cparam_conv2d_16_dma_flag_conds_2 : 
                                         (conv2d_16_row_select == 2)? (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)? 1 : cparam_conv2d_16_dma_flag_conds_1 : 1'd0;
  wire conv2d_16_mux_next_dma_flag_1;
  assign conv2d_16_mux_next_dma_flag_1 = (conv2d_16_row_select == 0)? (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)? 1 : cparam_conv2d_16_dma_flag_conds_1 : 
                                         (conv2d_16_row_select == 1)? (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)? 1 : cparam_conv2d_16_dma_flag_conds_0 : 
                                         (conv2d_16_row_select == 2)? (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)? 1 : cparam_conv2d_16_dma_flag_conds_2 : 1'd0;
  wire conv2d_16_mux_next_dma_flag_2;
  assign conv2d_16_mux_next_dma_flag_2 = (conv2d_16_row_select == 0)? (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)? 1 : cparam_conv2d_16_dma_flag_conds_2 : 
                                         (conv2d_16_row_select == 1)? (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)? 1 : cparam_conv2d_16_dma_flag_conds_1 : 
                                         (conv2d_16_row_select == 2)? (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)? 1 : cparam_conv2d_16_dma_flag_conds_0 : 1'd0;
  reg [32-1:0] max_pool_serial_18_objaddr;
  reg [32-1:0] max_pool_serial_18_arg_objaddr_0;
  reg [32-1:0] control_max_pool_serial_18;
  localparam control_max_pool_serial_18_init = 0;
  reg _control_max_pool_serial_18_called;
  wire signed [32-1:0] max_pool_serial_18_act_base_offset;
  reg signed [32-1:0] max_pool_serial_18_act_base_offset_row;
  reg signed [32-1:0] max_pool_serial_18_act_base_offset_bat;
  assign max_pool_serial_18_act_base_offset = max_pool_serial_18_act_base_offset_row + max_pool_serial_18_act_base_offset_bat;
  wire signed [32-1:0] max_pool_serial_18_out_base_offset;
  reg signed [32-1:0] max_pool_serial_18_out_base_offset_row;
  reg signed [32-1:0] max_pool_serial_18_out_base_offset_bat;
  assign max_pool_serial_18_out_base_offset = max_pool_serial_18_out_base_offset_row + max_pool_serial_18_out_base_offset_bat;
  reg [32-1:0] max_pool_serial_18_col_count;
  reg [32-1:0] max_pool_serial_18_row_count;
  reg [32-1:0] max_pool_serial_18_bat_count;
  reg [32-1:0] max_pool_serial_18_prev_row_count;
  reg [32-1:0] max_pool_serial_18_prev_bat_count;
  reg [32-1:0] max_pool_serial_18_stream_act_local;
  reg [32-1:0] max_pool_serial_18_stream_out_local;
  reg max_pool_serial_18_act_page;
  reg [32-1:0] max_pool_serial_18_act_page_comp_offset;
  reg [32-1:0] max_pool_serial_18_act_page_dma_offset;
  reg max_pool_serial_18_out_page;
  reg [32-1:0] max_pool_serial_18_out_page_comp_offset;
  reg [32-1:0] max_pool_serial_18_out_page_dma_offset;
  reg max_pool_serial_18_skip_read_act;
  reg max_pool_serial_18_skip_comp;
  reg max_pool_serial_18_skip_write_out;
  reg [32-1:0] max_pool_serial_18_comp_count;
  reg [32-1:0] max_pool_serial_18_out_count;
  wire max_pool_serial_18_dma_pad_mask_0;
  assign max_pool_serial_18_dma_pad_mask_0 = (max_pool_serial_18_row_count + 0 < cparam_max_pool_serial_18_pad_row_top) || (max_pool_serial_18_row_count + 0 >= cparam_max_pool_serial_18_act_num_row + cparam_max_pool_serial_18_pad_row_top);
  wire max_pool_serial_18_dma_pad_mask_1;
  assign max_pool_serial_18_dma_pad_mask_1 = (max_pool_serial_18_row_count + 1 < cparam_max_pool_serial_18_pad_row_top) || (max_pool_serial_18_row_count + 1 >= cparam_max_pool_serial_18_act_num_row + cparam_max_pool_serial_18_pad_row_top);
  reg axim_flag_1022;
  reg [32-1:0] _d1_control_max_pool_serial_18;
  reg _control_max_pool_serial_18_cond_5_0_1;
  reg axim_flag_1023;
  reg _control_max_pool_serial_18_cond_11_1_1;
  reg [32-1:0] max_pool_serial_18_comp_fsm;
  localparam max_pool_serial_18_comp_fsm_init = 0;
  reg [32-1:0] max_pool_serial_18_act_page_comp_offset_buf;
  reg [32-1:0] max_pool_serial_18_out_page_comp_offset_buf;
  reg [32-1:0] max_pool_serial_18_row_count_buf;
  wire max_pool_serial_18_stream_pad_mask_0_0;
  assign max_pool_serial_18_stream_pad_mask_0_0 = (max_pool_serial_18_col_count + 0 < cparam_max_pool_serial_18_pad_col_left) || (max_pool_serial_18_col_count + 0 >= cparam_max_pool_serial_18_act_num_col + cparam_max_pool_serial_18_pad_col_left) || (max_pool_serial_18_row_count_buf + 0 < cparam_max_pool_serial_18_pad_row_top) || (max_pool_serial_18_row_count_buf + 0 >= cparam_max_pool_serial_18_act_num_row + cparam_max_pool_serial_18_pad_row_top);
  wire max_pool_serial_18_stream_pad_mask_0_1;
  assign max_pool_serial_18_stream_pad_mask_0_1 = (max_pool_serial_18_col_count + 1 < cparam_max_pool_serial_18_pad_col_left) || (max_pool_serial_18_col_count + 1 >= cparam_max_pool_serial_18_act_num_col + cparam_max_pool_serial_18_pad_col_left) || (max_pool_serial_18_row_count_buf + 0 < cparam_max_pool_serial_18_pad_row_top) || (max_pool_serial_18_row_count_buf + 0 >= cparam_max_pool_serial_18_act_num_row + cparam_max_pool_serial_18_pad_row_top);
  wire max_pool_serial_18_stream_pad_mask_1_0;
  assign max_pool_serial_18_stream_pad_mask_1_0 = (max_pool_serial_18_col_count + 0 < cparam_max_pool_serial_18_pad_col_left) || (max_pool_serial_18_col_count + 0 >= cparam_max_pool_serial_18_act_num_col + cparam_max_pool_serial_18_pad_col_left) || (max_pool_serial_18_row_count_buf + 1 < cparam_max_pool_serial_18_pad_row_top) || (max_pool_serial_18_row_count_buf + 1 >= cparam_max_pool_serial_18_act_num_row + cparam_max_pool_serial_18_pad_row_top);
  wire max_pool_serial_18_stream_pad_mask_1_1;
  assign max_pool_serial_18_stream_pad_mask_1_1 = (max_pool_serial_18_col_count + 1 < cparam_max_pool_serial_18_pad_col_left) || (max_pool_serial_18_col_count + 1 >= cparam_max_pool_serial_18_act_num_col + cparam_max_pool_serial_18_pad_col_left) || (max_pool_serial_18_row_count_buf + 1 < cparam_max_pool_serial_18_pad_row_top) || (max_pool_serial_18_row_count_buf + 1 >= cparam_max_pool_serial_18_act_num_row + cparam_max_pool_serial_18_pad_row_top);
  reg [4-1:0] max_pool_serial_18_stream_pad_masks;
  wire [3-1:0] stream_max_pool_serial_18_constant_0_data;
  wire [8-1:0] stream_max_pool_serial_18_source_1_data;
  wire [4-1:0] stream_max_pool_serial_18_constant_2_data;
  reg [32-1:0] _counter_data_782;
  reg [32-1:0] _counter_count_782;
  wire [8-1:0] _reinterpretcast_src_789;
  assign _reinterpretcast_src_789 = stream_max_pool_serial_18_source_1_data;
  wire signed [8-1:0] _reinterpretcast_data_789;
  assign _reinterpretcast_data_789 = _reinterpretcast_src_789;
  reg [4-1:0] __delay_data_1411;
  reg signed [8-1:0] __delay_data_1412;
  reg [3-1:0] __delay_data_1414;
  reg [1-1:0] _pointer_data_784;
  reg signed [8-1:0] __delay_data_1413;
  reg [3-1:0] __delay_data_1415;
  reg signed [9-1:0] _cond_data_791;
  reg [3-1:0] __delay_data_1416;
  reg signed [8-1:0] __variable_wdata_207;
  assign _reduce_max_13_x_data = __variable_wdata_207;
  reg [8-1:0] __variable_wdata_208;
  assign _reduce_max_13_size_data = __variable_wdata_208;
  reg signed [8-1:0] __substreamoutput_data_793;
  reg [1-1:0] __substreamoutput_data_794;
  wire signed [8-1:0] _reinterpretcast_src_795;
  assign _reinterpretcast_src_795 = __substreamoutput_data_793;
  wire signed [8-1:0] _reinterpretcast_data_795;
  assign _reinterpretcast_data_795 = _reinterpretcast_src_795;
  wire [1-1:0] stream_max_pool_serial_18_sink_4_data;
  assign stream_max_pool_serial_18_sink_4_data = __substreamoutput_data_794;
  wire signed [8-1:0] stream_max_pool_serial_18_sink_3_data;
  assign stream_max_pool_serial_18_sink_3_data = _reinterpretcast_data_795;
  reg _set_flag_1024;
  reg [3-1:0] __variable_wdata_777;
  assign stream_max_pool_serial_18_constant_0_data = __variable_wdata_777;
  reg _set_flag_1025;
  reg [4-1:0] __variable_wdata_779;
  assign stream_max_pool_serial_18_constant_2_data = __variable_wdata_779;
  reg [32-1:0] _source_stream_max_pool_serial_18_source_1_pat_cur_offset_0;
  reg [32-1:0] _source_stream_max_pool_serial_18_source_1_pat_cur_offset_1;
  reg [32-1:0] _source_stream_max_pool_serial_18_source_1_pat_cur_offset_2;
  reg [32-1:0] _source_stream_max_pool_serial_18_source_1_pat_cur_offset_3;
  reg [33-1:0] _source_stream_max_pool_serial_18_source_1_pat_size_0;
  reg [33-1:0] _source_stream_max_pool_serial_18_source_1_pat_size_1;
  reg [33-1:0] _source_stream_max_pool_serial_18_source_1_pat_size_2;
  reg [33-1:0] _source_stream_max_pool_serial_18_source_1_pat_size_3;
  reg [32-1:0] _source_stream_max_pool_serial_18_source_1_pat_stride_0;
  reg [32-1:0] _source_stream_max_pool_serial_18_source_1_pat_stride_1;
  reg [32-1:0] _source_stream_max_pool_serial_18_source_1_pat_stride_2;
  reg [32-1:0] _source_stream_max_pool_serial_18_source_1_pat_stride_3;
  reg [33-1:0] _source_stream_max_pool_serial_18_source_1_pat_count_0;
  reg [33-1:0] _source_stream_max_pool_serial_18_source_1_pat_count_1;
  reg [33-1:0] _source_stream_max_pool_serial_18_source_1_pat_count_2;
  reg [33-1:0] _source_stream_max_pool_serial_18_source_1_pat_count_3;
  reg [33-1:0] _source_stream_max_pool_serial_18_source_1_pat_size_buf_0;
  reg [33-1:0] _source_stream_max_pool_serial_18_source_1_pat_size_buf_1;
  reg [33-1:0] _source_stream_max_pool_serial_18_source_1_pat_size_buf_2;
  reg [33-1:0] _source_stream_max_pool_serial_18_source_1_pat_size_buf_3;
  reg [32-1:0] _source_stream_max_pool_serial_18_source_1_pat_stride_buf_0;
  reg [32-1:0] _source_stream_max_pool_serial_18_source_1_pat_stride_buf_1;
  reg [32-1:0] _source_stream_max_pool_serial_18_source_1_pat_stride_buf_2;
  reg [32-1:0] _source_stream_max_pool_serial_18_source_1_pat_stride_buf_3;
  reg _set_flag_1026;
  wire [2-1:0] _tmp_1027;
  assign _tmp_1027 = _stream_max_pool_serial_18_source_1_source_ram_raddr;
  reg [2-1:0] __tmp_1027_1;
  reg [2-1:0] __tmp_1027_2;
  reg _tmp_1028;
  reg _ram_w8_l2048_id1_0_cond_3_1;
  reg _ram_w8_l2048_id1_0_cond_4_1;
  reg _ram_w8_l2048_id1_0_cond_4_2;
  reg _tmp_1029;
  reg _ram_w8_l2048_id1_1_cond_3_1;
  reg _ram_w8_l2048_id1_1_cond_4_1;
  reg _ram_w8_l2048_id1_1_cond_4_2;
  reg _tmp_1030;
  reg _ram_w8_l2048_id1_2_cond_3_1;
  reg _ram_w8_l2048_id1_2_cond_4_1;
  reg _ram_w8_l2048_id1_2_cond_4_2;
  reg _tmp_1031;
  reg _ram_w8_l2048_id1_3_cond_3_1;
  reg _ram_w8_l2048_id1_3_cond_4_1;
  reg _ram_w8_l2048_id1_3_cond_4_2;
  wire signed [8-1:0] _tmp_1032;
  wire _tmp_1033;
  assign _tmp_1032 = (__tmp_1027_2 == 0)? ram_w8_l2048_id1_0_0_rdata : 
                     (__tmp_1027_2 == 1)? ram_w8_l2048_id1_1_0_rdata : 
                     (__tmp_1027_2 == 2)? ram_w8_l2048_id1_2_0_rdata : 
                     (__tmp_1027_2 == 3)? ram_w8_l2048_id1_3_0_rdata : 0;
  assign _tmp_1033 = _tmp_1028;
  assign _stream_max_pool_serial_18_source_1_source_ram_rdata = (_stream_max_pool_serial_18_source_1_source_ram_sel == 1)? _tmp_1032 : 0;
  localparam _tmp_1034 = 1;
  wire [_tmp_1034-1:0] _tmp_1035;
  assign _tmp_1035 = _stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1);
  reg [_tmp_1034-1:0] __tmp_1035_1;
  reg [8-1:0] __variable_wdata_778;
  assign stream_max_pool_serial_18_source_1_data = __variable_wdata_778;
  reg [32-1:0] _stream_max_pool_serial_18_source_1_source_pat_fsm_0;
  localparam _stream_max_pool_serial_18_source_1_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_max_pool_serial_18_source_1_source_pat_all_offset;
  assign _stream_max_pool_serial_18_source_1_source_pat_all_offset = _stream_max_pool_serial_18_source_1_source_offset_buf + _source_stream_max_pool_serial_18_source_1_pat_cur_offset_0 + _source_stream_max_pool_serial_18_source_1_pat_cur_offset_1 + _source_stream_max_pool_serial_18_source_1_pat_cur_offset_2 + _source_stream_max_pool_serial_18_source_1_pat_cur_offset_3;
  reg _set_flag_1036;
  reg [32-1:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_1;
  reg [32-1:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_2;
  reg [32-1:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_3;
  reg [32-1:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_4;
  reg [32-1:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_5;
  reg [32-1:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_6;
  reg [32-1:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_7;
  reg [32-1:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_8;
  reg [32-1:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_9;
  reg [33-1:0] __stream_max_pool_serial_18_sink_3_sink_size_1_1;
  reg [33-1:0] __stream_max_pool_serial_18_sink_3_sink_size_1_2;
  reg [33-1:0] __stream_max_pool_serial_18_sink_3_sink_size_1_3;
  reg [33-1:0] __stream_max_pool_serial_18_sink_3_sink_size_1_4;
  reg [33-1:0] __stream_max_pool_serial_18_sink_3_sink_size_1_5;
  reg [33-1:0] __stream_max_pool_serial_18_sink_3_sink_size_1_6;
  reg [33-1:0] __stream_max_pool_serial_18_sink_3_sink_size_1_7;
  reg [33-1:0] __stream_max_pool_serial_18_sink_3_sink_size_1_8;
  reg [33-1:0] __stream_max_pool_serial_18_sink_3_sink_size_1_9;
  reg __stream_seq_15_cond_2_1;
  reg __stream_seq_15_cond_2_2;
  reg __stream_seq_15_cond_2_3;
  reg __stream_seq_15_cond_2_4;
  reg __stream_seq_15_cond_2_5;
  reg __stream_seq_15_cond_2_6;
  reg __stream_seq_15_cond_2_7;
  reg __stream_seq_15_cond_2_8;
  reg __stream_seq_15_cond_2_9;
  reg __set_flag_1036_1;
  reg __set_flag_1036_2;
  reg __set_flag_1036_3;
  reg __set_flag_1036_4;
  reg __set_flag_1036_5;
  reg __set_flag_1036_6;
  reg __set_flag_1036_7;
  reg __set_flag_1036_8;
  reg __set_flag_1036_9;
  wire [2-1:0] _tmp_1037;
  assign _tmp_1037 = _stream_max_pool_serial_18_sink_3_sink_waddr;
  reg _ram_w8_l2048_id0_0_cond_3_1;
  reg _ram_w8_l2048_id0_1_cond_3_1;
  reg _ram_w8_l2048_id0_2_cond_3_1;
  reg _ram_w8_l2048_id0_3_cond_3_1;
  reg __stream_max_pool_serial_18_start_1;
  reg __stream_max_pool_serial_18_start_2;
  reg __stream_max_pool_serial_18_start_3;
  reg __stream_max_pool_serial_18_start_4;
  reg __stream_max_pool_serial_18_start_5;
  reg __stream_max_pool_serial_18_start_6;
  reg __stream_max_pool_serial_18_start_7;
  reg __stream_max_pool_serial_18_start_8;
  reg __stream_max_pool_serial_18_start_9;
  reg __stream_max_pool_serial_18_start_10;
  reg [32-1:0] _stream_max_pool_serial_18_sink_3_sink_fsm_1;
  localparam _stream_max_pool_serial_18_sink_3_sink_fsm_1_init = 0;
  reg _set_flag_1038;
  assign _stream_max_pool_serial_18_start_flag = (_set_flag_1038)? 1 : 0;
  localparam _tmp_1039 = 1;
  wire [_tmp_1039-1:0] _tmp_1040;
  assign _tmp_1040 = (_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag;
  reg [_tmp_1039-1:0] __tmp_1040_1;
  reg [_tmp_1039-1:0] __tmp_1040_2;
  reg [_tmp_1039-1:0] __tmp_1040_3;
  reg [_tmp_1039-1:0] __tmp_1040_4;
  reg [_tmp_1039-1:0] __tmp_1040_5;
  localparam _tmp_1041 = 1;
  wire [_tmp_1041-1:0] _tmp_1042;
  assign _tmp_1042 = (_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag;
  reg [_tmp_1041-1:0] __tmp_1042_1;
  reg [_tmp_1041-1:0] __tmp_1042_2;
  reg [_tmp_1041-1:0] __tmp_1042_3;
  reg [_tmp_1041-1:0] __tmp_1042_4;
  reg [_tmp_1041-1:0] __tmp_1042_5;
  reg [_tmp_1041-1:0] __tmp_1042_6;
  reg [_tmp_1041-1:0] __tmp_1042_7;
  reg [_tmp_1041-1:0] __tmp_1042_8;
  reg [_tmp_1041-1:0] __tmp_1042_9;
  localparam _tmp_1043 = 1;
  wire [_tmp_1043-1:0] _tmp_1044;
  assign _tmp_1044 = (_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag;
  reg [_tmp_1043-1:0] __tmp_1044_1;
  reg [_tmp_1043-1:0] __tmp_1044_2;
  reg [_tmp_1043-1:0] __tmp_1044_3;
  reg [_tmp_1043-1:0] __tmp_1044_4;
  reg [_tmp_1043-1:0] __tmp_1044_5;
  reg [_tmp_1043-1:0] __tmp_1044_6;
  reg [_tmp_1043-1:0] __tmp_1044_7;
  localparam _tmp_1045 = 1;
  wire [_tmp_1045-1:0] _tmp_1046;
  assign _tmp_1046 = (_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag;
  reg [_tmp_1045-1:0] __tmp_1046_1;
  reg [_tmp_1045-1:0] __tmp_1046_2;
  reg [_tmp_1045-1:0] __tmp_1046_3;
  reg [_tmp_1045-1:0] __tmp_1046_4;
  reg [_tmp_1045-1:0] __tmp_1046_5;
  reg [_tmp_1045-1:0] __tmp_1046_6;
  reg [_tmp_1045-1:0] __tmp_1046_7;
  wire _stream_max_pool_serial_18_done;
  assign _stream_max_pool_serial_18_done = _stream_max_pool_serial_18_source_1_idle;
  localparam _tmp_1047 = 1;
  wire [_tmp_1047-1:0] _tmp_1048;
  assign _tmp_1048 = _stream_max_pool_serial_18_fsm == 3;
  reg [_tmp_1047-1:0] __tmp_1048_1;
  localparam _tmp_1049 = 1;
  wire [_tmp_1049-1:0] _tmp_1050;
  assign _tmp_1050 = _stream_max_pool_serial_18_fsm == 3;
  reg [_tmp_1049-1:0] __tmp_1050_1;
  reg [_tmp_1049-1:0] __tmp_1050_2;
  reg [_tmp_1049-1:0] __tmp_1050_3;
  reg [_tmp_1049-1:0] __tmp_1050_4;
  reg [_tmp_1049-1:0] __tmp_1050_5;
  localparam _tmp_1051 = 1;
  wire [_tmp_1051-1:0] _tmp_1052;
  assign _tmp_1052 = _stream_max_pool_serial_18_fsm == 3;
  reg [_tmp_1051-1:0] __tmp_1052_1;
  reg [_tmp_1051-1:0] __tmp_1052_2;
  reg [_tmp_1051-1:0] __tmp_1052_3;
  reg [_tmp_1051-1:0] __tmp_1052_4;
  localparam _tmp_1053 = 1;
  wire [_tmp_1053-1:0] _tmp_1054;
  assign _tmp_1054 = _stream_max_pool_serial_18_fsm == 3;
  reg [_tmp_1053-1:0] __tmp_1054_1;
  reg [_tmp_1053-1:0] __tmp_1054_2;
  reg [_tmp_1053-1:0] __tmp_1054_3;
  reg [_tmp_1053-1:0] __tmp_1054_4;
  reg [3-1:0] __reduce_max_13_sink_wait_count;
  localparam _tmp_1055 = 1;
  wire [_tmp_1055-1:0] _tmp_1056;
  assign _tmp_1056 = _stream_max_pool_serial_18_fsm == 3;
  reg [_tmp_1055-1:0] __tmp_1056_1;
  reg [_tmp_1055-1:0] __tmp_1056_2;
  reg [_tmp_1055-1:0] __tmp_1056_3;
  reg [_tmp_1055-1:0] __tmp_1056_4;
  reg [_tmp_1055-1:0] __tmp_1056_5;
  localparam _tmp_1057 = 1;
  wire [_tmp_1057-1:0] _tmp_1058;
  assign _tmp_1058 = _stream_max_pool_serial_18_fsm == 3;
  reg [_tmp_1057-1:0] __tmp_1058_1;
  reg [_tmp_1057-1:0] __tmp_1058_2;
  reg [_tmp_1057-1:0] __tmp_1058_3;
  reg [_tmp_1057-1:0] __tmp_1058_4;
  reg [_tmp_1057-1:0] __tmp_1058_5;
  localparam _tmp_1059 = 1;
  wire [_tmp_1059-1:0] _tmp_1060;
  assign _tmp_1060 = _stream_max_pool_serial_18_fsm == 3;
  reg [_tmp_1059-1:0] __tmp_1060_1;
  reg [_tmp_1059-1:0] __tmp_1060_2;
  reg [_tmp_1059-1:0] __tmp_1060_3;
  reg [_tmp_1059-1:0] __tmp_1060_4;
  reg [_tmp_1059-1:0] __tmp_1060_5;
  reg [4-1:0] _stream_max_pool_serial_18_sink_wait_count;
  localparam _tmp_1061 = 1;
  wire [_tmp_1061-1:0] _tmp_1062;
  assign _tmp_1062 = _stream_max_pool_serial_18_fsm == 3;
  reg [_tmp_1061-1:0] __tmp_1062_1;
  reg [_tmp_1061-1:0] __tmp_1062_2;
  reg [_tmp_1061-1:0] __tmp_1062_3;
  reg [_tmp_1061-1:0] __tmp_1062_4;
  reg [_tmp_1061-1:0] __tmp_1062_5;
  reg [_tmp_1061-1:0] __tmp_1062_6;
  reg [_tmp_1061-1:0] __tmp_1062_7;
  reg [_tmp_1061-1:0] __tmp_1062_8;
  reg [_tmp_1061-1:0] __tmp_1062_9;
  reg [_tmp_1061-1:0] __tmp_1062_10;
  localparam _tmp_1063 = 1;
  wire [_tmp_1063-1:0] _tmp_1064;
  assign _tmp_1064 = _stream_max_pool_serial_18_fsm == 3;
  reg [_tmp_1063-1:0] __tmp_1064_1;
  reg [_tmp_1063-1:0] __tmp_1064_2;
  reg [_tmp_1063-1:0] __tmp_1064_3;
  reg [_tmp_1063-1:0] __tmp_1064_4;
  reg [_tmp_1063-1:0] __tmp_1064_5;
  reg [_tmp_1063-1:0] __tmp_1064_6;
  reg [_tmp_1063-1:0] __tmp_1064_7;
  reg [_tmp_1063-1:0] __tmp_1064_8;
  reg [_tmp_1063-1:0] __tmp_1064_9;
  reg [_tmp_1063-1:0] __tmp_1064_10;
  localparam _tmp_1065 = 1;
  wire [_tmp_1065-1:0] _tmp_1066;
  assign _tmp_1066 = _stream_max_pool_serial_18_fsm == 3;
  reg [_tmp_1065-1:0] __tmp_1066_1;
  reg [_tmp_1065-1:0] __tmp_1066_2;
  reg [_tmp_1065-1:0] __tmp_1066_3;
  reg [_tmp_1065-1:0] __tmp_1066_4;
  reg [_tmp_1065-1:0] __tmp_1066_5;
  reg [_tmp_1065-1:0] __tmp_1066_6;
  reg [_tmp_1065-1:0] __tmp_1066_7;
  reg [_tmp_1065-1:0] __tmp_1066_8;
  reg [_tmp_1065-1:0] __tmp_1066_9;
  reg [_tmp_1065-1:0] __tmp_1066_10;
  localparam _tmp_1067 = 1;
  wire [_tmp_1067-1:0] _tmp_1068;
  assign _tmp_1068 = _stream_max_pool_serial_18_fsm == 3;
  reg [_tmp_1067-1:0] __tmp_1068_1;
  reg [_tmp_1067-1:0] __tmp_1068_2;
  reg [_tmp_1067-1:0] __tmp_1068_3;
  reg [_tmp_1067-1:0] __tmp_1068_4;
  reg [_tmp_1067-1:0] __tmp_1068_5;
  reg [_tmp_1067-1:0] __tmp_1068_6;
  reg [_tmp_1067-1:0] __tmp_1068_7;
  reg [_tmp_1067-1:0] __tmp_1068_8;
  reg [_tmp_1067-1:0] __tmp_1068_9;
  reg [_tmp_1067-1:0] __tmp_1068_10;
  localparam _tmp_1069 = 1;
  wire [_tmp_1069-1:0] _tmp_1070;
  assign _tmp_1070 = _stream_max_pool_serial_18_fsm == 3;
  reg [_tmp_1069-1:0] __tmp_1070_1;
  reg [_tmp_1069-1:0] __tmp_1070_2;
  reg [_tmp_1069-1:0] __tmp_1070_3;
  reg [_tmp_1069-1:0] __tmp_1070_4;
  reg [_tmp_1069-1:0] __tmp_1070_5;
  reg [_tmp_1069-1:0] __tmp_1070_6;
  reg axim_flag_1071;
  reg _control_max_pool_serial_18_cond_19_2_1;
  reg _maxi_ram_w8_l2048_id0_1_write_start;
  reg [8-1:0] _maxi_ram_w8_l2048_id0_1_write_op_sel;
  reg [32-1:0] _maxi_ram_w8_l2048_id0_1_write_local_addr;
  reg [32-1:0] _maxi_ram_w8_l2048_id0_1_write_global_addr;
  reg [33-1:0] _maxi_ram_w8_l2048_id0_1_write_size;
  reg [32-1:0] _maxi_ram_w8_l2048_id0_1_write_local_stride;
  reg _tmp_1072;
  reg _tmp_1073;
  wire _tmp_1074;
  wire _tmp_1075;
  assign _tmp_1075 = 1;
  localparam _tmp_1076 = 1;
  wire [_tmp_1076-1:0] _tmp_1077;
  assign _tmp_1077 = (_tmp_1074 || !_tmp_1072) && (_tmp_1075 || !_tmp_1073);
  reg [_tmp_1076-1:0] __tmp_1077_1;
  wire signed [8-1:0] _tmp_1078;
  reg signed [8-1:0] __tmp_1078_1;
  assign _tmp_1078 = (__tmp_1077_1)? ram_w8_l2048_id0_0_1_rdata : __tmp_1078_1;
  reg _tmp_1079;
  reg _tmp_1080;
  reg _tmp_1081;
  reg _tmp_1082;
  reg [34-1:0] _tmp_1083;
  reg _tmp_1084;
  reg _tmp_1085;
  wire _tmp_1086;
  wire _tmp_1087;
  assign _tmp_1087 = 1;
  localparam _tmp_1088 = 1;
  wire [_tmp_1088-1:0] _tmp_1089;
  assign _tmp_1089 = (_tmp_1086 || !_tmp_1084) && (_tmp_1087 || !_tmp_1085);
  reg [_tmp_1088-1:0] __tmp_1089_1;
  wire signed [8-1:0] _tmp_1090;
  reg signed [8-1:0] __tmp_1090_1;
  assign _tmp_1090 = (__tmp_1089_1)? ram_w8_l2048_id0_1_1_rdata : __tmp_1090_1;
  reg _tmp_1091;
  reg _tmp_1092;
  reg _tmp_1093;
  reg _tmp_1094;
  reg [34-1:0] _tmp_1095;
  reg _tmp_1096;
  reg _tmp_1097;
  wire _tmp_1098;
  wire _tmp_1099;
  assign _tmp_1099 = 1;
  localparam _tmp_1100 = 1;
  wire [_tmp_1100-1:0] _tmp_1101;
  assign _tmp_1101 = (_tmp_1098 || !_tmp_1096) && (_tmp_1099 || !_tmp_1097);
  reg [_tmp_1100-1:0] __tmp_1101_1;
  wire signed [8-1:0] _tmp_1102;
  reg signed [8-1:0] __tmp_1102_1;
  assign _tmp_1102 = (__tmp_1101_1)? ram_w8_l2048_id0_2_1_rdata : __tmp_1102_1;
  reg _tmp_1103;
  reg _tmp_1104;
  reg _tmp_1105;
  reg _tmp_1106;
  reg [34-1:0] _tmp_1107;
  reg _tmp_1108;
  reg _tmp_1109;
  wire _tmp_1110;
  wire _tmp_1111;
  assign _tmp_1111 = 1;
  localparam _tmp_1112 = 1;
  wire [_tmp_1112-1:0] _tmp_1113;
  assign _tmp_1113 = (_tmp_1110 || !_tmp_1108) && (_tmp_1111 || !_tmp_1109);
  reg [_tmp_1112-1:0] __tmp_1113_1;
  wire signed [8-1:0] _tmp_1114;
  reg signed [8-1:0] __tmp_1114_1;
  assign _tmp_1114 = (__tmp_1113_1)? ram_w8_l2048_id0_3_1_rdata : __tmp_1114_1;
  reg _tmp_1115;
  reg _tmp_1116;
  reg _tmp_1117;
  reg _tmp_1118;
  reg [34-1:0] _tmp_1119;
  reg _tmp_1120;
  wire [32-1:0] _dataflow_cat_odata_107;
  wire _dataflow_cat_ovalid_107;
  wire _dataflow_cat_oready_107;
  assign _dataflow_cat_oready_107 = (_maxi_write_fsm == 3) && (_maxi_write_op_sel == 2) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid));
  reg _maxi_cond_3_1;
  reg [32-1:0] matmul_29_objaddr;
  reg [32-1:0] matmul_29_arg_objaddr_0;
  reg [32-1:0] matmul_29_arg_objaddr_1;
  reg [32-1:0] matmul_29_arg_objaddr_2;
  reg [32-1:0] matmul_29_arg_objaddr_3;
  reg [32-1:0] control_matmul_29;
  localparam control_matmul_29_init = 0;
  reg _control_matmul_29_called;
  wire signed [32-1:0] matmul_29_act_base_offset;
  reg signed [32-1:0] matmul_29_act_base_offset_row;
  reg signed [32-1:0] matmul_29_act_base_offset_bat;
  assign matmul_29_act_base_offset = matmul_29_act_base_offset_row + matmul_29_act_base_offset_bat;
  reg signed [32-1:0] matmul_29_filter_base_offset;
  reg [32-1:0] matmul_29_next_stream_num_ops;
  wire signed [32-1:0] matmul_29_out_base_offset;
  reg signed [32-1:0] matmul_29_out_base_offset_val;
  reg signed [32-1:0] matmul_29_out_base_offset_col;
  reg signed [32-1:0] matmul_29_out_base_offset_row;
  reg signed [32-1:0] matmul_29_out_base_offset_bat;
  reg signed [32-1:0] matmul_29_out_base_offset_och;
  assign matmul_29_out_base_offset = matmul_29_out_base_offset_val + matmul_29_out_base_offset_col + matmul_29_out_base_offset_row + matmul_29_out_base_offset_bat + matmul_29_out_base_offset_och;
  reg matmul_29_dma_flag_0;
  reg [32-1:0] matmul_29_sync_comp_count;
  reg [32-1:0] matmul_29_sync_out_count;
  reg [32-1:0] matmul_29_write_count;
  reg [32-1:0] matmul_29_next_out_write_size;
  reg [32-1:0] matmul_29_col_count;
  reg [32-1:0] matmul_29_row_count;
  reg [32-1:0] matmul_29_bat_count;
  reg [32-1:0] matmul_29_och_count;
  reg [1-1:0] matmul_29_col_select;
  reg [1-1:0] matmul_29_row_select;
  reg [32-1:0] matmul_29_out_col_count;
  reg [32-1:0] matmul_29_out_row_count;
  reg [32-1:0] matmul_29_out_ram_select;
  reg [32-1:0] matmul_29_prev_col_count;
  reg [32-1:0] matmul_29_prev_row_count;
  reg [32-1:0] matmul_29_prev_bat_count;
  reg [32-1:0] matmul_29_prev_och_count;
  reg [1-1:0] matmul_29_prev_row_select;
  reg [32-1:0] matmul_29_stream_act_local_0;
  reg [32-1:0] matmul_29_stream_out_local_val;
  reg [32-1:0] matmul_29_stream_out_local_col;
  wire [32-1:0] matmul_29_stream_out_local;
  assign matmul_29_stream_out_local = matmul_29_stream_out_local_val + matmul_29_stream_out_local_col;
  reg [32-1:0] matmul_29_act_page_comp_offset_0;
  reg [32-1:0] matmul_29_act_page_dma_offset_0;
  reg [32-1:0] matmul_29_filter_page_comp_offset;
  reg [32-1:0] matmul_29_filter_page_dma_offset;
  reg matmul_29_out_page;
  reg [32-1:0] matmul_29_out_page_comp_offset;
  reg [32-1:0] matmul_29_out_page_dma_offset;
  reg [32-1:0] matmul_29_out_laddr_offset;
  reg matmul_29_skip_read_filter;
  reg matmul_29_skip_read_act;
  reg matmul_29_skip_comp;
  reg matmul_29_skip_write_out;
  reg axim_flag_1121;
  reg [32-1:0] _d1_control_matmul_29;
  reg _control_matmul_29_cond_3_0_1;
  reg _maxi_ram_w8_l2048_id2_1_read_start;
  reg [8-1:0] _maxi_ram_w8_l2048_id2_1_read_op_sel;
  reg [32-1:0] _maxi_ram_w8_l2048_id2_1_read_local_addr;
  reg [32-1:0] _maxi_ram_w8_l2048_id2_1_read_global_addr;
  reg [33-1:0] _maxi_ram_w8_l2048_id2_1_read_size;
  reg [32-1:0] _maxi_ram_w8_l2048_id2_1_read_local_stride;
  reg [32-1:0] _wdata_1122;
  reg _wvalid_1123;
  reg [34-1:0] _tmp_1124;
  reg _tmp_1125;
  wire [8-1:0] _dataflow_slice_odata_111;
  wire _dataflow_slice_ovalid_111;
  wire _dataflow_slice_oready_111;
  assign _dataflow_slice_oready_111 = (_tmp_1124 > 0) && !_tmp_1125;
  reg _ram_w8_l2048_id2_0_cond_4_1;
  reg [34-1:0] _tmp_1126;
  reg _tmp_1127;
  wire [8-1:0] _dataflow_slice_odata_114;
  wire _dataflow_slice_ovalid_114;
  wire _dataflow_slice_oready_114;
  assign _dataflow_slice_oready_114 = (_tmp_1126 > 0) && !_tmp_1127;
  reg _ram_w8_l2048_id2_1_cond_4_1;
  reg [34-1:0] _tmp_1128;
  reg _tmp_1129;
  wire [8-1:0] _dataflow_slice_odata_117;
  wire _dataflow_slice_ovalid_117;
  wire _dataflow_slice_oready_117;
  assign _dataflow_slice_oready_117 = (_tmp_1128 > 0) && !_tmp_1129;
  reg _ram_w8_l2048_id2_2_cond_4_1;
  reg [34-1:0] _tmp_1130;
  reg _tmp_1131;
  wire [8-1:0] _dataflow_slice_odata_120;
  wire _dataflow_slice_ovalid_120;
  wire _dataflow_slice_oready_120;
  assign _dataflow_slice_oready_120 = (_tmp_1130 > 0) && !_tmp_1131;
  reg _ram_w8_l2048_id2_3_cond_4_1;
  reg __maxi_read_fsm_cond_3_7_1;
  reg axim_flag_1132;
  reg _control_matmul_29_cond_8_1_1;
  reg axim_flag_1133;
  reg _control_matmul_29_cond_14_2_1;
  reg _maxi_ram_w4_l8192_id0_1_read_start;
  reg [8-1:0] _maxi_ram_w4_l8192_id0_1_read_op_sel;
  reg [32-1:0] _maxi_ram_w4_l8192_id0_1_read_local_addr;
  reg [32-1:0] _maxi_ram_w4_l8192_id0_1_read_global_addr;
  reg [33-1:0] _maxi_ram_w4_l8192_id0_1_read_size;
  reg [32-1:0] _maxi_ram_w4_l8192_id0_1_read_local_stride;
  reg [32-1:0] _wdata_1134;
  reg _wvalid_1135;
  reg [34-1:0] _tmp_1136;
  reg _tmp_1137;
  wire [4-1:0] _dataflow_slice_odata_124;
  wire _dataflow_slice_ovalid_124;
  wire _dataflow_slice_oready_124;
  assign _dataflow_slice_oready_124 = (_tmp_1136 > 0) && !_tmp_1137;
  reg _ram_w4_l8192_id0_0_cond_4_1;
  reg [34-1:0] _tmp_1138;
  reg _tmp_1139;
  wire [4-1:0] _dataflow_slice_odata_127;
  wire _dataflow_slice_ovalid_127;
  wire _dataflow_slice_oready_127;
  assign _dataflow_slice_oready_127 = (_tmp_1138 > 0) && !_tmp_1139;
  reg _ram_w4_l8192_id0_1_cond_4_1;
  reg [34-1:0] _tmp_1140;
  reg _tmp_1141;
  wire [4-1:0] _dataflow_slice_odata_130;
  wire _dataflow_slice_ovalid_130;
  wire _dataflow_slice_oready_130;
  assign _dataflow_slice_oready_130 = (_tmp_1140 > 0) && !_tmp_1141;
  reg _ram_w4_l8192_id0_2_cond_4_1;
  reg [34-1:0] _tmp_1142;
  reg _tmp_1143;
  wire [4-1:0] _dataflow_slice_odata_133;
  wire _dataflow_slice_ovalid_133;
  wire _dataflow_slice_oready_133;
  assign _dataflow_slice_oready_133 = (_tmp_1142 > 0) && !_tmp_1143;
  reg _ram_w4_l8192_id0_3_cond_4_1;
  reg [34-1:0] _tmp_1144;
  reg _tmp_1145;
  wire [4-1:0] _dataflow_slice_odata_136;
  wire _dataflow_slice_ovalid_136;
  wire _dataflow_slice_oready_136;
  assign _dataflow_slice_oready_136 = (_tmp_1144 > 0) && !_tmp_1145;
  reg _ram_w4_l8192_id0_4_cond_4_1;
  reg [34-1:0] _tmp_1146;
  reg _tmp_1147;
  wire [4-1:0] _dataflow_slice_odata_139;
  wire _dataflow_slice_ovalid_139;
  wire _dataflow_slice_oready_139;
  assign _dataflow_slice_oready_139 = (_tmp_1146 > 0) && !_tmp_1147;
  reg _ram_w4_l8192_id0_5_cond_4_1;
  reg [34-1:0] _tmp_1148;
  reg _tmp_1149;
  wire [4-1:0] _dataflow_slice_odata_142;
  wire _dataflow_slice_ovalid_142;
  wire _dataflow_slice_oready_142;
  assign _dataflow_slice_oready_142 = (_tmp_1148 > 0) && !_tmp_1149;
  reg _ram_w4_l8192_id0_6_cond_4_1;
  reg [34-1:0] _tmp_1150;
  reg _tmp_1151;
  wire [4-1:0] _dataflow_slice_odata_145;
  wire _dataflow_slice_ovalid_145;
  wire _dataflow_slice_oready_145;
  assign _dataflow_slice_oready_145 = (_tmp_1150 > 0) && !_tmp_1151;
  reg _ram_w4_l8192_id0_7_cond_4_1;
  reg __maxi_read_fsm_cond_3_8_1;
  wire [32-1:0] matmul_29_mux_act_gaddr_0;
  assign matmul_29_mux_act_gaddr_0 = (matmul_29_row_select == 0)? matmul_29_arg_objaddr_0 + (matmul_29_act_base_offset + cparam_matmul_29_act_offset_values_0) : 1'd0;
  wire matmul_29_dma_pad_mask_0;
  assign matmul_29_dma_pad_mask_0 = (matmul_29_row_count + 0 < cparam_matmul_29_pad_row_top) || (matmul_29_row_count + 0 >= cparam_matmul_29_act_num_row + cparam_matmul_29_pad_row_top);
  wire matmul_29_mux_dma_pad_mask_0;
  assign matmul_29_mux_dma_pad_mask_0 = (matmul_29_row_select == 0)? matmul_29_dma_pad_mask_0 : 1'd0;
  wire matmul_29_mux_dma_flag_0;
  assign matmul_29_mux_dma_flag_0 = (matmul_29_prev_row_select == 0)? matmul_29_dma_flag_0 : 1'd0;
  reg axim_flag_1152;
  reg _control_matmul_29_cond_22_3_1;
  reg _maxi_ram_w8_l2048_id3_1_read_start;
  reg [8-1:0] _maxi_ram_w8_l2048_id3_1_read_op_sel;
  reg [32-1:0] _maxi_ram_w8_l2048_id3_1_read_local_addr;
  reg [32-1:0] _maxi_ram_w8_l2048_id3_1_read_global_addr;
  reg [33-1:0] _maxi_ram_w8_l2048_id3_1_read_size;
  reg [32-1:0] _maxi_ram_w8_l2048_id3_1_read_local_stride;
  reg [32-1:0] _wdata_1153;
  reg _wvalid_1154;
  reg [34-1:0] _tmp_1155;
  reg _tmp_1156;
  wire [8-1:0] _dataflow_slice_odata_149;
  wire _dataflow_slice_ovalid_149;
  wire _dataflow_slice_oready_149;
  assign _dataflow_slice_oready_149 = (_tmp_1155 > 0) && !_tmp_1156;
  reg _ram_w8_l2048_id3_0_cond_3_1;
  reg [34-1:0] _tmp_1157;
  reg _tmp_1158;
  wire [8-1:0] _dataflow_slice_odata_152;
  wire _dataflow_slice_ovalid_152;
  wire _dataflow_slice_oready_152;
  assign _dataflow_slice_oready_152 = (_tmp_1157 > 0) && !_tmp_1158;
  reg _ram_w8_l2048_id3_1_cond_3_1;
  reg [34-1:0] _tmp_1159;
  reg _tmp_1160;
  wire [8-1:0] _dataflow_slice_odata_155;
  wire _dataflow_slice_ovalid_155;
  wire _dataflow_slice_oready_155;
  assign _dataflow_slice_oready_155 = (_tmp_1159 > 0) && !_tmp_1160;
  reg _ram_w8_l2048_id3_2_cond_3_1;
  reg [34-1:0] _tmp_1161;
  reg _tmp_1162;
  wire [8-1:0] _dataflow_slice_odata_158;
  wire _dataflow_slice_ovalid_158;
  wire _dataflow_slice_oready_158;
  assign _dataflow_slice_oready_158 = (_tmp_1161 > 0) && !_tmp_1162;
  reg _ram_w8_l2048_id3_3_cond_3_1;
  reg __maxi_read_fsm_cond_3_9_1;
  reg [32-1:0] matmul_29_comp_fsm;
  localparam matmul_29_comp_fsm_init = 0;
  reg [32-1:0] matmul_29_filter_page_comp_offset_buf;
  reg [32-1:0] matmul_29_act_page_comp_offset_buf_0;
  reg [32-1:0] matmul_29_out_page_comp_offset_buf;
  reg [32-1:0] matmul_29_row_count_buf;
  reg [1-1:0] matmul_29_row_select_buf;
  reg [32-1:0] matmul_29_och_count_buf;
  wire matmul_29_stream_pad_mask_0_0;
  assign matmul_29_stream_pad_mask_0_0 = (matmul_29_col_count + 0 < cparam_matmul_29_pad_col_left) || (matmul_29_col_count + 0 >= cparam_matmul_29_act_num_col + cparam_matmul_29_pad_col_left) || (matmul_29_row_count_buf + 0 < cparam_matmul_29_pad_row_top) || (matmul_29_row_count_buf + 0 >= cparam_matmul_29_act_num_row + cparam_matmul_29_pad_row_top);
  reg [1-1:0] matmul_29_stream_pad_masks;
  wire [11-1:0] stream_matmul_29_constant_0_data;
  wire [1-1:0] stream_matmul_29_constant_1_data;
  wire [1-1:0] stream_matmul_29_constant_2_data;
  wire [1-1:0] stream_matmul_29_constant_3_data;
  wire [1-1:0] stream_matmul_29_constant_4_data;
  wire [1-1:0] stream_matmul_29_constant_5_data;
  wire [8-1:0] stream_matmul_29_source_6_data;
  wire [1-1:0] stream_matmul_29_constant_7_data;
  wire [8-1:0] stream_matmul_29_source_8_data;
  wire [1-1:0] stream_matmul_29_constant_9_data;
  wire [8-1:0] stream_matmul_29_source_10_data;
  wire [1-1:0] stream_matmul_29_constant_11_data;
  wire [8-1:0] stream_matmul_29_source_12_data;
  wire [1-1:0] stream_matmul_29_constant_13_data;
  wire [8-1:0] stream_matmul_29_source_14_data;
  wire [1-1:0] stream_matmul_29_constant_15_data;
  wire [1-1:0] stream_matmul_29_constant_16_data;
  wire [4-1:0] stream_matmul_29_constant_17_data;
  wire [2-1:0] stream_matmul_29_constant_18_data;
  wire [8-1:0] stream_matmul_29_source_19_data;
  wire [4-1:0] stream_matmul_29_source_20_data;
  wire [8-1:0] _slice_data_815;
  assign _slice_data_815 = stream_matmul_29_source_6_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_816;
  assign _reinterpretcast_src_816 = _slice_data_815;
  wire signed [8-1:0] _reinterpretcast_data_816;
  assign _reinterpretcast_data_816 = _reinterpretcast_src_816;
  reg signed [8-1:0] _cond_data_817;
  wire [8-1:0] _slice_data_822;
  assign _slice_data_822 = stream_matmul_29_source_8_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_823;
  assign _reinterpretcast_src_823 = _slice_data_822;
  wire signed [8-1:0] _reinterpretcast_data_823;
  assign _reinterpretcast_data_823 = _reinterpretcast_src_823;
  reg signed [8-1:0] _cond_data_824;
  wire [8-1:0] _slice_data_829;
  assign _slice_data_829 = stream_matmul_29_source_10_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_830;
  assign _reinterpretcast_src_830 = _slice_data_829;
  wire [8-1:0] _reinterpretcast_data_830;
  assign _reinterpretcast_data_830 = _reinterpretcast_src_830;
  reg [8-1:0] _cond_data_831;
  wire [8-1:0] _slice_data_836;
  assign _slice_data_836 = stream_matmul_29_source_12_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_837;
  assign _reinterpretcast_src_837 = _slice_data_836;
  wire [8-1:0] _reinterpretcast_data_837;
  assign _reinterpretcast_data_837 = _reinterpretcast_src_837;
  reg [8-1:0] _cond_data_838;
  wire [8-1:0] _slice_data_843;
  assign _slice_data_843 = stream_matmul_29_source_14_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_844;
  assign _reinterpretcast_src_844 = _slice_data_843;
  wire [8-1:0] _reinterpretcast_data_844;
  assign _reinterpretcast_data_844 = _reinterpretcast_src_844;
  reg [8-1:0] _cond_data_845;
  reg [1-1:0] _eq_data_851;
  reg [1-1:0] _eq_data_855;
  wire [4-1:0] _reinterpretcast_src_869;
  assign _reinterpretcast_src_869 = stream_matmul_29_source_20_data;
  wire signed [4-1:0] _reinterpretcast_data_869;
  assign _reinterpretcast_data_869 = _reinterpretcast_src_869;
  wire [1-1:0] _pointer_data_870;
  assign _pointer_data_870 = stream_matmul_29_constant_3_data[1'sd0];
  reg [1-1:0] _eq_data_891;
  reg [1-1:0] _eq_data_894;
  reg [8-1:0] __delay_data_1417;
  reg [1-1:0] __delay_data_1419;
  reg [1-1:0] __delay_data_1422;
  reg signed [4-1:0] __delay_data_1423;
  reg [1-1:0] __delay_data_1429;
  reg [11-1:0] __delay_data_1444;
  reg [4-1:0] __delay_data_1482;
  reg signed [8-1:0] _cond_data_853;
  reg [8-1:0] _plus_data_875;
  reg [8-1:0] _plus_data_880;
  reg [8-1:0] _plus_data_885;
  reg [1-1:0] __delay_data_1418;
  reg [1-1:0] __delay_data_1420;
  reg signed [4-1:0] __delay_data_1424;
  reg [11-1:0] __delay_data_1445;
  reg signed [8-1:0] __delay_data_1460;
  reg signed [8-1:0] __delay_data_1483;
  reg [1-1:0] __delay_data_1529;
  reg [1-1:0] __delay_data_1565;
  reg signed [8-1:0] _cond_data_857;
  reg [1-1:0] __delay_data_1421;
  reg signed [4-1:0] __delay_data_1425;
  reg [8-1:0] __delay_data_1427;
  reg [8-1:0] __delay_data_1430;
  reg [11-1:0] __delay_data_1446;
  reg signed [8-1:0] __delay_data_1461;
  reg signed [8-1:0] __delay_data_1484;
  reg [8-1:0] __delay_data_1506;
  reg [1-1:0] __delay_data_1530;
  reg [1-1:0] __delay_data_1566;
  wire signed [8-1:0] _reinterpretcast_src_863;
  assign _reinterpretcast_src_863 = _cond_data_857;
  wire signed [8-1:0] _reinterpretcast_data_863;
  assign _reinterpretcast_data_863 = _reinterpretcast_src_863;
  reg signed [8-1:0] _cond_data_873;
  reg signed [4-1:0] __delay_data_1426;
  reg [8-1:0] __delay_data_1428;
  reg [8-1:0] __delay_data_1431;
  reg [11-1:0] __delay_data_1447;
  reg signed [8-1:0] __delay_data_1462;
  reg signed [8-1:0] __delay_data_1485;
  reg [8-1:0] __delay_data_1507;
  reg [1-1:0] __delay_data_1531;
  reg [1-1:0] __delay_data_1567;
  reg [8-1:0] __delay_data_1432;
  reg [11-1:0] __delay_data_1448;
  reg signed [8-1:0] __delay_data_1463;
  reg signed [8-1:0] __delay_data_1486;
  reg [8-1:0] __delay_data_1508;
  reg [1-1:0] __delay_data_1532;
  reg [1-1:0] __delay_data_1568;
  reg [8-1:0] __delay_data_1433;
  reg [11-1:0] __delay_data_1449;
  reg signed [8-1:0] __delay_data_1464;
  reg signed [8-1:0] __delay_data_1487;
  reg [8-1:0] __delay_data_1509;
  reg [1-1:0] __delay_data_1533;
  reg [1-1:0] __delay_data_1569;
  reg [8-1:0] __delay_data_1434;
  reg [11-1:0] __delay_data_1450;
  reg signed [8-1:0] __delay_data_1465;
  reg signed [8-1:0] __delay_data_1488;
  reg [8-1:0] __delay_data_1510;
  reg [1-1:0] __delay_data_1534;
  reg [1-1:0] __delay_data_1570;
  reg [8-1:0] __delay_data_1435;
  reg [11-1:0] __delay_data_1451;
  reg signed [8-1:0] __delay_data_1466;
  reg signed [8-1:0] __delay_data_1489;
  reg [8-1:0] __delay_data_1511;
  reg [1-1:0] __delay_data_1535;
  reg [1-1:0] __delay_data_1571;
  reg [8-1:0] __delay_data_1436;
  reg [11-1:0] __delay_data_1452;
  reg signed [8-1:0] __delay_data_1467;
  reg signed [8-1:0] __delay_data_1490;
  reg [8-1:0] __delay_data_1512;
  reg [1-1:0] __delay_data_1536;
  reg [1-1:0] __delay_data_1572;
  reg [8-1:0] __delay_data_1437;
  reg [11-1:0] __delay_data_1453;
  reg signed [8-1:0] __delay_data_1468;
  reg signed [8-1:0] __delay_data_1491;
  reg [8-1:0] __delay_data_1513;
  reg [1-1:0] __delay_data_1537;
  reg [1-1:0] __delay_data_1573;
  reg [8-1:0] __delay_data_1438;
  reg [11-1:0] __delay_data_1454;
  reg signed [8-1:0] __delay_data_1469;
  reg signed [8-1:0] __delay_data_1492;
  reg [8-1:0] __delay_data_1514;
  reg [1-1:0] __delay_data_1538;
  reg [1-1:0] __delay_data_1574;
  reg [8-1:0] __delay_data_1439;
  reg [11-1:0] __delay_data_1455;
  reg signed [8-1:0] __delay_data_1470;
  reg signed [8-1:0] __delay_data_1493;
  reg [8-1:0] __delay_data_1515;
  reg [1-1:0] __delay_data_1539;
  reg [1-1:0] __delay_data_1575;
  reg [8-1:0] __delay_data_1440;
  reg [11-1:0] __delay_data_1456;
  reg signed [8-1:0] __delay_data_1471;
  reg signed [8-1:0] __delay_data_1494;
  reg [8-1:0] __delay_data_1516;
  reg [1-1:0] __delay_data_1540;
  reg [1-1:0] __delay_data_1576;
  reg signed [12-1:0] __substreamoutput_data_876;
  reg [8-1:0] __delay_data_1441;
  reg [11-1:0] __delay_data_1457;
  reg signed [8-1:0] __delay_data_1472;
  reg signed [8-1:0] __delay_data_1495;
  reg [8-1:0] __delay_data_1517;
  reg [1-1:0] __delay_data_1541;
  reg [1-1:0] __delay_data_1577;
  reg signed [32-1:0] __variable_wdata_22;
  assign add_tree_1_var0_data = __variable_wdata_22;
  reg [8-1:0] __delay_data_1442;
  reg [11-1:0] __delay_data_1458;
  reg signed [8-1:0] __delay_data_1473;
  reg signed [8-1:0] __delay_data_1496;
  reg [8-1:0] __delay_data_1518;
  reg [1-1:0] __delay_data_1542;
  reg [1-1:0] __delay_data_1578;
  reg signed [32-1:0] __substreamoutput_data_878;
  reg [8-1:0] __delay_data_1443;
  reg [11-1:0] __delay_data_1459;
  reg signed [8-1:0] __delay_data_1474;
  reg signed [8-1:0] __delay_data_1497;
  reg [8-1:0] __delay_data_1519;
  reg [1-1:0] __delay_data_1543;
  reg [1-1:0] __delay_data_1579;
  reg signed [8-1:0] __delay_data_1475;
  reg signed [8-1:0] __delay_data_1498;
  reg [8-1:0] __delay_data_1520;
  reg [1-1:0] __delay_data_1544;
  reg [1-1:0] __delay_data_1580;
  reg signed [8-1:0] __delay_data_1476;
  reg signed [8-1:0] __delay_data_1499;
  reg [8-1:0] __delay_data_1521;
  reg [1-1:0] __delay_data_1545;
  reg [1-1:0] __delay_data_1581;
  reg signed [8-1:0] __delay_data_1477;
  reg signed [8-1:0] __delay_data_1500;
  reg [8-1:0] __delay_data_1522;
  reg [1-1:0] __delay_data_1546;
  reg [1-1:0] __delay_data_1582;
  reg signed [8-1:0] __delay_data_1478;
  reg signed [8-1:0] __delay_data_1501;
  reg [8-1:0] __delay_data_1523;
  reg [1-1:0] __delay_data_1547;
  reg [1-1:0] __delay_data_1583;
  reg signed [8-1:0] __delay_data_1479;
  reg signed [8-1:0] __delay_data_1502;
  reg [8-1:0] __delay_data_1524;
  reg [1-1:0] __delay_data_1548;
  reg [1-1:0] __delay_data_1584;
  reg signed [8-1:0] __delay_data_1480;
  reg signed [8-1:0] __delay_data_1503;
  reg [8-1:0] __delay_data_1525;
  reg [1-1:0] __delay_data_1549;
  reg [1-1:0] __delay_data_1585;
  reg signed [32-1:0] __substreamoutput_data_881;
  reg [1-1:0] __substreamoutput_data_882;
  reg signed [8-1:0] __delay_data_1481;
  reg signed [8-1:0] __delay_data_1504;
  reg [8-1:0] __delay_data_1526;
  reg [1-1:0] __delay_data_1550;
  reg [1-1:0] __delay_data_1586;
  reg signed [32-1:0] _plus_data_883;
  reg signed [8-1:0] __delay_data_1505;
  reg [8-1:0] __delay_data_1527;
  reg [1-1:0] __delay_data_1551;
  reg [1-1:0] __delay_data_1587;
  reg [1-1:0] __delay_data_1602;
  reg [1-1:0] __delay_data_1552;
  reg [1-1:0] __delay_data_1588;
  reg [1-1:0] __delay_data_1603;
  reg [1-1:0] __delay_data_1553;
  reg [1-1:0] __delay_data_1589;
  reg [1-1:0] __delay_data_1604;
  reg [1-1:0] __delay_data_1554;
  reg [1-1:0] __delay_data_1590;
  reg [1-1:0] __delay_data_1605;
  reg [1-1:0] __delay_data_1555;
  reg [1-1:0] __delay_data_1591;
  reg [1-1:0] __delay_data_1606;
  reg [1-1:0] __delay_data_1556;
  reg [1-1:0] __delay_data_1592;
  reg [1-1:0] __delay_data_1607;
  reg [1-1:0] __delay_data_1557;
  reg [1-1:0] __delay_data_1593;
  reg [1-1:0] __delay_data_1608;
  reg [1-1:0] __delay_data_1558;
  reg [1-1:0] __delay_data_1594;
  reg [1-1:0] __delay_data_1609;
  reg [1-1:0] __delay_data_1559;
  reg [1-1:0] __delay_data_1595;
  reg [1-1:0] __delay_data_1610;
  reg [1-1:0] __delay_data_1560;
  reg [1-1:0] __delay_data_1596;
  reg [1-1:0] __delay_data_1611;
  reg signed [8-1:0] __substreamoutput_data_886;
  reg [1-1:0] __delay_data_1561;
  reg [1-1:0] __delay_data_1597;
  reg [1-1:0] __delay_data_1612;
  reg [1-1:0] _greaterthan_data_888;
  reg signed [8-1:0] __delay_data_1528;
  reg [1-1:0] __delay_data_1562;
  reg [1-1:0] __delay_data_1598;
  reg [1-1:0] __delay_data_1613;
  reg signed [8-1:0] _cond_data_890;
  reg [1-1:0] __delay_data_1563;
  reg signed [8-1:0] __delay_data_1564;
  reg [1-1:0] __delay_data_1599;
  reg [1-1:0] __delay_data_1614;
  reg signed [8-1:0] _cond_data_893;
  reg [1-1:0] __delay_data_1600;
  reg signed [8-1:0] __delay_data_1601;
  reg [1-1:0] __delay_data_1615;
  reg signed [8-1:0] _cond_data_896;
  reg [1-1:0] __delay_data_1616;
  wire signed [8-1:0] _reinterpretcast_src_897;
  assign _reinterpretcast_src_897 = _cond_data_896;
  wire signed [8-1:0] _reinterpretcast_data_897;
  assign _reinterpretcast_data_897 = _reinterpretcast_src_897;
  wire signed [8-1:0] stream_matmul_29_sink_21_data;
  assign stream_matmul_29_sink_21_data = _reinterpretcast_data_897;
  wire [1-1:0] stream_matmul_29_sink_22_data;
  assign stream_matmul_29_sink_22_data = __delay_data_1616;
  reg _set_flag_1163;
  reg [11-1:0] __variable_wdata_796;
  assign stream_matmul_29_constant_0_data = __variable_wdata_796;
  reg _set_flag_1164;
  reg [1-1:0] __variable_wdata_797;
  assign stream_matmul_29_constant_1_data = __variable_wdata_797;
  reg _set_flag_1165;
  reg [1-1:0] __variable_wdata_798;
  assign stream_matmul_29_constant_2_data = __variable_wdata_798;
  reg _set_flag_1166;
  reg [1-1:0] __variable_wdata_799;
  assign stream_matmul_29_constant_3_data = __variable_wdata_799;
  reg _set_flag_1167;
  reg [1-1:0] __variable_wdata_800;
  assign stream_matmul_29_constant_4_data = __variable_wdata_800;
  reg _set_flag_1168;
  reg [1-1:0] __variable_wdata_811;
  assign stream_matmul_29_constant_5_data = __variable_wdata_811;
  reg [32-1:0] _source_stream_matmul_29_source_6_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_29_source_6_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_29_source_6_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_29_source_6_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_29_source_6_pat_size_0;
  reg [33-1:0] _source_stream_matmul_29_source_6_pat_size_1;
  reg [33-1:0] _source_stream_matmul_29_source_6_pat_size_2;
  reg [33-1:0] _source_stream_matmul_29_source_6_pat_size_3;
  reg [32-1:0] _source_stream_matmul_29_source_6_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_29_source_6_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_29_source_6_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_29_source_6_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_29_source_6_pat_count_0;
  reg [33-1:0] _source_stream_matmul_29_source_6_pat_count_1;
  reg [33-1:0] _source_stream_matmul_29_source_6_pat_count_2;
  reg [33-1:0] _source_stream_matmul_29_source_6_pat_count_3;
  reg [33-1:0] _source_stream_matmul_29_source_6_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_29_source_6_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_29_source_6_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_29_source_6_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_29_source_6_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_29_source_6_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_29_source_6_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_29_source_6_pat_stride_buf_3;
  reg _set_flag_1169;
  wire [2-1:0] _tmp_1170;
  assign _tmp_1170 = _stream_matmul_29_source_6_source_ram_raddr;
  reg [2-1:0] __tmp_1170_1;
  reg [2-1:0] __tmp_1170_2;
  reg _tmp_1171;
  reg _ram_w8_l2048_id2_0_cond_5_1;
  reg _ram_w8_l2048_id2_0_cond_6_1;
  reg _ram_w8_l2048_id2_0_cond_6_2;
  reg _tmp_1172;
  reg _ram_w8_l2048_id2_1_cond_5_1;
  reg _ram_w8_l2048_id2_1_cond_6_1;
  reg _ram_w8_l2048_id2_1_cond_6_2;
  reg _tmp_1173;
  reg _ram_w8_l2048_id2_2_cond_5_1;
  reg _ram_w8_l2048_id2_2_cond_6_1;
  reg _ram_w8_l2048_id2_2_cond_6_2;
  reg _tmp_1174;
  reg _ram_w8_l2048_id2_3_cond_5_1;
  reg _ram_w8_l2048_id2_3_cond_6_1;
  reg _ram_w8_l2048_id2_3_cond_6_2;
  wire signed [8-1:0] _tmp_1175;
  wire _tmp_1176;
  assign _tmp_1175 = (__tmp_1170_2 == 0)? ram_w8_l2048_id2_0_0_rdata : 
                     (__tmp_1170_2 == 1)? ram_w8_l2048_id2_1_0_rdata : 
                     (__tmp_1170_2 == 2)? ram_w8_l2048_id2_2_0_rdata : 
                     (__tmp_1170_2 == 3)? ram_w8_l2048_id2_3_0_rdata : 0;
  assign _tmp_1176 = _tmp_1171;
  assign _stream_matmul_29_source_6_source_ram_rdata = (_stream_matmul_29_source_6_source_ram_sel == 1)? _tmp_1175 : 0;
  localparam _tmp_1177 = 1;
  wire [_tmp_1177-1:0] _tmp_1178;
  assign _tmp_1178 = _stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1);
  reg [_tmp_1177-1:0] __tmp_1178_1;
  reg [8-1:0] __variable_wdata_812;
  assign stream_matmul_29_source_6_data = __variable_wdata_812;
  reg [32-1:0] _stream_matmul_29_source_6_source_pat_fsm_0;
  localparam _stream_matmul_29_source_6_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_matmul_29_source_6_source_pat_all_offset;
  assign _stream_matmul_29_source_6_source_pat_all_offset = _stream_matmul_29_source_6_source_offset_buf + _source_stream_matmul_29_source_6_pat_cur_offset_0 + _source_stream_matmul_29_source_6_pat_cur_offset_1 + _source_stream_matmul_29_source_6_pat_cur_offset_2 + _source_stream_matmul_29_source_6_pat_cur_offset_3;
  reg _set_flag_1179;
  reg [1-1:0] __variable_wdata_818;
  assign stream_matmul_29_constant_7_data = __variable_wdata_818;
  reg [32-1:0] _source_stream_matmul_29_source_8_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_29_source_8_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_29_source_8_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_29_source_8_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_29_source_8_pat_size_0;
  reg [33-1:0] _source_stream_matmul_29_source_8_pat_size_1;
  reg [33-1:0] _source_stream_matmul_29_source_8_pat_size_2;
  reg [33-1:0] _source_stream_matmul_29_source_8_pat_size_3;
  reg [32-1:0] _source_stream_matmul_29_source_8_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_29_source_8_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_29_source_8_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_29_source_8_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_29_source_8_pat_count_0;
  reg [33-1:0] _source_stream_matmul_29_source_8_pat_count_1;
  reg [33-1:0] _source_stream_matmul_29_source_8_pat_count_2;
  reg [33-1:0] _source_stream_matmul_29_source_8_pat_count_3;
  reg [33-1:0] _source_stream_matmul_29_source_8_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_29_source_8_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_29_source_8_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_29_source_8_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_29_source_8_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_29_source_8_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_29_source_8_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_29_source_8_pat_stride_buf_3;
  reg _set_flag_1180;
  wire [2-1:0] _tmp_1181;
  assign _tmp_1181 = _stream_matmul_29_source_8_source_ram_raddr;
  reg [2-1:0] __tmp_1181_1;
  reg [2-1:0] __tmp_1181_2;
  reg _tmp_1182;
  reg _ram_w8_l2048_id0_0_cond_4_1;
  reg _ram_w8_l2048_id0_0_cond_5_1;
  reg _ram_w8_l2048_id0_0_cond_5_2;
  reg _tmp_1183;
  reg _ram_w8_l2048_id0_1_cond_4_1;
  reg _ram_w8_l2048_id0_1_cond_5_1;
  reg _ram_w8_l2048_id0_1_cond_5_2;
  reg _tmp_1184;
  reg _ram_w8_l2048_id0_2_cond_4_1;
  reg _ram_w8_l2048_id0_2_cond_5_1;
  reg _ram_w8_l2048_id0_2_cond_5_2;
  reg _tmp_1185;
  reg _ram_w8_l2048_id0_3_cond_4_1;
  reg _ram_w8_l2048_id0_3_cond_5_1;
  reg _ram_w8_l2048_id0_3_cond_5_2;
  wire signed [8-1:0] _tmp_1186;
  wire _tmp_1187;
  assign _tmp_1186 = (__tmp_1181_2 == 0)? ram_w8_l2048_id0_0_0_rdata : 
                     (__tmp_1181_2 == 1)? ram_w8_l2048_id0_1_0_rdata : 
                     (__tmp_1181_2 == 2)? ram_w8_l2048_id0_2_0_rdata : 
                     (__tmp_1181_2 == 3)? ram_w8_l2048_id0_3_0_rdata : 0;
  assign _tmp_1187 = _tmp_1182;
  assign _stream_matmul_29_source_8_source_ram_rdata = (_stream_matmul_29_source_8_source_ram_sel == 2)? _tmp_1186 : 0;
  localparam _tmp_1188 = 1;
  wire [_tmp_1188-1:0] _tmp_1189;
  assign _tmp_1189 = _stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2);
  reg [_tmp_1188-1:0] __tmp_1189_1;
  reg [8-1:0] __variable_wdata_819;
  assign stream_matmul_29_source_8_data = __variable_wdata_819;
  reg [32-1:0] _stream_matmul_29_source_8_source_pat_fsm_1;
  localparam _stream_matmul_29_source_8_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_matmul_29_source_8_source_pat_all_offset;
  assign _stream_matmul_29_source_8_source_pat_all_offset = _stream_matmul_29_source_8_source_offset_buf + _source_stream_matmul_29_source_8_pat_cur_offset_0 + _source_stream_matmul_29_source_8_pat_cur_offset_1 + _source_stream_matmul_29_source_8_pat_cur_offset_2 + _source_stream_matmul_29_source_8_pat_cur_offset_3;
  reg _set_flag_1190;
  reg [1-1:0] __variable_wdata_825;
  assign stream_matmul_29_constant_9_data = __variable_wdata_825;
  reg _set_flag_1191;
  reg [8-1:0] __variable_wdata_826;
  assign stream_matmul_29_source_10_data = __variable_wdata_826;
  reg _set_flag_1192;
  reg [1-1:0] __variable_wdata_832;
  assign stream_matmul_29_constant_11_data = __variable_wdata_832;
  reg _set_flag_1193;
  reg [8-1:0] __variable_wdata_833;
  assign stream_matmul_29_source_12_data = __variable_wdata_833;
  reg _set_flag_1194;
  reg [1-1:0] __variable_wdata_839;
  assign stream_matmul_29_constant_13_data = __variable_wdata_839;
  reg _set_flag_1195;
  reg [8-1:0] __variable_wdata_840;
  assign stream_matmul_29_source_14_data = __variable_wdata_840;
  reg _set_flag_1196;
  reg [1-1:0] __variable_wdata_846;
  assign stream_matmul_29_constant_15_data = __variable_wdata_846;
  reg _set_flag_1197;
  reg [1-1:0] __variable_wdata_847;
  assign stream_matmul_29_constant_16_data = __variable_wdata_847;
  reg _set_flag_1198;
  reg [4-1:0] __variable_wdata_848;
  assign stream_matmul_29_constant_17_data = __variable_wdata_848;
  reg _set_flag_1199;
  reg [2-1:0] __variable_wdata_849;
  assign stream_matmul_29_constant_18_data = __variable_wdata_849;
  reg [32-1:0] _source_stream_matmul_29_source_19_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_29_source_19_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_29_source_19_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_29_source_19_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_29_source_19_pat_size_0;
  reg [33-1:0] _source_stream_matmul_29_source_19_pat_size_1;
  reg [33-1:0] _source_stream_matmul_29_source_19_pat_size_2;
  reg [33-1:0] _source_stream_matmul_29_source_19_pat_size_3;
  reg [32-1:0] _source_stream_matmul_29_source_19_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_29_source_19_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_29_source_19_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_29_source_19_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_29_source_19_pat_count_0;
  reg [33-1:0] _source_stream_matmul_29_source_19_pat_count_1;
  reg [33-1:0] _source_stream_matmul_29_source_19_pat_count_2;
  reg [33-1:0] _source_stream_matmul_29_source_19_pat_count_3;
  reg [33-1:0] _source_stream_matmul_29_source_19_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_29_source_19_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_29_source_19_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_29_source_19_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_29_source_19_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_29_source_19_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_29_source_19_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_29_source_19_pat_stride_buf_3;
  reg _set_flag_1200;
  wire [2-1:0] _tmp_1201;
  assign _tmp_1201 = _stream_matmul_29_source_19_source_ram_raddr;
  reg [2-1:0] __tmp_1201_1;
  reg [2-1:0] __tmp_1201_2;
  reg _tmp_1202;
  reg _ram_w8_l2048_id3_0_cond_4_1;
  reg _ram_w8_l2048_id3_0_cond_5_1;
  reg _ram_w8_l2048_id3_0_cond_5_2;
  reg _tmp_1203;
  reg _ram_w8_l2048_id3_1_cond_4_1;
  reg _ram_w8_l2048_id3_1_cond_5_1;
  reg _ram_w8_l2048_id3_1_cond_5_2;
  reg _tmp_1204;
  reg _ram_w8_l2048_id3_2_cond_4_1;
  reg _ram_w8_l2048_id3_2_cond_5_1;
  reg _ram_w8_l2048_id3_2_cond_5_2;
  reg _tmp_1205;
  reg _ram_w8_l2048_id3_3_cond_4_1;
  reg _ram_w8_l2048_id3_3_cond_5_1;
  reg _ram_w8_l2048_id3_3_cond_5_2;
  wire signed [8-1:0] _tmp_1206;
  wire _tmp_1207;
  assign _tmp_1206 = (__tmp_1201_2 == 0)? ram_w8_l2048_id3_0_0_rdata : 
                     (__tmp_1201_2 == 1)? ram_w8_l2048_id3_1_0_rdata : 
                     (__tmp_1201_2 == 2)? ram_w8_l2048_id3_2_0_rdata : 
                     (__tmp_1201_2 == 3)? ram_w8_l2048_id3_3_0_rdata : 0;
  assign _tmp_1207 = _tmp_1202;
  assign _stream_matmul_29_source_19_source_ram_rdata = (_stream_matmul_29_source_19_source_ram_sel == 3)? _tmp_1206 : 0;
  localparam _tmp_1208 = 1;
  wire [_tmp_1208-1:0] _tmp_1209;
  assign _tmp_1209 = _stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3);
  reg [_tmp_1208-1:0] __tmp_1209_1;
  reg [8-1:0] __variable_wdata_850;
  assign stream_matmul_29_source_19_data = __variable_wdata_850;
  reg [32-1:0] _stream_matmul_29_source_19_source_pat_fsm_2;
  localparam _stream_matmul_29_source_19_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_matmul_29_source_19_source_pat_all_offset;
  assign _stream_matmul_29_source_19_source_pat_all_offset = _stream_matmul_29_source_19_source_offset_buf + _source_stream_matmul_29_source_19_pat_cur_offset_0 + _source_stream_matmul_29_source_19_pat_cur_offset_1 + _source_stream_matmul_29_source_19_pat_cur_offset_2 + _source_stream_matmul_29_source_19_pat_cur_offset_3;
  reg [32-1:0] _source_stream_matmul_29_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_29_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_29_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_29_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_29_source_20_pat_size_0;
  reg [33-1:0] _source_stream_matmul_29_source_20_pat_size_1;
  reg [33-1:0] _source_stream_matmul_29_source_20_pat_size_2;
  reg [33-1:0] _source_stream_matmul_29_source_20_pat_size_3;
  reg [32-1:0] _source_stream_matmul_29_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_29_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_29_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_29_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_29_source_20_pat_count_0;
  reg [33-1:0] _source_stream_matmul_29_source_20_pat_count_1;
  reg [33-1:0] _source_stream_matmul_29_source_20_pat_count_2;
  reg [33-1:0] _source_stream_matmul_29_source_20_pat_count_3;
  reg [33-1:0] _source_stream_matmul_29_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_29_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_29_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_29_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_29_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_29_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_29_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_29_source_20_pat_stride_buf_3;
  reg _set_flag_1210;
  wire [3-1:0] _tmp_1211;
  assign _tmp_1211 = _stream_matmul_29_source_20_source_ram_raddr;
  reg [3-1:0] __tmp_1211_1;
  reg [3-1:0] __tmp_1211_2;
  reg _tmp_1212;
  reg _ram_w4_l8192_id0_0_cond_5_1;
  reg _ram_w4_l8192_id0_0_cond_6_1;
  reg _ram_w4_l8192_id0_0_cond_6_2;
  reg _tmp_1213;
  reg _ram_w4_l8192_id0_1_cond_5_1;
  reg _ram_w4_l8192_id0_1_cond_6_1;
  reg _ram_w4_l8192_id0_1_cond_6_2;
  reg _tmp_1214;
  reg _ram_w4_l8192_id0_2_cond_5_1;
  reg _ram_w4_l8192_id0_2_cond_6_1;
  reg _ram_w4_l8192_id0_2_cond_6_2;
  reg _tmp_1215;
  reg _ram_w4_l8192_id0_3_cond_5_1;
  reg _ram_w4_l8192_id0_3_cond_6_1;
  reg _ram_w4_l8192_id0_3_cond_6_2;
  reg _tmp_1216;
  reg _ram_w4_l8192_id0_4_cond_5_1;
  reg _ram_w4_l8192_id0_4_cond_6_1;
  reg _ram_w4_l8192_id0_4_cond_6_2;
  reg _tmp_1217;
  reg _ram_w4_l8192_id0_5_cond_5_1;
  reg _ram_w4_l8192_id0_5_cond_6_1;
  reg _ram_w4_l8192_id0_5_cond_6_2;
  reg _tmp_1218;
  reg _ram_w4_l8192_id0_6_cond_5_1;
  reg _ram_w4_l8192_id0_6_cond_6_1;
  reg _ram_w4_l8192_id0_6_cond_6_2;
  reg _tmp_1219;
  reg _ram_w4_l8192_id0_7_cond_5_1;
  reg _ram_w4_l8192_id0_7_cond_6_1;
  reg _ram_w4_l8192_id0_7_cond_6_2;
  wire signed [4-1:0] _tmp_1220;
  wire _tmp_1221;
  assign _tmp_1220 = (__tmp_1211_2 == 0)? ram_w4_l8192_id0_0_0_rdata : 
                     (__tmp_1211_2 == 1)? ram_w4_l8192_id0_1_0_rdata : 
                     (__tmp_1211_2 == 2)? ram_w4_l8192_id0_2_0_rdata : 
                     (__tmp_1211_2 == 3)? ram_w4_l8192_id0_3_0_rdata : 
                     (__tmp_1211_2 == 4)? ram_w4_l8192_id0_4_0_rdata : 
                     (__tmp_1211_2 == 5)? ram_w4_l8192_id0_5_0_rdata : 
                     (__tmp_1211_2 == 6)? ram_w4_l8192_id0_6_0_rdata : 
                     (__tmp_1211_2 == 7)? ram_w4_l8192_id0_7_0_rdata : 0;
  assign _tmp_1221 = _tmp_1212;
  assign _stream_matmul_29_source_20_source_ram_rdata = (_stream_matmul_29_source_20_source_ram_sel == 4)? _tmp_1220 : 0;
  localparam _tmp_1222 = 1;
  wire [_tmp_1222-1:0] _tmp_1223;
  assign _tmp_1223 = _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
  reg [_tmp_1222-1:0] __tmp_1223_1;
  reg [4-1:0] __variable_wdata_864;
  assign stream_matmul_29_source_20_data = __variable_wdata_864;
  reg [32-1:0] _stream_matmul_29_source_20_source_pat_fsm_3;
  localparam _stream_matmul_29_source_20_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_matmul_29_source_20_source_pat_all_offset;
  assign _stream_matmul_29_source_20_source_pat_all_offset = _stream_matmul_29_source_20_source_offset_buf + _source_stream_matmul_29_source_20_pat_cur_offset_0 + _source_stream_matmul_29_source_20_pat_cur_offset_1 + _source_stream_matmul_29_source_20_pat_cur_offset_2 + _source_stream_matmul_29_source_20_pat_cur_offset_3;
  reg _set_flag_1224;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_1;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_2;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_3;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_4;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_5;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_6;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_7;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_8;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_9;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_10;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_11;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_12;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_13;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_14;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_15;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_16;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_17;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_18;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_19;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_20;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_21;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_22;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_23;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_24;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_25;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_26;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_27;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_28;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_29;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_30;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_31;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_32;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_33;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_34;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_35;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_36;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_37;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_38;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_39;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_40;
  reg [32-1:0] __stream_matmul_29_sink_21_sink_offset_0_41;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_1;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_2;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_3;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_4;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_5;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_6;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_7;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_8;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_9;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_10;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_11;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_12;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_13;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_14;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_15;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_16;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_17;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_18;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_19;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_20;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_21;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_22;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_23;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_24;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_25;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_26;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_27;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_28;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_29;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_30;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_31;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_32;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_33;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_34;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_35;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_36;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_37;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_38;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_39;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_40;
  reg [33-1:0] __stream_matmul_29_sink_21_sink_size_1_41;
  reg __stream_seq_16_cond_2_1;
  reg __stream_seq_16_cond_2_2;
  reg __stream_seq_16_cond_2_3;
  reg __stream_seq_16_cond_2_4;
  reg __stream_seq_16_cond_2_5;
  reg __stream_seq_16_cond_2_6;
  reg __stream_seq_16_cond_2_7;
  reg __stream_seq_16_cond_2_8;
  reg __stream_seq_16_cond_2_9;
  reg __stream_seq_16_cond_2_10;
  reg __stream_seq_16_cond_2_11;
  reg __stream_seq_16_cond_2_12;
  reg __stream_seq_16_cond_2_13;
  reg __stream_seq_16_cond_2_14;
  reg __stream_seq_16_cond_2_15;
  reg __stream_seq_16_cond_2_16;
  reg __stream_seq_16_cond_2_17;
  reg __stream_seq_16_cond_2_18;
  reg __stream_seq_16_cond_2_19;
  reg __stream_seq_16_cond_2_20;
  reg __stream_seq_16_cond_2_21;
  reg __stream_seq_16_cond_2_22;
  reg __stream_seq_16_cond_2_23;
  reg __stream_seq_16_cond_2_24;
  reg __stream_seq_16_cond_2_25;
  reg __stream_seq_16_cond_2_26;
  reg __stream_seq_16_cond_2_27;
  reg __stream_seq_16_cond_2_28;
  reg __stream_seq_16_cond_2_29;
  reg __stream_seq_16_cond_2_30;
  reg __stream_seq_16_cond_2_31;
  reg __stream_seq_16_cond_2_32;
  reg __stream_seq_16_cond_2_33;
  reg __stream_seq_16_cond_2_34;
  reg __stream_seq_16_cond_2_35;
  reg __stream_seq_16_cond_2_36;
  reg __stream_seq_16_cond_2_37;
  reg __stream_seq_16_cond_2_38;
  reg __stream_seq_16_cond_2_39;
  reg __stream_seq_16_cond_2_40;
  reg __stream_seq_16_cond_2_41;
  reg __set_flag_1224_1;
  reg __set_flag_1224_2;
  reg __set_flag_1224_3;
  reg __set_flag_1224_4;
  reg __set_flag_1224_5;
  reg __set_flag_1224_6;
  reg __set_flag_1224_7;
  reg __set_flag_1224_8;
  reg __set_flag_1224_9;
  reg __set_flag_1224_10;
  reg __set_flag_1224_11;
  reg __set_flag_1224_12;
  reg __set_flag_1224_13;
  reg __set_flag_1224_14;
  reg __set_flag_1224_15;
  reg __set_flag_1224_16;
  reg __set_flag_1224_17;
  reg __set_flag_1224_18;
  reg __set_flag_1224_19;
  reg __set_flag_1224_20;
  reg __set_flag_1224_21;
  reg __set_flag_1224_22;
  reg __set_flag_1224_23;
  reg __set_flag_1224_24;
  reg __set_flag_1224_25;
  reg __set_flag_1224_26;
  reg __set_flag_1224_27;
  reg __set_flag_1224_28;
  reg __set_flag_1224_29;
  reg __set_flag_1224_30;
  reg __set_flag_1224_31;
  reg __set_flag_1224_32;
  reg __set_flag_1224_33;
  reg __set_flag_1224_34;
  reg __set_flag_1224_35;
  reg __set_flag_1224_36;
  reg __set_flag_1224_37;
  reg __set_flag_1224_38;
  reg __set_flag_1224_39;
  reg __set_flag_1224_40;
  reg __set_flag_1224_41;
  wire [2-1:0] _tmp_1225;
  assign _tmp_1225 = _stream_matmul_29_sink_21_sink_waddr;
  reg _ram_w8_l2048_id1_0_cond_5_1;
  reg _ram_w8_l2048_id1_1_cond_5_1;
  reg _ram_w8_l2048_id1_2_cond_5_1;
  reg _ram_w8_l2048_id1_3_cond_5_1;
  reg __stream_matmul_29_start_1;
  reg __stream_matmul_29_start_2;
  reg __stream_matmul_29_start_3;
  reg __stream_matmul_29_start_4;
  reg __stream_matmul_29_start_5;
  reg __stream_matmul_29_start_6;
  reg __stream_matmul_29_start_7;
  reg __stream_matmul_29_start_8;
  reg __stream_matmul_29_start_9;
  reg __stream_matmul_29_start_10;
  reg __stream_matmul_29_start_11;
  reg __stream_matmul_29_start_12;
  reg __stream_matmul_29_start_13;
  reg __stream_matmul_29_start_14;
  reg __stream_matmul_29_start_15;
  reg __stream_matmul_29_start_16;
  reg __stream_matmul_29_start_17;
  reg __stream_matmul_29_start_18;
  reg __stream_matmul_29_start_19;
  reg __stream_matmul_29_start_20;
  reg __stream_matmul_29_start_21;
  reg __stream_matmul_29_start_22;
  reg __stream_matmul_29_start_23;
  reg __stream_matmul_29_start_24;
  reg __stream_matmul_29_start_25;
  reg __stream_matmul_29_start_26;
  reg __stream_matmul_29_start_27;
  reg __stream_matmul_29_start_28;
  reg __stream_matmul_29_start_29;
  reg __stream_matmul_29_start_30;
  reg __stream_matmul_29_start_31;
  reg __stream_matmul_29_start_32;
  reg __stream_matmul_29_start_33;
  reg __stream_matmul_29_start_34;
  reg __stream_matmul_29_start_35;
  reg __stream_matmul_29_start_36;
  reg __stream_matmul_29_start_37;
  reg __stream_matmul_29_start_38;
  reg __stream_matmul_29_start_39;
  reg __stream_matmul_29_start_40;
  reg __stream_matmul_29_start_41;
  reg __stream_matmul_29_start_42;
  reg [32-1:0] _stream_matmul_29_sink_21_sink_fsm_4;
  localparam _stream_matmul_29_sink_21_sink_fsm_4_init = 0;
  assign _stream_matmul_29_start_flag = ((matmul_29_comp_fsm == 4) && !_stream_matmul_29_source_busy)? 1 : 0;
  localparam _tmp_1226 = 1;
  wire [_tmp_1226-1:0] _tmp_1227;
  assign _tmp_1227 = (_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag;
  reg [_tmp_1226-1:0] __tmp_1227_1;
  reg [_tmp_1226-1:0] __tmp_1227_2;
  reg [_tmp_1226-1:0] __tmp_1227_3;
  reg [_tmp_1226-1:0] __tmp_1227_4;
  reg [_tmp_1226-1:0] __tmp_1227_5;
  localparam _tmp_1228 = 1;
  wire [_tmp_1228-1:0] _tmp_1229;
  assign _tmp_1229 = (_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag;
  reg [_tmp_1228-1:0] __tmp_1229_1;
  reg [_tmp_1228-1:0] __tmp_1229_2;
  reg [_tmp_1228-1:0] __tmp_1229_3;
  reg [_tmp_1228-1:0] __tmp_1229_4;
  reg [_tmp_1228-1:0] __tmp_1229_5;
  reg [_tmp_1228-1:0] __tmp_1229_6;
  reg [_tmp_1228-1:0] __tmp_1229_7;
  reg [_tmp_1228-1:0] __tmp_1229_8;
  localparam _tmp_1230 = 1;
  wire [_tmp_1230-1:0] _tmp_1231;
  assign _tmp_1231 = (_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag;
  reg [_tmp_1230-1:0] __tmp_1231_1;
  reg [_tmp_1230-1:0] __tmp_1231_2;
  reg [_tmp_1230-1:0] __tmp_1231_3;
  reg [_tmp_1230-1:0] __tmp_1231_4;
  reg [_tmp_1230-1:0] __tmp_1231_5;
  reg [_tmp_1230-1:0] __tmp_1231_6;
  reg [_tmp_1230-1:0] __tmp_1231_7;
  reg [_tmp_1230-1:0] __tmp_1231_8;
  localparam _tmp_1232 = 1;
  wire [_tmp_1232-1:0] _tmp_1233;
  assign _tmp_1233 = (_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag;
  reg [_tmp_1232-1:0] __tmp_1233_1;
  reg [_tmp_1232-1:0] __tmp_1233_2;
  reg [_tmp_1232-1:0] __tmp_1233_3;
  reg [_tmp_1232-1:0] __tmp_1233_4;
  reg [_tmp_1232-1:0] __tmp_1233_5;
  reg [_tmp_1232-1:0] __tmp_1233_6;
  reg [_tmp_1232-1:0] __tmp_1233_7;
  reg [_tmp_1232-1:0] __tmp_1233_8;
  localparam _tmp_1234 = 1;
  wire [_tmp_1234-1:0] _tmp_1235;
  assign _tmp_1235 = (_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag;
  reg [_tmp_1234-1:0] __tmp_1235_1;
  reg [_tmp_1234-1:0] __tmp_1235_2;
  reg [_tmp_1234-1:0] __tmp_1235_3;
  reg [_tmp_1234-1:0] __tmp_1235_4;
  reg [_tmp_1234-1:0] __tmp_1235_5;
  reg [_tmp_1234-1:0] __tmp_1235_6;
  reg [_tmp_1234-1:0] __tmp_1235_7;
  reg [_tmp_1234-1:0] __tmp_1235_8;
  reg [_tmp_1234-1:0] __tmp_1235_9;
  reg [_tmp_1234-1:0] __tmp_1235_10;
  reg [_tmp_1234-1:0] __tmp_1235_11;
  reg [_tmp_1234-1:0] __tmp_1235_12;
  reg [_tmp_1234-1:0] __tmp_1235_13;
  reg [_tmp_1234-1:0] __tmp_1235_14;
  reg [_tmp_1234-1:0] __tmp_1235_15;
  reg [_tmp_1234-1:0] __tmp_1235_16;
  reg [_tmp_1234-1:0] __tmp_1235_17;
  reg [_tmp_1234-1:0] __tmp_1235_18;
  localparam _tmp_1236 = 1;
  wire [_tmp_1236-1:0] _tmp_1237;
  assign _tmp_1237 = (_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag;
  reg [_tmp_1236-1:0] __tmp_1237_1;
  reg [_tmp_1236-1:0] __tmp_1237_2;
  reg [_tmp_1236-1:0] __tmp_1237_3;
  reg [_tmp_1236-1:0] __tmp_1237_4;
  reg [_tmp_1236-1:0] __tmp_1237_5;
  reg [_tmp_1236-1:0] __tmp_1237_6;
  reg [_tmp_1236-1:0] __tmp_1237_7;
  reg [_tmp_1236-1:0] __tmp_1237_8;
  reg [_tmp_1236-1:0] __tmp_1237_9;
  reg [_tmp_1236-1:0] __tmp_1237_10;
  reg [_tmp_1236-1:0] __tmp_1237_11;
  reg [_tmp_1236-1:0] __tmp_1237_12;
  reg [_tmp_1236-1:0] __tmp_1237_13;
  reg [_tmp_1236-1:0] __tmp_1237_14;
  reg [_tmp_1236-1:0] __tmp_1237_15;
  reg [_tmp_1236-1:0] __tmp_1237_16;
  reg [_tmp_1236-1:0] __tmp_1237_17;
  reg [_tmp_1236-1:0] __tmp_1237_18;
  reg [_tmp_1236-1:0] __tmp_1237_19;
  reg [_tmp_1236-1:0] __tmp_1237_20;
  reg [_tmp_1236-1:0] __tmp_1237_21;
  reg [_tmp_1236-1:0] __tmp_1237_22;
  localparam _tmp_1238 = 1;
  wire [_tmp_1238-1:0] _tmp_1239;
  assign _tmp_1239 = (_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag;
  reg [_tmp_1238-1:0] __tmp_1239_1;
  reg [_tmp_1238-1:0] __tmp_1239_2;
  reg [_tmp_1238-1:0] __tmp_1239_3;
  reg [_tmp_1238-1:0] __tmp_1239_4;
  reg [_tmp_1238-1:0] __tmp_1239_5;
  reg [_tmp_1238-1:0] __tmp_1239_6;
  reg [_tmp_1238-1:0] __tmp_1239_7;
  reg [_tmp_1238-1:0] __tmp_1239_8;
  reg [_tmp_1238-1:0] __tmp_1239_9;
  reg [_tmp_1238-1:0] __tmp_1239_10;
  reg [_tmp_1238-1:0] __tmp_1239_11;
  reg [_tmp_1238-1:0] __tmp_1239_12;
  reg [_tmp_1238-1:0] __tmp_1239_13;
  reg [_tmp_1238-1:0] __tmp_1239_14;
  reg [_tmp_1238-1:0] __tmp_1239_15;
  reg [_tmp_1238-1:0] __tmp_1239_16;
  reg [_tmp_1238-1:0] __tmp_1239_17;
  reg [_tmp_1238-1:0] __tmp_1239_18;
  reg [_tmp_1238-1:0] __tmp_1239_19;
  reg [_tmp_1238-1:0] __tmp_1239_20;
  localparam _tmp_1240 = 1;
  wire [_tmp_1240-1:0] _tmp_1241;
  assign _tmp_1241 = (_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag;
  reg [_tmp_1240-1:0] __tmp_1241_1;
  reg [_tmp_1240-1:0] __tmp_1241_2;
  reg [_tmp_1240-1:0] __tmp_1241_3;
  reg [_tmp_1240-1:0] __tmp_1241_4;
  reg [_tmp_1240-1:0] __tmp_1241_5;
  reg [_tmp_1240-1:0] __tmp_1241_6;
  reg [_tmp_1240-1:0] __tmp_1241_7;
  reg [_tmp_1240-1:0] __tmp_1241_8;
  reg [_tmp_1240-1:0] __tmp_1241_9;
  reg [_tmp_1240-1:0] __tmp_1241_10;
  reg [_tmp_1240-1:0] __tmp_1241_11;
  reg [_tmp_1240-1:0] __tmp_1241_12;
  reg [_tmp_1240-1:0] __tmp_1241_13;
  reg [_tmp_1240-1:0] __tmp_1241_14;
  reg [_tmp_1240-1:0] __tmp_1241_15;
  reg [_tmp_1240-1:0] __tmp_1241_16;
  reg [_tmp_1240-1:0] __tmp_1241_17;
  reg [_tmp_1240-1:0] __tmp_1241_18;
  reg [_tmp_1240-1:0] __tmp_1241_19;
  reg [_tmp_1240-1:0] __tmp_1241_20;
  localparam _tmp_1242 = 1;
  wire [_tmp_1242-1:0] _tmp_1243;
  assign _tmp_1243 = (_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag;
  reg [_tmp_1242-1:0] __tmp_1243_1;
  reg [_tmp_1242-1:0] __tmp_1243_2;
  reg [_tmp_1242-1:0] __tmp_1243_3;
  reg [_tmp_1242-1:0] __tmp_1243_4;
  reg [_tmp_1242-1:0] __tmp_1243_5;
  reg [_tmp_1242-1:0] __tmp_1243_6;
  reg [_tmp_1242-1:0] __tmp_1243_7;
  reg [_tmp_1242-1:0] __tmp_1243_8;
  reg [_tmp_1242-1:0] __tmp_1243_9;
  reg [_tmp_1242-1:0] __tmp_1243_10;
  reg [_tmp_1242-1:0] __tmp_1243_11;
  reg [_tmp_1242-1:0] __tmp_1243_12;
  reg [_tmp_1242-1:0] __tmp_1243_13;
  reg [_tmp_1242-1:0] __tmp_1243_14;
  reg [_tmp_1242-1:0] __tmp_1243_15;
  reg [_tmp_1242-1:0] __tmp_1243_16;
  reg [_tmp_1242-1:0] __tmp_1243_17;
  reg [_tmp_1242-1:0] __tmp_1243_18;
  reg [_tmp_1242-1:0] __tmp_1243_19;
  reg [_tmp_1242-1:0] __tmp_1243_20;
  localparam _tmp_1244 = 1;
  wire [_tmp_1244-1:0] _tmp_1245;
  assign _tmp_1245 = (_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag;
  reg [_tmp_1244-1:0] __tmp_1245_1;
  reg [_tmp_1244-1:0] __tmp_1245_2;
  reg [_tmp_1244-1:0] __tmp_1245_3;
  reg [_tmp_1244-1:0] __tmp_1245_4;
  reg [_tmp_1244-1:0] __tmp_1245_5;
  reg [_tmp_1244-1:0] __tmp_1245_6;
  reg [_tmp_1244-1:0] __tmp_1245_7;
  reg [_tmp_1244-1:0] __tmp_1245_8;
  reg [_tmp_1244-1:0] __tmp_1245_9;
  reg [_tmp_1244-1:0] __tmp_1245_10;
  reg [_tmp_1244-1:0] __tmp_1245_11;
  reg [_tmp_1244-1:0] __tmp_1245_12;
  reg [_tmp_1244-1:0] __tmp_1245_13;
  reg [_tmp_1244-1:0] __tmp_1245_14;
  reg [_tmp_1244-1:0] __tmp_1245_15;
  reg [_tmp_1244-1:0] __tmp_1245_16;
  reg [_tmp_1244-1:0] __tmp_1245_17;
  reg [_tmp_1244-1:0] __tmp_1245_18;
  reg [_tmp_1244-1:0] __tmp_1245_19;
  reg [_tmp_1244-1:0] __tmp_1245_20;
  reg [_tmp_1244-1:0] __tmp_1245_21;
  reg [_tmp_1244-1:0] __tmp_1245_22;
  reg [_tmp_1244-1:0] __tmp_1245_23;
  reg [_tmp_1244-1:0] __tmp_1245_24;
  reg [_tmp_1244-1:0] __tmp_1245_25;
  reg [_tmp_1244-1:0] __tmp_1245_26;
  reg [_tmp_1244-1:0] __tmp_1245_27;
  reg [_tmp_1244-1:0] __tmp_1245_28;
  localparam _tmp_1246 = 1;
  wire [_tmp_1246-1:0] _tmp_1247;
  assign _tmp_1247 = (_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag;
  reg [_tmp_1246-1:0] __tmp_1247_1;
  reg [_tmp_1246-1:0] __tmp_1247_2;
  reg [_tmp_1246-1:0] __tmp_1247_3;
  reg [_tmp_1246-1:0] __tmp_1247_4;
  reg [_tmp_1246-1:0] __tmp_1247_5;
  reg [_tmp_1246-1:0] __tmp_1247_6;
  reg [_tmp_1246-1:0] __tmp_1247_7;
  reg [_tmp_1246-1:0] __tmp_1247_8;
  reg [_tmp_1246-1:0] __tmp_1247_9;
  reg [_tmp_1246-1:0] __tmp_1247_10;
  reg [_tmp_1246-1:0] __tmp_1247_11;
  reg [_tmp_1246-1:0] __tmp_1247_12;
  reg [_tmp_1246-1:0] __tmp_1247_13;
  reg [_tmp_1246-1:0] __tmp_1247_14;
  reg [_tmp_1246-1:0] __tmp_1247_15;
  reg [_tmp_1246-1:0] __tmp_1247_16;
  reg [_tmp_1246-1:0] __tmp_1247_17;
  reg [_tmp_1246-1:0] __tmp_1247_18;
  reg [_tmp_1246-1:0] __tmp_1247_19;
  reg [_tmp_1246-1:0] __tmp_1247_20;
  reg [_tmp_1246-1:0] __tmp_1247_21;
  reg [_tmp_1246-1:0] __tmp_1247_22;
  reg [_tmp_1246-1:0] __tmp_1247_23;
  reg [_tmp_1246-1:0] __tmp_1247_24;
  reg [_tmp_1246-1:0] __tmp_1247_25;
  reg [_tmp_1246-1:0] __tmp_1247_26;
  reg [_tmp_1246-1:0] __tmp_1247_27;
  reg [_tmp_1246-1:0] __tmp_1247_28;
  localparam _tmp_1248 = 1;
  wire [_tmp_1248-1:0] _tmp_1249;
  assign _tmp_1249 = (_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag;
  reg [_tmp_1248-1:0] __tmp_1249_1;
  reg [_tmp_1248-1:0] __tmp_1249_2;
  reg [_tmp_1248-1:0] __tmp_1249_3;
  reg [_tmp_1248-1:0] __tmp_1249_4;
  reg [_tmp_1248-1:0] __tmp_1249_5;
  reg [_tmp_1248-1:0] __tmp_1249_6;
  reg [_tmp_1248-1:0] __tmp_1249_7;
  reg [_tmp_1248-1:0] __tmp_1249_8;
  reg [_tmp_1248-1:0] __tmp_1249_9;
  reg [_tmp_1248-1:0] __tmp_1249_10;
  reg [_tmp_1248-1:0] __tmp_1249_11;
  reg [_tmp_1248-1:0] __tmp_1249_12;
  reg [_tmp_1248-1:0] __tmp_1249_13;
  reg [_tmp_1248-1:0] __tmp_1249_14;
  reg [_tmp_1248-1:0] __tmp_1249_15;
  reg [_tmp_1248-1:0] __tmp_1249_16;
  reg [_tmp_1248-1:0] __tmp_1249_17;
  reg [_tmp_1248-1:0] __tmp_1249_18;
  reg [_tmp_1248-1:0] __tmp_1249_19;
  reg [_tmp_1248-1:0] __tmp_1249_20;
  reg [_tmp_1248-1:0] __tmp_1249_21;
  reg [_tmp_1248-1:0] __tmp_1249_22;
  reg [_tmp_1248-1:0] __tmp_1249_23;
  reg [_tmp_1248-1:0] __tmp_1249_24;
  reg [_tmp_1248-1:0] __tmp_1249_25;
  reg [_tmp_1248-1:0] __tmp_1249_26;
  reg [_tmp_1248-1:0] __tmp_1249_27;
  reg [_tmp_1248-1:0] __tmp_1249_28;
  wire _stream_matmul_29_done;
  assign _stream_matmul_29_done = _stream_matmul_29_source_10_idle && _stream_matmul_29_source_12_idle && _stream_matmul_29_source_14_idle && _stream_matmul_29_source_19_idle && _stream_matmul_29_source_20_idle && _stream_matmul_29_source_6_idle && _stream_matmul_29_source_8_idle;
  localparam _tmp_1250 = 1;
  wire [_tmp_1250-1:0] _tmp_1251;
  assign _tmp_1251 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1250-1:0] __tmp_1251_1;
  localparam _tmp_1252 = 1;
  wire [_tmp_1252-1:0] _tmp_1253;
  assign _tmp_1253 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1252-1:0] __tmp_1253_1;
  reg [_tmp_1252-1:0] __tmp_1253_2;
  reg [_tmp_1252-1:0] __tmp_1253_3;
  reg [_tmp_1252-1:0] __tmp_1253_4;
  reg [_tmp_1252-1:0] __tmp_1253_5;
  localparam _tmp_1254 = 1;
  wire [_tmp_1254-1:0] _tmp_1255;
  assign _tmp_1255 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1254-1:0] __tmp_1255_1;
  reg [_tmp_1254-1:0] __tmp_1255_2;
  reg [_tmp_1254-1:0] __tmp_1255_3;
  reg [_tmp_1254-1:0] __tmp_1255_4;
  reg [_tmp_1254-1:0] __tmp_1255_5;
  localparam _tmp_1256 = 1;
  wire [_tmp_1256-1:0] _tmp_1257;
  assign _tmp_1257 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1256-1:0] __tmp_1257_1;
  reg [_tmp_1256-1:0] __tmp_1257_2;
  reg [_tmp_1256-1:0] __tmp_1257_3;
  reg [_tmp_1256-1:0] __tmp_1257_4;
  reg [_tmp_1256-1:0] __tmp_1257_5;
  localparam _tmp_1258 = 1;
  wire [_tmp_1258-1:0] _tmp_1259;
  assign _tmp_1259 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1258-1:0] __tmp_1259_1;
  reg [_tmp_1258-1:0] __tmp_1259_2;
  reg [_tmp_1258-1:0] __tmp_1259_3;
  reg [_tmp_1258-1:0] __tmp_1259_4;
  reg [_tmp_1258-1:0] __tmp_1259_5;
  reg [_tmp_1258-1:0] __tmp_1259_6;
  reg [_tmp_1258-1:0] __tmp_1259_7;
  reg [_tmp_1258-1:0] __tmp_1259_8;
  reg [_tmp_1258-1:0] __tmp_1259_9;
  reg [_tmp_1258-1:0] __tmp_1259_10;
  reg [_tmp_1258-1:0] __tmp_1259_11;
  reg [_tmp_1258-1:0] __tmp_1259_12;
  localparam _tmp_1260 = 1;
  wire [_tmp_1260-1:0] _tmp_1261;
  assign _tmp_1261 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1260-1:0] __tmp_1261_1;
  reg [_tmp_1260-1:0] __tmp_1261_2;
  reg [_tmp_1260-1:0] __tmp_1261_3;
  reg [_tmp_1260-1:0] __tmp_1261_4;
  reg [_tmp_1260-1:0] __tmp_1261_5;
  reg [_tmp_1260-1:0] __tmp_1261_6;
  reg [_tmp_1260-1:0] __tmp_1261_7;
  reg [_tmp_1260-1:0] __tmp_1261_8;
  reg [_tmp_1260-1:0] __tmp_1261_9;
  reg [_tmp_1260-1:0] __tmp_1261_10;
  reg [_tmp_1260-1:0] __tmp_1261_11;
  reg [_tmp_1260-1:0] __tmp_1261_12;
  localparam _tmp_1262 = 1;
  wire [_tmp_1262-1:0] _tmp_1263;
  assign _tmp_1263 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1262-1:0] __tmp_1263_1;
  reg [_tmp_1262-1:0] __tmp_1263_2;
  reg [_tmp_1262-1:0] __tmp_1263_3;
  reg [_tmp_1262-1:0] __tmp_1263_4;
  reg [_tmp_1262-1:0] __tmp_1263_5;
  reg [_tmp_1262-1:0] __tmp_1263_6;
  reg [_tmp_1262-1:0] __tmp_1263_7;
  reg [_tmp_1262-1:0] __tmp_1263_8;
  reg [_tmp_1262-1:0] __tmp_1263_9;
  reg [_tmp_1262-1:0] __tmp_1263_10;
  reg [_tmp_1262-1:0] __tmp_1263_11;
  reg [_tmp_1262-1:0] __tmp_1263_12;
  localparam _tmp_1264 = 1;
  wire [_tmp_1264-1:0] _tmp_1265;
  assign _tmp_1265 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1264-1:0] __tmp_1265_1;
  reg [_tmp_1264-1:0] __tmp_1265_2;
  reg [_tmp_1264-1:0] __tmp_1265_3;
  reg [_tmp_1264-1:0] __tmp_1265_4;
  reg [_tmp_1264-1:0] __tmp_1265_5;
  reg [_tmp_1264-1:0] __tmp_1265_6;
  reg [_tmp_1264-1:0] __tmp_1265_7;
  reg [_tmp_1264-1:0] __tmp_1265_8;
  reg [_tmp_1264-1:0] __tmp_1265_9;
  reg [_tmp_1264-1:0] __tmp_1265_10;
  reg [_tmp_1264-1:0] __tmp_1265_11;
  reg [_tmp_1264-1:0] __tmp_1265_12;
  reg [_tmp_1264-1:0] __tmp_1265_13;
  reg [_tmp_1264-1:0] __tmp_1265_14;
  reg [_tmp_1264-1:0] __tmp_1265_15;
  reg [2-1:0] _add_tree_1_sink_wait_count;
  localparam _tmp_1266 = 1;
  wire [_tmp_1266-1:0] _tmp_1267;
  assign _tmp_1267 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1266-1:0] __tmp_1267_1;
  reg [_tmp_1266-1:0] __tmp_1267_2;
  reg [_tmp_1266-1:0] __tmp_1267_3;
  reg [_tmp_1266-1:0] __tmp_1267_4;
  localparam _tmp_1268 = 1;
  wire [_tmp_1268-1:0] _tmp_1269;
  assign _tmp_1269 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1268-1:0] __tmp_1269_1;
  reg [_tmp_1268-1:0] __tmp_1269_2;
  reg [_tmp_1268-1:0] __tmp_1269_3;
  reg [_tmp_1268-1:0] __tmp_1269_4;
  localparam _tmp_1270 = 1;
  wire [_tmp_1270-1:0] _tmp_1271;
  assign _tmp_1271 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1270-1:0] __tmp_1271_1;
  reg [_tmp_1270-1:0] __tmp_1271_2;
  reg [_tmp_1270-1:0] __tmp_1271_3;
  reg [_tmp_1270-1:0] __tmp_1271_4;
  localparam _tmp_1272 = 1;
  wire [_tmp_1272-1:0] _tmp_1273;
  assign _tmp_1273 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1272-1:0] __tmp_1273_1;
  reg [_tmp_1272-1:0] __tmp_1273_2;
  reg [_tmp_1272-1:0] __tmp_1273_3;
  reg [_tmp_1272-1:0] __tmp_1273_4;
  reg [_tmp_1272-1:0] __tmp_1273_5;
  reg [_tmp_1272-1:0] __tmp_1273_6;
  reg [_tmp_1272-1:0] __tmp_1273_7;
  reg [_tmp_1272-1:0] __tmp_1273_8;
  reg [_tmp_1272-1:0] __tmp_1273_9;
  reg [_tmp_1272-1:0] __tmp_1273_10;
  reg [_tmp_1272-1:0] __tmp_1273_11;
  reg [_tmp_1272-1:0] __tmp_1273_12;
  reg [_tmp_1272-1:0] __tmp_1273_13;
  reg [_tmp_1272-1:0] __tmp_1273_14;
  reg [_tmp_1272-1:0] __tmp_1273_15;
  reg [_tmp_1272-1:0] __tmp_1273_16;
  reg [_tmp_1272-1:0] __tmp_1273_17;
  reg [_tmp_1272-1:0] __tmp_1273_18;
  localparam _tmp_1274 = 1;
  wire [_tmp_1274-1:0] _tmp_1275;
  assign _tmp_1275 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1274-1:0] __tmp_1275_1;
  reg [_tmp_1274-1:0] __tmp_1275_2;
  reg [_tmp_1274-1:0] __tmp_1275_3;
  reg [_tmp_1274-1:0] __tmp_1275_4;
  reg [_tmp_1274-1:0] __tmp_1275_5;
  reg [_tmp_1274-1:0] __tmp_1275_6;
  reg [_tmp_1274-1:0] __tmp_1275_7;
  reg [_tmp_1274-1:0] __tmp_1275_8;
  reg [_tmp_1274-1:0] __tmp_1275_9;
  reg [_tmp_1274-1:0] __tmp_1275_10;
  reg [_tmp_1274-1:0] __tmp_1275_11;
  reg [_tmp_1274-1:0] __tmp_1275_12;
  reg [_tmp_1274-1:0] __tmp_1275_13;
  reg [_tmp_1274-1:0] __tmp_1275_14;
  reg [_tmp_1274-1:0] __tmp_1275_15;
  reg [_tmp_1274-1:0] __tmp_1275_16;
  reg [_tmp_1274-1:0] __tmp_1275_17;
  localparam _tmp_1276 = 1;
  wire [_tmp_1276-1:0] _tmp_1277;
  assign _tmp_1277 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1276-1:0] __tmp_1277_1;
  reg [_tmp_1276-1:0] __tmp_1277_2;
  reg [_tmp_1276-1:0] __tmp_1277_3;
  reg [_tmp_1276-1:0] __tmp_1277_4;
  reg [_tmp_1276-1:0] __tmp_1277_5;
  reg [_tmp_1276-1:0] __tmp_1277_6;
  reg [_tmp_1276-1:0] __tmp_1277_7;
  reg [_tmp_1276-1:0] __tmp_1277_8;
  reg [_tmp_1276-1:0] __tmp_1277_9;
  reg [_tmp_1276-1:0] __tmp_1277_10;
  reg [_tmp_1276-1:0] __tmp_1277_11;
  reg [_tmp_1276-1:0] __tmp_1277_12;
  reg [_tmp_1276-1:0] __tmp_1277_13;
  reg [_tmp_1276-1:0] __tmp_1277_14;
  reg [_tmp_1276-1:0] __tmp_1277_15;
  reg [_tmp_1276-1:0] __tmp_1277_16;
  reg [_tmp_1276-1:0] __tmp_1277_17;
  localparam _tmp_1278 = 1;
  wire [_tmp_1278-1:0] _tmp_1279;
  assign _tmp_1279 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1278-1:0] __tmp_1279_1;
  reg [_tmp_1278-1:0] __tmp_1279_2;
  reg [_tmp_1278-1:0] __tmp_1279_3;
  reg [_tmp_1278-1:0] __tmp_1279_4;
  reg [_tmp_1278-1:0] __tmp_1279_5;
  reg [_tmp_1278-1:0] __tmp_1279_6;
  reg [_tmp_1278-1:0] __tmp_1279_7;
  reg [_tmp_1278-1:0] __tmp_1279_8;
  reg [_tmp_1278-1:0] __tmp_1279_9;
  reg [_tmp_1278-1:0] __tmp_1279_10;
  reg [_tmp_1278-1:0] __tmp_1279_11;
  reg [_tmp_1278-1:0] __tmp_1279_12;
  reg [_tmp_1278-1:0] __tmp_1279_13;
  reg [_tmp_1278-1:0] __tmp_1279_14;
  reg [_tmp_1278-1:0] __tmp_1279_15;
  reg [_tmp_1278-1:0] __tmp_1279_16;
  reg [_tmp_1278-1:0] __tmp_1279_17;
  localparam _tmp_1280 = 1;
  wire [_tmp_1280-1:0] _tmp_1281;
  assign _tmp_1281 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1280-1:0] __tmp_1281_1;
  reg [_tmp_1280-1:0] __tmp_1281_2;
  reg [_tmp_1280-1:0] __tmp_1281_3;
  reg [_tmp_1280-1:0] __tmp_1281_4;
  reg [_tmp_1280-1:0] __tmp_1281_5;
  reg [_tmp_1280-1:0] __tmp_1281_6;
  reg [_tmp_1280-1:0] __tmp_1281_7;
  reg [_tmp_1280-1:0] __tmp_1281_8;
  reg [_tmp_1280-1:0] __tmp_1281_9;
  localparam _tmp_1282 = 1;
  wire [_tmp_1282-1:0] _tmp_1283;
  assign _tmp_1283 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1282-1:0] __tmp_1283_1;
  reg [_tmp_1282-1:0] __tmp_1283_2;
  reg [_tmp_1282-1:0] __tmp_1283_3;
  reg [_tmp_1282-1:0] __tmp_1283_4;
  reg [_tmp_1282-1:0] __tmp_1283_5;
  reg [_tmp_1282-1:0] __tmp_1283_6;
  reg [_tmp_1282-1:0] __tmp_1283_7;
  reg [_tmp_1282-1:0] __tmp_1283_8;
  reg [_tmp_1282-1:0] __tmp_1283_9;
  localparam _tmp_1284 = 1;
  wire [_tmp_1284-1:0] _tmp_1285;
  assign _tmp_1285 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1284-1:0] __tmp_1285_1;
  reg [_tmp_1284-1:0] __tmp_1285_2;
  reg [_tmp_1284-1:0] __tmp_1285_3;
  reg [_tmp_1284-1:0] __tmp_1285_4;
  reg [_tmp_1284-1:0] __tmp_1285_5;
  reg [_tmp_1284-1:0] __tmp_1285_6;
  reg [_tmp_1284-1:0] __tmp_1285_7;
  reg [_tmp_1284-1:0] __tmp_1285_8;
  reg [_tmp_1284-1:0] __tmp_1285_9;
  localparam _tmp_1286 = 1;
  wire [_tmp_1286-1:0] _tmp_1287;
  assign _tmp_1287 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1286-1:0] __tmp_1287_1;
  reg [_tmp_1286-1:0] __tmp_1287_2;
  reg [_tmp_1286-1:0] __tmp_1287_3;
  reg [_tmp_1286-1:0] __tmp_1287_4;
  reg [_tmp_1286-1:0] __tmp_1287_5;
  reg [_tmp_1286-1:0] __tmp_1287_6;
  reg [_tmp_1286-1:0] __tmp_1287_7;
  reg [_tmp_1286-1:0] __tmp_1287_8;
  reg [_tmp_1286-1:0] __tmp_1287_9;
  reg [_tmp_1286-1:0] __tmp_1287_10;
  reg [_tmp_1286-1:0] __tmp_1287_11;
  reg [_tmp_1286-1:0] __tmp_1287_12;
  reg [_tmp_1286-1:0] __tmp_1287_13;
  reg [_tmp_1286-1:0] __tmp_1287_14;
  reg [_tmp_1286-1:0] __tmp_1287_15;
  reg [_tmp_1286-1:0] __tmp_1287_16;
  reg [_tmp_1286-1:0] __tmp_1287_17;
  reg [_tmp_1286-1:0] __tmp_1287_18;
  reg [_tmp_1286-1:0] __tmp_1287_19;
  reg [_tmp_1286-1:0] __tmp_1287_20;
  reg [_tmp_1286-1:0] __tmp_1287_21;
  reg [_tmp_1286-1:0] __tmp_1287_22;
  reg [_tmp_1286-1:0] __tmp_1287_23;
  reg [_tmp_1286-1:0] __tmp_1287_24;
  reg [_tmp_1286-1:0] __tmp_1287_25;
  localparam _tmp_1288 = 1;
  wire [_tmp_1288-1:0] _tmp_1289;
  assign _tmp_1289 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1288-1:0] __tmp_1289_1;
  reg [_tmp_1288-1:0] __tmp_1289_2;
  reg [_tmp_1288-1:0] __tmp_1289_3;
  reg [_tmp_1288-1:0] __tmp_1289_4;
  reg [_tmp_1288-1:0] __tmp_1289_5;
  reg [_tmp_1288-1:0] __tmp_1289_6;
  reg [_tmp_1288-1:0] __tmp_1289_7;
  reg [_tmp_1288-1:0] __tmp_1289_8;
  reg [_tmp_1288-1:0] __tmp_1289_9;
  reg [_tmp_1288-1:0] __tmp_1289_10;
  reg [_tmp_1288-1:0] __tmp_1289_11;
  reg [_tmp_1288-1:0] __tmp_1289_12;
  reg [_tmp_1288-1:0] __tmp_1289_13;
  reg [_tmp_1288-1:0] __tmp_1289_14;
  reg [_tmp_1288-1:0] __tmp_1289_15;
  reg [_tmp_1288-1:0] __tmp_1289_16;
  reg [_tmp_1288-1:0] __tmp_1289_17;
  reg [_tmp_1288-1:0] __tmp_1289_18;
  reg [_tmp_1288-1:0] __tmp_1289_19;
  reg [_tmp_1288-1:0] __tmp_1289_20;
  reg [_tmp_1288-1:0] __tmp_1289_21;
  reg [_tmp_1288-1:0] __tmp_1289_22;
  reg [_tmp_1288-1:0] __tmp_1289_23;
  reg [_tmp_1288-1:0] __tmp_1289_24;
  reg [_tmp_1288-1:0] __tmp_1289_25;
  localparam _tmp_1290 = 1;
  wire [_tmp_1290-1:0] _tmp_1291;
  assign _tmp_1291 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1290-1:0] __tmp_1291_1;
  reg [_tmp_1290-1:0] __tmp_1291_2;
  reg [_tmp_1290-1:0] __tmp_1291_3;
  reg [_tmp_1290-1:0] __tmp_1291_4;
  reg [_tmp_1290-1:0] __tmp_1291_5;
  reg [_tmp_1290-1:0] __tmp_1291_6;
  reg [_tmp_1290-1:0] __tmp_1291_7;
  reg [_tmp_1290-1:0] __tmp_1291_8;
  reg [_tmp_1290-1:0] __tmp_1291_9;
  reg [_tmp_1290-1:0] __tmp_1291_10;
  reg [_tmp_1290-1:0] __tmp_1291_11;
  reg [_tmp_1290-1:0] __tmp_1291_12;
  reg [_tmp_1290-1:0] __tmp_1291_13;
  reg [_tmp_1290-1:0] __tmp_1291_14;
  reg [_tmp_1290-1:0] __tmp_1291_15;
  reg [_tmp_1290-1:0] __tmp_1291_16;
  reg [_tmp_1290-1:0] __tmp_1291_17;
  reg [_tmp_1290-1:0] __tmp_1291_18;
  reg [_tmp_1290-1:0] __tmp_1291_19;
  reg [_tmp_1290-1:0] __tmp_1291_20;
  reg [_tmp_1290-1:0] __tmp_1291_21;
  reg [_tmp_1290-1:0] __tmp_1291_22;
  reg [_tmp_1290-1:0] __tmp_1291_23;
  reg [_tmp_1290-1:0] __tmp_1291_24;
  reg [_tmp_1290-1:0] __tmp_1291_25;
  localparam _tmp_1292 = 1;
  wire [_tmp_1292-1:0] _tmp_1293;
  assign _tmp_1293 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1292-1:0] __tmp_1293_1;
  reg [_tmp_1292-1:0] __tmp_1293_2;
  reg [_tmp_1292-1:0] __tmp_1293_3;
  reg [_tmp_1292-1:0] __tmp_1293_4;
  reg [_tmp_1292-1:0] __tmp_1293_5;
  reg [_tmp_1292-1:0] __tmp_1293_6;
  reg [_tmp_1292-1:0] __tmp_1293_7;
  reg [_tmp_1292-1:0] __tmp_1293_8;
  reg [_tmp_1292-1:0] __tmp_1293_9;
  reg [_tmp_1292-1:0] __tmp_1293_10;
  reg [_tmp_1292-1:0] __tmp_1293_11;
  reg [_tmp_1292-1:0] __tmp_1293_12;
  localparam _tmp_1294 = 1;
  wire [_tmp_1294-1:0] _tmp_1295;
  assign _tmp_1295 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1294-1:0] __tmp_1295_1;
  reg [_tmp_1294-1:0] __tmp_1295_2;
  reg [_tmp_1294-1:0] __tmp_1295_3;
  reg [_tmp_1294-1:0] __tmp_1295_4;
  reg [_tmp_1294-1:0] __tmp_1295_5;
  reg [_tmp_1294-1:0] __tmp_1295_6;
  reg [_tmp_1294-1:0] __tmp_1295_7;
  reg [_tmp_1294-1:0] __tmp_1295_8;
  reg [_tmp_1294-1:0] __tmp_1295_9;
  reg [_tmp_1294-1:0] __tmp_1295_10;
  reg [_tmp_1294-1:0] __tmp_1295_11;
  reg [_tmp_1294-1:0] __tmp_1295_12;
  localparam _tmp_1296 = 1;
  wire [_tmp_1296-1:0] _tmp_1297;
  assign _tmp_1297 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1296-1:0] __tmp_1297_1;
  reg [_tmp_1296-1:0] __tmp_1297_2;
  reg [_tmp_1296-1:0] __tmp_1297_3;
  reg [_tmp_1296-1:0] __tmp_1297_4;
  reg [_tmp_1296-1:0] __tmp_1297_5;
  reg [_tmp_1296-1:0] __tmp_1297_6;
  reg [_tmp_1296-1:0] __tmp_1297_7;
  reg [_tmp_1296-1:0] __tmp_1297_8;
  reg [_tmp_1296-1:0] __tmp_1297_9;
  reg [_tmp_1296-1:0] __tmp_1297_10;
  reg [_tmp_1296-1:0] __tmp_1297_11;
  reg [_tmp_1296-1:0] __tmp_1297_12;
  reg [6-1:0] _stream_matmul_29_sink_wait_count;
  localparam _tmp_1298 = 1;
  wire [_tmp_1298-1:0] _tmp_1299;
  assign _tmp_1299 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1298-1:0] __tmp_1299_1;
  reg [_tmp_1298-1:0] __tmp_1299_2;
  reg [_tmp_1298-1:0] __tmp_1299_3;
  reg [_tmp_1298-1:0] __tmp_1299_4;
  reg [_tmp_1298-1:0] __tmp_1299_5;
  reg [_tmp_1298-1:0] __tmp_1299_6;
  reg [_tmp_1298-1:0] __tmp_1299_7;
  reg [_tmp_1298-1:0] __tmp_1299_8;
  reg [_tmp_1298-1:0] __tmp_1299_9;
  reg [_tmp_1298-1:0] __tmp_1299_10;
  reg [_tmp_1298-1:0] __tmp_1299_11;
  reg [_tmp_1298-1:0] __tmp_1299_12;
  reg [_tmp_1298-1:0] __tmp_1299_13;
  reg [_tmp_1298-1:0] __tmp_1299_14;
  reg [_tmp_1298-1:0] __tmp_1299_15;
  reg [_tmp_1298-1:0] __tmp_1299_16;
  reg [_tmp_1298-1:0] __tmp_1299_17;
  reg [_tmp_1298-1:0] __tmp_1299_18;
  reg [_tmp_1298-1:0] __tmp_1299_19;
  reg [_tmp_1298-1:0] __tmp_1299_20;
  reg [_tmp_1298-1:0] __tmp_1299_21;
  reg [_tmp_1298-1:0] __tmp_1299_22;
  reg [_tmp_1298-1:0] __tmp_1299_23;
  reg [_tmp_1298-1:0] __tmp_1299_24;
  reg [_tmp_1298-1:0] __tmp_1299_25;
  reg [_tmp_1298-1:0] __tmp_1299_26;
  reg [_tmp_1298-1:0] __tmp_1299_27;
  reg [_tmp_1298-1:0] __tmp_1299_28;
  reg [_tmp_1298-1:0] __tmp_1299_29;
  reg [_tmp_1298-1:0] __tmp_1299_30;
  reg [_tmp_1298-1:0] __tmp_1299_31;
  reg [_tmp_1298-1:0] __tmp_1299_32;
  reg [_tmp_1298-1:0] __tmp_1299_33;
  reg [_tmp_1298-1:0] __tmp_1299_34;
  reg [_tmp_1298-1:0] __tmp_1299_35;
  reg [_tmp_1298-1:0] __tmp_1299_36;
  reg [_tmp_1298-1:0] __tmp_1299_37;
  reg [_tmp_1298-1:0] __tmp_1299_38;
  reg [_tmp_1298-1:0] __tmp_1299_39;
  reg [_tmp_1298-1:0] __tmp_1299_40;
  reg [_tmp_1298-1:0] __tmp_1299_41;
  reg [_tmp_1298-1:0] __tmp_1299_42;
  localparam _tmp_1300 = 1;
  wire [_tmp_1300-1:0] _tmp_1301;
  assign _tmp_1301 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1300-1:0] __tmp_1301_1;
  reg [_tmp_1300-1:0] __tmp_1301_2;
  reg [_tmp_1300-1:0] __tmp_1301_3;
  reg [_tmp_1300-1:0] __tmp_1301_4;
  reg [_tmp_1300-1:0] __tmp_1301_5;
  reg [_tmp_1300-1:0] __tmp_1301_6;
  reg [_tmp_1300-1:0] __tmp_1301_7;
  reg [_tmp_1300-1:0] __tmp_1301_8;
  reg [_tmp_1300-1:0] __tmp_1301_9;
  reg [_tmp_1300-1:0] __tmp_1301_10;
  reg [_tmp_1300-1:0] __tmp_1301_11;
  reg [_tmp_1300-1:0] __tmp_1301_12;
  reg [_tmp_1300-1:0] __tmp_1301_13;
  reg [_tmp_1300-1:0] __tmp_1301_14;
  reg [_tmp_1300-1:0] __tmp_1301_15;
  reg [_tmp_1300-1:0] __tmp_1301_16;
  reg [_tmp_1300-1:0] __tmp_1301_17;
  reg [_tmp_1300-1:0] __tmp_1301_18;
  reg [_tmp_1300-1:0] __tmp_1301_19;
  reg [_tmp_1300-1:0] __tmp_1301_20;
  reg [_tmp_1300-1:0] __tmp_1301_21;
  reg [_tmp_1300-1:0] __tmp_1301_22;
  reg [_tmp_1300-1:0] __tmp_1301_23;
  reg [_tmp_1300-1:0] __tmp_1301_24;
  reg [_tmp_1300-1:0] __tmp_1301_25;
  reg [_tmp_1300-1:0] __tmp_1301_26;
  reg [_tmp_1300-1:0] __tmp_1301_27;
  reg [_tmp_1300-1:0] __tmp_1301_28;
  reg [_tmp_1300-1:0] __tmp_1301_29;
  reg [_tmp_1300-1:0] __tmp_1301_30;
  reg [_tmp_1300-1:0] __tmp_1301_31;
  reg [_tmp_1300-1:0] __tmp_1301_32;
  reg [_tmp_1300-1:0] __tmp_1301_33;
  reg [_tmp_1300-1:0] __tmp_1301_34;
  reg [_tmp_1300-1:0] __tmp_1301_35;
  reg [_tmp_1300-1:0] __tmp_1301_36;
  reg [_tmp_1300-1:0] __tmp_1301_37;
  reg [_tmp_1300-1:0] __tmp_1301_38;
  reg [_tmp_1300-1:0] __tmp_1301_39;
  reg [_tmp_1300-1:0] __tmp_1301_40;
  reg [_tmp_1300-1:0] __tmp_1301_41;
  reg [_tmp_1300-1:0] __tmp_1301_42;
  localparam _tmp_1302 = 1;
  wire [_tmp_1302-1:0] _tmp_1303;
  assign _tmp_1303 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1302-1:0] __tmp_1303_1;
  reg [_tmp_1302-1:0] __tmp_1303_2;
  reg [_tmp_1302-1:0] __tmp_1303_3;
  reg [_tmp_1302-1:0] __tmp_1303_4;
  reg [_tmp_1302-1:0] __tmp_1303_5;
  reg [_tmp_1302-1:0] __tmp_1303_6;
  reg [_tmp_1302-1:0] __tmp_1303_7;
  reg [_tmp_1302-1:0] __tmp_1303_8;
  reg [_tmp_1302-1:0] __tmp_1303_9;
  reg [_tmp_1302-1:0] __tmp_1303_10;
  reg [_tmp_1302-1:0] __tmp_1303_11;
  reg [_tmp_1302-1:0] __tmp_1303_12;
  reg [_tmp_1302-1:0] __tmp_1303_13;
  reg [_tmp_1302-1:0] __tmp_1303_14;
  reg [_tmp_1302-1:0] __tmp_1303_15;
  reg [_tmp_1302-1:0] __tmp_1303_16;
  reg [_tmp_1302-1:0] __tmp_1303_17;
  reg [_tmp_1302-1:0] __tmp_1303_18;
  reg [_tmp_1302-1:0] __tmp_1303_19;
  reg [_tmp_1302-1:0] __tmp_1303_20;
  reg [_tmp_1302-1:0] __tmp_1303_21;
  reg [_tmp_1302-1:0] __tmp_1303_22;
  reg [_tmp_1302-1:0] __tmp_1303_23;
  reg [_tmp_1302-1:0] __tmp_1303_24;
  reg [_tmp_1302-1:0] __tmp_1303_25;
  reg [_tmp_1302-1:0] __tmp_1303_26;
  reg [_tmp_1302-1:0] __tmp_1303_27;
  reg [_tmp_1302-1:0] __tmp_1303_28;
  reg [_tmp_1302-1:0] __tmp_1303_29;
  reg [_tmp_1302-1:0] __tmp_1303_30;
  reg [_tmp_1302-1:0] __tmp_1303_31;
  reg [_tmp_1302-1:0] __tmp_1303_32;
  reg [_tmp_1302-1:0] __tmp_1303_33;
  reg [_tmp_1302-1:0] __tmp_1303_34;
  reg [_tmp_1302-1:0] __tmp_1303_35;
  reg [_tmp_1302-1:0] __tmp_1303_36;
  reg [_tmp_1302-1:0] __tmp_1303_37;
  reg [_tmp_1302-1:0] __tmp_1303_38;
  reg [_tmp_1302-1:0] __tmp_1303_39;
  reg [_tmp_1302-1:0] __tmp_1303_40;
  reg [_tmp_1302-1:0] __tmp_1303_41;
  reg [_tmp_1302-1:0] __tmp_1303_42;
  localparam _tmp_1304 = 1;
  wire [_tmp_1304-1:0] _tmp_1305;
  assign _tmp_1305 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1304-1:0] __tmp_1305_1;
  reg [_tmp_1304-1:0] __tmp_1305_2;
  reg [_tmp_1304-1:0] __tmp_1305_3;
  reg [_tmp_1304-1:0] __tmp_1305_4;
  reg [_tmp_1304-1:0] __tmp_1305_5;
  reg [_tmp_1304-1:0] __tmp_1305_6;
  reg [_tmp_1304-1:0] __tmp_1305_7;
  reg [_tmp_1304-1:0] __tmp_1305_8;
  reg [_tmp_1304-1:0] __tmp_1305_9;
  reg [_tmp_1304-1:0] __tmp_1305_10;
  reg [_tmp_1304-1:0] __tmp_1305_11;
  reg [_tmp_1304-1:0] __tmp_1305_12;
  reg [_tmp_1304-1:0] __tmp_1305_13;
  reg [_tmp_1304-1:0] __tmp_1305_14;
  reg [_tmp_1304-1:0] __tmp_1305_15;
  reg [_tmp_1304-1:0] __tmp_1305_16;
  reg [_tmp_1304-1:0] __tmp_1305_17;
  reg [_tmp_1304-1:0] __tmp_1305_18;
  reg [_tmp_1304-1:0] __tmp_1305_19;
  reg [_tmp_1304-1:0] __tmp_1305_20;
  reg [_tmp_1304-1:0] __tmp_1305_21;
  reg [_tmp_1304-1:0] __tmp_1305_22;
  reg [_tmp_1304-1:0] __tmp_1305_23;
  reg [_tmp_1304-1:0] __tmp_1305_24;
  reg [_tmp_1304-1:0] __tmp_1305_25;
  reg [_tmp_1304-1:0] __tmp_1305_26;
  reg [_tmp_1304-1:0] __tmp_1305_27;
  reg [_tmp_1304-1:0] __tmp_1305_28;
  reg [_tmp_1304-1:0] __tmp_1305_29;
  reg [_tmp_1304-1:0] __tmp_1305_30;
  reg [_tmp_1304-1:0] __tmp_1305_31;
  reg [_tmp_1304-1:0] __tmp_1305_32;
  reg [_tmp_1304-1:0] __tmp_1305_33;
  reg [_tmp_1304-1:0] __tmp_1305_34;
  reg [_tmp_1304-1:0] __tmp_1305_35;
  reg [_tmp_1304-1:0] __tmp_1305_36;
  reg [_tmp_1304-1:0] __tmp_1305_37;
  reg [_tmp_1304-1:0] __tmp_1305_38;
  reg [_tmp_1304-1:0] __tmp_1305_39;
  reg [_tmp_1304-1:0] __tmp_1305_40;
  reg [_tmp_1304-1:0] __tmp_1305_41;
  reg [_tmp_1304-1:0] __tmp_1305_42;
  localparam _tmp_1306 = 1;
  wire [_tmp_1306-1:0] _tmp_1307;
  assign _tmp_1307 = _stream_matmul_29_fsm == 3;
  reg [_tmp_1306-1:0] __tmp_1307_1;
  reg [_tmp_1306-1:0] __tmp_1307_2;
  reg [_tmp_1306-1:0] __tmp_1307_3;
  reg [_tmp_1306-1:0] __tmp_1307_4;
  reg [_tmp_1306-1:0] __tmp_1307_5;
  reg [_tmp_1306-1:0] __tmp_1307_6;
  reg [_tmp_1306-1:0] __tmp_1307_7;
  reg [_tmp_1306-1:0] __tmp_1307_8;
  reg [_tmp_1306-1:0] __tmp_1307_9;
  reg [_tmp_1306-1:0] __tmp_1307_10;
  reg [_tmp_1306-1:0] __tmp_1307_11;
  reg [_tmp_1306-1:0] __tmp_1307_12;
  reg [_tmp_1306-1:0] __tmp_1307_13;
  reg [_tmp_1306-1:0] __tmp_1307_14;
  reg [_tmp_1306-1:0] __tmp_1307_15;
  reg [_tmp_1306-1:0] __tmp_1307_16;
  reg [_tmp_1306-1:0] __tmp_1307_17;
  reg [_tmp_1306-1:0] __tmp_1307_18;
  reg [_tmp_1306-1:0] __tmp_1307_19;
  reg [_tmp_1306-1:0] __tmp_1307_20;
  reg [_tmp_1306-1:0] __tmp_1307_21;
  reg [_tmp_1306-1:0] __tmp_1307_22;
  reg [_tmp_1306-1:0] __tmp_1307_23;
  reg [_tmp_1306-1:0] __tmp_1307_24;
  reg [_tmp_1306-1:0] __tmp_1307_25;
  reg [_tmp_1306-1:0] __tmp_1307_26;
  reg [_tmp_1306-1:0] __tmp_1307_27;
  reg [_tmp_1306-1:0] __tmp_1307_28;
  reg [_tmp_1306-1:0] __tmp_1307_29;
  reg [_tmp_1306-1:0] __tmp_1307_30;
  reg [_tmp_1306-1:0] __tmp_1307_31;
  reg [_tmp_1306-1:0] __tmp_1307_32;
  reg [_tmp_1306-1:0] __tmp_1307_33;
  reg [_tmp_1306-1:0] __tmp_1307_34;
  reg [_tmp_1306-1:0] __tmp_1307_35;
  reg [_tmp_1306-1:0] __tmp_1307_36;
  reg [_tmp_1306-1:0] __tmp_1307_37;
  reg [_tmp_1306-1:0] __tmp_1307_38;
  wire matmul_29_dma_out_mask_0;
  assign matmul_29_dma_out_mask_0 = matmul_29_out_row_count + 0 >= cparam_matmul_29_out_num_row;
  reg axim_flag_1308;
  reg _control_matmul_29_cond_32_4_1;
  reg _maxi_ram_w8_l2048_id1_1_write_start;
  reg [8-1:0] _maxi_ram_w8_l2048_id1_1_write_op_sel;
  reg [32-1:0] _maxi_ram_w8_l2048_id1_1_write_local_addr;
  reg [32-1:0] _maxi_ram_w8_l2048_id1_1_write_global_addr;
  reg [33-1:0] _maxi_ram_w8_l2048_id1_1_write_size;
  reg [32-1:0] _maxi_ram_w8_l2048_id1_1_write_local_stride;
  reg _tmp_1309;
  reg _tmp_1310;
  wire _tmp_1311;
  wire _tmp_1312;
  assign _tmp_1312 = 1;
  localparam _tmp_1313 = 1;
  wire [_tmp_1313-1:0] _tmp_1314;
  assign _tmp_1314 = (_tmp_1311 || !_tmp_1309) && (_tmp_1312 || !_tmp_1310);
  reg [_tmp_1313-1:0] __tmp_1314_1;
  wire signed [8-1:0] _tmp_1315;
  reg signed [8-1:0] __tmp_1315_1;
  assign _tmp_1315 = (__tmp_1314_1)? ram_w8_l2048_id1_0_1_rdata : __tmp_1315_1;
  reg _tmp_1316;
  reg _tmp_1317;
  reg _tmp_1318;
  reg _tmp_1319;
  reg [34-1:0] _tmp_1320;
  reg _tmp_1321;
  reg _tmp_1322;
  wire _tmp_1323;
  wire _tmp_1324;
  assign _tmp_1324 = 1;
  localparam _tmp_1325 = 1;
  wire [_tmp_1325-1:0] _tmp_1326;
  assign _tmp_1326 = (_tmp_1323 || !_tmp_1321) && (_tmp_1324 || !_tmp_1322);
  reg [_tmp_1325-1:0] __tmp_1326_1;
  wire signed [8-1:0] _tmp_1327;
  reg signed [8-1:0] __tmp_1327_1;
  assign _tmp_1327 = (__tmp_1326_1)? ram_w8_l2048_id1_1_1_rdata : __tmp_1327_1;
  reg _tmp_1328;
  reg _tmp_1329;
  reg _tmp_1330;
  reg _tmp_1331;
  reg [34-1:0] _tmp_1332;
  reg _tmp_1333;
  reg _tmp_1334;
  wire _tmp_1335;
  wire _tmp_1336;
  assign _tmp_1336 = 1;
  localparam _tmp_1337 = 1;
  wire [_tmp_1337-1:0] _tmp_1338;
  assign _tmp_1338 = (_tmp_1335 || !_tmp_1333) && (_tmp_1336 || !_tmp_1334);
  reg [_tmp_1337-1:0] __tmp_1338_1;
  wire signed [8-1:0] _tmp_1339;
  reg signed [8-1:0] __tmp_1339_1;
  assign _tmp_1339 = (__tmp_1338_1)? ram_w8_l2048_id1_2_1_rdata : __tmp_1339_1;
  reg _tmp_1340;
  reg _tmp_1341;
  reg _tmp_1342;
  reg _tmp_1343;
  reg [34-1:0] _tmp_1344;
  reg _tmp_1345;
  reg _tmp_1346;
  wire _tmp_1347;
  wire _tmp_1348;
  assign _tmp_1348 = 1;
  localparam _tmp_1349 = 1;
  wire [_tmp_1349-1:0] _tmp_1350;
  assign _tmp_1350 = (_tmp_1347 || !_tmp_1345) && (_tmp_1348 || !_tmp_1346);
  reg [_tmp_1349-1:0] __tmp_1350_1;
  wire signed [8-1:0] _tmp_1351;
  reg signed [8-1:0] __tmp_1351_1;
  assign _tmp_1351 = (__tmp_1350_1)? ram_w8_l2048_id1_3_1_rdata : __tmp_1351_1;
  reg _tmp_1352;
  reg _tmp_1353;
  reg _tmp_1354;
  reg _tmp_1355;
  reg [34-1:0] _tmp_1356;
  reg _tmp_1357;
  wire [32-1:0] _dataflow_cat_odata_167;
  wire _dataflow_cat_ovalid_167;
  wire _dataflow_cat_oready_167;
  assign _dataflow_cat_oready_167 = (_maxi_write_fsm == 3) && (_maxi_write_op_sel == 3) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid));
  reg _maxi_cond_4_1;
  assign _maxi_write_data_done = (_tmp_1357 && maxi_wvalid && maxi_wready)? 1 : 
                                 (_tmp_1120 && maxi_wvalid && maxi_wready)? 1 : 
                                 (_tmp_1020 && maxi_wvalid && maxi_wready)? 1 : 0;
  wire matmul_29_update_filter;
  assign matmul_29_update_filter = (cparam_matmul_29_data_stationary == 0) && (matmul_29_row_count >= cparam_matmul_29_max_row_count) && (matmul_29_bat_count >= cparam_matmul_29_max_bat_count) || (cparam_matmul_29_data_stationary == 1) && !cparam_matmul_29_keep_filter;
  wire matmul_29_update_act;
  assign matmul_29_update_act = (cparam_matmul_29_data_stationary == 1) && (matmul_29_och_count >= cparam_matmul_29_max_och_count) || (cparam_matmul_29_data_stationary == 0);
  wire matmul_29_mux_next_dma_flag_0;
  assign matmul_29_mux_next_dma_flag_0 = (matmul_29_row_select == 0)? (matmul_29_row_count >= cparam_matmul_29_max_row_count)? 1 : cparam_matmul_29_dma_flag_conds_0 : 1'd0;

  always @(posedge CLK) begin
    _RESETN_inv_1 <= RESETN_inv;
    _RESETN_inv_2 <= _RESETN_inv_1;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= 0;
      _maxi_ram_w8_l2048_id1_1_read_start <= 0;
      _maxi_ram_w8_l2048_id1_1_read_op_sel <= 0;
      _maxi_ram_w8_l2048_id1_1_read_local_addr <= 0;
      _maxi_ram_w8_l2048_id1_1_read_global_addr <= 0;
      _maxi_ram_w8_l2048_id1_1_read_size <= 0;
      _maxi_ram_w8_l2048_id1_1_read_local_stride <= 0;
      _maxi_read_idle <= 1;
      _maxi_read_op_sel <= 0;
      _maxi_read_local_addr <= 0;
      _maxi_read_global_addr <= 0;
      _maxi_read_size <= 0;
      _maxi_read_local_stride <= 0;
      maxi_araddr <= 0;
      maxi_arlen <= 0;
      maxi_arvalid <= 0;
      _tmp_20 <= 0;
      _maxi_cond_0_1 <= 0;
      _maxi_ram_w8_l2048_id0_1_read_start <= 0;
      _maxi_ram_w8_l2048_id0_1_read_op_sel <= 0;
      _maxi_ram_w8_l2048_id0_1_read_local_addr <= 0;
      _maxi_ram_w8_l2048_id0_1_read_global_addr <= 0;
      _maxi_ram_w8_l2048_id0_1_read_size <= 0;
      _maxi_ram_w8_l2048_id0_1_read_local_stride <= 0;
      _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start <= 0;
      _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_op_sel <= 0;
      _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_addr <= 0;
      _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_global_addr <= 0;
      _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_size <= 0;
      _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_stride <= 0;
      _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start <= 0;
      _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_op_sel <= 0;
      _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_addr <= 0;
      _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_global_addr <= 0;
      _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_size <= 0;
      _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_stride <= 0;
      _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start <= 0;
      _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_op_sel <= 0;
      _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_addr <= 0;
      _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_global_addr <= 0;
      _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_size <= 0;
      _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_stride <= 0;
      _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start <= 0;
      _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_op_sel <= 0;
      _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_addr <= 0;
      _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_global_addr <= 0;
      _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_size <= 0;
      _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_stride <= 0;
      _maxi_ram_w8_l2048_id11_1_write_start <= 0;
      _maxi_ram_w8_l2048_id11_1_write_op_sel <= 0;
      _maxi_ram_w8_l2048_id11_1_write_local_addr <= 0;
      _maxi_ram_w8_l2048_id11_1_write_global_addr <= 0;
      _maxi_ram_w8_l2048_id11_1_write_size <= 0;
      _maxi_ram_w8_l2048_id11_1_write_local_stride <= 0;
      _maxi_write_idle <= 1;
      _maxi_write_op_sel <= 0;
      _maxi_write_local_addr <= 0;
      _maxi_write_global_addr <= 0;
      _maxi_write_size <= 0;
      _maxi_write_local_stride <= 0;
      maxi_awaddr <= 0;
      maxi_awlen <= 0;
      maxi_awvalid <= 0;
      _tmp_1019 <= 0;
      _maxi_cond_1_1 <= 0;
      maxi_wdata <= 0;
      maxi_wvalid <= 0;
      maxi_wlast <= 0;
      maxi_wstrb <= 0;
      _tmp_1020 <= 0;
      _maxi_cond_2_1 <= 0;
      _maxi_ram_w8_l2048_id0_1_write_start <= 0;
      _maxi_ram_w8_l2048_id0_1_write_op_sel <= 0;
      _maxi_ram_w8_l2048_id0_1_write_local_addr <= 0;
      _maxi_ram_w8_l2048_id0_1_write_global_addr <= 0;
      _maxi_ram_w8_l2048_id0_1_write_size <= 0;
      _maxi_ram_w8_l2048_id0_1_write_local_stride <= 0;
      _tmp_1120 <= 0;
      _maxi_cond_3_1 <= 0;
      _maxi_ram_w8_l2048_id2_1_read_start <= 0;
      _maxi_ram_w8_l2048_id2_1_read_op_sel <= 0;
      _maxi_ram_w8_l2048_id2_1_read_local_addr <= 0;
      _maxi_ram_w8_l2048_id2_1_read_global_addr <= 0;
      _maxi_ram_w8_l2048_id2_1_read_size <= 0;
      _maxi_ram_w8_l2048_id2_1_read_local_stride <= 0;
      _maxi_ram_w4_l8192_id0_1_read_start <= 0;
      _maxi_ram_w4_l8192_id0_1_read_op_sel <= 0;
      _maxi_ram_w4_l8192_id0_1_read_local_addr <= 0;
      _maxi_ram_w4_l8192_id0_1_read_global_addr <= 0;
      _maxi_ram_w4_l8192_id0_1_read_size <= 0;
      _maxi_ram_w4_l8192_id0_1_read_local_stride <= 0;
      _maxi_ram_w8_l2048_id3_1_read_start <= 0;
      _maxi_ram_w8_l2048_id3_1_read_op_sel <= 0;
      _maxi_ram_w8_l2048_id3_1_read_local_addr <= 0;
      _maxi_ram_w8_l2048_id3_1_read_global_addr <= 0;
      _maxi_ram_w8_l2048_id3_1_read_size <= 0;
      _maxi_ram_w8_l2048_id3_1_read_local_stride <= 0;
      _maxi_ram_w8_l2048_id1_1_write_start <= 0;
      _maxi_ram_w8_l2048_id1_1_write_op_sel <= 0;
      _maxi_ram_w8_l2048_id1_1_write_local_addr <= 0;
      _maxi_ram_w8_l2048_id1_1_write_global_addr <= 0;
      _maxi_ram_w8_l2048_id1_1_write_size <= 0;
      _maxi_ram_w8_l2048_id1_1_write_local_stride <= 0;
      _tmp_1357 <= 0;
      _maxi_cond_4_1 <= 0;
    end else begin
      if(_maxi_cond_0_1) begin
        maxi_arvalid <= 0;
      end 
      if(_maxi_cond_1_1) begin
        maxi_awvalid <= 0;
      end 
      if(_maxi_cond_2_1) begin
        maxi_wvalid <= 0;
        maxi_wlast <= 0;
        _tmp_1020 <= 0;
      end 
      if(_maxi_cond_3_1) begin
        maxi_wvalid <= 0;
        maxi_wlast <= 0;
        _tmp_1120 <= 0;
      end 
      if(_maxi_cond_4_1) begin
        maxi_wvalid <= 0;
        maxi_wlast <= 0;
        _tmp_1357 <= 0;
      end 
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= _saxi_register_9;
      _maxi_ram_w8_l2048_id1_1_read_start <= 0;
      if(axim_flag_9) begin
        _maxi_ram_w8_l2048_id1_1_read_start <= 1;
        _maxi_ram_w8_l2048_id1_1_read_op_sel <= 1;
        _maxi_ram_w8_l2048_id1_1_read_local_addr <= 0;
        _maxi_ram_w8_l2048_id1_1_read_global_addr <= conv2d_16_arg_objaddr_2;
        _maxi_ram_w8_l2048_id1_1_read_size <= (cparam_conv2d_16_bias_num >> 2) + (((cparam_conv2d_16_bias_num & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id1_1_read_local_stride <= 1;
      end 
      if(_maxi_ram_w8_l2048_id1_1_read_start) begin
        _maxi_read_idle <= 0;
      end 
      if(_maxi_ram_w8_l2048_id1_1_read_start) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= _maxi_ram_w8_l2048_id1_1_read_op_sel;
        _maxi_read_local_addr <= _maxi_ram_w8_l2048_id1_1_read_local_addr;
        _maxi_read_global_addr <= _maxi_ram_w8_l2048_id1_1_read_global_addr;
        _maxi_read_size <= _maxi_ram_w8_l2048_id1_1_read_size;
        _maxi_read_local_stride <= _maxi_ram_w8_l2048_id1_1_read_local_stride;
      end 
      if((_maxi_read_fsm == 2) && ((maxi_arready || !maxi_arvalid) && (_tmp_20 == 0))) begin
        maxi_araddr <= _maxi_read_cur_global_addr;
        maxi_arlen <= _maxi_read_cur_size - 1;
        maxi_arvalid <= 1;
        _tmp_20 <= _maxi_read_cur_size;
      end 
      _maxi_cond_0_1 <= 1;
      if(maxi_arvalid && !maxi_arready) begin
        maxi_arvalid <= maxi_arvalid;
      end 
      if(maxi_rready && maxi_rvalid && (_tmp_20 > 0)) begin
        _tmp_20 <= _tmp_20 - 1;
      end 
      if(axim_flag_21) begin
        _maxi_read_idle <= 1;
      end 
      _maxi_ram_w8_l2048_id0_1_read_start <= 0;
      if(axim_flag_22) begin
        _maxi_ram_w8_l2048_id0_1_read_start <= 1;
        _maxi_ram_w8_l2048_id0_1_read_op_sel <= 2;
        _maxi_ram_w8_l2048_id0_1_read_local_addr <= 0;
        _maxi_ram_w8_l2048_id0_1_read_global_addr <= conv2d_16_arg_objaddr_3;
        _maxi_ram_w8_l2048_id0_1_read_size <= (cparam_conv2d_16_scale_num >> 2) + (((cparam_conv2d_16_scale_num & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id0_1_read_local_stride <= 1;
      end 
      if(_maxi_ram_w8_l2048_id0_1_read_start) begin
        _maxi_read_idle <= 0;
      end 
      if(_maxi_ram_w8_l2048_id0_1_read_start) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= _maxi_ram_w8_l2048_id0_1_read_op_sel;
        _maxi_read_local_addr <= _maxi_ram_w8_l2048_id0_1_read_local_addr;
        _maxi_read_global_addr <= _maxi_ram_w8_l2048_id0_1_read_global_addr;
        _maxi_read_size <= _maxi_ram_w8_l2048_id0_1_read_size;
        _maxi_read_local_stride <= _maxi_ram_w8_l2048_id0_1_read_local_stride;
      end 
      _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start <= 0;
      if(axim_flag_35) begin
        _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start <= 1;
        _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_op_sel <= 3;
        _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_addr <= conv2d_16_filter_page_dma_offset >> 3;
        _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_global_addr <= conv2d_16_arg_objaddr_1 + conv2d_16_filter_base_offset;
        _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_size <= (cparam_conv2d_16_filter_read_size >> 3) + (((cparam_conv2d_16_filter_read_size & { 3{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_stride <= 1;
      end 
      if(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start) begin
        _maxi_read_idle <= 0;
      end 
      if(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_op_sel;
        _maxi_read_local_addr <= _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_addr;
        _maxi_read_global_addr <= _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_global_addr;
        _maxi_read_size <= _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_size;
        _maxi_read_local_stride <= _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_stride;
      end 
      _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start <= 0;
      if(axim_flag_288) begin
        _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start <= 1;
        _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_op_sel <= 4;
        _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_addr <= conv2d_16_act_page_dma_offset_0 >> 2;
        _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_global_addr <= conv2d_16_mux_act_gaddr_0;
        _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_size <= (cparam_conv2d_16_act_read_size >> 2) + (((cparam_conv2d_16_act_read_size & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_stride <= 1;
      end 
      if(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start) begin
        _maxi_read_idle <= 0;
      end 
      if(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_op_sel;
        _maxi_read_local_addr <= _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_addr;
        _maxi_read_global_addr <= _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_global_addr;
        _maxi_read_size <= _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_size;
        _maxi_read_local_stride <= _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_stride;
      end 
      _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start <= 0;
      if(axim_flag_345) begin
        _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start <= 1;
        _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_op_sel <= 5;
        _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_addr <= conv2d_16_act_page_dma_offset_1 >> 2;
        _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_global_addr <= conv2d_16_mux_act_gaddr_1;
        _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_size <= (cparam_conv2d_16_act_read_size >> 2) + (((cparam_conv2d_16_act_read_size & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_stride <= 1;
      end 
      if(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start) begin
        _maxi_read_idle <= 0;
      end 
      if(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_op_sel;
        _maxi_read_local_addr <= _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_addr;
        _maxi_read_global_addr <= _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_global_addr;
        _maxi_read_size <= _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_size;
        _maxi_read_local_stride <= _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_stride;
      end 
      _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start <= 0;
      if(axim_flag_402) begin
        _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start <= 1;
        _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_op_sel <= 6;
        _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_addr <= conv2d_16_act_page_dma_offset_2 >> 2;
        _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_global_addr <= conv2d_16_mux_act_gaddr_2;
        _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_size <= (cparam_conv2d_16_act_read_size >> 2) + (((cparam_conv2d_16_act_read_size & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_stride <= 1;
      end 
      if(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start) begin
        _maxi_read_idle <= 0;
      end 
      if(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_op_sel;
        _maxi_read_local_addr <= _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_addr;
        _maxi_read_global_addr <= _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_global_addr;
        _maxi_read_size <= _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_size;
        _maxi_read_local_stride <= _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_stride;
      end 
      _maxi_ram_w8_l2048_id11_1_write_start <= 0;
      if(axim_flag_970) begin
        _maxi_ram_w8_l2048_id11_1_write_start <= 1;
        _maxi_ram_w8_l2048_id11_1_write_op_sel <= 1;
        _maxi_ram_w8_l2048_id11_1_write_local_addr <= conv2d_16_out_laddr_offset + conv2d_16_out_page_dma_offset >> 2;
        _maxi_ram_w8_l2048_id11_1_write_global_addr <= conv2d_16_objaddr + (conv2d_16_out_base_offset + cparam_conv2d_16_out_offset_values_0);
        _maxi_ram_w8_l2048_id11_1_write_size <= (conv2d_16_next_out_write_size >> 2) + (((conv2d_16_next_out_write_size & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id11_1_write_local_stride <= 1;
      end 
      if(_maxi_ram_w8_l2048_id11_1_write_start) begin
        _maxi_write_idle <= 0;
      end 
      if(_maxi_ram_w8_l2048_id11_1_write_start) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= _maxi_ram_w8_l2048_id11_1_write_op_sel;
        _maxi_write_local_addr <= _maxi_ram_w8_l2048_id11_1_write_local_addr;
        _maxi_write_global_addr <= _maxi_ram_w8_l2048_id11_1_write_global_addr;
        _maxi_write_size <= _maxi_ram_w8_l2048_id11_1_write_size;
        _maxi_write_local_stride <= _maxi_ram_w8_l2048_id11_1_write_local_stride;
      end 
      if((_maxi_write_fsm == 2) && ((maxi_awready || !maxi_awvalid) && (_tmp_1019 == 0))) begin
        maxi_awaddr <= _maxi_write_cur_global_addr;
        maxi_awlen <= _maxi_write_cur_size - 1;
        maxi_awvalid <= 1;
        _tmp_1019 <= _maxi_write_cur_size;
      end 
      if((_maxi_write_fsm == 2) && ((maxi_awready || !maxi_awvalid) && (_tmp_1019 == 0)) && (_maxi_write_cur_size == 0)) begin
        maxi_awvalid <= 0;
      end 
      _maxi_cond_1_1 <= 1;
      if(maxi_awvalid && !maxi_awready) begin
        maxi_awvalid <= maxi_awvalid;
      end 
      if(_dataflow_cat_ovalid_98 && ((_maxi_write_fsm == 3) && (_maxi_write_op_sel == 1) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid))) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid) && (_tmp_1019 > 0))) begin
        maxi_wdata <= _dataflow_cat_odata_98;
        maxi_wvalid <= 1;
        maxi_wlast <= 0;
        maxi_wstrb <= { 4{ 1'd1 } };
        _tmp_1019 <= _tmp_1019 - 1;
      end 
      if(_dataflow_cat_ovalid_98 && ((_maxi_write_fsm == 3) && (_maxi_write_op_sel == 1) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid))) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid) && (_tmp_1019 > 0)) && (_tmp_1019 == 1)) begin
        maxi_wlast <= 1;
        _tmp_1020 <= 1;
      end 
      _maxi_cond_2_1 <= 1;
      if(maxi_wvalid && !maxi_wready) begin
        maxi_wvalid <= maxi_wvalid;
        maxi_wlast <= maxi_wlast;
        _tmp_1020 <= _tmp_1020;
      end 
      if(axim_flag_1021) begin
        _maxi_write_idle <= 1;
      end 
      if(axim_flag_1022) begin
        _maxi_ram_w8_l2048_id1_1_read_start <= 1;
        _maxi_ram_w8_l2048_id1_1_read_op_sel <= 1;
        _maxi_ram_w8_l2048_id1_1_read_local_addr <= max_pool_serial_18_act_page_dma_offset >> 2;
        _maxi_ram_w8_l2048_id1_1_read_global_addr <= max_pool_serial_18_arg_objaddr_0 + (max_pool_serial_18_act_base_offset + cparam_max_pool_serial_18_act_offset_values_0);
        _maxi_ram_w8_l2048_id1_1_read_size <= (cparam_max_pool_serial_18_act_read_size >> 2) + (((cparam_max_pool_serial_18_act_read_size & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id1_1_read_local_stride <= 1;
      end 
      if(axim_flag_1023) begin
        _maxi_ram_w8_l2048_id1_1_read_start <= 1;
        _maxi_ram_w8_l2048_id1_1_read_op_sel <= 1;
        _maxi_ram_w8_l2048_id1_1_read_local_addr <= max_pool_serial_18_act_page_dma_offset + cparam_max_pool_serial_18_act_read_size >> 2;
        _maxi_ram_w8_l2048_id1_1_read_global_addr <= max_pool_serial_18_arg_objaddr_0 + (max_pool_serial_18_act_base_offset + cparam_max_pool_serial_18_act_offset_values_1);
        _maxi_ram_w8_l2048_id1_1_read_size <= (cparam_max_pool_serial_18_act_read_size >> 2) + (((cparam_max_pool_serial_18_act_read_size & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id1_1_read_local_stride <= 1;
      end 
      _maxi_ram_w8_l2048_id0_1_write_start <= 0;
      if(axim_flag_1071) begin
        _maxi_ram_w8_l2048_id0_1_write_start <= 1;
        _maxi_ram_w8_l2048_id0_1_write_op_sel <= 2;
        _maxi_ram_w8_l2048_id0_1_write_local_addr <= max_pool_serial_18_out_page_dma_offset >> 2;
        _maxi_ram_w8_l2048_id0_1_write_global_addr <= max_pool_serial_18_objaddr + max_pool_serial_18_out_base_offset;
        _maxi_ram_w8_l2048_id0_1_write_size <= (cparam_max_pool_serial_18_out_write_size >> 2) + (((cparam_max_pool_serial_18_out_write_size & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id0_1_write_local_stride <= 1;
      end 
      if(_maxi_ram_w8_l2048_id0_1_write_start) begin
        _maxi_write_idle <= 0;
      end 
      if(_maxi_ram_w8_l2048_id0_1_write_start) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= _maxi_ram_w8_l2048_id0_1_write_op_sel;
        _maxi_write_local_addr <= _maxi_ram_w8_l2048_id0_1_write_local_addr;
        _maxi_write_global_addr <= _maxi_ram_w8_l2048_id0_1_write_global_addr;
        _maxi_write_size <= _maxi_ram_w8_l2048_id0_1_write_size;
        _maxi_write_local_stride <= _maxi_ram_w8_l2048_id0_1_write_local_stride;
      end 
      if(_dataflow_cat_ovalid_107 && ((_maxi_write_fsm == 3) && (_maxi_write_op_sel == 2) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid))) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid) && (_tmp_1019 > 0))) begin
        maxi_wdata <= _dataflow_cat_odata_107;
        maxi_wvalid <= 1;
        maxi_wlast <= 0;
        maxi_wstrb <= { 4{ 1'd1 } };
        _tmp_1019 <= _tmp_1019 - 1;
      end 
      if(_dataflow_cat_ovalid_107 && ((_maxi_write_fsm == 3) && (_maxi_write_op_sel == 2) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid))) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid) && (_tmp_1019 > 0)) && (_tmp_1019 == 1)) begin
        maxi_wlast <= 1;
        _tmp_1120 <= 1;
      end 
      _maxi_cond_3_1 <= 1;
      if(maxi_wvalid && !maxi_wready) begin
        maxi_wvalid <= maxi_wvalid;
        maxi_wlast <= maxi_wlast;
        _tmp_1120 <= _tmp_1120;
      end 
      _maxi_ram_w8_l2048_id2_1_read_start <= 0;
      if(axim_flag_1121) begin
        _maxi_ram_w8_l2048_id2_1_read_start <= 1;
        _maxi_ram_w8_l2048_id2_1_read_op_sel <= 7;
        _maxi_ram_w8_l2048_id2_1_read_local_addr <= 0;
        _maxi_ram_w8_l2048_id2_1_read_global_addr <= matmul_29_arg_objaddr_2;
        _maxi_ram_w8_l2048_id2_1_read_size <= (cparam_matmul_29_bias_num >> 2) + (((cparam_matmul_29_bias_num & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id2_1_read_local_stride <= 1;
      end 
      if(_maxi_ram_w8_l2048_id2_1_read_start) begin
        _maxi_read_idle <= 0;
      end 
      if(_maxi_ram_w8_l2048_id2_1_read_start) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= _maxi_ram_w8_l2048_id2_1_read_op_sel;
        _maxi_read_local_addr <= _maxi_ram_w8_l2048_id2_1_read_local_addr;
        _maxi_read_global_addr <= _maxi_ram_w8_l2048_id2_1_read_global_addr;
        _maxi_read_size <= _maxi_ram_w8_l2048_id2_1_read_size;
        _maxi_read_local_stride <= _maxi_ram_w8_l2048_id2_1_read_local_stride;
      end 
      if(axim_flag_1132) begin
        _maxi_ram_w8_l2048_id0_1_read_start <= 1;
        _maxi_ram_w8_l2048_id0_1_read_op_sel <= 2;
        _maxi_ram_w8_l2048_id0_1_read_local_addr <= 0;
        _maxi_ram_w8_l2048_id0_1_read_global_addr <= matmul_29_arg_objaddr_3;
        _maxi_ram_w8_l2048_id0_1_read_size <= (cparam_matmul_29_scale_num >> 2) + (((cparam_matmul_29_scale_num & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id0_1_read_local_stride <= 1;
      end 
      _maxi_ram_w4_l8192_id0_1_read_start <= 0;
      if(axim_flag_1133) begin
        _maxi_ram_w4_l8192_id0_1_read_start <= 1;
        _maxi_ram_w4_l8192_id0_1_read_op_sel <= 8;
        _maxi_ram_w4_l8192_id0_1_read_local_addr <= matmul_29_filter_page_dma_offset >> 3;
        _maxi_ram_w4_l8192_id0_1_read_global_addr <= matmul_29_arg_objaddr_1 + matmul_29_filter_base_offset;
        _maxi_ram_w4_l8192_id0_1_read_size <= (cparam_matmul_29_filter_read_size >> 3) + (((cparam_matmul_29_filter_read_size & { 3{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w4_l8192_id0_1_read_local_stride <= 1;
      end 
      if(_maxi_ram_w4_l8192_id0_1_read_start) begin
        _maxi_read_idle <= 0;
      end 
      if(_maxi_ram_w4_l8192_id0_1_read_start) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= _maxi_ram_w4_l8192_id0_1_read_op_sel;
        _maxi_read_local_addr <= _maxi_ram_w4_l8192_id0_1_read_local_addr;
        _maxi_read_global_addr <= _maxi_ram_w4_l8192_id0_1_read_global_addr;
        _maxi_read_size <= _maxi_ram_w4_l8192_id0_1_read_size;
        _maxi_read_local_stride <= _maxi_ram_w4_l8192_id0_1_read_local_stride;
      end 
      _maxi_ram_w8_l2048_id3_1_read_start <= 0;
      if(axim_flag_1152) begin
        _maxi_ram_w8_l2048_id3_1_read_start <= 1;
        _maxi_ram_w8_l2048_id3_1_read_op_sel <= 9;
        _maxi_ram_w8_l2048_id3_1_read_local_addr <= matmul_29_act_page_dma_offset_0 >> 2;
        _maxi_ram_w8_l2048_id3_1_read_global_addr <= matmul_29_mux_act_gaddr_0;
        _maxi_ram_w8_l2048_id3_1_read_size <= (cparam_matmul_29_act_read_size >> 2) + (((cparam_matmul_29_act_read_size & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id3_1_read_local_stride <= 1;
      end 
      if(_maxi_ram_w8_l2048_id3_1_read_start) begin
        _maxi_read_idle <= 0;
      end 
      if(_maxi_ram_w8_l2048_id3_1_read_start) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= _maxi_ram_w8_l2048_id3_1_read_op_sel;
        _maxi_read_local_addr <= _maxi_ram_w8_l2048_id3_1_read_local_addr;
        _maxi_read_global_addr <= _maxi_ram_w8_l2048_id3_1_read_global_addr;
        _maxi_read_size <= _maxi_ram_w8_l2048_id3_1_read_size;
        _maxi_read_local_stride <= _maxi_ram_w8_l2048_id3_1_read_local_stride;
      end 
      _maxi_ram_w8_l2048_id1_1_write_start <= 0;
      if(axim_flag_1308) begin
        _maxi_ram_w8_l2048_id1_1_write_start <= 1;
        _maxi_ram_w8_l2048_id1_1_write_op_sel <= 3;
        _maxi_ram_w8_l2048_id1_1_write_local_addr <= matmul_29_out_laddr_offset + matmul_29_out_page_dma_offset >> 2;
        _maxi_ram_w8_l2048_id1_1_write_global_addr <= matmul_29_objaddr + (matmul_29_out_base_offset + cparam_matmul_29_out_offset_values_0);
        _maxi_ram_w8_l2048_id1_1_write_size <= (matmul_29_next_out_write_size >> 2) + (((matmul_29_next_out_write_size & { 2{ 1'd1 } }) > 0)? 1 : 0);
        _maxi_ram_w8_l2048_id1_1_write_local_stride <= 1;
      end 
      if(_maxi_ram_w8_l2048_id1_1_write_start) begin
        _maxi_write_idle <= 0;
      end 
      if(_maxi_ram_w8_l2048_id1_1_write_start) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= _maxi_ram_w8_l2048_id1_1_write_op_sel;
        _maxi_write_local_addr <= _maxi_ram_w8_l2048_id1_1_write_local_addr;
        _maxi_write_global_addr <= _maxi_ram_w8_l2048_id1_1_write_global_addr;
        _maxi_write_size <= _maxi_ram_w8_l2048_id1_1_write_size;
        _maxi_write_local_stride <= _maxi_ram_w8_l2048_id1_1_write_local_stride;
      end 
      if(_dataflow_cat_ovalid_167 && ((_maxi_write_fsm == 3) && (_maxi_write_op_sel == 3) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid))) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid) && (_tmp_1019 > 0))) begin
        maxi_wdata <= _dataflow_cat_odata_167;
        maxi_wvalid <= 1;
        maxi_wlast <= 0;
        maxi_wstrb <= { 4{ 1'd1 } };
        _tmp_1019 <= _tmp_1019 - 1;
      end 
      if(_dataflow_cat_ovalid_167 && ((_maxi_write_fsm == 3) && (_maxi_write_op_sel == 3) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid))) && ((_tmp_1019 > 0) && (maxi_wready || !maxi_wvalid) && (_tmp_1019 > 0)) && (_tmp_1019 == 1)) begin
        maxi_wlast <= 1;
        _tmp_1357 <= 1;
      end 
      _maxi_cond_4_1 <= 1;
      if(maxi_wvalid && !maxi_wready) begin
        maxi_wvalid <= maxi_wvalid;
        maxi_wlast <= maxi_wlast;
        _tmp_1357 <= _tmp_1357;
      end 
    end
  end

  reg [8-1:0] _dataflow_slice_data_3;
  reg _dataflow_slice_valid_3;
  wire _dataflow_slice_ready_3;
  reg [8-1:0] _dataflow_slice_data_6;
  reg _dataflow_slice_valid_6;
  wire _dataflow_slice_ready_6;
  reg [8-1:0] _dataflow_slice_data_9;
  reg _dataflow_slice_valid_9;
  wire _dataflow_slice_ready_9;
  reg [8-1:0] _dataflow_slice_data_12;
  reg _dataflow_slice_valid_12;
  wire _dataflow_slice_ready_12;
  reg [8-1:0] _dataflow_slice_data_16;
  reg _dataflow_slice_valid_16;
  wire _dataflow_slice_ready_16;
  reg [8-1:0] _dataflow_slice_data_19;
  reg _dataflow_slice_valid_19;
  wire _dataflow_slice_ready_19;
  reg [8-1:0] _dataflow_slice_data_22;
  reg _dataflow_slice_valid_22;
  wire _dataflow_slice_ready_22;
  reg [8-1:0] _dataflow_slice_data_25;
  reg _dataflow_slice_valid_25;
  wire _dataflow_slice_ready_25;
  reg [4-1:0] _dataflow_slice_data_29;
  reg _dataflow_slice_valid_29;
  wire _dataflow_slice_ready_29;
  reg [4-1:0] _dataflow_slice_data_32;
  reg _dataflow_slice_valid_32;
  wire _dataflow_slice_ready_32;
  reg [4-1:0] _dataflow_slice_data_35;
  reg _dataflow_slice_valid_35;
  wire _dataflow_slice_ready_35;
  reg [4-1:0] _dataflow_slice_data_38;
  reg _dataflow_slice_valid_38;
  wire _dataflow_slice_ready_38;
  reg [4-1:0] _dataflow_slice_data_41;
  reg _dataflow_slice_valid_41;
  wire _dataflow_slice_ready_41;
  reg [4-1:0] _dataflow_slice_data_44;
  reg _dataflow_slice_valid_44;
  wire _dataflow_slice_ready_44;
  reg [4-1:0] _dataflow_slice_data_47;
  reg _dataflow_slice_valid_47;
  wire _dataflow_slice_ready_47;
  reg [4-1:0] _dataflow_slice_data_50;
  reg _dataflow_slice_valid_50;
  wire _dataflow_slice_ready_50;
  reg [8-1:0] _dataflow_slice_data_54;
  reg _dataflow_slice_valid_54;
  wire _dataflow_slice_ready_54;
  reg [8-1:0] _dataflow_slice_data_57;
  reg _dataflow_slice_valid_57;
  wire _dataflow_slice_ready_57;
  reg [8-1:0] _dataflow_slice_data_60;
  reg _dataflow_slice_valid_60;
  wire _dataflow_slice_ready_60;
  reg [8-1:0] _dataflow_slice_data_63;
  reg _dataflow_slice_valid_63;
  wire _dataflow_slice_ready_63;
  reg [8-1:0] _dataflow_slice_data_67;
  reg _dataflow_slice_valid_67;
  wire _dataflow_slice_ready_67;
  reg [8-1:0] _dataflow_slice_data_70;
  reg _dataflow_slice_valid_70;
  wire _dataflow_slice_ready_70;
  reg [8-1:0] _dataflow_slice_data_73;
  reg _dataflow_slice_valid_73;
  wire _dataflow_slice_ready_73;
  reg [8-1:0] _dataflow_slice_data_76;
  reg _dataflow_slice_valid_76;
  wire _dataflow_slice_ready_76;
  reg [8-1:0] _dataflow_slice_data_80;
  reg _dataflow_slice_valid_80;
  wire _dataflow_slice_ready_80;
  reg [8-1:0] _dataflow_slice_data_83;
  reg _dataflow_slice_valid_83;
  wire _dataflow_slice_ready_83;
  reg [8-1:0] _dataflow_slice_data_86;
  reg _dataflow_slice_valid_86;
  wire _dataflow_slice_ready_86;
  reg [8-1:0] _dataflow_slice_data_89;
  reg _dataflow_slice_valid_89;
  wire _dataflow_slice_ready_89;
  reg [8-1:0] _dataflow_slice_data_111;
  reg _dataflow_slice_valid_111;
  wire _dataflow_slice_ready_111;
  reg [8-1:0] _dataflow_slice_data_114;
  reg _dataflow_slice_valid_114;
  wire _dataflow_slice_ready_114;
  reg [8-1:0] _dataflow_slice_data_117;
  reg _dataflow_slice_valid_117;
  wire _dataflow_slice_ready_117;
  reg [8-1:0] _dataflow_slice_data_120;
  reg _dataflow_slice_valid_120;
  wire _dataflow_slice_ready_120;
  reg [4-1:0] _dataflow_slice_data_124;
  reg _dataflow_slice_valid_124;
  wire _dataflow_slice_ready_124;
  reg [4-1:0] _dataflow_slice_data_127;
  reg _dataflow_slice_valid_127;
  wire _dataflow_slice_ready_127;
  reg [4-1:0] _dataflow_slice_data_130;
  reg _dataflow_slice_valid_130;
  wire _dataflow_slice_ready_130;
  reg [4-1:0] _dataflow_slice_data_133;
  reg _dataflow_slice_valid_133;
  wire _dataflow_slice_ready_133;
  reg [4-1:0] _dataflow_slice_data_136;
  reg _dataflow_slice_valid_136;
  wire _dataflow_slice_ready_136;
  reg [4-1:0] _dataflow_slice_data_139;
  reg _dataflow_slice_valid_139;
  wire _dataflow_slice_ready_139;
  reg [4-1:0] _dataflow_slice_data_142;
  reg _dataflow_slice_valid_142;
  wire _dataflow_slice_ready_142;
  reg [4-1:0] _dataflow_slice_data_145;
  reg _dataflow_slice_valid_145;
  wire _dataflow_slice_ready_145;
  reg [8-1:0] _dataflow_slice_data_149;
  reg _dataflow_slice_valid_149;
  wire _dataflow_slice_ready_149;
  reg [8-1:0] _dataflow_slice_data_152;
  reg _dataflow_slice_valid_152;
  wire _dataflow_slice_ready_152;
  reg [8-1:0] _dataflow_slice_data_155;
  reg _dataflow_slice_valid_155;
  wire _dataflow_slice_ready_155;
  reg [8-1:0] _dataflow_slice_data_158;
  reg _dataflow_slice_valid_158;
  wire _dataflow_slice_ready_158;
  assign _dataflow_slice_odata_3 = _dataflow_slice_data_3;
  assign _dataflow_slice_ovalid_3 = _dataflow_slice_valid_3;
  assign _dataflow_slice_ready_3 = _dataflow_slice_oready_3;
  assign _dataflow_slice_odata_6 = _dataflow_slice_data_6;
  assign _dataflow_slice_ovalid_6 = _dataflow_slice_valid_6;
  assign _dataflow_slice_ready_6 = _dataflow_slice_oready_6;
  assign _dataflow_slice_odata_9 = _dataflow_slice_data_9;
  assign _dataflow_slice_ovalid_9 = _dataflow_slice_valid_9;
  assign _dataflow_slice_ready_9 = _dataflow_slice_oready_9;
  assign _dataflow_slice_odata_12 = _dataflow_slice_data_12;
  assign _dataflow_slice_ovalid_12 = _dataflow_slice_valid_12;
  assign _dataflow_slice_ready_12 = _dataflow_slice_oready_12;
  assign _dataflow_slice_odata_16 = _dataflow_slice_data_16;
  assign _dataflow_slice_ovalid_16 = _dataflow_slice_valid_16;
  assign _dataflow_slice_ready_16 = _dataflow_slice_oready_16;
  assign _dataflow_slice_odata_19 = _dataflow_slice_data_19;
  assign _dataflow_slice_ovalid_19 = _dataflow_slice_valid_19;
  assign _dataflow_slice_ready_19 = _dataflow_slice_oready_19;
  assign _dataflow_slice_odata_22 = _dataflow_slice_data_22;
  assign _dataflow_slice_ovalid_22 = _dataflow_slice_valid_22;
  assign _dataflow_slice_ready_22 = _dataflow_slice_oready_22;
  assign _dataflow_slice_odata_25 = _dataflow_slice_data_25;
  assign _dataflow_slice_ovalid_25 = _dataflow_slice_valid_25;
  assign _dataflow_slice_ready_25 = _dataflow_slice_oready_25;
  assign _dataflow_slice_odata_29 = _dataflow_slice_data_29;
  assign _dataflow_slice_ovalid_29 = _dataflow_slice_valid_29;
  assign _dataflow_slice_ready_29 = _dataflow_slice_oready_29;
  assign _dataflow_slice_odata_32 = _dataflow_slice_data_32;
  assign _dataflow_slice_ovalid_32 = _dataflow_slice_valid_32;
  assign _dataflow_slice_ready_32 = _dataflow_slice_oready_32;
  assign _dataflow_slice_odata_35 = _dataflow_slice_data_35;
  assign _dataflow_slice_ovalid_35 = _dataflow_slice_valid_35;
  assign _dataflow_slice_ready_35 = _dataflow_slice_oready_35;
  assign _dataflow_slice_odata_38 = _dataflow_slice_data_38;
  assign _dataflow_slice_ovalid_38 = _dataflow_slice_valid_38;
  assign _dataflow_slice_ready_38 = _dataflow_slice_oready_38;
  assign _dataflow_slice_odata_41 = _dataflow_slice_data_41;
  assign _dataflow_slice_ovalid_41 = _dataflow_slice_valid_41;
  assign _dataflow_slice_ready_41 = _dataflow_slice_oready_41;
  assign _dataflow_slice_odata_44 = _dataflow_slice_data_44;
  assign _dataflow_slice_ovalid_44 = _dataflow_slice_valid_44;
  assign _dataflow_slice_ready_44 = _dataflow_slice_oready_44;
  assign _dataflow_slice_odata_47 = _dataflow_slice_data_47;
  assign _dataflow_slice_ovalid_47 = _dataflow_slice_valid_47;
  assign _dataflow_slice_ready_47 = _dataflow_slice_oready_47;
  assign _dataflow_slice_odata_50 = _dataflow_slice_data_50;
  assign _dataflow_slice_ovalid_50 = _dataflow_slice_valid_50;
  assign _dataflow_slice_ready_50 = _dataflow_slice_oready_50;
  assign _dataflow_slice_odata_54 = _dataflow_slice_data_54;
  assign _dataflow_slice_ovalid_54 = _dataflow_slice_valid_54;
  assign _dataflow_slice_ready_54 = _dataflow_slice_oready_54;
  assign _dataflow_slice_odata_57 = _dataflow_slice_data_57;
  assign _dataflow_slice_ovalid_57 = _dataflow_slice_valid_57;
  assign _dataflow_slice_ready_57 = _dataflow_slice_oready_57;
  assign _dataflow_slice_odata_60 = _dataflow_slice_data_60;
  assign _dataflow_slice_ovalid_60 = _dataflow_slice_valid_60;
  assign _dataflow_slice_ready_60 = _dataflow_slice_oready_60;
  assign _dataflow_slice_odata_63 = _dataflow_slice_data_63;
  assign _dataflow_slice_ovalid_63 = _dataflow_slice_valid_63;
  assign _dataflow_slice_ready_63 = _dataflow_slice_oready_63;
  assign _dataflow_slice_odata_67 = _dataflow_slice_data_67;
  assign _dataflow_slice_ovalid_67 = _dataflow_slice_valid_67;
  assign _dataflow_slice_ready_67 = _dataflow_slice_oready_67;
  assign _dataflow_slice_odata_70 = _dataflow_slice_data_70;
  assign _dataflow_slice_ovalid_70 = _dataflow_slice_valid_70;
  assign _dataflow_slice_ready_70 = _dataflow_slice_oready_70;
  assign _dataflow_slice_odata_73 = _dataflow_slice_data_73;
  assign _dataflow_slice_ovalid_73 = _dataflow_slice_valid_73;
  assign _dataflow_slice_ready_73 = _dataflow_slice_oready_73;
  assign _dataflow_slice_odata_76 = _dataflow_slice_data_76;
  assign _dataflow_slice_ovalid_76 = _dataflow_slice_valid_76;
  assign _dataflow_slice_ready_76 = _dataflow_slice_oready_76;
  assign _dataflow_slice_odata_80 = _dataflow_slice_data_80;
  assign _dataflow_slice_ovalid_80 = _dataflow_slice_valid_80;
  assign _dataflow_slice_ready_80 = _dataflow_slice_oready_80;
  assign _dataflow_slice_odata_83 = _dataflow_slice_data_83;
  assign _dataflow_slice_ovalid_83 = _dataflow_slice_valid_83;
  assign _dataflow_slice_ready_83 = _dataflow_slice_oready_83;
  assign _dataflow_slice_odata_86 = _dataflow_slice_data_86;
  assign _dataflow_slice_ovalid_86 = _dataflow_slice_valid_86;
  assign _dataflow_slice_ready_86 = _dataflow_slice_oready_86;
  assign _dataflow_slice_odata_89 = _dataflow_slice_data_89;
  assign _dataflow_slice_ovalid_89 = _dataflow_slice_valid_89;
  assign _dataflow_slice_ready_89 = _dataflow_slice_oready_89;
  assign _dataflow_slice_odata_111 = _dataflow_slice_data_111;
  assign _dataflow_slice_ovalid_111 = _dataflow_slice_valid_111;
  assign _dataflow_slice_ready_111 = _dataflow_slice_oready_111;
  assign _dataflow_slice_odata_114 = _dataflow_slice_data_114;
  assign _dataflow_slice_ovalid_114 = _dataflow_slice_valid_114;
  assign _dataflow_slice_ready_114 = _dataflow_slice_oready_114;
  assign _dataflow_slice_odata_117 = _dataflow_slice_data_117;
  assign _dataflow_slice_ovalid_117 = _dataflow_slice_valid_117;
  assign _dataflow_slice_ready_117 = _dataflow_slice_oready_117;
  assign _dataflow_slice_odata_120 = _dataflow_slice_data_120;
  assign _dataflow_slice_ovalid_120 = _dataflow_slice_valid_120;
  assign _dataflow_slice_ready_120 = _dataflow_slice_oready_120;
  assign _dataflow_slice_odata_124 = _dataflow_slice_data_124;
  assign _dataflow_slice_ovalid_124 = _dataflow_slice_valid_124;
  assign _dataflow_slice_ready_124 = _dataflow_slice_oready_124;
  assign _dataflow_slice_odata_127 = _dataflow_slice_data_127;
  assign _dataflow_slice_ovalid_127 = _dataflow_slice_valid_127;
  assign _dataflow_slice_ready_127 = _dataflow_slice_oready_127;
  assign _dataflow_slice_odata_130 = _dataflow_slice_data_130;
  assign _dataflow_slice_ovalid_130 = _dataflow_slice_valid_130;
  assign _dataflow_slice_ready_130 = _dataflow_slice_oready_130;
  assign _dataflow_slice_odata_133 = _dataflow_slice_data_133;
  assign _dataflow_slice_ovalid_133 = _dataflow_slice_valid_133;
  assign _dataflow_slice_ready_133 = _dataflow_slice_oready_133;
  assign _dataflow_slice_odata_136 = _dataflow_slice_data_136;
  assign _dataflow_slice_ovalid_136 = _dataflow_slice_valid_136;
  assign _dataflow_slice_ready_136 = _dataflow_slice_oready_136;
  assign _dataflow_slice_odata_139 = _dataflow_slice_data_139;
  assign _dataflow_slice_ovalid_139 = _dataflow_slice_valid_139;
  assign _dataflow_slice_ready_139 = _dataflow_slice_oready_139;
  assign _dataflow_slice_odata_142 = _dataflow_slice_data_142;
  assign _dataflow_slice_ovalid_142 = _dataflow_slice_valid_142;
  assign _dataflow_slice_ready_142 = _dataflow_slice_oready_142;
  assign _dataflow_slice_odata_145 = _dataflow_slice_data_145;
  assign _dataflow_slice_ovalid_145 = _dataflow_slice_valid_145;
  assign _dataflow_slice_ready_145 = _dataflow_slice_oready_145;
  assign _dataflow_slice_odata_149 = _dataflow_slice_data_149;
  assign _dataflow_slice_ovalid_149 = _dataflow_slice_valid_149;
  assign _dataflow_slice_ready_149 = _dataflow_slice_oready_149;
  assign _dataflow_slice_odata_152 = _dataflow_slice_data_152;
  assign _dataflow_slice_ovalid_152 = _dataflow_slice_valid_152;
  assign _dataflow_slice_ready_152 = _dataflow_slice_oready_152;
  assign _dataflow_slice_odata_155 = _dataflow_slice_data_155;
  assign _dataflow_slice_ovalid_155 = _dataflow_slice_valid_155;
  assign _dataflow_slice_ready_155 = _dataflow_slice_oready_155;
  assign _dataflow_slice_odata_158 = _dataflow_slice_data_158;
  assign _dataflow_slice_ovalid_158 = _dataflow_slice_valid_158;
  assign _dataflow_slice_ready_158 = _dataflow_slice_oready_158;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _dataflow_slice_data_3 <= 0;
      _dataflow_slice_valid_3 <= 0;
      _dataflow_slice_data_6 <= 0;
      _dataflow_slice_valid_6 <= 0;
      _dataflow_slice_data_9 <= 0;
      _dataflow_slice_valid_9 <= 0;
      _dataflow_slice_data_12 <= 0;
      _dataflow_slice_valid_12 <= 0;
      _dataflow_slice_data_16 <= 0;
      _dataflow_slice_valid_16 <= 0;
      _dataflow_slice_data_19 <= 0;
      _dataflow_slice_valid_19 <= 0;
      _dataflow_slice_data_22 <= 0;
      _dataflow_slice_valid_22 <= 0;
      _dataflow_slice_data_25 <= 0;
      _dataflow_slice_valid_25 <= 0;
      _dataflow_slice_data_29 <= 0;
      _dataflow_slice_valid_29 <= 0;
      _dataflow_slice_data_32 <= 0;
      _dataflow_slice_valid_32 <= 0;
      _dataflow_slice_data_35 <= 0;
      _dataflow_slice_valid_35 <= 0;
      _dataflow_slice_data_38 <= 0;
      _dataflow_slice_valid_38 <= 0;
      _dataflow_slice_data_41 <= 0;
      _dataflow_slice_valid_41 <= 0;
      _dataflow_slice_data_44 <= 0;
      _dataflow_slice_valid_44 <= 0;
      _dataflow_slice_data_47 <= 0;
      _dataflow_slice_valid_47 <= 0;
      _dataflow_slice_data_50 <= 0;
      _dataflow_slice_valid_50 <= 0;
      _dataflow_slice_data_54 <= 0;
      _dataflow_slice_valid_54 <= 0;
      _dataflow_slice_data_57 <= 0;
      _dataflow_slice_valid_57 <= 0;
      _dataflow_slice_data_60 <= 0;
      _dataflow_slice_valid_60 <= 0;
      _dataflow_slice_data_63 <= 0;
      _dataflow_slice_valid_63 <= 0;
      _dataflow_slice_data_67 <= 0;
      _dataflow_slice_valid_67 <= 0;
      _dataflow_slice_data_70 <= 0;
      _dataflow_slice_valid_70 <= 0;
      _dataflow_slice_data_73 <= 0;
      _dataflow_slice_valid_73 <= 0;
      _dataflow_slice_data_76 <= 0;
      _dataflow_slice_valid_76 <= 0;
      _dataflow_slice_data_80 <= 0;
      _dataflow_slice_valid_80 <= 0;
      _dataflow_slice_data_83 <= 0;
      _dataflow_slice_valid_83 <= 0;
      _dataflow_slice_data_86 <= 0;
      _dataflow_slice_valid_86 <= 0;
      _dataflow_slice_data_89 <= 0;
      _dataflow_slice_valid_89 <= 0;
      _dataflow_slice_data_111 <= 0;
      _dataflow_slice_valid_111 <= 0;
      _dataflow_slice_data_114 <= 0;
      _dataflow_slice_valid_114 <= 0;
      _dataflow_slice_data_117 <= 0;
      _dataflow_slice_valid_117 <= 0;
      _dataflow_slice_data_120 <= 0;
      _dataflow_slice_valid_120 <= 0;
      _dataflow_slice_data_124 <= 0;
      _dataflow_slice_valid_124 <= 0;
      _dataflow_slice_data_127 <= 0;
      _dataflow_slice_valid_127 <= 0;
      _dataflow_slice_data_130 <= 0;
      _dataflow_slice_valid_130 <= 0;
      _dataflow_slice_data_133 <= 0;
      _dataflow_slice_valid_133 <= 0;
      _dataflow_slice_data_136 <= 0;
      _dataflow_slice_valid_136 <= 0;
      _dataflow_slice_data_139 <= 0;
      _dataflow_slice_valid_139 <= 0;
      _dataflow_slice_data_142 <= 0;
      _dataflow_slice_valid_142 <= 0;
      _dataflow_slice_data_145 <= 0;
      _dataflow_slice_valid_145 <= 0;
      _dataflow_slice_data_149 <= 0;
      _dataflow_slice_valid_149 <= 0;
      _dataflow_slice_data_152 <= 0;
      _dataflow_slice_valid_152 <= 0;
      _dataflow_slice_data_155 <= 0;
      _dataflow_slice_valid_155 <= 0;
      _dataflow_slice_data_158 <= 0;
      _dataflow_slice_valid_158 <= 0;
    end else begin
      if((_dataflow_slice_ready_3 || !_dataflow_slice_valid_3) && 1 && _wvalid_11) begin
        _dataflow_slice_data_3 <= _wdata_10[4'd7:1'd0];
      end 
      if(_dataflow_slice_valid_3 && _dataflow_slice_ready_3) begin
        _dataflow_slice_valid_3 <= 0;
      end 
      if((_dataflow_slice_ready_3 || !_dataflow_slice_valid_3) && 1) begin
        _dataflow_slice_valid_3 <= _wvalid_11;
      end 
      if((_dataflow_slice_ready_6 || !_dataflow_slice_valid_6) && 1 && _wvalid_11) begin
        _dataflow_slice_data_6 <= _wdata_10[5'd15:5'd8];
      end 
      if(_dataflow_slice_valid_6 && _dataflow_slice_ready_6) begin
        _dataflow_slice_valid_6 <= 0;
      end 
      if((_dataflow_slice_ready_6 || !_dataflow_slice_valid_6) && 1) begin
        _dataflow_slice_valid_6 <= _wvalid_11;
      end 
      if((_dataflow_slice_ready_9 || !_dataflow_slice_valid_9) && 1 && _wvalid_11) begin
        _dataflow_slice_data_9 <= _wdata_10[6'd23:6'd16];
      end 
      if(_dataflow_slice_valid_9 && _dataflow_slice_ready_9) begin
        _dataflow_slice_valid_9 <= 0;
      end 
      if((_dataflow_slice_ready_9 || !_dataflow_slice_valid_9) && 1) begin
        _dataflow_slice_valid_9 <= _wvalid_11;
      end 
      if((_dataflow_slice_ready_12 || !_dataflow_slice_valid_12) && 1 && _wvalid_11) begin
        _dataflow_slice_data_12 <= _wdata_10[6'd31:6'd24];
      end 
      if(_dataflow_slice_valid_12 && _dataflow_slice_ready_12) begin
        _dataflow_slice_valid_12 <= 0;
      end 
      if((_dataflow_slice_ready_12 || !_dataflow_slice_valid_12) && 1) begin
        _dataflow_slice_valid_12 <= _wvalid_11;
      end 
      if((_dataflow_slice_ready_16 || !_dataflow_slice_valid_16) && 1 && _wvalid_24) begin
        _dataflow_slice_data_16 <= _wdata_23[4'd7:1'd0];
      end 
      if(_dataflow_slice_valid_16 && _dataflow_slice_ready_16) begin
        _dataflow_slice_valid_16 <= 0;
      end 
      if((_dataflow_slice_ready_16 || !_dataflow_slice_valid_16) && 1) begin
        _dataflow_slice_valid_16 <= _wvalid_24;
      end 
      if((_dataflow_slice_ready_19 || !_dataflow_slice_valid_19) && 1 && _wvalid_24) begin
        _dataflow_slice_data_19 <= _wdata_23[5'd15:5'd8];
      end 
      if(_dataflow_slice_valid_19 && _dataflow_slice_ready_19) begin
        _dataflow_slice_valid_19 <= 0;
      end 
      if((_dataflow_slice_ready_19 || !_dataflow_slice_valid_19) && 1) begin
        _dataflow_slice_valid_19 <= _wvalid_24;
      end 
      if((_dataflow_slice_ready_22 || !_dataflow_slice_valid_22) && 1 && _wvalid_24) begin
        _dataflow_slice_data_22 <= _wdata_23[6'd23:6'd16];
      end 
      if(_dataflow_slice_valid_22 && _dataflow_slice_ready_22) begin
        _dataflow_slice_valid_22 <= 0;
      end 
      if((_dataflow_slice_ready_22 || !_dataflow_slice_valid_22) && 1) begin
        _dataflow_slice_valid_22 <= _wvalid_24;
      end 
      if((_dataflow_slice_ready_25 || !_dataflow_slice_valid_25) && 1 && _wvalid_24) begin
        _dataflow_slice_data_25 <= _wdata_23[6'd31:6'd24];
      end 
      if(_dataflow_slice_valid_25 && _dataflow_slice_ready_25) begin
        _dataflow_slice_valid_25 <= 0;
      end 
      if((_dataflow_slice_ready_25 || !_dataflow_slice_valid_25) && 1) begin
        _dataflow_slice_valid_25 <= _wvalid_24;
      end 
      if((_dataflow_slice_ready_29 || !_dataflow_slice_valid_29) && 1 && _wvalid_37) begin
        _dataflow_slice_data_29 <= _wdata_36[3'd3:1'd0];
      end 
      if(_dataflow_slice_valid_29 && _dataflow_slice_ready_29) begin
        _dataflow_slice_valid_29 <= 0;
      end 
      if((_dataflow_slice_ready_29 || !_dataflow_slice_valid_29) && 1) begin
        _dataflow_slice_valid_29 <= _wvalid_37;
      end 
      if((_dataflow_slice_ready_32 || !_dataflow_slice_valid_32) && 1 && _wvalid_37) begin
        _dataflow_slice_data_32 <= _wdata_36[4'd7:4'd4];
      end 
      if(_dataflow_slice_valid_32 && _dataflow_slice_ready_32) begin
        _dataflow_slice_valid_32 <= 0;
      end 
      if((_dataflow_slice_ready_32 || !_dataflow_slice_valid_32) && 1) begin
        _dataflow_slice_valid_32 <= _wvalid_37;
      end 
      if((_dataflow_slice_ready_35 || !_dataflow_slice_valid_35) && 1 && _wvalid_37) begin
        _dataflow_slice_data_35 <= _wdata_36[5'd11:5'd8];
      end 
      if(_dataflow_slice_valid_35 && _dataflow_slice_ready_35) begin
        _dataflow_slice_valid_35 <= 0;
      end 
      if((_dataflow_slice_ready_35 || !_dataflow_slice_valid_35) && 1) begin
        _dataflow_slice_valid_35 <= _wvalid_37;
      end 
      if((_dataflow_slice_ready_38 || !_dataflow_slice_valid_38) && 1 && _wvalid_37) begin
        _dataflow_slice_data_38 <= _wdata_36[5'd15:5'd12];
      end 
      if(_dataflow_slice_valid_38 && _dataflow_slice_ready_38) begin
        _dataflow_slice_valid_38 <= 0;
      end 
      if((_dataflow_slice_ready_38 || !_dataflow_slice_valid_38) && 1) begin
        _dataflow_slice_valid_38 <= _wvalid_37;
      end 
      if((_dataflow_slice_ready_41 || !_dataflow_slice_valid_41) && 1 && _wvalid_37) begin
        _dataflow_slice_data_41 <= _wdata_36[6'd19:6'd16];
      end 
      if(_dataflow_slice_valid_41 && _dataflow_slice_ready_41) begin
        _dataflow_slice_valid_41 <= 0;
      end 
      if((_dataflow_slice_ready_41 || !_dataflow_slice_valid_41) && 1) begin
        _dataflow_slice_valid_41 <= _wvalid_37;
      end 
      if((_dataflow_slice_ready_44 || !_dataflow_slice_valid_44) && 1 && _wvalid_37) begin
        _dataflow_slice_data_44 <= _wdata_36[6'd23:6'd20];
      end 
      if(_dataflow_slice_valid_44 && _dataflow_slice_ready_44) begin
        _dataflow_slice_valid_44 <= 0;
      end 
      if((_dataflow_slice_ready_44 || !_dataflow_slice_valid_44) && 1) begin
        _dataflow_slice_valid_44 <= _wvalid_37;
      end 
      if((_dataflow_slice_ready_47 || !_dataflow_slice_valid_47) && 1 && _wvalid_37) begin
        _dataflow_slice_data_47 <= _wdata_36[6'd27:6'd24];
      end 
      if(_dataflow_slice_valid_47 && _dataflow_slice_ready_47) begin
        _dataflow_slice_valid_47 <= 0;
      end 
      if((_dataflow_slice_ready_47 || !_dataflow_slice_valid_47) && 1) begin
        _dataflow_slice_valid_47 <= _wvalid_37;
      end 
      if((_dataflow_slice_ready_50 || !_dataflow_slice_valid_50) && 1 && _wvalid_37) begin
        _dataflow_slice_data_50 <= _wdata_36[6'd31:6'd28];
      end 
      if(_dataflow_slice_valid_50 && _dataflow_slice_ready_50) begin
        _dataflow_slice_valid_50 <= 0;
      end 
      if((_dataflow_slice_ready_50 || !_dataflow_slice_valid_50) && 1) begin
        _dataflow_slice_valid_50 <= _wvalid_37;
      end 
      if((_dataflow_slice_ready_54 || !_dataflow_slice_valid_54) && 1 && _wvalid_290) begin
        _dataflow_slice_data_54 <= _wdata_289[4'd7:1'd0];
      end 
      if(_dataflow_slice_valid_54 && _dataflow_slice_ready_54) begin
        _dataflow_slice_valid_54 <= 0;
      end 
      if((_dataflow_slice_ready_54 || !_dataflow_slice_valid_54) && 1) begin
        _dataflow_slice_valid_54 <= _wvalid_290;
      end 
      if((_dataflow_slice_ready_57 || !_dataflow_slice_valid_57) && 1 && _wvalid_290) begin
        _dataflow_slice_data_57 <= _wdata_289[5'd15:5'd8];
      end 
      if(_dataflow_slice_valid_57 && _dataflow_slice_ready_57) begin
        _dataflow_slice_valid_57 <= 0;
      end 
      if((_dataflow_slice_ready_57 || !_dataflow_slice_valid_57) && 1) begin
        _dataflow_slice_valid_57 <= _wvalid_290;
      end 
      if((_dataflow_slice_ready_60 || !_dataflow_slice_valid_60) && 1 && _wvalid_290) begin
        _dataflow_slice_data_60 <= _wdata_289[6'd23:6'd16];
      end 
      if(_dataflow_slice_valid_60 && _dataflow_slice_ready_60) begin
        _dataflow_slice_valid_60 <= 0;
      end 
      if((_dataflow_slice_ready_60 || !_dataflow_slice_valid_60) && 1) begin
        _dataflow_slice_valid_60 <= _wvalid_290;
      end 
      if((_dataflow_slice_ready_63 || !_dataflow_slice_valid_63) && 1 && _wvalid_290) begin
        _dataflow_slice_data_63 <= _wdata_289[6'd31:6'd24];
      end 
      if(_dataflow_slice_valid_63 && _dataflow_slice_ready_63) begin
        _dataflow_slice_valid_63 <= 0;
      end 
      if((_dataflow_slice_ready_63 || !_dataflow_slice_valid_63) && 1) begin
        _dataflow_slice_valid_63 <= _wvalid_290;
      end 
      if((_dataflow_slice_ready_67 || !_dataflow_slice_valid_67) && 1 && _wvalid_347) begin
        _dataflow_slice_data_67 <= _wdata_346[4'd7:1'd0];
      end 
      if(_dataflow_slice_valid_67 && _dataflow_slice_ready_67) begin
        _dataflow_slice_valid_67 <= 0;
      end 
      if((_dataflow_slice_ready_67 || !_dataflow_slice_valid_67) && 1) begin
        _dataflow_slice_valid_67 <= _wvalid_347;
      end 
      if((_dataflow_slice_ready_70 || !_dataflow_slice_valid_70) && 1 && _wvalid_347) begin
        _dataflow_slice_data_70 <= _wdata_346[5'd15:5'd8];
      end 
      if(_dataflow_slice_valid_70 && _dataflow_slice_ready_70) begin
        _dataflow_slice_valid_70 <= 0;
      end 
      if((_dataflow_slice_ready_70 || !_dataflow_slice_valid_70) && 1) begin
        _dataflow_slice_valid_70 <= _wvalid_347;
      end 
      if((_dataflow_slice_ready_73 || !_dataflow_slice_valid_73) && 1 && _wvalid_347) begin
        _dataflow_slice_data_73 <= _wdata_346[6'd23:6'd16];
      end 
      if(_dataflow_slice_valid_73 && _dataflow_slice_ready_73) begin
        _dataflow_slice_valid_73 <= 0;
      end 
      if((_dataflow_slice_ready_73 || !_dataflow_slice_valid_73) && 1) begin
        _dataflow_slice_valid_73 <= _wvalid_347;
      end 
      if((_dataflow_slice_ready_76 || !_dataflow_slice_valid_76) && 1 && _wvalid_347) begin
        _dataflow_slice_data_76 <= _wdata_346[6'd31:6'd24];
      end 
      if(_dataflow_slice_valid_76 && _dataflow_slice_ready_76) begin
        _dataflow_slice_valid_76 <= 0;
      end 
      if((_dataflow_slice_ready_76 || !_dataflow_slice_valid_76) && 1) begin
        _dataflow_slice_valid_76 <= _wvalid_347;
      end 
      if((_dataflow_slice_ready_80 || !_dataflow_slice_valid_80) && 1 && _wvalid_404) begin
        _dataflow_slice_data_80 <= _wdata_403[4'd7:1'd0];
      end 
      if(_dataflow_slice_valid_80 && _dataflow_slice_ready_80) begin
        _dataflow_slice_valid_80 <= 0;
      end 
      if((_dataflow_slice_ready_80 || !_dataflow_slice_valid_80) && 1) begin
        _dataflow_slice_valid_80 <= _wvalid_404;
      end 
      if((_dataflow_slice_ready_83 || !_dataflow_slice_valid_83) && 1 && _wvalid_404) begin
        _dataflow_slice_data_83 <= _wdata_403[5'd15:5'd8];
      end 
      if(_dataflow_slice_valid_83 && _dataflow_slice_ready_83) begin
        _dataflow_slice_valid_83 <= 0;
      end 
      if((_dataflow_slice_ready_83 || !_dataflow_slice_valid_83) && 1) begin
        _dataflow_slice_valid_83 <= _wvalid_404;
      end 
      if((_dataflow_slice_ready_86 || !_dataflow_slice_valid_86) && 1 && _wvalid_404) begin
        _dataflow_slice_data_86 <= _wdata_403[6'd23:6'd16];
      end 
      if(_dataflow_slice_valid_86 && _dataflow_slice_ready_86) begin
        _dataflow_slice_valid_86 <= 0;
      end 
      if((_dataflow_slice_ready_86 || !_dataflow_slice_valid_86) && 1) begin
        _dataflow_slice_valid_86 <= _wvalid_404;
      end 
      if((_dataflow_slice_ready_89 || !_dataflow_slice_valid_89) && 1 && _wvalid_404) begin
        _dataflow_slice_data_89 <= _wdata_403[6'd31:6'd24];
      end 
      if(_dataflow_slice_valid_89 && _dataflow_slice_ready_89) begin
        _dataflow_slice_valid_89 <= 0;
      end 
      if((_dataflow_slice_ready_89 || !_dataflow_slice_valid_89) && 1) begin
        _dataflow_slice_valid_89 <= _wvalid_404;
      end 
      if((_dataflow_slice_ready_111 || !_dataflow_slice_valid_111) && 1 && _wvalid_1123) begin
        _dataflow_slice_data_111 <= _wdata_1122[4'd7:1'd0];
      end 
      if(_dataflow_slice_valid_111 && _dataflow_slice_ready_111) begin
        _dataflow_slice_valid_111 <= 0;
      end 
      if((_dataflow_slice_ready_111 || !_dataflow_slice_valid_111) && 1) begin
        _dataflow_slice_valid_111 <= _wvalid_1123;
      end 
      if((_dataflow_slice_ready_114 || !_dataflow_slice_valid_114) && 1 && _wvalid_1123) begin
        _dataflow_slice_data_114 <= _wdata_1122[5'd15:5'd8];
      end 
      if(_dataflow_slice_valid_114 && _dataflow_slice_ready_114) begin
        _dataflow_slice_valid_114 <= 0;
      end 
      if((_dataflow_slice_ready_114 || !_dataflow_slice_valid_114) && 1) begin
        _dataflow_slice_valid_114 <= _wvalid_1123;
      end 
      if((_dataflow_slice_ready_117 || !_dataflow_slice_valid_117) && 1 && _wvalid_1123) begin
        _dataflow_slice_data_117 <= _wdata_1122[6'd23:6'd16];
      end 
      if(_dataflow_slice_valid_117 && _dataflow_slice_ready_117) begin
        _dataflow_slice_valid_117 <= 0;
      end 
      if((_dataflow_slice_ready_117 || !_dataflow_slice_valid_117) && 1) begin
        _dataflow_slice_valid_117 <= _wvalid_1123;
      end 
      if((_dataflow_slice_ready_120 || !_dataflow_slice_valid_120) && 1 && _wvalid_1123) begin
        _dataflow_slice_data_120 <= _wdata_1122[6'd31:6'd24];
      end 
      if(_dataflow_slice_valid_120 && _dataflow_slice_ready_120) begin
        _dataflow_slice_valid_120 <= 0;
      end 
      if((_dataflow_slice_ready_120 || !_dataflow_slice_valid_120) && 1) begin
        _dataflow_slice_valid_120 <= _wvalid_1123;
      end 
      if((_dataflow_slice_ready_124 || !_dataflow_slice_valid_124) && 1 && _wvalid_1135) begin
        _dataflow_slice_data_124 <= _wdata_1134[3'd3:1'd0];
      end 
      if(_dataflow_slice_valid_124 && _dataflow_slice_ready_124) begin
        _dataflow_slice_valid_124 <= 0;
      end 
      if((_dataflow_slice_ready_124 || !_dataflow_slice_valid_124) && 1) begin
        _dataflow_slice_valid_124 <= _wvalid_1135;
      end 
      if((_dataflow_slice_ready_127 || !_dataflow_slice_valid_127) && 1 && _wvalid_1135) begin
        _dataflow_slice_data_127 <= _wdata_1134[4'd7:4'd4];
      end 
      if(_dataflow_slice_valid_127 && _dataflow_slice_ready_127) begin
        _dataflow_slice_valid_127 <= 0;
      end 
      if((_dataflow_slice_ready_127 || !_dataflow_slice_valid_127) && 1) begin
        _dataflow_slice_valid_127 <= _wvalid_1135;
      end 
      if((_dataflow_slice_ready_130 || !_dataflow_slice_valid_130) && 1 && _wvalid_1135) begin
        _dataflow_slice_data_130 <= _wdata_1134[5'd11:5'd8];
      end 
      if(_dataflow_slice_valid_130 && _dataflow_slice_ready_130) begin
        _dataflow_slice_valid_130 <= 0;
      end 
      if((_dataflow_slice_ready_130 || !_dataflow_slice_valid_130) && 1) begin
        _dataflow_slice_valid_130 <= _wvalid_1135;
      end 
      if((_dataflow_slice_ready_133 || !_dataflow_slice_valid_133) && 1 && _wvalid_1135) begin
        _dataflow_slice_data_133 <= _wdata_1134[5'd15:5'd12];
      end 
      if(_dataflow_slice_valid_133 && _dataflow_slice_ready_133) begin
        _dataflow_slice_valid_133 <= 0;
      end 
      if((_dataflow_slice_ready_133 || !_dataflow_slice_valid_133) && 1) begin
        _dataflow_slice_valid_133 <= _wvalid_1135;
      end 
      if((_dataflow_slice_ready_136 || !_dataflow_slice_valid_136) && 1 && _wvalid_1135) begin
        _dataflow_slice_data_136 <= _wdata_1134[6'd19:6'd16];
      end 
      if(_dataflow_slice_valid_136 && _dataflow_slice_ready_136) begin
        _dataflow_slice_valid_136 <= 0;
      end 
      if((_dataflow_slice_ready_136 || !_dataflow_slice_valid_136) && 1) begin
        _dataflow_slice_valid_136 <= _wvalid_1135;
      end 
      if((_dataflow_slice_ready_139 || !_dataflow_slice_valid_139) && 1 && _wvalid_1135) begin
        _dataflow_slice_data_139 <= _wdata_1134[6'd23:6'd20];
      end 
      if(_dataflow_slice_valid_139 && _dataflow_slice_ready_139) begin
        _dataflow_slice_valid_139 <= 0;
      end 
      if((_dataflow_slice_ready_139 || !_dataflow_slice_valid_139) && 1) begin
        _dataflow_slice_valid_139 <= _wvalid_1135;
      end 
      if((_dataflow_slice_ready_142 || !_dataflow_slice_valid_142) && 1 && _wvalid_1135) begin
        _dataflow_slice_data_142 <= _wdata_1134[6'd27:6'd24];
      end 
      if(_dataflow_slice_valid_142 && _dataflow_slice_ready_142) begin
        _dataflow_slice_valid_142 <= 0;
      end 
      if((_dataflow_slice_ready_142 || !_dataflow_slice_valid_142) && 1) begin
        _dataflow_slice_valid_142 <= _wvalid_1135;
      end 
      if((_dataflow_slice_ready_145 || !_dataflow_slice_valid_145) && 1 && _wvalid_1135) begin
        _dataflow_slice_data_145 <= _wdata_1134[6'd31:6'd28];
      end 
      if(_dataflow_slice_valid_145 && _dataflow_slice_ready_145) begin
        _dataflow_slice_valid_145 <= 0;
      end 
      if((_dataflow_slice_ready_145 || !_dataflow_slice_valid_145) && 1) begin
        _dataflow_slice_valid_145 <= _wvalid_1135;
      end 
      if((_dataflow_slice_ready_149 || !_dataflow_slice_valid_149) && 1 && _wvalid_1154) begin
        _dataflow_slice_data_149 <= _wdata_1153[4'd7:1'd0];
      end 
      if(_dataflow_slice_valid_149 && _dataflow_slice_ready_149) begin
        _dataflow_slice_valid_149 <= 0;
      end 
      if((_dataflow_slice_ready_149 || !_dataflow_slice_valid_149) && 1) begin
        _dataflow_slice_valid_149 <= _wvalid_1154;
      end 
      if((_dataflow_slice_ready_152 || !_dataflow_slice_valid_152) && 1 && _wvalid_1154) begin
        _dataflow_slice_data_152 <= _wdata_1153[5'd15:5'd8];
      end 
      if(_dataflow_slice_valid_152 && _dataflow_slice_ready_152) begin
        _dataflow_slice_valid_152 <= 0;
      end 
      if((_dataflow_slice_ready_152 || !_dataflow_slice_valid_152) && 1) begin
        _dataflow_slice_valid_152 <= _wvalid_1154;
      end 
      if((_dataflow_slice_ready_155 || !_dataflow_slice_valid_155) && 1 && _wvalid_1154) begin
        _dataflow_slice_data_155 <= _wdata_1153[6'd23:6'd16];
      end 
      if(_dataflow_slice_valid_155 && _dataflow_slice_ready_155) begin
        _dataflow_slice_valid_155 <= 0;
      end 
      if((_dataflow_slice_ready_155 || !_dataflow_slice_valid_155) && 1) begin
        _dataflow_slice_valid_155 <= _wvalid_1154;
      end 
      if((_dataflow_slice_ready_158 || !_dataflow_slice_valid_158) && 1 && _wvalid_1154) begin
        _dataflow_slice_data_158 <= _wdata_1153[6'd31:6'd24];
      end 
      if(_dataflow_slice_valid_158 && _dataflow_slice_ready_158) begin
        _dataflow_slice_valid_158 <= 0;
      end 
      if((_dataflow_slice_ready_158 || !_dataflow_slice_valid_158) && 1) begin
        _dataflow_slice_valid_158 <= _wvalid_1154;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      saxi_bvalid <= 0;
      _tmp_3 <= 0;
      _tmp_4 <= 0;
      _tmp_1 <= 0;
      _tmp_2 <= 0;
      _tmp_0 <= 0;
      saxi_rdata <= 0;
      saxi_rvalid <= 0;
      _saxi_cond_0_1 <= 0;
      _saxi_register_0 <= 0;
      _saxi_flag_0 <= 0;
      _saxi_register_1 <= 0;
      _saxi_flag_1 <= 0;
      _saxi_register_2 <= 0;
      _saxi_flag_2 <= 0;
      _saxi_register_3 <= 0;
      _saxi_flag_3 <= 0;
      _saxi_register_4 <= 0;
      _saxi_flag_4 <= 0;
      _saxi_register_5 <= 0;
      _saxi_flag_5 <= 0;
      _saxi_register_6 <= 0;
      _saxi_flag_6 <= 0;
      _saxi_register_7 <= 0;
      _saxi_flag_7 <= 0;
      _saxi_register_8 <= 0;
      _saxi_flag_8 <= 0;
      _saxi_register_9 <= 0;
      _saxi_flag_9 <= 0;
      _saxi_register_10 <= 165376;
      _saxi_flag_10 <= 0;
      _saxi_register_11 <= 0;
      _saxi_flag_11 <= 0;
      _saxi_register_12 <= 64;
      _saxi_flag_12 <= 0;
      _saxi_register_13 <= 4160;
      _saxi_flag_13 <= 0;
    end else begin
      if(_saxi_cond_0_1) begin
        saxi_rvalid <= 0;
      end 
      if(saxi_bvalid && saxi_bready) begin
        saxi_bvalid <= 0;
      end 
      if(saxi_wvalid && saxi_wready) begin
        saxi_bvalid <= 1;
      end 
      _tmp_3 <= saxi_awvalid;
      _tmp_4 <= saxi_arvalid;
      _tmp_1 <= 0;
      _tmp_2 <= 0;
      if(saxi_awready && saxi_awvalid && !saxi_bvalid) begin
        _tmp_0 <= saxi_awaddr;
        _tmp_1 <= 1;
      end else if(saxi_arready && saxi_arvalid) begin
        _tmp_0 <= saxi_araddr;
        _tmp_2 <= 1;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid)) begin
        saxi_rdata <= _tmp_6;
        saxi_rvalid <= 1;
      end 
      _saxi_cond_0_1 <= 1;
      if(saxi_rvalid && !saxi_rready) begin
        saxi_rvalid <= saxi_rvalid;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 0)) begin
        _saxi_register_0 <= _tmp_8;
        _saxi_flag_0 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 1)) begin
        _saxi_register_1 <= _tmp_8;
        _saxi_flag_1 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 2)) begin
        _saxi_register_2 <= _tmp_8;
        _saxi_flag_2 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 3)) begin
        _saxi_register_3 <= _tmp_8;
        _saxi_flag_3 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 4)) begin
        _saxi_register_4 <= _tmp_8;
        _saxi_flag_4 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 5)) begin
        _saxi_register_5 <= _tmp_8;
        _saxi_flag_5 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 6)) begin
        _saxi_register_6 <= _tmp_8;
        _saxi_flag_6 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 7)) begin
        _saxi_register_7 <= _tmp_8;
        _saxi_flag_7 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 8)) begin
        _saxi_register_8 <= _tmp_8;
        _saxi_flag_8 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 9)) begin
        _saxi_register_9 <= _tmp_8;
        _saxi_flag_9 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 10)) begin
        _saxi_register_10 <= _tmp_8;
        _saxi_flag_10 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 11)) begin
        _saxi_register_11 <= _tmp_8;
        _saxi_flag_11 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 12)) begin
        _saxi_register_12 <= _tmp_8;
        _saxi_flag_12 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && _tmp_7 && (_tmp_5 == 13)) begin
        _saxi_register_13 <= _tmp_8;
        _saxi_flag_13 <= 0;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 0)) begin
        _saxi_register_0 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 1)) begin
        _saxi_register_1 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 2)) begin
        _saxi_register_2 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 3)) begin
        _saxi_register_3 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 4)) begin
        _saxi_register_4 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 5)) begin
        _saxi_register_5 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 6)) begin
        _saxi_register_6 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 7)) begin
        _saxi_register_7 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 8)) begin
        _saxi_register_8 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 9)) begin
        _saxi_register_9 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 10)) begin
        _saxi_register_10 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 11)) begin
        _saxi_register_11 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 12)) begin
        _saxi_register_12 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && (saxi_wready && saxi_wvalid) && (_tmp_5 == 13)) begin
        _saxi_register_13 <= saxi_wdata;
      end 
      if(main_fsm == 0) begin
        _saxi_register_5 <= 0;
        _saxi_register_6 <= 0;
        _saxi_register_7 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_0 <= 1;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_1 <= 1;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_2 <= 1;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_3 <= 1;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_4 <= 1;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 1) && 1) begin
        _saxi_register_5 <= 1;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_6 <= 1;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_7 <= 1;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_8 <= 1;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_9 <= 1;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_10 <= 1;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_11 <= 1;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_12 <= 1;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_13 <= 1;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 2) && 1) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 89) && 1) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 89) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
    end
  end

  localparam _saxi_register_fsm_1 = 1;
  localparam _saxi_register_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _saxi_register_fsm <= _saxi_register_fsm_init;
    end else begin
      case(_saxi_register_fsm)
        _saxi_register_fsm_init: begin
          if(_tmp_2 || _tmp_1) begin
            _tmp_5 <= (_tmp_0 >> _saxi_shift) & _saxi_mask;
          end 
          if(_tmp_2) begin
            _saxi_register_fsm <= _saxi_register_fsm_1;
          end 
          if(_tmp_1) begin
            _saxi_register_fsm <= _saxi_register_fsm_2;
          end 
        end
        _saxi_register_fsm_1: begin
          if(saxi_rready || !saxi_rvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
        _saxi_register_fsm_2: begin
          _saxi_register_fsm <= _saxi_register_fsm_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    _rst_logic_1 <= rst_logic;
    _rst_logic_2 <= _rst_logic_1;
    RST <= rst_logic | _rst_logic_1 | _rst_logic_2;
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_68 <= 0;
      _tmp_38 <= 0;
      _tmp_39 <= 0;
      _tmp_41 <= 0;
      _tmp_42 <= 0;
      _tmp_43 <= 0;
      _tmp_44 <= 0;
      _tmp_45 <= 0;
      _tmp_46 <= 0;
      _tmp_47 <= 0;
      _tmp_48 <= 0;
      _tmp_49 <= 0;
      ram_w4_l8192_id0_0_1_addr <= 0;
      ram_w4_l8192_id0_0_1_wdata <= 0;
      ram_w4_l8192_id0_0_1_wenable <= 0;
      _tmp_40 <= 0;
      _ram_w4_l8192_id0_0_cond_0_1 <= 0;
      _ram_w4_l8192_id0_0_cond_1_1 <= 0;
      ram_w4_l8192_id0_0_0_addr <= 0;
      _ram_w4_l8192_id0_0_cond_2_1 <= 0;
      _tmp_586 <= 0;
      _ram_w4_l8192_id0_0_cond_3_1 <= 0;
      _ram_w4_l8192_id0_0_cond_3_2 <= 0;
      _tmp_1136 <= 0;
      _tmp_1137 <= 0;
      _ram_w4_l8192_id0_0_cond_4_1 <= 0;
      _ram_w4_l8192_id0_0_cond_5_1 <= 0;
      _tmp_1212 <= 0;
      _ram_w4_l8192_id0_0_cond_6_1 <= 0;
      _ram_w4_l8192_id0_0_cond_6_2 <= 0;
      ram_w4_l8192_id0_0_0_wdata <= 0;
      ram_w4_l8192_id0_0_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id0_0_cond_3_2) begin
        _tmp_586 <= 0;
      end 
      if(_ram_w4_l8192_id0_0_cond_6_2) begin
        _tmp_1212 <= 0;
      end 
      if(_ram_w4_l8192_id0_0_cond_0_1) begin
        _tmp_40 <= 0;
      end 
      if(_ram_w4_l8192_id0_0_cond_1_1) begin
        ram_w4_l8192_id0_0_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id0_0_cond_2_1) begin
        _tmp_586 <= 1;
      end 
      _ram_w4_l8192_id0_0_cond_3_2 <= _ram_w4_l8192_id0_0_cond_3_1;
      if(_ram_w4_l8192_id0_0_cond_4_1) begin
        ram_w4_l8192_id0_0_1_wenable <= 0;
        _tmp_1137 <= 0;
      end 
      if(_ram_w4_l8192_id0_0_cond_5_1) begin
        _tmp_1212 <= 1;
      end 
      _ram_w4_l8192_id0_0_cond_6_2 <= _ram_w4_l8192_id0_0_cond_6_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_39 == 0)) begin
        _tmp_68 <= 0;
        _tmp_38 <= req_block_size_33 - 1;
        _tmp_39 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_39 == 0)) begin
        _tmp_41 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_39 == 0)) begin
        _tmp_42 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_39 == 0)) begin
        _tmp_43 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_39 == 0)) begin
        _tmp_44 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_39 == 0)) begin
        _tmp_45 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_39 == 0)) begin
        _tmp_46 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_39 == 0)) begin
        _tmp_47 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_39 == 0)) begin
        _tmp_48 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_39 == 0)) begin
        _tmp_49 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0)) begin
        _tmp_38 <= _tmp_38 - 1;
        _tmp_39 <= _tmp_39 - 1;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0) && (_tmp_38 == 0)) begin
        _tmp_38 <= req_block_size_33 - 1;
        _tmp_68 <= _tmp_68 + 1;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0) && (_tmp_38 == 0) && (_tmp_68 == 8)) begin
        _tmp_68 <= 0;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0) && (_tmp_68 == 0)) begin
        _tmp_41 <= _tmp_50;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0) && (_tmp_68 == 1)) begin
        _tmp_42 <= _tmp_51;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0) && (_tmp_68 == 2)) begin
        _tmp_43 <= _tmp_52;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0) && (_tmp_68 == 3)) begin
        _tmp_44 <= _tmp_53;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0) && (_tmp_68 == 4)) begin
        _tmp_45 <= _tmp_54;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0) && (_tmp_68 == 5)) begin
        _tmp_46 <= _tmp_55;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0) && (_tmp_68 == 6)) begin
        _tmp_47 <= _tmp_56;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0) && (_tmp_68 == 7)) begin
        _tmp_48 <= _tmp_57;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0) && (_tmp_68 == 8)) begin
        _tmp_49 <= _tmp_58;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0)) begin
        ram_w4_l8192_id0_0_1_addr <= _tmp_59;
        ram_w4_l8192_id0_0_1_wdata <= _dataflow_slice_odata_29;
        ram_w4_l8192_id0_0_1_wenable <= _tmp_68 == 0;
      end 
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 == 1)) begin
        _tmp_40 <= 1;
      end 
      _ram_w4_l8192_id0_0_cond_0_1 <= 1;
      _ram_w4_l8192_id0_0_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12)) begin
        ram_w4_l8192_id0_0_0_addr <= _stream_conv2d_16_source_28_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_0_cond_2_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      _ram_w4_l8192_id0_0_cond_3_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      if(_maxi_read_start && (_maxi_read_op_sel == 8) && (_tmp_1136 == 0)) begin
        ram_w4_l8192_id0_0_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1136 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_124 && ((_tmp_1136 > 0) && !_tmp_1137) && (_tmp_1136 > 0)) begin
        ram_w4_l8192_id0_0_1_addr <= ram_w4_l8192_id0_0_1_addr + _maxi_read_local_stride;
        ram_w4_l8192_id0_0_1_wdata <= _dataflow_slice_odata_124;
        ram_w4_l8192_id0_0_1_wenable <= 1;
        _tmp_1136 <= _tmp_1136 - 1;
      end 
      if(_dataflow_slice_ovalid_124 && ((_tmp_1136 > 0) && !_tmp_1137) && (_tmp_1136 == 1)) begin
        _tmp_1137 <= 1;
      end 
      _ram_w4_l8192_id0_0_cond_4_1 <= 1;
      if(_stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4)) begin
        ram_w4_l8192_id0_0_0_addr <= _stream_matmul_29_source_20_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_0_cond_5_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      _ram_w4_l8192_id0_0_cond_6_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      ram_w4_l8192_id0_0_0_wdata <= 0;
      ram_w4_l8192_id0_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_99 <= 0;
      _tmp_69 <= 0;
      _tmp_70 <= 0;
      _tmp_72 <= 0;
      _tmp_73 <= 0;
      _tmp_74 <= 0;
      _tmp_75 <= 0;
      _tmp_76 <= 0;
      _tmp_77 <= 0;
      _tmp_78 <= 0;
      _tmp_79 <= 0;
      _tmp_80 <= 0;
      ram_w4_l8192_id0_1_1_addr <= 0;
      ram_w4_l8192_id0_1_1_wdata <= 0;
      ram_w4_l8192_id0_1_1_wenable <= 0;
      _tmp_71 <= 0;
      _ram_w4_l8192_id0_1_cond_0_1 <= 0;
      _ram_w4_l8192_id0_1_cond_1_1 <= 0;
      ram_w4_l8192_id0_1_0_addr <= 0;
      _ram_w4_l8192_id0_1_cond_2_1 <= 0;
      _tmp_587 <= 0;
      _ram_w4_l8192_id0_1_cond_3_1 <= 0;
      _ram_w4_l8192_id0_1_cond_3_2 <= 0;
      _tmp_1138 <= 0;
      _tmp_1139 <= 0;
      _ram_w4_l8192_id0_1_cond_4_1 <= 0;
      _ram_w4_l8192_id0_1_cond_5_1 <= 0;
      _tmp_1213 <= 0;
      _ram_w4_l8192_id0_1_cond_6_1 <= 0;
      _ram_w4_l8192_id0_1_cond_6_2 <= 0;
      ram_w4_l8192_id0_1_0_wdata <= 0;
      ram_w4_l8192_id0_1_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id0_1_cond_3_2) begin
        _tmp_587 <= 0;
      end 
      if(_ram_w4_l8192_id0_1_cond_6_2) begin
        _tmp_1213 <= 0;
      end 
      if(_ram_w4_l8192_id0_1_cond_0_1) begin
        _tmp_71 <= 0;
      end 
      if(_ram_w4_l8192_id0_1_cond_1_1) begin
        ram_w4_l8192_id0_1_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id0_1_cond_2_1) begin
        _tmp_587 <= 1;
      end 
      _ram_w4_l8192_id0_1_cond_3_2 <= _ram_w4_l8192_id0_1_cond_3_1;
      if(_ram_w4_l8192_id0_1_cond_4_1) begin
        ram_w4_l8192_id0_1_1_wenable <= 0;
        _tmp_1139 <= 0;
      end 
      if(_ram_w4_l8192_id0_1_cond_5_1) begin
        _tmp_1213 <= 1;
      end 
      _ram_w4_l8192_id0_1_cond_6_2 <= _ram_w4_l8192_id0_1_cond_6_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_70 == 0)) begin
        _tmp_99 <= 0;
        _tmp_69 <= req_block_size_33 - 1;
        _tmp_70 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_70 == 0)) begin
        _tmp_72 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_70 == 0)) begin
        _tmp_73 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_70 == 0)) begin
        _tmp_74 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_70 == 0)) begin
        _tmp_75 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_70 == 0)) begin
        _tmp_76 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_70 == 0)) begin
        _tmp_77 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_70 == 0)) begin
        _tmp_78 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_70 == 0)) begin
        _tmp_79 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_70 == 0)) begin
        _tmp_80 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0)) begin
        _tmp_69 <= _tmp_69 - 1;
        _tmp_70 <= _tmp_70 - 1;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0) && (_tmp_69 == 0)) begin
        _tmp_69 <= req_block_size_33 - 1;
        _tmp_99 <= _tmp_99 + 1;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0) && (_tmp_69 == 0) && (_tmp_99 == 8)) begin
        _tmp_99 <= 0;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0) && (_tmp_99 == 0)) begin
        _tmp_72 <= _tmp_81;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0) && (_tmp_99 == 1)) begin
        _tmp_73 <= _tmp_82;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0) && (_tmp_99 == 2)) begin
        _tmp_74 <= _tmp_83;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0) && (_tmp_99 == 3)) begin
        _tmp_75 <= _tmp_84;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0) && (_tmp_99 == 4)) begin
        _tmp_76 <= _tmp_85;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0) && (_tmp_99 == 5)) begin
        _tmp_77 <= _tmp_86;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0) && (_tmp_99 == 6)) begin
        _tmp_78 <= _tmp_87;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0) && (_tmp_99 == 7)) begin
        _tmp_79 <= _tmp_88;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0) && (_tmp_99 == 8)) begin
        _tmp_80 <= _tmp_89;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0)) begin
        ram_w4_l8192_id0_1_1_addr <= _tmp_90;
        ram_w4_l8192_id0_1_1_wdata <= _dataflow_slice_odata_32;
        ram_w4_l8192_id0_1_1_wenable <= _tmp_99 == 0;
      end 
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 == 1)) begin
        _tmp_71 <= 1;
      end 
      _ram_w4_l8192_id0_1_cond_0_1 <= 1;
      _ram_w4_l8192_id0_1_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12)) begin
        ram_w4_l8192_id0_1_0_addr <= _stream_conv2d_16_source_28_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_1_cond_2_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      _ram_w4_l8192_id0_1_cond_3_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      if(_maxi_read_start && (_maxi_read_op_sel == 8) && (_tmp_1138 == 0)) begin
        ram_w4_l8192_id0_1_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1138 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_127 && ((_tmp_1138 > 0) && !_tmp_1139) && (_tmp_1138 > 0)) begin
        ram_w4_l8192_id0_1_1_addr <= ram_w4_l8192_id0_1_1_addr + _maxi_read_local_stride;
        ram_w4_l8192_id0_1_1_wdata <= _dataflow_slice_odata_127;
        ram_w4_l8192_id0_1_1_wenable <= 1;
        _tmp_1138 <= _tmp_1138 - 1;
      end 
      if(_dataflow_slice_ovalid_127 && ((_tmp_1138 > 0) && !_tmp_1139) && (_tmp_1138 == 1)) begin
        _tmp_1139 <= 1;
      end 
      _ram_w4_l8192_id0_1_cond_4_1 <= 1;
      if(_stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4)) begin
        ram_w4_l8192_id0_1_0_addr <= _stream_matmul_29_source_20_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_1_cond_5_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      _ram_w4_l8192_id0_1_cond_6_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      ram_w4_l8192_id0_1_0_wdata <= 0;
      ram_w4_l8192_id0_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_130 <= 0;
      _tmp_100 <= 0;
      _tmp_101 <= 0;
      _tmp_103 <= 0;
      _tmp_104 <= 0;
      _tmp_105 <= 0;
      _tmp_106 <= 0;
      _tmp_107 <= 0;
      _tmp_108 <= 0;
      _tmp_109 <= 0;
      _tmp_110 <= 0;
      _tmp_111 <= 0;
      ram_w4_l8192_id0_2_1_addr <= 0;
      ram_w4_l8192_id0_2_1_wdata <= 0;
      ram_w4_l8192_id0_2_1_wenable <= 0;
      _tmp_102 <= 0;
      _ram_w4_l8192_id0_2_cond_0_1 <= 0;
      _ram_w4_l8192_id0_2_cond_1_1 <= 0;
      ram_w4_l8192_id0_2_0_addr <= 0;
      _ram_w4_l8192_id0_2_cond_2_1 <= 0;
      _tmp_588 <= 0;
      _ram_w4_l8192_id0_2_cond_3_1 <= 0;
      _ram_w4_l8192_id0_2_cond_3_2 <= 0;
      _tmp_1140 <= 0;
      _tmp_1141 <= 0;
      _ram_w4_l8192_id0_2_cond_4_1 <= 0;
      _ram_w4_l8192_id0_2_cond_5_1 <= 0;
      _tmp_1214 <= 0;
      _ram_w4_l8192_id0_2_cond_6_1 <= 0;
      _ram_w4_l8192_id0_2_cond_6_2 <= 0;
      ram_w4_l8192_id0_2_0_wdata <= 0;
      ram_w4_l8192_id0_2_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id0_2_cond_3_2) begin
        _tmp_588 <= 0;
      end 
      if(_ram_w4_l8192_id0_2_cond_6_2) begin
        _tmp_1214 <= 0;
      end 
      if(_ram_w4_l8192_id0_2_cond_0_1) begin
        _tmp_102 <= 0;
      end 
      if(_ram_w4_l8192_id0_2_cond_1_1) begin
        ram_w4_l8192_id0_2_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id0_2_cond_2_1) begin
        _tmp_588 <= 1;
      end 
      _ram_w4_l8192_id0_2_cond_3_2 <= _ram_w4_l8192_id0_2_cond_3_1;
      if(_ram_w4_l8192_id0_2_cond_4_1) begin
        ram_w4_l8192_id0_2_1_wenable <= 0;
        _tmp_1141 <= 0;
      end 
      if(_ram_w4_l8192_id0_2_cond_5_1) begin
        _tmp_1214 <= 1;
      end 
      _ram_w4_l8192_id0_2_cond_6_2 <= _ram_w4_l8192_id0_2_cond_6_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_101 == 0)) begin
        _tmp_130 <= 0;
        _tmp_100 <= req_block_size_33 - 1;
        _tmp_101 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_101 == 0)) begin
        _tmp_103 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_101 == 0)) begin
        _tmp_104 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_101 == 0)) begin
        _tmp_105 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_101 == 0)) begin
        _tmp_106 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_101 == 0)) begin
        _tmp_107 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_101 == 0)) begin
        _tmp_108 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_101 == 0)) begin
        _tmp_109 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_101 == 0)) begin
        _tmp_110 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_101 == 0)) begin
        _tmp_111 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0)) begin
        _tmp_100 <= _tmp_100 - 1;
        _tmp_101 <= _tmp_101 - 1;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0) && (_tmp_100 == 0)) begin
        _tmp_100 <= req_block_size_33 - 1;
        _tmp_130 <= _tmp_130 + 1;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0) && (_tmp_100 == 0) && (_tmp_130 == 8)) begin
        _tmp_130 <= 0;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0) && (_tmp_130 == 0)) begin
        _tmp_103 <= _tmp_112;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0) && (_tmp_130 == 1)) begin
        _tmp_104 <= _tmp_113;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0) && (_tmp_130 == 2)) begin
        _tmp_105 <= _tmp_114;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0) && (_tmp_130 == 3)) begin
        _tmp_106 <= _tmp_115;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0) && (_tmp_130 == 4)) begin
        _tmp_107 <= _tmp_116;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0) && (_tmp_130 == 5)) begin
        _tmp_108 <= _tmp_117;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0) && (_tmp_130 == 6)) begin
        _tmp_109 <= _tmp_118;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0) && (_tmp_130 == 7)) begin
        _tmp_110 <= _tmp_119;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0) && (_tmp_130 == 8)) begin
        _tmp_111 <= _tmp_120;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0)) begin
        ram_w4_l8192_id0_2_1_addr <= _tmp_121;
        ram_w4_l8192_id0_2_1_wdata <= _dataflow_slice_odata_35;
        ram_w4_l8192_id0_2_1_wenable <= _tmp_130 == 0;
      end 
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 == 1)) begin
        _tmp_102 <= 1;
      end 
      _ram_w4_l8192_id0_2_cond_0_1 <= 1;
      _ram_w4_l8192_id0_2_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12)) begin
        ram_w4_l8192_id0_2_0_addr <= _stream_conv2d_16_source_28_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_2_cond_2_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      _ram_w4_l8192_id0_2_cond_3_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      if(_maxi_read_start && (_maxi_read_op_sel == 8) && (_tmp_1140 == 0)) begin
        ram_w4_l8192_id0_2_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1140 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_130 && ((_tmp_1140 > 0) && !_tmp_1141) && (_tmp_1140 > 0)) begin
        ram_w4_l8192_id0_2_1_addr <= ram_w4_l8192_id0_2_1_addr + _maxi_read_local_stride;
        ram_w4_l8192_id0_2_1_wdata <= _dataflow_slice_odata_130;
        ram_w4_l8192_id0_2_1_wenable <= 1;
        _tmp_1140 <= _tmp_1140 - 1;
      end 
      if(_dataflow_slice_ovalid_130 && ((_tmp_1140 > 0) && !_tmp_1141) && (_tmp_1140 == 1)) begin
        _tmp_1141 <= 1;
      end 
      _ram_w4_l8192_id0_2_cond_4_1 <= 1;
      if(_stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4)) begin
        ram_w4_l8192_id0_2_0_addr <= _stream_matmul_29_source_20_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_2_cond_5_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      _ram_w4_l8192_id0_2_cond_6_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      ram_w4_l8192_id0_2_0_wdata <= 0;
      ram_w4_l8192_id0_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_161 <= 0;
      _tmp_131 <= 0;
      _tmp_132 <= 0;
      _tmp_134 <= 0;
      _tmp_135 <= 0;
      _tmp_136 <= 0;
      _tmp_137 <= 0;
      _tmp_138 <= 0;
      _tmp_139 <= 0;
      _tmp_140 <= 0;
      _tmp_141 <= 0;
      _tmp_142 <= 0;
      ram_w4_l8192_id0_3_1_addr <= 0;
      ram_w4_l8192_id0_3_1_wdata <= 0;
      ram_w4_l8192_id0_3_1_wenable <= 0;
      _tmp_133 <= 0;
      _ram_w4_l8192_id0_3_cond_0_1 <= 0;
      _ram_w4_l8192_id0_3_cond_1_1 <= 0;
      ram_w4_l8192_id0_3_0_addr <= 0;
      _ram_w4_l8192_id0_3_cond_2_1 <= 0;
      _tmp_589 <= 0;
      _ram_w4_l8192_id0_3_cond_3_1 <= 0;
      _ram_w4_l8192_id0_3_cond_3_2 <= 0;
      _tmp_1142 <= 0;
      _tmp_1143 <= 0;
      _ram_w4_l8192_id0_3_cond_4_1 <= 0;
      _ram_w4_l8192_id0_3_cond_5_1 <= 0;
      _tmp_1215 <= 0;
      _ram_w4_l8192_id0_3_cond_6_1 <= 0;
      _ram_w4_l8192_id0_3_cond_6_2 <= 0;
      ram_w4_l8192_id0_3_0_wdata <= 0;
      ram_w4_l8192_id0_3_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id0_3_cond_3_2) begin
        _tmp_589 <= 0;
      end 
      if(_ram_w4_l8192_id0_3_cond_6_2) begin
        _tmp_1215 <= 0;
      end 
      if(_ram_w4_l8192_id0_3_cond_0_1) begin
        _tmp_133 <= 0;
      end 
      if(_ram_w4_l8192_id0_3_cond_1_1) begin
        ram_w4_l8192_id0_3_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id0_3_cond_2_1) begin
        _tmp_589 <= 1;
      end 
      _ram_w4_l8192_id0_3_cond_3_2 <= _ram_w4_l8192_id0_3_cond_3_1;
      if(_ram_w4_l8192_id0_3_cond_4_1) begin
        ram_w4_l8192_id0_3_1_wenable <= 0;
        _tmp_1143 <= 0;
      end 
      if(_ram_w4_l8192_id0_3_cond_5_1) begin
        _tmp_1215 <= 1;
      end 
      _ram_w4_l8192_id0_3_cond_6_2 <= _ram_w4_l8192_id0_3_cond_6_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_132 == 0)) begin
        _tmp_161 <= 0;
        _tmp_131 <= req_block_size_33 - 1;
        _tmp_132 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_132 == 0)) begin
        _tmp_134 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_132 == 0)) begin
        _tmp_135 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_132 == 0)) begin
        _tmp_136 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_132 == 0)) begin
        _tmp_137 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_132 == 0)) begin
        _tmp_138 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_132 == 0)) begin
        _tmp_139 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_132 == 0)) begin
        _tmp_140 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_132 == 0)) begin
        _tmp_141 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_132 == 0)) begin
        _tmp_142 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0)) begin
        _tmp_131 <= _tmp_131 - 1;
        _tmp_132 <= _tmp_132 - 1;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0) && (_tmp_131 == 0)) begin
        _tmp_131 <= req_block_size_33 - 1;
        _tmp_161 <= _tmp_161 + 1;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0) && (_tmp_131 == 0) && (_tmp_161 == 8)) begin
        _tmp_161 <= 0;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0) && (_tmp_161 == 0)) begin
        _tmp_134 <= _tmp_143;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0) && (_tmp_161 == 1)) begin
        _tmp_135 <= _tmp_144;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0) && (_tmp_161 == 2)) begin
        _tmp_136 <= _tmp_145;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0) && (_tmp_161 == 3)) begin
        _tmp_137 <= _tmp_146;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0) && (_tmp_161 == 4)) begin
        _tmp_138 <= _tmp_147;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0) && (_tmp_161 == 5)) begin
        _tmp_139 <= _tmp_148;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0) && (_tmp_161 == 6)) begin
        _tmp_140 <= _tmp_149;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0) && (_tmp_161 == 7)) begin
        _tmp_141 <= _tmp_150;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0) && (_tmp_161 == 8)) begin
        _tmp_142 <= _tmp_151;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0)) begin
        ram_w4_l8192_id0_3_1_addr <= _tmp_152;
        ram_w4_l8192_id0_3_1_wdata <= _dataflow_slice_odata_38;
        ram_w4_l8192_id0_3_1_wenable <= _tmp_161 == 0;
      end 
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 == 1)) begin
        _tmp_133 <= 1;
      end 
      _ram_w4_l8192_id0_3_cond_0_1 <= 1;
      _ram_w4_l8192_id0_3_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12)) begin
        ram_w4_l8192_id0_3_0_addr <= _stream_conv2d_16_source_28_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_3_cond_2_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      _ram_w4_l8192_id0_3_cond_3_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      if(_maxi_read_start && (_maxi_read_op_sel == 8) && (_tmp_1142 == 0)) begin
        ram_w4_l8192_id0_3_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1142 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_133 && ((_tmp_1142 > 0) && !_tmp_1143) && (_tmp_1142 > 0)) begin
        ram_w4_l8192_id0_3_1_addr <= ram_w4_l8192_id0_3_1_addr + _maxi_read_local_stride;
        ram_w4_l8192_id0_3_1_wdata <= _dataflow_slice_odata_133;
        ram_w4_l8192_id0_3_1_wenable <= 1;
        _tmp_1142 <= _tmp_1142 - 1;
      end 
      if(_dataflow_slice_ovalid_133 && ((_tmp_1142 > 0) && !_tmp_1143) && (_tmp_1142 == 1)) begin
        _tmp_1143 <= 1;
      end 
      _ram_w4_l8192_id0_3_cond_4_1 <= 1;
      if(_stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4)) begin
        ram_w4_l8192_id0_3_0_addr <= _stream_matmul_29_source_20_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_3_cond_5_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      _ram_w4_l8192_id0_3_cond_6_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      ram_w4_l8192_id0_3_0_wdata <= 0;
      ram_w4_l8192_id0_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_192 <= 0;
      _tmp_162 <= 0;
      _tmp_163 <= 0;
      _tmp_165 <= 0;
      _tmp_166 <= 0;
      _tmp_167 <= 0;
      _tmp_168 <= 0;
      _tmp_169 <= 0;
      _tmp_170 <= 0;
      _tmp_171 <= 0;
      _tmp_172 <= 0;
      _tmp_173 <= 0;
      ram_w4_l8192_id0_4_1_addr <= 0;
      ram_w4_l8192_id0_4_1_wdata <= 0;
      ram_w4_l8192_id0_4_1_wenable <= 0;
      _tmp_164 <= 0;
      _ram_w4_l8192_id0_4_cond_0_1 <= 0;
      _ram_w4_l8192_id0_4_cond_1_1 <= 0;
      ram_w4_l8192_id0_4_0_addr <= 0;
      _ram_w4_l8192_id0_4_cond_2_1 <= 0;
      _tmp_590 <= 0;
      _ram_w4_l8192_id0_4_cond_3_1 <= 0;
      _ram_w4_l8192_id0_4_cond_3_2 <= 0;
      _tmp_1144 <= 0;
      _tmp_1145 <= 0;
      _ram_w4_l8192_id0_4_cond_4_1 <= 0;
      _ram_w4_l8192_id0_4_cond_5_1 <= 0;
      _tmp_1216 <= 0;
      _ram_w4_l8192_id0_4_cond_6_1 <= 0;
      _ram_w4_l8192_id0_4_cond_6_2 <= 0;
      ram_w4_l8192_id0_4_0_wdata <= 0;
      ram_w4_l8192_id0_4_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id0_4_cond_3_2) begin
        _tmp_590 <= 0;
      end 
      if(_ram_w4_l8192_id0_4_cond_6_2) begin
        _tmp_1216 <= 0;
      end 
      if(_ram_w4_l8192_id0_4_cond_0_1) begin
        _tmp_164 <= 0;
      end 
      if(_ram_w4_l8192_id0_4_cond_1_1) begin
        ram_w4_l8192_id0_4_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id0_4_cond_2_1) begin
        _tmp_590 <= 1;
      end 
      _ram_w4_l8192_id0_4_cond_3_2 <= _ram_w4_l8192_id0_4_cond_3_1;
      if(_ram_w4_l8192_id0_4_cond_4_1) begin
        ram_w4_l8192_id0_4_1_wenable <= 0;
        _tmp_1145 <= 0;
      end 
      if(_ram_w4_l8192_id0_4_cond_5_1) begin
        _tmp_1216 <= 1;
      end 
      _ram_w4_l8192_id0_4_cond_6_2 <= _ram_w4_l8192_id0_4_cond_6_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_163 == 0)) begin
        _tmp_192 <= 0;
        _tmp_162 <= req_block_size_33 - 1;
        _tmp_163 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_163 == 0)) begin
        _tmp_165 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_163 == 0)) begin
        _tmp_166 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_163 == 0)) begin
        _tmp_167 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_163 == 0)) begin
        _tmp_168 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_163 == 0)) begin
        _tmp_169 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_163 == 0)) begin
        _tmp_170 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_163 == 0)) begin
        _tmp_171 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_163 == 0)) begin
        _tmp_172 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_163 == 0)) begin
        _tmp_173 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0)) begin
        _tmp_162 <= _tmp_162 - 1;
        _tmp_163 <= _tmp_163 - 1;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0) && (_tmp_162 == 0)) begin
        _tmp_162 <= req_block_size_33 - 1;
        _tmp_192 <= _tmp_192 + 1;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0) && (_tmp_162 == 0) && (_tmp_192 == 8)) begin
        _tmp_192 <= 0;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0) && (_tmp_192 == 0)) begin
        _tmp_165 <= _tmp_174;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0) && (_tmp_192 == 1)) begin
        _tmp_166 <= _tmp_175;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0) && (_tmp_192 == 2)) begin
        _tmp_167 <= _tmp_176;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0) && (_tmp_192 == 3)) begin
        _tmp_168 <= _tmp_177;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0) && (_tmp_192 == 4)) begin
        _tmp_169 <= _tmp_178;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0) && (_tmp_192 == 5)) begin
        _tmp_170 <= _tmp_179;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0) && (_tmp_192 == 6)) begin
        _tmp_171 <= _tmp_180;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0) && (_tmp_192 == 7)) begin
        _tmp_172 <= _tmp_181;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0) && (_tmp_192 == 8)) begin
        _tmp_173 <= _tmp_182;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0)) begin
        ram_w4_l8192_id0_4_1_addr <= _tmp_183;
        ram_w4_l8192_id0_4_1_wdata <= _dataflow_slice_odata_41;
        ram_w4_l8192_id0_4_1_wenable <= _tmp_192 == 0;
      end 
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 == 1)) begin
        _tmp_164 <= 1;
      end 
      _ram_w4_l8192_id0_4_cond_0_1 <= 1;
      _ram_w4_l8192_id0_4_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12)) begin
        ram_w4_l8192_id0_4_0_addr <= _stream_conv2d_16_source_28_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_4_cond_2_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      _ram_w4_l8192_id0_4_cond_3_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      if(_maxi_read_start && (_maxi_read_op_sel == 8) && (_tmp_1144 == 0)) begin
        ram_w4_l8192_id0_4_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1144 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_136 && ((_tmp_1144 > 0) && !_tmp_1145) && (_tmp_1144 > 0)) begin
        ram_w4_l8192_id0_4_1_addr <= ram_w4_l8192_id0_4_1_addr + _maxi_read_local_stride;
        ram_w4_l8192_id0_4_1_wdata <= _dataflow_slice_odata_136;
        ram_w4_l8192_id0_4_1_wenable <= 1;
        _tmp_1144 <= _tmp_1144 - 1;
      end 
      if(_dataflow_slice_ovalid_136 && ((_tmp_1144 > 0) && !_tmp_1145) && (_tmp_1144 == 1)) begin
        _tmp_1145 <= 1;
      end 
      _ram_w4_l8192_id0_4_cond_4_1 <= 1;
      if(_stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4)) begin
        ram_w4_l8192_id0_4_0_addr <= _stream_matmul_29_source_20_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_4_cond_5_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      _ram_w4_l8192_id0_4_cond_6_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      ram_w4_l8192_id0_4_0_wdata <= 0;
      ram_w4_l8192_id0_4_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_223 <= 0;
      _tmp_193 <= 0;
      _tmp_194 <= 0;
      _tmp_196 <= 0;
      _tmp_197 <= 0;
      _tmp_198 <= 0;
      _tmp_199 <= 0;
      _tmp_200 <= 0;
      _tmp_201 <= 0;
      _tmp_202 <= 0;
      _tmp_203 <= 0;
      _tmp_204 <= 0;
      ram_w4_l8192_id0_5_1_addr <= 0;
      ram_w4_l8192_id0_5_1_wdata <= 0;
      ram_w4_l8192_id0_5_1_wenable <= 0;
      _tmp_195 <= 0;
      _ram_w4_l8192_id0_5_cond_0_1 <= 0;
      _ram_w4_l8192_id0_5_cond_1_1 <= 0;
      ram_w4_l8192_id0_5_0_addr <= 0;
      _ram_w4_l8192_id0_5_cond_2_1 <= 0;
      _tmp_591 <= 0;
      _ram_w4_l8192_id0_5_cond_3_1 <= 0;
      _ram_w4_l8192_id0_5_cond_3_2 <= 0;
      _tmp_1146 <= 0;
      _tmp_1147 <= 0;
      _ram_w4_l8192_id0_5_cond_4_1 <= 0;
      _ram_w4_l8192_id0_5_cond_5_1 <= 0;
      _tmp_1217 <= 0;
      _ram_w4_l8192_id0_5_cond_6_1 <= 0;
      _ram_w4_l8192_id0_5_cond_6_2 <= 0;
      ram_w4_l8192_id0_5_0_wdata <= 0;
      ram_w4_l8192_id0_5_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id0_5_cond_3_2) begin
        _tmp_591 <= 0;
      end 
      if(_ram_w4_l8192_id0_5_cond_6_2) begin
        _tmp_1217 <= 0;
      end 
      if(_ram_w4_l8192_id0_5_cond_0_1) begin
        _tmp_195 <= 0;
      end 
      if(_ram_w4_l8192_id0_5_cond_1_1) begin
        ram_w4_l8192_id0_5_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id0_5_cond_2_1) begin
        _tmp_591 <= 1;
      end 
      _ram_w4_l8192_id0_5_cond_3_2 <= _ram_w4_l8192_id0_5_cond_3_1;
      if(_ram_w4_l8192_id0_5_cond_4_1) begin
        ram_w4_l8192_id0_5_1_wenable <= 0;
        _tmp_1147 <= 0;
      end 
      if(_ram_w4_l8192_id0_5_cond_5_1) begin
        _tmp_1217 <= 1;
      end 
      _ram_w4_l8192_id0_5_cond_6_2 <= _ram_w4_l8192_id0_5_cond_6_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_194 == 0)) begin
        _tmp_223 <= 0;
        _tmp_193 <= req_block_size_33 - 1;
        _tmp_194 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_194 == 0)) begin
        _tmp_196 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_194 == 0)) begin
        _tmp_197 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_194 == 0)) begin
        _tmp_198 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_194 == 0)) begin
        _tmp_199 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_194 == 0)) begin
        _tmp_200 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_194 == 0)) begin
        _tmp_201 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_194 == 0)) begin
        _tmp_202 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_194 == 0)) begin
        _tmp_203 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_194 == 0)) begin
        _tmp_204 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0)) begin
        _tmp_193 <= _tmp_193 - 1;
        _tmp_194 <= _tmp_194 - 1;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0) && (_tmp_193 == 0)) begin
        _tmp_193 <= req_block_size_33 - 1;
        _tmp_223 <= _tmp_223 + 1;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0) && (_tmp_193 == 0) && (_tmp_223 == 8)) begin
        _tmp_223 <= 0;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0) && (_tmp_223 == 0)) begin
        _tmp_196 <= _tmp_205;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0) && (_tmp_223 == 1)) begin
        _tmp_197 <= _tmp_206;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0) && (_tmp_223 == 2)) begin
        _tmp_198 <= _tmp_207;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0) && (_tmp_223 == 3)) begin
        _tmp_199 <= _tmp_208;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0) && (_tmp_223 == 4)) begin
        _tmp_200 <= _tmp_209;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0) && (_tmp_223 == 5)) begin
        _tmp_201 <= _tmp_210;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0) && (_tmp_223 == 6)) begin
        _tmp_202 <= _tmp_211;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0) && (_tmp_223 == 7)) begin
        _tmp_203 <= _tmp_212;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0) && (_tmp_223 == 8)) begin
        _tmp_204 <= _tmp_213;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0)) begin
        ram_w4_l8192_id0_5_1_addr <= _tmp_214;
        ram_w4_l8192_id0_5_1_wdata <= _dataflow_slice_odata_44;
        ram_w4_l8192_id0_5_1_wenable <= _tmp_223 == 0;
      end 
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 == 1)) begin
        _tmp_195 <= 1;
      end 
      _ram_w4_l8192_id0_5_cond_0_1 <= 1;
      _ram_w4_l8192_id0_5_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12)) begin
        ram_w4_l8192_id0_5_0_addr <= _stream_conv2d_16_source_28_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_5_cond_2_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      _ram_w4_l8192_id0_5_cond_3_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      if(_maxi_read_start && (_maxi_read_op_sel == 8) && (_tmp_1146 == 0)) begin
        ram_w4_l8192_id0_5_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1146 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_139 && ((_tmp_1146 > 0) && !_tmp_1147) && (_tmp_1146 > 0)) begin
        ram_w4_l8192_id0_5_1_addr <= ram_w4_l8192_id0_5_1_addr + _maxi_read_local_stride;
        ram_w4_l8192_id0_5_1_wdata <= _dataflow_slice_odata_139;
        ram_w4_l8192_id0_5_1_wenable <= 1;
        _tmp_1146 <= _tmp_1146 - 1;
      end 
      if(_dataflow_slice_ovalid_139 && ((_tmp_1146 > 0) && !_tmp_1147) && (_tmp_1146 == 1)) begin
        _tmp_1147 <= 1;
      end 
      _ram_w4_l8192_id0_5_cond_4_1 <= 1;
      if(_stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4)) begin
        ram_w4_l8192_id0_5_0_addr <= _stream_matmul_29_source_20_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_5_cond_5_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      _ram_w4_l8192_id0_5_cond_6_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      ram_w4_l8192_id0_5_0_wdata <= 0;
      ram_w4_l8192_id0_5_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_254 <= 0;
      _tmp_224 <= 0;
      _tmp_225 <= 0;
      _tmp_227 <= 0;
      _tmp_228 <= 0;
      _tmp_229 <= 0;
      _tmp_230 <= 0;
      _tmp_231 <= 0;
      _tmp_232 <= 0;
      _tmp_233 <= 0;
      _tmp_234 <= 0;
      _tmp_235 <= 0;
      ram_w4_l8192_id0_6_1_addr <= 0;
      ram_w4_l8192_id0_6_1_wdata <= 0;
      ram_w4_l8192_id0_6_1_wenable <= 0;
      _tmp_226 <= 0;
      _ram_w4_l8192_id0_6_cond_0_1 <= 0;
      _ram_w4_l8192_id0_6_cond_1_1 <= 0;
      ram_w4_l8192_id0_6_0_addr <= 0;
      _ram_w4_l8192_id0_6_cond_2_1 <= 0;
      _tmp_592 <= 0;
      _ram_w4_l8192_id0_6_cond_3_1 <= 0;
      _ram_w4_l8192_id0_6_cond_3_2 <= 0;
      _tmp_1148 <= 0;
      _tmp_1149 <= 0;
      _ram_w4_l8192_id0_6_cond_4_1 <= 0;
      _ram_w4_l8192_id0_6_cond_5_1 <= 0;
      _tmp_1218 <= 0;
      _ram_w4_l8192_id0_6_cond_6_1 <= 0;
      _ram_w4_l8192_id0_6_cond_6_2 <= 0;
      ram_w4_l8192_id0_6_0_wdata <= 0;
      ram_w4_l8192_id0_6_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id0_6_cond_3_2) begin
        _tmp_592 <= 0;
      end 
      if(_ram_w4_l8192_id0_6_cond_6_2) begin
        _tmp_1218 <= 0;
      end 
      if(_ram_w4_l8192_id0_6_cond_0_1) begin
        _tmp_226 <= 0;
      end 
      if(_ram_w4_l8192_id0_6_cond_1_1) begin
        ram_w4_l8192_id0_6_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id0_6_cond_2_1) begin
        _tmp_592 <= 1;
      end 
      _ram_w4_l8192_id0_6_cond_3_2 <= _ram_w4_l8192_id0_6_cond_3_1;
      if(_ram_w4_l8192_id0_6_cond_4_1) begin
        ram_w4_l8192_id0_6_1_wenable <= 0;
        _tmp_1149 <= 0;
      end 
      if(_ram_w4_l8192_id0_6_cond_5_1) begin
        _tmp_1218 <= 1;
      end 
      _ram_w4_l8192_id0_6_cond_6_2 <= _ram_w4_l8192_id0_6_cond_6_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_225 == 0)) begin
        _tmp_254 <= 0;
        _tmp_224 <= req_block_size_33 - 1;
        _tmp_225 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_225 == 0)) begin
        _tmp_227 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_225 == 0)) begin
        _tmp_228 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_225 == 0)) begin
        _tmp_229 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_225 == 0)) begin
        _tmp_230 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_225 == 0)) begin
        _tmp_231 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_225 == 0)) begin
        _tmp_232 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_225 == 0)) begin
        _tmp_233 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_225 == 0)) begin
        _tmp_234 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_225 == 0)) begin
        _tmp_235 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0)) begin
        _tmp_224 <= _tmp_224 - 1;
        _tmp_225 <= _tmp_225 - 1;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0) && (_tmp_224 == 0)) begin
        _tmp_224 <= req_block_size_33 - 1;
        _tmp_254 <= _tmp_254 + 1;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0) && (_tmp_224 == 0) && (_tmp_254 == 8)) begin
        _tmp_254 <= 0;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0) && (_tmp_254 == 0)) begin
        _tmp_227 <= _tmp_236;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0) && (_tmp_254 == 1)) begin
        _tmp_228 <= _tmp_237;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0) && (_tmp_254 == 2)) begin
        _tmp_229 <= _tmp_238;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0) && (_tmp_254 == 3)) begin
        _tmp_230 <= _tmp_239;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0) && (_tmp_254 == 4)) begin
        _tmp_231 <= _tmp_240;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0) && (_tmp_254 == 5)) begin
        _tmp_232 <= _tmp_241;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0) && (_tmp_254 == 6)) begin
        _tmp_233 <= _tmp_242;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0) && (_tmp_254 == 7)) begin
        _tmp_234 <= _tmp_243;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0) && (_tmp_254 == 8)) begin
        _tmp_235 <= _tmp_244;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0)) begin
        ram_w4_l8192_id0_6_1_addr <= _tmp_245;
        ram_w4_l8192_id0_6_1_wdata <= _dataflow_slice_odata_47;
        ram_w4_l8192_id0_6_1_wenable <= _tmp_254 == 0;
      end 
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 == 1)) begin
        _tmp_226 <= 1;
      end 
      _ram_w4_l8192_id0_6_cond_0_1 <= 1;
      _ram_w4_l8192_id0_6_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12)) begin
        ram_w4_l8192_id0_6_0_addr <= _stream_conv2d_16_source_28_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_6_cond_2_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      _ram_w4_l8192_id0_6_cond_3_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      if(_maxi_read_start && (_maxi_read_op_sel == 8) && (_tmp_1148 == 0)) begin
        ram_w4_l8192_id0_6_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1148 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_142 && ((_tmp_1148 > 0) && !_tmp_1149) && (_tmp_1148 > 0)) begin
        ram_w4_l8192_id0_6_1_addr <= ram_w4_l8192_id0_6_1_addr + _maxi_read_local_stride;
        ram_w4_l8192_id0_6_1_wdata <= _dataflow_slice_odata_142;
        ram_w4_l8192_id0_6_1_wenable <= 1;
        _tmp_1148 <= _tmp_1148 - 1;
      end 
      if(_dataflow_slice_ovalid_142 && ((_tmp_1148 > 0) && !_tmp_1149) && (_tmp_1148 == 1)) begin
        _tmp_1149 <= 1;
      end 
      _ram_w4_l8192_id0_6_cond_4_1 <= 1;
      if(_stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4)) begin
        ram_w4_l8192_id0_6_0_addr <= _stream_matmul_29_source_20_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_6_cond_5_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      _ram_w4_l8192_id0_6_cond_6_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      ram_w4_l8192_id0_6_0_wdata <= 0;
      ram_w4_l8192_id0_6_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_285 <= 0;
      _tmp_255 <= 0;
      _tmp_256 <= 0;
      _tmp_258 <= 0;
      _tmp_259 <= 0;
      _tmp_260 <= 0;
      _tmp_261 <= 0;
      _tmp_262 <= 0;
      _tmp_263 <= 0;
      _tmp_264 <= 0;
      _tmp_265 <= 0;
      _tmp_266 <= 0;
      ram_w4_l8192_id0_7_1_addr <= 0;
      ram_w4_l8192_id0_7_1_wdata <= 0;
      ram_w4_l8192_id0_7_1_wenable <= 0;
      _tmp_257 <= 0;
      _ram_w4_l8192_id0_7_cond_0_1 <= 0;
      _ram_w4_l8192_id0_7_cond_1_1 <= 0;
      ram_w4_l8192_id0_7_0_addr <= 0;
      _ram_w4_l8192_id0_7_cond_2_1 <= 0;
      _tmp_593 <= 0;
      _ram_w4_l8192_id0_7_cond_3_1 <= 0;
      _ram_w4_l8192_id0_7_cond_3_2 <= 0;
      _tmp_1150 <= 0;
      _tmp_1151 <= 0;
      _ram_w4_l8192_id0_7_cond_4_1 <= 0;
      _ram_w4_l8192_id0_7_cond_5_1 <= 0;
      _tmp_1219 <= 0;
      _ram_w4_l8192_id0_7_cond_6_1 <= 0;
      _ram_w4_l8192_id0_7_cond_6_2 <= 0;
      ram_w4_l8192_id0_7_0_wdata <= 0;
      ram_w4_l8192_id0_7_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id0_7_cond_3_2) begin
        _tmp_593 <= 0;
      end 
      if(_ram_w4_l8192_id0_7_cond_6_2) begin
        _tmp_1219 <= 0;
      end 
      if(_ram_w4_l8192_id0_7_cond_0_1) begin
        _tmp_257 <= 0;
      end 
      if(_ram_w4_l8192_id0_7_cond_1_1) begin
        ram_w4_l8192_id0_7_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id0_7_cond_2_1) begin
        _tmp_593 <= 1;
      end 
      _ram_w4_l8192_id0_7_cond_3_2 <= _ram_w4_l8192_id0_7_cond_3_1;
      if(_ram_w4_l8192_id0_7_cond_4_1) begin
        ram_w4_l8192_id0_7_1_wenable <= 0;
        _tmp_1151 <= 0;
      end 
      if(_ram_w4_l8192_id0_7_cond_5_1) begin
        _tmp_1219 <= 1;
      end 
      _ram_w4_l8192_id0_7_cond_6_2 <= _ram_w4_l8192_id0_7_cond_6_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_256 == 0)) begin
        _tmp_285 <= 0;
        _tmp_255 <= req_block_size_33 - 1;
        _tmp_256 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_256 == 0)) begin
        _tmp_258 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_256 == 0)) begin
        _tmp_259 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_256 == 0)) begin
        _tmp_260 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_256 == 0)) begin
        _tmp_261 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_256 == 0)) begin
        _tmp_262 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_256 == 0)) begin
        _tmp_263 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_256 == 0)) begin
        _tmp_264 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_256 == 0)) begin
        _tmp_265 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 3) && (_tmp_256 == 0)) begin
        _tmp_266 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0)) begin
        _tmp_255 <= _tmp_255 - 1;
        _tmp_256 <= _tmp_256 - 1;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0) && (_tmp_255 == 0)) begin
        _tmp_255 <= req_block_size_33 - 1;
        _tmp_285 <= _tmp_285 + 1;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0) && (_tmp_255 == 0) && (_tmp_285 == 8)) begin
        _tmp_285 <= 0;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0) && (_tmp_285 == 0)) begin
        _tmp_258 <= _tmp_267;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0) && (_tmp_285 == 1)) begin
        _tmp_259 <= _tmp_268;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0) && (_tmp_285 == 2)) begin
        _tmp_260 <= _tmp_269;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0) && (_tmp_285 == 3)) begin
        _tmp_261 <= _tmp_270;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0) && (_tmp_285 == 4)) begin
        _tmp_262 <= _tmp_271;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0) && (_tmp_285 == 5)) begin
        _tmp_263 <= _tmp_272;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0) && (_tmp_285 == 6)) begin
        _tmp_264 <= _tmp_273;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0) && (_tmp_285 == 7)) begin
        _tmp_265 <= _tmp_274;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0) && (_tmp_285 == 8)) begin
        _tmp_266 <= _tmp_275;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0)) begin
        ram_w4_l8192_id0_7_1_addr <= _tmp_276;
        ram_w4_l8192_id0_7_1_wdata <= _dataflow_slice_odata_50;
        ram_w4_l8192_id0_7_1_wenable <= _tmp_285 == 0;
      end 
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 == 1)) begin
        _tmp_257 <= 1;
      end 
      _ram_w4_l8192_id0_7_cond_0_1 <= 1;
      _ram_w4_l8192_id0_7_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12)) begin
        ram_w4_l8192_id0_7_0_addr <= _stream_conv2d_16_source_28_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_7_cond_2_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      _ram_w4_l8192_id0_7_cond_3_1 <= _stream_conv2d_16_source_28_source_ram_renable && (_stream_conv2d_16_source_28_source_ram_sel == 12);
      if(_maxi_read_start && (_maxi_read_op_sel == 8) && (_tmp_1150 == 0)) begin
        ram_w4_l8192_id0_7_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1150 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_145 && ((_tmp_1150 > 0) && !_tmp_1151) && (_tmp_1150 > 0)) begin
        ram_w4_l8192_id0_7_1_addr <= ram_w4_l8192_id0_7_1_addr + _maxi_read_local_stride;
        ram_w4_l8192_id0_7_1_wdata <= _dataflow_slice_odata_145;
        ram_w4_l8192_id0_7_1_wenable <= 1;
        _tmp_1150 <= _tmp_1150 - 1;
      end 
      if(_dataflow_slice_ovalid_145 && ((_tmp_1150 > 0) && !_tmp_1151) && (_tmp_1150 == 1)) begin
        _tmp_1151 <= 1;
      end 
      _ram_w4_l8192_id0_7_cond_4_1 <= 1;
      if(_stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4)) begin
        ram_w4_l8192_id0_7_0_addr <= _stream_matmul_29_source_20_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id0_7_cond_5_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      _ram_w4_l8192_id0_7_cond_6_1 <= _stream_matmul_29_source_20_source_ram_renable && (_stream_matmul_29_source_20_source_ram_sel == 4);
      ram_w4_l8192_id0_7_0_wdata <= 0;
      ram_w4_l8192_id0_7_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id1_0_1_addr <= 0;
      ram_w4_l8192_id1_0_1_wdata <= 0;
      ram_w4_l8192_id1_0_1_wenable <= 0;
      _ram_w4_l8192_id1_0_cond_0_1 <= 0;
      ram_w4_l8192_id1_0_0_addr <= 0;
      _ram_w4_l8192_id1_0_cond_1_1 <= 0;
      _tmp_600 <= 0;
      _ram_w4_l8192_id1_0_cond_2_1 <= 0;
      _ram_w4_l8192_id1_0_cond_2_2 <= 0;
      ram_w4_l8192_id1_0_0_wdata <= 0;
      ram_w4_l8192_id1_0_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id1_0_cond_2_2) begin
        _tmp_600 <= 0;
      end 
      if(_ram_w4_l8192_id1_0_cond_0_1) begin
        ram_w4_l8192_id1_0_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id1_0_cond_1_1) begin
        _tmp_600 <= 1;
      end 
      _ram_w4_l8192_id1_0_cond_2_2 <= _ram_w4_l8192_id1_0_cond_2_1;
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0)) begin
        ram_w4_l8192_id1_0_1_addr <= _tmp_60;
        ram_w4_l8192_id1_0_1_wdata <= _dataflow_slice_odata_29;
        ram_w4_l8192_id1_0_1_wenable <= _tmp_68 == 1;
      end 
      _ram_w4_l8192_id1_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13)) begin
        ram_w4_l8192_id1_0_0_addr <= _stream_conv2d_16_source_29_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id1_0_cond_1_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      _ram_w4_l8192_id1_0_cond_2_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      ram_w4_l8192_id1_0_0_wdata <= 0;
      ram_w4_l8192_id1_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id1_1_1_addr <= 0;
      ram_w4_l8192_id1_1_1_wdata <= 0;
      ram_w4_l8192_id1_1_1_wenable <= 0;
      _ram_w4_l8192_id1_1_cond_0_1 <= 0;
      ram_w4_l8192_id1_1_0_addr <= 0;
      _ram_w4_l8192_id1_1_cond_1_1 <= 0;
      _tmp_601 <= 0;
      _ram_w4_l8192_id1_1_cond_2_1 <= 0;
      _ram_w4_l8192_id1_1_cond_2_2 <= 0;
      ram_w4_l8192_id1_1_0_wdata <= 0;
      ram_w4_l8192_id1_1_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id1_1_cond_2_2) begin
        _tmp_601 <= 0;
      end 
      if(_ram_w4_l8192_id1_1_cond_0_1) begin
        ram_w4_l8192_id1_1_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id1_1_cond_1_1) begin
        _tmp_601 <= 1;
      end 
      _ram_w4_l8192_id1_1_cond_2_2 <= _ram_w4_l8192_id1_1_cond_2_1;
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0)) begin
        ram_w4_l8192_id1_1_1_addr <= _tmp_91;
        ram_w4_l8192_id1_1_1_wdata <= _dataflow_slice_odata_32;
        ram_w4_l8192_id1_1_1_wenable <= _tmp_99 == 1;
      end 
      _ram_w4_l8192_id1_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13)) begin
        ram_w4_l8192_id1_1_0_addr <= _stream_conv2d_16_source_29_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id1_1_cond_1_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      _ram_w4_l8192_id1_1_cond_2_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      ram_w4_l8192_id1_1_0_wdata <= 0;
      ram_w4_l8192_id1_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id1_2_1_addr <= 0;
      ram_w4_l8192_id1_2_1_wdata <= 0;
      ram_w4_l8192_id1_2_1_wenable <= 0;
      _ram_w4_l8192_id1_2_cond_0_1 <= 0;
      ram_w4_l8192_id1_2_0_addr <= 0;
      _ram_w4_l8192_id1_2_cond_1_1 <= 0;
      _tmp_602 <= 0;
      _ram_w4_l8192_id1_2_cond_2_1 <= 0;
      _ram_w4_l8192_id1_2_cond_2_2 <= 0;
      ram_w4_l8192_id1_2_0_wdata <= 0;
      ram_w4_l8192_id1_2_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id1_2_cond_2_2) begin
        _tmp_602 <= 0;
      end 
      if(_ram_w4_l8192_id1_2_cond_0_1) begin
        ram_w4_l8192_id1_2_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id1_2_cond_1_1) begin
        _tmp_602 <= 1;
      end 
      _ram_w4_l8192_id1_2_cond_2_2 <= _ram_w4_l8192_id1_2_cond_2_1;
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0)) begin
        ram_w4_l8192_id1_2_1_addr <= _tmp_122;
        ram_w4_l8192_id1_2_1_wdata <= _dataflow_slice_odata_35;
        ram_w4_l8192_id1_2_1_wenable <= _tmp_130 == 1;
      end 
      _ram_w4_l8192_id1_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13)) begin
        ram_w4_l8192_id1_2_0_addr <= _stream_conv2d_16_source_29_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id1_2_cond_1_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      _ram_w4_l8192_id1_2_cond_2_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      ram_w4_l8192_id1_2_0_wdata <= 0;
      ram_w4_l8192_id1_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id1_3_1_addr <= 0;
      ram_w4_l8192_id1_3_1_wdata <= 0;
      ram_w4_l8192_id1_3_1_wenable <= 0;
      _ram_w4_l8192_id1_3_cond_0_1 <= 0;
      ram_w4_l8192_id1_3_0_addr <= 0;
      _ram_w4_l8192_id1_3_cond_1_1 <= 0;
      _tmp_603 <= 0;
      _ram_w4_l8192_id1_3_cond_2_1 <= 0;
      _ram_w4_l8192_id1_3_cond_2_2 <= 0;
      ram_w4_l8192_id1_3_0_wdata <= 0;
      ram_w4_l8192_id1_3_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id1_3_cond_2_2) begin
        _tmp_603 <= 0;
      end 
      if(_ram_w4_l8192_id1_3_cond_0_1) begin
        ram_w4_l8192_id1_3_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id1_3_cond_1_1) begin
        _tmp_603 <= 1;
      end 
      _ram_w4_l8192_id1_3_cond_2_2 <= _ram_w4_l8192_id1_3_cond_2_1;
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0)) begin
        ram_w4_l8192_id1_3_1_addr <= _tmp_153;
        ram_w4_l8192_id1_3_1_wdata <= _dataflow_slice_odata_38;
        ram_w4_l8192_id1_3_1_wenable <= _tmp_161 == 1;
      end 
      _ram_w4_l8192_id1_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13)) begin
        ram_w4_l8192_id1_3_0_addr <= _stream_conv2d_16_source_29_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id1_3_cond_1_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      _ram_w4_l8192_id1_3_cond_2_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      ram_w4_l8192_id1_3_0_wdata <= 0;
      ram_w4_l8192_id1_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id1_4_1_addr <= 0;
      ram_w4_l8192_id1_4_1_wdata <= 0;
      ram_w4_l8192_id1_4_1_wenable <= 0;
      _ram_w4_l8192_id1_4_cond_0_1 <= 0;
      ram_w4_l8192_id1_4_0_addr <= 0;
      _ram_w4_l8192_id1_4_cond_1_1 <= 0;
      _tmp_604 <= 0;
      _ram_w4_l8192_id1_4_cond_2_1 <= 0;
      _ram_w4_l8192_id1_4_cond_2_2 <= 0;
      ram_w4_l8192_id1_4_0_wdata <= 0;
      ram_w4_l8192_id1_4_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id1_4_cond_2_2) begin
        _tmp_604 <= 0;
      end 
      if(_ram_w4_l8192_id1_4_cond_0_1) begin
        ram_w4_l8192_id1_4_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id1_4_cond_1_1) begin
        _tmp_604 <= 1;
      end 
      _ram_w4_l8192_id1_4_cond_2_2 <= _ram_w4_l8192_id1_4_cond_2_1;
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0)) begin
        ram_w4_l8192_id1_4_1_addr <= _tmp_184;
        ram_w4_l8192_id1_4_1_wdata <= _dataflow_slice_odata_41;
        ram_w4_l8192_id1_4_1_wenable <= _tmp_192 == 1;
      end 
      _ram_w4_l8192_id1_4_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13)) begin
        ram_w4_l8192_id1_4_0_addr <= _stream_conv2d_16_source_29_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id1_4_cond_1_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      _ram_w4_l8192_id1_4_cond_2_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      ram_w4_l8192_id1_4_0_wdata <= 0;
      ram_w4_l8192_id1_4_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id1_5_1_addr <= 0;
      ram_w4_l8192_id1_5_1_wdata <= 0;
      ram_w4_l8192_id1_5_1_wenable <= 0;
      _ram_w4_l8192_id1_5_cond_0_1 <= 0;
      ram_w4_l8192_id1_5_0_addr <= 0;
      _ram_w4_l8192_id1_5_cond_1_1 <= 0;
      _tmp_605 <= 0;
      _ram_w4_l8192_id1_5_cond_2_1 <= 0;
      _ram_w4_l8192_id1_5_cond_2_2 <= 0;
      ram_w4_l8192_id1_5_0_wdata <= 0;
      ram_w4_l8192_id1_5_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id1_5_cond_2_2) begin
        _tmp_605 <= 0;
      end 
      if(_ram_w4_l8192_id1_5_cond_0_1) begin
        ram_w4_l8192_id1_5_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id1_5_cond_1_1) begin
        _tmp_605 <= 1;
      end 
      _ram_w4_l8192_id1_5_cond_2_2 <= _ram_w4_l8192_id1_5_cond_2_1;
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0)) begin
        ram_w4_l8192_id1_5_1_addr <= _tmp_215;
        ram_w4_l8192_id1_5_1_wdata <= _dataflow_slice_odata_44;
        ram_w4_l8192_id1_5_1_wenable <= _tmp_223 == 1;
      end 
      _ram_w4_l8192_id1_5_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13)) begin
        ram_w4_l8192_id1_5_0_addr <= _stream_conv2d_16_source_29_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id1_5_cond_1_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      _ram_w4_l8192_id1_5_cond_2_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      ram_w4_l8192_id1_5_0_wdata <= 0;
      ram_w4_l8192_id1_5_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id1_6_1_addr <= 0;
      ram_w4_l8192_id1_6_1_wdata <= 0;
      ram_w4_l8192_id1_6_1_wenable <= 0;
      _ram_w4_l8192_id1_6_cond_0_1 <= 0;
      ram_w4_l8192_id1_6_0_addr <= 0;
      _ram_w4_l8192_id1_6_cond_1_1 <= 0;
      _tmp_606 <= 0;
      _ram_w4_l8192_id1_6_cond_2_1 <= 0;
      _ram_w4_l8192_id1_6_cond_2_2 <= 0;
      ram_w4_l8192_id1_6_0_wdata <= 0;
      ram_w4_l8192_id1_6_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id1_6_cond_2_2) begin
        _tmp_606 <= 0;
      end 
      if(_ram_w4_l8192_id1_6_cond_0_1) begin
        ram_w4_l8192_id1_6_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id1_6_cond_1_1) begin
        _tmp_606 <= 1;
      end 
      _ram_w4_l8192_id1_6_cond_2_2 <= _ram_w4_l8192_id1_6_cond_2_1;
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0)) begin
        ram_w4_l8192_id1_6_1_addr <= _tmp_246;
        ram_w4_l8192_id1_6_1_wdata <= _dataflow_slice_odata_47;
        ram_w4_l8192_id1_6_1_wenable <= _tmp_254 == 1;
      end 
      _ram_w4_l8192_id1_6_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13)) begin
        ram_w4_l8192_id1_6_0_addr <= _stream_conv2d_16_source_29_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id1_6_cond_1_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      _ram_w4_l8192_id1_6_cond_2_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      ram_w4_l8192_id1_6_0_wdata <= 0;
      ram_w4_l8192_id1_6_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id1_7_1_addr <= 0;
      ram_w4_l8192_id1_7_1_wdata <= 0;
      ram_w4_l8192_id1_7_1_wenable <= 0;
      _ram_w4_l8192_id1_7_cond_0_1 <= 0;
      ram_w4_l8192_id1_7_0_addr <= 0;
      _ram_w4_l8192_id1_7_cond_1_1 <= 0;
      _tmp_607 <= 0;
      _ram_w4_l8192_id1_7_cond_2_1 <= 0;
      _ram_w4_l8192_id1_7_cond_2_2 <= 0;
      ram_w4_l8192_id1_7_0_wdata <= 0;
      ram_w4_l8192_id1_7_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id1_7_cond_2_2) begin
        _tmp_607 <= 0;
      end 
      if(_ram_w4_l8192_id1_7_cond_0_1) begin
        ram_w4_l8192_id1_7_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id1_7_cond_1_1) begin
        _tmp_607 <= 1;
      end 
      _ram_w4_l8192_id1_7_cond_2_2 <= _ram_w4_l8192_id1_7_cond_2_1;
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0)) begin
        ram_w4_l8192_id1_7_1_addr <= _tmp_277;
        ram_w4_l8192_id1_7_1_wdata <= _dataflow_slice_odata_50;
        ram_w4_l8192_id1_7_1_wenable <= _tmp_285 == 1;
      end 
      _ram_w4_l8192_id1_7_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13)) begin
        ram_w4_l8192_id1_7_0_addr <= _stream_conv2d_16_source_29_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id1_7_cond_1_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      _ram_w4_l8192_id1_7_cond_2_1 <= _stream_conv2d_16_source_29_source_ram_renable && (_stream_conv2d_16_source_29_source_ram_sel == 13);
      ram_w4_l8192_id1_7_0_wdata <= 0;
      ram_w4_l8192_id1_7_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id2_0_1_addr <= 0;
      ram_w4_l8192_id2_0_1_wdata <= 0;
      ram_w4_l8192_id2_0_1_wenable <= 0;
      _ram_w4_l8192_id2_0_cond_0_1 <= 0;
      ram_w4_l8192_id2_0_0_addr <= 0;
      _ram_w4_l8192_id2_0_cond_1_1 <= 0;
      _tmp_614 <= 0;
      _ram_w4_l8192_id2_0_cond_2_1 <= 0;
      _ram_w4_l8192_id2_0_cond_2_2 <= 0;
      ram_w4_l8192_id2_0_0_wdata <= 0;
      ram_w4_l8192_id2_0_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id2_0_cond_2_2) begin
        _tmp_614 <= 0;
      end 
      if(_ram_w4_l8192_id2_0_cond_0_1) begin
        ram_w4_l8192_id2_0_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id2_0_cond_1_1) begin
        _tmp_614 <= 1;
      end 
      _ram_w4_l8192_id2_0_cond_2_2 <= _ram_w4_l8192_id2_0_cond_2_1;
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0)) begin
        ram_w4_l8192_id2_0_1_addr <= _tmp_61;
        ram_w4_l8192_id2_0_1_wdata <= _dataflow_slice_odata_29;
        ram_w4_l8192_id2_0_1_wenable <= _tmp_68 == 2;
      end 
      _ram_w4_l8192_id2_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14)) begin
        ram_w4_l8192_id2_0_0_addr <= _stream_conv2d_16_source_30_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id2_0_cond_1_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      _ram_w4_l8192_id2_0_cond_2_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      ram_w4_l8192_id2_0_0_wdata <= 0;
      ram_w4_l8192_id2_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id2_1_1_addr <= 0;
      ram_w4_l8192_id2_1_1_wdata <= 0;
      ram_w4_l8192_id2_1_1_wenable <= 0;
      _ram_w4_l8192_id2_1_cond_0_1 <= 0;
      ram_w4_l8192_id2_1_0_addr <= 0;
      _ram_w4_l8192_id2_1_cond_1_1 <= 0;
      _tmp_615 <= 0;
      _ram_w4_l8192_id2_1_cond_2_1 <= 0;
      _ram_w4_l8192_id2_1_cond_2_2 <= 0;
      ram_w4_l8192_id2_1_0_wdata <= 0;
      ram_w4_l8192_id2_1_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id2_1_cond_2_2) begin
        _tmp_615 <= 0;
      end 
      if(_ram_w4_l8192_id2_1_cond_0_1) begin
        ram_w4_l8192_id2_1_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id2_1_cond_1_1) begin
        _tmp_615 <= 1;
      end 
      _ram_w4_l8192_id2_1_cond_2_2 <= _ram_w4_l8192_id2_1_cond_2_1;
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0)) begin
        ram_w4_l8192_id2_1_1_addr <= _tmp_92;
        ram_w4_l8192_id2_1_1_wdata <= _dataflow_slice_odata_32;
        ram_w4_l8192_id2_1_1_wenable <= _tmp_99 == 2;
      end 
      _ram_w4_l8192_id2_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14)) begin
        ram_w4_l8192_id2_1_0_addr <= _stream_conv2d_16_source_30_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id2_1_cond_1_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      _ram_w4_l8192_id2_1_cond_2_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      ram_w4_l8192_id2_1_0_wdata <= 0;
      ram_w4_l8192_id2_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id2_2_1_addr <= 0;
      ram_w4_l8192_id2_2_1_wdata <= 0;
      ram_w4_l8192_id2_2_1_wenable <= 0;
      _ram_w4_l8192_id2_2_cond_0_1 <= 0;
      ram_w4_l8192_id2_2_0_addr <= 0;
      _ram_w4_l8192_id2_2_cond_1_1 <= 0;
      _tmp_616 <= 0;
      _ram_w4_l8192_id2_2_cond_2_1 <= 0;
      _ram_w4_l8192_id2_2_cond_2_2 <= 0;
      ram_w4_l8192_id2_2_0_wdata <= 0;
      ram_w4_l8192_id2_2_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id2_2_cond_2_2) begin
        _tmp_616 <= 0;
      end 
      if(_ram_w4_l8192_id2_2_cond_0_1) begin
        ram_w4_l8192_id2_2_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id2_2_cond_1_1) begin
        _tmp_616 <= 1;
      end 
      _ram_w4_l8192_id2_2_cond_2_2 <= _ram_w4_l8192_id2_2_cond_2_1;
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0)) begin
        ram_w4_l8192_id2_2_1_addr <= _tmp_123;
        ram_w4_l8192_id2_2_1_wdata <= _dataflow_slice_odata_35;
        ram_w4_l8192_id2_2_1_wenable <= _tmp_130 == 2;
      end 
      _ram_w4_l8192_id2_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14)) begin
        ram_w4_l8192_id2_2_0_addr <= _stream_conv2d_16_source_30_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id2_2_cond_1_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      _ram_w4_l8192_id2_2_cond_2_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      ram_w4_l8192_id2_2_0_wdata <= 0;
      ram_w4_l8192_id2_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id2_3_1_addr <= 0;
      ram_w4_l8192_id2_3_1_wdata <= 0;
      ram_w4_l8192_id2_3_1_wenable <= 0;
      _ram_w4_l8192_id2_3_cond_0_1 <= 0;
      ram_w4_l8192_id2_3_0_addr <= 0;
      _ram_w4_l8192_id2_3_cond_1_1 <= 0;
      _tmp_617 <= 0;
      _ram_w4_l8192_id2_3_cond_2_1 <= 0;
      _ram_w4_l8192_id2_3_cond_2_2 <= 0;
      ram_w4_l8192_id2_3_0_wdata <= 0;
      ram_w4_l8192_id2_3_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id2_3_cond_2_2) begin
        _tmp_617 <= 0;
      end 
      if(_ram_w4_l8192_id2_3_cond_0_1) begin
        ram_w4_l8192_id2_3_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id2_3_cond_1_1) begin
        _tmp_617 <= 1;
      end 
      _ram_w4_l8192_id2_3_cond_2_2 <= _ram_w4_l8192_id2_3_cond_2_1;
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0)) begin
        ram_w4_l8192_id2_3_1_addr <= _tmp_154;
        ram_w4_l8192_id2_3_1_wdata <= _dataflow_slice_odata_38;
        ram_w4_l8192_id2_3_1_wenable <= _tmp_161 == 2;
      end 
      _ram_w4_l8192_id2_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14)) begin
        ram_w4_l8192_id2_3_0_addr <= _stream_conv2d_16_source_30_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id2_3_cond_1_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      _ram_w4_l8192_id2_3_cond_2_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      ram_w4_l8192_id2_3_0_wdata <= 0;
      ram_w4_l8192_id2_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id2_4_1_addr <= 0;
      ram_w4_l8192_id2_4_1_wdata <= 0;
      ram_w4_l8192_id2_4_1_wenable <= 0;
      _ram_w4_l8192_id2_4_cond_0_1 <= 0;
      ram_w4_l8192_id2_4_0_addr <= 0;
      _ram_w4_l8192_id2_4_cond_1_1 <= 0;
      _tmp_618 <= 0;
      _ram_w4_l8192_id2_4_cond_2_1 <= 0;
      _ram_w4_l8192_id2_4_cond_2_2 <= 0;
      ram_w4_l8192_id2_4_0_wdata <= 0;
      ram_w4_l8192_id2_4_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id2_4_cond_2_2) begin
        _tmp_618 <= 0;
      end 
      if(_ram_w4_l8192_id2_4_cond_0_1) begin
        ram_w4_l8192_id2_4_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id2_4_cond_1_1) begin
        _tmp_618 <= 1;
      end 
      _ram_w4_l8192_id2_4_cond_2_2 <= _ram_w4_l8192_id2_4_cond_2_1;
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0)) begin
        ram_w4_l8192_id2_4_1_addr <= _tmp_185;
        ram_w4_l8192_id2_4_1_wdata <= _dataflow_slice_odata_41;
        ram_w4_l8192_id2_4_1_wenable <= _tmp_192 == 2;
      end 
      _ram_w4_l8192_id2_4_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14)) begin
        ram_w4_l8192_id2_4_0_addr <= _stream_conv2d_16_source_30_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id2_4_cond_1_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      _ram_w4_l8192_id2_4_cond_2_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      ram_w4_l8192_id2_4_0_wdata <= 0;
      ram_w4_l8192_id2_4_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id2_5_1_addr <= 0;
      ram_w4_l8192_id2_5_1_wdata <= 0;
      ram_w4_l8192_id2_5_1_wenable <= 0;
      _ram_w4_l8192_id2_5_cond_0_1 <= 0;
      ram_w4_l8192_id2_5_0_addr <= 0;
      _ram_w4_l8192_id2_5_cond_1_1 <= 0;
      _tmp_619 <= 0;
      _ram_w4_l8192_id2_5_cond_2_1 <= 0;
      _ram_w4_l8192_id2_5_cond_2_2 <= 0;
      ram_w4_l8192_id2_5_0_wdata <= 0;
      ram_w4_l8192_id2_5_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id2_5_cond_2_2) begin
        _tmp_619 <= 0;
      end 
      if(_ram_w4_l8192_id2_5_cond_0_1) begin
        ram_w4_l8192_id2_5_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id2_5_cond_1_1) begin
        _tmp_619 <= 1;
      end 
      _ram_w4_l8192_id2_5_cond_2_2 <= _ram_w4_l8192_id2_5_cond_2_1;
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0)) begin
        ram_w4_l8192_id2_5_1_addr <= _tmp_216;
        ram_w4_l8192_id2_5_1_wdata <= _dataflow_slice_odata_44;
        ram_w4_l8192_id2_5_1_wenable <= _tmp_223 == 2;
      end 
      _ram_w4_l8192_id2_5_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14)) begin
        ram_w4_l8192_id2_5_0_addr <= _stream_conv2d_16_source_30_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id2_5_cond_1_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      _ram_w4_l8192_id2_5_cond_2_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      ram_w4_l8192_id2_5_0_wdata <= 0;
      ram_w4_l8192_id2_5_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id2_6_1_addr <= 0;
      ram_w4_l8192_id2_6_1_wdata <= 0;
      ram_w4_l8192_id2_6_1_wenable <= 0;
      _ram_w4_l8192_id2_6_cond_0_1 <= 0;
      ram_w4_l8192_id2_6_0_addr <= 0;
      _ram_w4_l8192_id2_6_cond_1_1 <= 0;
      _tmp_620 <= 0;
      _ram_w4_l8192_id2_6_cond_2_1 <= 0;
      _ram_w4_l8192_id2_6_cond_2_2 <= 0;
      ram_w4_l8192_id2_6_0_wdata <= 0;
      ram_w4_l8192_id2_6_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id2_6_cond_2_2) begin
        _tmp_620 <= 0;
      end 
      if(_ram_w4_l8192_id2_6_cond_0_1) begin
        ram_w4_l8192_id2_6_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id2_6_cond_1_1) begin
        _tmp_620 <= 1;
      end 
      _ram_w4_l8192_id2_6_cond_2_2 <= _ram_w4_l8192_id2_6_cond_2_1;
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0)) begin
        ram_w4_l8192_id2_6_1_addr <= _tmp_247;
        ram_w4_l8192_id2_6_1_wdata <= _dataflow_slice_odata_47;
        ram_w4_l8192_id2_6_1_wenable <= _tmp_254 == 2;
      end 
      _ram_w4_l8192_id2_6_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14)) begin
        ram_w4_l8192_id2_6_0_addr <= _stream_conv2d_16_source_30_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id2_6_cond_1_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      _ram_w4_l8192_id2_6_cond_2_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      ram_w4_l8192_id2_6_0_wdata <= 0;
      ram_w4_l8192_id2_6_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id2_7_1_addr <= 0;
      ram_w4_l8192_id2_7_1_wdata <= 0;
      ram_w4_l8192_id2_7_1_wenable <= 0;
      _ram_w4_l8192_id2_7_cond_0_1 <= 0;
      ram_w4_l8192_id2_7_0_addr <= 0;
      _ram_w4_l8192_id2_7_cond_1_1 <= 0;
      _tmp_621 <= 0;
      _ram_w4_l8192_id2_7_cond_2_1 <= 0;
      _ram_w4_l8192_id2_7_cond_2_2 <= 0;
      ram_w4_l8192_id2_7_0_wdata <= 0;
      ram_w4_l8192_id2_7_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id2_7_cond_2_2) begin
        _tmp_621 <= 0;
      end 
      if(_ram_w4_l8192_id2_7_cond_0_1) begin
        ram_w4_l8192_id2_7_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id2_7_cond_1_1) begin
        _tmp_621 <= 1;
      end 
      _ram_w4_l8192_id2_7_cond_2_2 <= _ram_w4_l8192_id2_7_cond_2_1;
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0)) begin
        ram_w4_l8192_id2_7_1_addr <= _tmp_278;
        ram_w4_l8192_id2_7_1_wdata <= _dataflow_slice_odata_50;
        ram_w4_l8192_id2_7_1_wenable <= _tmp_285 == 2;
      end 
      _ram_w4_l8192_id2_7_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14)) begin
        ram_w4_l8192_id2_7_0_addr <= _stream_conv2d_16_source_30_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id2_7_cond_1_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      _ram_w4_l8192_id2_7_cond_2_1 <= _stream_conv2d_16_source_30_source_ram_renable && (_stream_conv2d_16_source_30_source_ram_sel == 14);
      ram_w4_l8192_id2_7_0_wdata <= 0;
      ram_w4_l8192_id2_7_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id3_0_1_addr <= 0;
      ram_w4_l8192_id3_0_1_wdata <= 0;
      ram_w4_l8192_id3_0_1_wenable <= 0;
      _ram_w4_l8192_id3_0_cond_0_1 <= 0;
      ram_w4_l8192_id3_0_0_addr <= 0;
      _ram_w4_l8192_id3_0_cond_1_1 <= 0;
      _tmp_628 <= 0;
      _ram_w4_l8192_id3_0_cond_2_1 <= 0;
      _ram_w4_l8192_id3_0_cond_2_2 <= 0;
      ram_w4_l8192_id3_0_0_wdata <= 0;
      ram_w4_l8192_id3_0_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id3_0_cond_2_2) begin
        _tmp_628 <= 0;
      end 
      if(_ram_w4_l8192_id3_0_cond_0_1) begin
        ram_w4_l8192_id3_0_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id3_0_cond_1_1) begin
        _tmp_628 <= 1;
      end 
      _ram_w4_l8192_id3_0_cond_2_2 <= _ram_w4_l8192_id3_0_cond_2_1;
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0)) begin
        ram_w4_l8192_id3_0_1_addr <= _tmp_62;
        ram_w4_l8192_id3_0_1_wdata <= _dataflow_slice_odata_29;
        ram_w4_l8192_id3_0_1_wenable <= _tmp_68 == 3;
      end 
      _ram_w4_l8192_id3_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15)) begin
        ram_w4_l8192_id3_0_0_addr <= _stream_conv2d_16_source_31_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id3_0_cond_1_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      _ram_w4_l8192_id3_0_cond_2_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      ram_w4_l8192_id3_0_0_wdata <= 0;
      ram_w4_l8192_id3_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id3_1_1_addr <= 0;
      ram_w4_l8192_id3_1_1_wdata <= 0;
      ram_w4_l8192_id3_1_1_wenable <= 0;
      _ram_w4_l8192_id3_1_cond_0_1 <= 0;
      ram_w4_l8192_id3_1_0_addr <= 0;
      _ram_w4_l8192_id3_1_cond_1_1 <= 0;
      _tmp_629 <= 0;
      _ram_w4_l8192_id3_1_cond_2_1 <= 0;
      _ram_w4_l8192_id3_1_cond_2_2 <= 0;
      ram_w4_l8192_id3_1_0_wdata <= 0;
      ram_w4_l8192_id3_1_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id3_1_cond_2_2) begin
        _tmp_629 <= 0;
      end 
      if(_ram_w4_l8192_id3_1_cond_0_1) begin
        ram_w4_l8192_id3_1_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id3_1_cond_1_1) begin
        _tmp_629 <= 1;
      end 
      _ram_w4_l8192_id3_1_cond_2_2 <= _ram_w4_l8192_id3_1_cond_2_1;
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0)) begin
        ram_w4_l8192_id3_1_1_addr <= _tmp_93;
        ram_w4_l8192_id3_1_1_wdata <= _dataflow_slice_odata_32;
        ram_w4_l8192_id3_1_1_wenable <= _tmp_99 == 3;
      end 
      _ram_w4_l8192_id3_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15)) begin
        ram_w4_l8192_id3_1_0_addr <= _stream_conv2d_16_source_31_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id3_1_cond_1_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      _ram_w4_l8192_id3_1_cond_2_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      ram_w4_l8192_id3_1_0_wdata <= 0;
      ram_w4_l8192_id3_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id3_2_1_addr <= 0;
      ram_w4_l8192_id3_2_1_wdata <= 0;
      ram_w4_l8192_id3_2_1_wenable <= 0;
      _ram_w4_l8192_id3_2_cond_0_1 <= 0;
      ram_w4_l8192_id3_2_0_addr <= 0;
      _ram_w4_l8192_id3_2_cond_1_1 <= 0;
      _tmp_630 <= 0;
      _ram_w4_l8192_id3_2_cond_2_1 <= 0;
      _ram_w4_l8192_id3_2_cond_2_2 <= 0;
      ram_w4_l8192_id3_2_0_wdata <= 0;
      ram_w4_l8192_id3_2_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id3_2_cond_2_2) begin
        _tmp_630 <= 0;
      end 
      if(_ram_w4_l8192_id3_2_cond_0_1) begin
        ram_w4_l8192_id3_2_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id3_2_cond_1_1) begin
        _tmp_630 <= 1;
      end 
      _ram_w4_l8192_id3_2_cond_2_2 <= _ram_w4_l8192_id3_2_cond_2_1;
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0)) begin
        ram_w4_l8192_id3_2_1_addr <= _tmp_124;
        ram_w4_l8192_id3_2_1_wdata <= _dataflow_slice_odata_35;
        ram_w4_l8192_id3_2_1_wenable <= _tmp_130 == 3;
      end 
      _ram_w4_l8192_id3_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15)) begin
        ram_w4_l8192_id3_2_0_addr <= _stream_conv2d_16_source_31_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id3_2_cond_1_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      _ram_w4_l8192_id3_2_cond_2_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      ram_w4_l8192_id3_2_0_wdata <= 0;
      ram_w4_l8192_id3_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id3_3_1_addr <= 0;
      ram_w4_l8192_id3_3_1_wdata <= 0;
      ram_w4_l8192_id3_3_1_wenable <= 0;
      _ram_w4_l8192_id3_3_cond_0_1 <= 0;
      ram_w4_l8192_id3_3_0_addr <= 0;
      _ram_w4_l8192_id3_3_cond_1_1 <= 0;
      _tmp_631 <= 0;
      _ram_w4_l8192_id3_3_cond_2_1 <= 0;
      _ram_w4_l8192_id3_3_cond_2_2 <= 0;
      ram_w4_l8192_id3_3_0_wdata <= 0;
      ram_w4_l8192_id3_3_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id3_3_cond_2_2) begin
        _tmp_631 <= 0;
      end 
      if(_ram_w4_l8192_id3_3_cond_0_1) begin
        ram_w4_l8192_id3_3_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id3_3_cond_1_1) begin
        _tmp_631 <= 1;
      end 
      _ram_w4_l8192_id3_3_cond_2_2 <= _ram_w4_l8192_id3_3_cond_2_1;
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0)) begin
        ram_w4_l8192_id3_3_1_addr <= _tmp_155;
        ram_w4_l8192_id3_3_1_wdata <= _dataflow_slice_odata_38;
        ram_w4_l8192_id3_3_1_wenable <= _tmp_161 == 3;
      end 
      _ram_w4_l8192_id3_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15)) begin
        ram_w4_l8192_id3_3_0_addr <= _stream_conv2d_16_source_31_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id3_3_cond_1_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      _ram_w4_l8192_id3_3_cond_2_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      ram_w4_l8192_id3_3_0_wdata <= 0;
      ram_w4_l8192_id3_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id3_4_1_addr <= 0;
      ram_w4_l8192_id3_4_1_wdata <= 0;
      ram_w4_l8192_id3_4_1_wenable <= 0;
      _ram_w4_l8192_id3_4_cond_0_1 <= 0;
      ram_w4_l8192_id3_4_0_addr <= 0;
      _ram_w4_l8192_id3_4_cond_1_1 <= 0;
      _tmp_632 <= 0;
      _ram_w4_l8192_id3_4_cond_2_1 <= 0;
      _ram_w4_l8192_id3_4_cond_2_2 <= 0;
      ram_w4_l8192_id3_4_0_wdata <= 0;
      ram_w4_l8192_id3_4_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id3_4_cond_2_2) begin
        _tmp_632 <= 0;
      end 
      if(_ram_w4_l8192_id3_4_cond_0_1) begin
        ram_w4_l8192_id3_4_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id3_4_cond_1_1) begin
        _tmp_632 <= 1;
      end 
      _ram_w4_l8192_id3_4_cond_2_2 <= _ram_w4_l8192_id3_4_cond_2_1;
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0)) begin
        ram_w4_l8192_id3_4_1_addr <= _tmp_186;
        ram_w4_l8192_id3_4_1_wdata <= _dataflow_slice_odata_41;
        ram_w4_l8192_id3_4_1_wenable <= _tmp_192 == 3;
      end 
      _ram_w4_l8192_id3_4_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15)) begin
        ram_w4_l8192_id3_4_0_addr <= _stream_conv2d_16_source_31_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id3_4_cond_1_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      _ram_w4_l8192_id3_4_cond_2_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      ram_w4_l8192_id3_4_0_wdata <= 0;
      ram_w4_l8192_id3_4_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id3_5_1_addr <= 0;
      ram_w4_l8192_id3_5_1_wdata <= 0;
      ram_w4_l8192_id3_5_1_wenable <= 0;
      _ram_w4_l8192_id3_5_cond_0_1 <= 0;
      ram_w4_l8192_id3_5_0_addr <= 0;
      _ram_w4_l8192_id3_5_cond_1_1 <= 0;
      _tmp_633 <= 0;
      _ram_w4_l8192_id3_5_cond_2_1 <= 0;
      _ram_w4_l8192_id3_5_cond_2_2 <= 0;
      ram_w4_l8192_id3_5_0_wdata <= 0;
      ram_w4_l8192_id3_5_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id3_5_cond_2_2) begin
        _tmp_633 <= 0;
      end 
      if(_ram_w4_l8192_id3_5_cond_0_1) begin
        ram_w4_l8192_id3_5_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id3_5_cond_1_1) begin
        _tmp_633 <= 1;
      end 
      _ram_w4_l8192_id3_5_cond_2_2 <= _ram_w4_l8192_id3_5_cond_2_1;
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0)) begin
        ram_w4_l8192_id3_5_1_addr <= _tmp_217;
        ram_w4_l8192_id3_5_1_wdata <= _dataflow_slice_odata_44;
        ram_w4_l8192_id3_5_1_wenable <= _tmp_223 == 3;
      end 
      _ram_w4_l8192_id3_5_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15)) begin
        ram_w4_l8192_id3_5_0_addr <= _stream_conv2d_16_source_31_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id3_5_cond_1_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      _ram_w4_l8192_id3_5_cond_2_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      ram_w4_l8192_id3_5_0_wdata <= 0;
      ram_w4_l8192_id3_5_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id3_6_1_addr <= 0;
      ram_w4_l8192_id3_6_1_wdata <= 0;
      ram_w4_l8192_id3_6_1_wenable <= 0;
      _ram_w4_l8192_id3_6_cond_0_1 <= 0;
      ram_w4_l8192_id3_6_0_addr <= 0;
      _ram_w4_l8192_id3_6_cond_1_1 <= 0;
      _tmp_634 <= 0;
      _ram_w4_l8192_id3_6_cond_2_1 <= 0;
      _ram_w4_l8192_id3_6_cond_2_2 <= 0;
      ram_w4_l8192_id3_6_0_wdata <= 0;
      ram_w4_l8192_id3_6_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id3_6_cond_2_2) begin
        _tmp_634 <= 0;
      end 
      if(_ram_w4_l8192_id3_6_cond_0_1) begin
        ram_w4_l8192_id3_6_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id3_6_cond_1_1) begin
        _tmp_634 <= 1;
      end 
      _ram_w4_l8192_id3_6_cond_2_2 <= _ram_w4_l8192_id3_6_cond_2_1;
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0)) begin
        ram_w4_l8192_id3_6_1_addr <= _tmp_248;
        ram_w4_l8192_id3_6_1_wdata <= _dataflow_slice_odata_47;
        ram_w4_l8192_id3_6_1_wenable <= _tmp_254 == 3;
      end 
      _ram_w4_l8192_id3_6_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15)) begin
        ram_w4_l8192_id3_6_0_addr <= _stream_conv2d_16_source_31_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id3_6_cond_1_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      _ram_w4_l8192_id3_6_cond_2_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      ram_w4_l8192_id3_6_0_wdata <= 0;
      ram_w4_l8192_id3_6_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id3_7_1_addr <= 0;
      ram_w4_l8192_id3_7_1_wdata <= 0;
      ram_w4_l8192_id3_7_1_wenable <= 0;
      _ram_w4_l8192_id3_7_cond_0_1 <= 0;
      ram_w4_l8192_id3_7_0_addr <= 0;
      _ram_w4_l8192_id3_7_cond_1_1 <= 0;
      _tmp_635 <= 0;
      _ram_w4_l8192_id3_7_cond_2_1 <= 0;
      _ram_w4_l8192_id3_7_cond_2_2 <= 0;
      ram_w4_l8192_id3_7_0_wdata <= 0;
      ram_w4_l8192_id3_7_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id3_7_cond_2_2) begin
        _tmp_635 <= 0;
      end 
      if(_ram_w4_l8192_id3_7_cond_0_1) begin
        ram_w4_l8192_id3_7_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id3_7_cond_1_1) begin
        _tmp_635 <= 1;
      end 
      _ram_w4_l8192_id3_7_cond_2_2 <= _ram_w4_l8192_id3_7_cond_2_1;
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0)) begin
        ram_w4_l8192_id3_7_1_addr <= _tmp_279;
        ram_w4_l8192_id3_7_1_wdata <= _dataflow_slice_odata_50;
        ram_w4_l8192_id3_7_1_wenable <= _tmp_285 == 3;
      end 
      _ram_w4_l8192_id3_7_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15)) begin
        ram_w4_l8192_id3_7_0_addr <= _stream_conv2d_16_source_31_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id3_7_cond_1_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      _ram_w4_l8192_id3_7_cond_2_1 <= _stream_conv2d_16_source_31_source_ram_renable && (_stream_conv2d_16_source_31_source_ram_sel == 15);
      ram_w4_l8192_id3_7_0_wdata <= 0;
      ram_w4_l8192_id3_7_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id4_0_1_addr <= 0;
      ram_w4_l8192_id4_0_1_wdata <= 0;
      ram_w4_l8192_id4_0_1_wenable <= 0;
      _ram_w4_l8192_id4_0_cond_0_1 <= 0;
      ram_w4_l8192_id4_0_0_addr <= 0;
      _ram_w4_l8192_id4_0_cond_1_1 <= 0;
      _tmp_642 <= 0;
      _ram_w4_l8192_id4_0_cond_2_1 <= 0;
      _ram_w4_l8192_id4_0_cond_2_2 <= 0;
      ram_w4_l8192_id4_0_0_wdata <= 0;
      ram_w4_l8192_id4_0_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id4_0_cond_2_2) begin
        _tmp_642 <= 0;
      end 
      if(_ram_w4_l8192_id4_0_cond_0_1) begin
        ram_w4_l8192_id4_0_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id4_0_cond_1_1) begin
        _tmp_642 <= 1;
      end 
      _ram_w4_l8192_id4_0_cond_2_2 <= _ram_w4_l8192_id4_0_cond_2_1;
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0)) begin
        ram_w4_l8192_id4_0_1_addr <= _tmp_63;
        ram_w4_l8192_id4_0_1_wdata <= _dataflow_slice_odata_29;
        ram_w4_l8192_id4_0_1_wenable <= _tmp_68 == 4;
      end 
      _ram_w4_l8192_id4_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16)) begin
        ram_w4_l8192_id4_0_0_addr <= _stream_conv2d_16_source_32_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id4_0_cond_1_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      _ram_w4_l8192_id4_0_cond_2_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      ram_w4_l8192_id4_0_0_wdata <= 0;
      ram_w4_l8192_id4_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id4_1_1_addr <= 0;
      ram_w4_l8192_id4_1_1_wdata <= 0;
      ram_w4_l8192_id4_1_1_wenable <= 0;
      _ram_w4_l8192_id4_1_cond_0_1 <= 0;
      ram_w4_l8192_id4_1_0_addr <= 0;
      _ram_w4_l8192_id4_1_cond_1_1 <= 0;
      _tmp_643 <= 0;
      _ram_w4_l8192_id4_1_cond_2_1 <= 0;
      _ram_w4_l8192_id4_1_cond_2_2 <= 0;
      ram_w4_l8192_id4_1_0_wdata <= 0;
      ram_w4_l8192_id4_1_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id4_1_cond_2_2) begin
        _tmp_643 <= 0;
      end 
      if(_ram_w4_l8192_id4_1_cond_0_1) begin
        ram_w4_l8192_id4_1_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id4_1_cond_1_1) begin
        _tmp_643 <= 1;
      end 
      _ram_w4_l8192_id4_1_cond_2_2 <= _ram_w4_l8192_id4_1_cond_2_1;
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0)) begin
        ram_w4_l8192_id4_1_1_addr <= _tmp_94;
        ram_w4_l8192_id4_1_1_wdata <= _dataflow_slice_odata_32;
        ram_w4_l8192_id4_1_1_wenable <= _tmp_99 == 4;
      end 
      _ram_w4_l8192_id4_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16)) begin
        ram_w4_l8192_id4_1_0_addr <= _stream_conv2d_16_source_32_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id4_1_cond_1_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      _ram_w4_l8192_id4_1_cond_2_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      ram_w4_l8192_id4_1_0_wdata <= 0;
      ram_w4_l8192_id4_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id4_2_1_addr <= 0;
      ram_w4_l8192_id4_2_1_wdata <= 0;
      ram_w4_l8192_id4_2_1_wenable <= 0;
      _ram_w4_l8192_id4_2_cond_0_1 <= 0;
      ram_w4_l8192_id4_2_0_addr <= 0;
      _ram_w4_l8192_id4_2_cond_1_1 <= 0;
      _tmp_644 <= 0;
      _ram_w4_l8192_id4_2_cond_2_1 <= 0;
      _ram_w4_l8192_id4_2_cond_2_2 <= 0;
      ram_w4_l8192_id4_2_0_wdata <= 0;
      ram_w4_l8192_id4_2_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id4_2_cond_2_2) begin
        _tmp_644 <= 0;
      end 
      if(_ram_w4_l8192_id4_2_cond_0_1) begin
        ram_w4_l8192_id4_2_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id4_2_cond_1_1) begin
        _tmp_644 <= 1;
      end 
      _ram_w4_l8192_id4_2_cond_2_2 <= _ram_w4_l8192_id4_2_cond_2_1;
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0)) begin
        ram_w4_l8192_id4_2_1_addr <= _tmp_125;
        ram_w4_l8192_id4_2_1_wdata <= _dataflow_slice_odata_35;
        ram_w4_l8192_id4_2_1_wenable <= _tmp_130 == 4;
      end 
      _ram_w4_l8192_id4_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16)) begin
        ram_w4_l8192_id4_2_0_addr <= _stream_conv2d_16_source_32_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id4_2_cond_1_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      _ram_w4_l8192_id4_2_cond_2_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      ram_w4_l8192_id4_2_0_wdata <= 0;
      ram_w4_l8192_id4_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id4_3_1_addr <= 0;
      ram_w4_l8192_id4_3_1_wdata <= 0;
      ram_w4_l8192_id4_3_1_wenable <= 0;
      _ram_w4_l8192_id4_3_cond_0_1 <= 0;
      ram_w4_l8192_id4_3_0_addr <= 0;
      _ram_w4_l8192_id4_3_cond_1_1 <= 0;
      _tmp_645 <= 0;
      _ram_w4_l8192_id4_3_cond_2_1 <= 0;
      _ram_w4_l8192_id4_3_cond_2_2 <= 0;
      ram_w4_l8192_id4_3_0_wdata <= 0;
      ram_w4_l8192_id4_3_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id4_3_cond_2_2) begin
        _tmp_645 <= 0;
      end 
      if(_ram_w4_l8192_id4_3_cond_0_1) begin
        ram_w4_l8192_id4_3_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id4_3_cond_1_1) begin
        _tmp_645 <= 1;
      end 
      _ram_w4_l8192_id4_3_cond_2_2 <= _ram_w4_l8192_id4_3_cond_2_1;
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0)) begin
        ram_w4_l8192_id4_3_1_addr <= _tmp_156;
        ram_w4_l8192_id4_3_1_wdata <= _dataflow_slice_odata_38;
        ram_w4_l8192_id4_3_1_wenable <= _tmp_161 == 4;
      end 
      _ram_w4_l8192_id4_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16)) begin
        ram_w4_l8192_id4_3_0_addr <= _stream_conv2d_16_source_32_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id4_3_cond_1_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      _ram_w4_l8192_id4_3_cond_2_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      ram_w4_l8192_id4_3_0_wdata <= 0;
      ram_w4_l8192_id4_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id4_4_1_addr <= 0;
      ram_w4_l8192_id4_4_1_wdata <= 0;
      ram_w4_l8192_id4_4_1_wenable <= 0;
      _ram_w4_l8192_id4_4_cond_0_1 <= 0;
      ram_w4_l8192_id4_4_0_addr <= 0;
      _ram_w4_l8192_id4_4_cond_1_1 <= 0;
      _tmp_646 <= 0;
      _ram_w4_l8192_id4_4_cond_2_1 <= 0;
      _ram_w4_l8192_id4_4_cond_2_2 <= 0;
      ram_w4_l8192_id4_4_0_wdata <= 0;
      ram_w4_l8192_id4_4_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id4_4_cond_2_2) begin
        _tmp_646 <= 0;
      end 
      if(_ram_w4_l8192_id4_4_cond_0_1) begin
        ram_w4_l8192_id4_4_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id4_4_cond_1_1) begin
        _tmp_646 <= 1;
      end 
      _ram_w4_l8192_id4_4_cond_2_2 <= _ram_w4_l8192_id4_4_cond_2_1;
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0)) begin
        ram_w4_l8192_id4_4_1_addr <= _tmp_187;
        ram_w4_l8192_id4_4_1_wdata <= _dataflow_slice_odata_41;
        ram_w4_l8192_id4_4_1_wenable <= _tmp_192 == 4;
      end 
      _ram_w4_l8192_id4_4_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16)) begin
        ram_w4_l8192_id4_4_0_addr <= _stream_conv2d_16_source_32_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id4_4_cond_1_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      _ram_w4_l8192_id4_4_cond_2_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      ram_w4_l8192_id4_4_0_wdata <= 0;
      ram_w4_l8192_id4_4_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id4_5_1_addr <= 0;
      ram_w4_l8192_id4_5_1_wdata <= 0;
      ram_w4_l8192_id4_5_1_wenable <= 0;
      _ram_w4_l8192_id4_5_cond_0_1 <= 0;
      ram_w4_l8192_id4_5_0_addr <= 0;
      _ram_w4_l8192_id4_5_cond_1_1 <= 0;
      _tmp_647 <= 0;
      _ram_w4_l8192_id4_5_cond_2_1 <= 0;
      _ram_w4_l8192_id4_5_cond_2_2 <= 0;
      ram_w4_l8192_id4_5_0_wdata <= 0;
      ram_w4_l8192_id4_5_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id4_5_cond_2_2) begin
        _tmp_647 <= 0;
      end 
      if(_ram_w4_l8192_id4_5_cond_0_1) begin
        ram_w4_l8192_id4_5_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id4_5_cond_1_1) begin
        _tmp_647 <= 1;
      end 
      _ram_w4_l8192_id4_5_cond_2_2 <= _ram_w4_l8192_id4_5_cond_2_1;
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0)) begin
        ram_w4_l8192_id4_5_1_addr <= _tmp_218;
        ram_w4_l8192_id4_5_1_wdata <= _dataflow_slice_odata_44;
        ram_w4_l8192_id4_5_1_wenable <= _tmp_223 == 4;
      end 
      _ram_w4_l8192_id4_5_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16)) begin
        ram_w4_l8192_id4_5_0_addr <= _stream_conv2d_16_source_32_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id4_5_cond_1_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      _ram_w4_l8192_id4_5_cond_2_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      ram_w4_l8192_id4_5_0_wdata <= 0;
      ram_w4_l8192_id4_5_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id4_6_1_addr <= 0;
      ram_w4_l8192_id4_6_1_wdata <= 0;
      ram_w4_l8192_id4_6_1_wenable <= 0;
      _ram_w4_l8192_id4_6_cond_0_1 <= 0;
      ram_w4_l8192_id4_6_0_addr <= 0;
      _ram_w4_l8192_id4_6_cond_1_1 <= 0;
      _tmp_648 <= 0;
      _ram_w4_l8192_id4_6_cond_2_1 <= 0;
      _ram_w4_l8192_id4_6_cond_2_2 <= 0;
      ram_w4_l8192_id4_6_0_wdata <= 0;
      ram_w4_l8192_id4_6_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id4_6_cond_2_2) begin
        _tmp_648 <= 0;
      end 
      if(_ram_w4_l8192_id4_6_cond_0_1) begin
        ram_w4_l8192_id4_6_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id4_6_cond_1_1) begin
        _tmp_648 <= 1;
      end 
      _ram_w4_l8192_id4_6_cond_2_2 <= _ram_w4_l8192_id4_6_cond_2_1;
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0)) begin
        ram_w4_l8192_id4_6_1_addr <= _tmp_249;
        ram_w4_l8192_id4_6_1_wdata <= _dataflow_slice_odata_47;
        ram_w4_l8192_id4_6_1_wenable <= _tmp_254 == 4;
      end 
      _ram_w4_l8192_id4_6_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16)) begin
        ram_w4_l8192_id4_6_0_addr <= _stream_conv2d_16_source_32_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id4_6_cond_1_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      _ram_w4_l8192_id4_6_cond_2_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      ram_w4_l8192_id4_6_0_wdata <= 0;
      ram_w4_l8192_id4_6_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id4_7_1_addr <= 0;
      ram_w4_l8192_id4_7_1_wdata <= 0;
      ram_w4_l8192_id4_7_1_wenable <= 0;
      _ram_w4_l8192_id4_7_cond_0_1 <= 0;
      ram_w4_l8192_id4_7_0_addr <= 0;
      _ram_w4_l8192_id4_7_cond_1_1 <= 0;
      _tmp_649 <= 0;
      _ram_w4_l8192_id4_7_cond_2_1 <= 0;
      _ram_w4_l8192_id4_7_cond_2_2 <= 0;
      ram_w4_l8192_id4_7_0_wdata <= 0;
      ram_w4_l8192_id4_7_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id4_7_cond_2_2) begin
        _tmp_649 <= 0;
      end 
      if(_ram_w4_l8192_id4_7_cond_0_1) begin
        ram_w4_l8192_id4_7_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id4_7_cond_1_1) begin
        _tmp_649 <= 1;
      end 
      _ram_w4_l8192_id4_7_cond_2_2 <= _ram_w4_l8192_id4_7_cond_2_1;
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0)) begin
        ram_w4_l8192_id4_7_1_addr <= _tmp_280;
        ram_w4_l8192_id4_7_1_wdata <= _dataflow_slice_odata_50;
        ram_w4_l8192_id4_7_1_wenable <= _tmp_285 == 4;
      end 
      _ram_w4_l8192_id4_7_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16)) begin
        ram_w4_l8192_id4_7_0_addr <= _stream_conv2d_16_source_32_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id4_7_cond_1_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      _ram_w4_l8192_id4_7_cond_2_1 <= _stream_conv2d_16_source_32_source_ram_renable && (_stream_conv2d_16_source_32_source_ram_sel == 16);
      ram_w4_l8192_id4_7_0_wdata <= 0;
      ram_w4_l8192_id4_7_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id5_0_1_addr <= 0;
      ram_w4_l8192_id5_0_1_wdata <= 0;
      ram_w4_l8192_id5_0_1_wenable <= 0;
      _ram_w4_l8192_id5_0_cond_0_1 <= 0;
      ram_w4_l8192_id5_0_0_addr <= 0;
      _ram_w4_l8192_id5_0_cond_1_1 <= 0;
      _tmp_656 <= 0;
      _ram_w4_l8192_id5_0_cond_2_1 <= 0;
      _ram_w4_l8192_id5_0_cond_2_2 <= 0;
      ram_w4_l8192_id5_0_0_wdata <= 0;
      ram_w4_l8192_id5_0_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id5_0_cond_2_2) begin
        _tmp_656 <= 0;
      end 
      if(_ram_w4_l8192_id5_0_cond_0_1) begin
        ram_w4_l8192_id5_0_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id5_0_cond_1_1) begin
        _tmp_656 <= 1;
      end 
      _ram_w4_l8192_id5_0_cond_2_2 <= _ram_w4_l8192_id5_0_cond_2_1;
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0)) begin
        ram_w4_l8192_id5_0_1_addr <= _tmp_64;
        ram_w4_l8192_id5_0_1_wdata <= _dataflow_slice_odata_29;
        ram_w4_l8192_id5_0_1_wenable <= _tmp_68 == 5;
      end 
      _ram_w4_l8192_id5_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17)) begin
        ram_w4_l8192_id5_0_0_addr <= _stream_conv2d_16_source_33_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id5_0_cond_1_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      _ram_w4_l8192_id5_0_cond_2_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      ram_w4_l8192_id5_0_0_wdata <= 0;
      ram_w4_l8192_id5_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id5_1_1_addr <= 0;
      ram_w4_l8192_id5_1_1_wdata <= 0;
      ram_w4_l8192_id5_1_1_wenable <= 0;
      _ram_w4_l8192_id5_1_cond_0_1 <= 0;
      ram_w4_l8192_id5_1_0_addr <= 0;
      _ram_w4_l8192_id5_1_cond_1_1 <= 0;
      _tmp_657 <= 0;
      _ram_w4_l8192_id5_1_cond_2_1 <= 0;
      _ram_w4_l8192_id5_1_cond_2_2 <= 0;
      ram_w4_l8192_id5_1_0_wdata <= 0;
      ram_w4_l8192_id5_1_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id5_1_cond_2_2) begin
        _tmp_657 <= 0;
      end 
      if(_ram_w4_l8192_id5_1_cond_0_1) begin
        ram_w4_l8192_id5_1_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id5_1_cond_1_1) begin
        _tmp_657 <= 1;
      end 
      _ram_w4_l8192_id5_1_cond_2_2 <= _ram_w4_l8192_id5_1_cond_2_1;
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0)) begin
        ram_w4_l8192_id5_1_1_addr <= _tmp_95;
        ram_w4_l8192_id5_1_1_wdata <= _dataflow_slice_odata_32;
        ram_w4_l8192_id5_1_1_wenable <= _tmp_99 == 5;
      end 
      _ram_w4_l8192_id5_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17)) begin
        ram_w4_l8192_id5_1_0_addr <= _stream_conv2d_16_source_33_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id5_1_cond_1_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      _ram_w4_l8192_id5_1_cond_2_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      ram_w4_l8192_id5_1_0_wdata <= 0;
      ram_w4_l8192_id5_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id5_2_1_addr <= 0;
      ram_w4_l8192_id5_2_1_wdata <= 0;
      ram_w4_l8192_id5_2_1_wenable <= 0;
      _ram_w4_l8192_id5_2_cond_0_1 <= 0;
      ram_w4_l8192_id5_2_0_addr <= 0;
      _ram_w4_l8192_id5_2_cond_1_1 <= 0;
      _tmp_658 <= 0;
      _ram_w4_l8192_id5_2_cond_2_1 <= 0;
      _ram_w4_l8192_id5_2_cond_2_2 <= 0;
      ram_w4_l8192_id5_2_0_wdata <= 0;
      ram_w4_l8192_id5_2_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id5_2_cond_2_2) begin
        _tmp_658 <= 0;
      end 
      if(_ram_w4_l8192_id5_2_cond_0_1) begin
        ram_w4_l8192_id5_2_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id5_2_cond_1_1) begin
        _tmp_658 <= 1;
      end 
      _ram_w4_l8192_id5_2_cond_2_2 <= _ram_w4_l8192_id5_2_cond_2_1;
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0)) begin
        ram_w4_l8192_id5_2_1_addr <= _tmp_126;
        ram_w4_l8192_id5_2_1_wdata <= _dataflow_slice_odata_35;
        ram_w4_l8192_id5_2_1_wenable <= _tmp_130 == 5;
      end 
      _ram_w4_l8192_id5_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17)) begin
        ram_w4_l8192_id5_2_0_addr <= _stream_conv2d_16_source_33_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id5_2_cond_1_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      _ram_w4_l8192_id5_2_cond_2_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      ram_w4_l8192_id5_2_0_wdata <= 0;
      ram_w4_l8192_id5_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id5_3_1_addr <= 0;
      ram_w4_l8192_id5_3_1_wdata <= 0;
      ram_w4_l8192_id5_3_1_wenable <= 0;
      _ram_w4_l8192_id5_3_cond_0_1 <= 0;
      ram_w4_l8192_id5_3_0_addr <= 0;
      _ram_w4_l8192_id5_3_cond_1_1 <= 0;
      _tmp_659 <= 0;
      _ram_w4_l8192_id5_3_cond_2_1 <= 0;
      _ram_w4_l8192_id5_3_cond_2_2 <= 0;
      ram_w4_l8192_id5_3_0_wdata <= 0;
      ram_w4_l8192_id5_3_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id5_3_cond_2_2) begin
        _tmp_659 <= 0;
      end 
      if(_ram_w4_l8192_id5_3_cond_0_1) begin
        ram_w4_l8192_id5_3_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id5_3_cond_1_1) begin
        _tmp_659 <= 1;
      end 
      _ram_w4_l8192_id5_3_cond_2_2 <= _ram_w4_l8192_id5_3_cond_2_1;
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0)) begin
        ram_w4_l8192_id5_3_1_addr <= _tmp_157;
        ram_w4_l8192_id5_3_1_wdata <= _dataflow_slice_odata_38;
        ram_w4_l8192_id5_3_1_wenable <= _tmp_161 == 5;
      end 
      _ram_w4_l8192_id5_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17)) begin
        ram_w4_l8192_id5_3_0_addr <= _stream_conv2d_16_source_33_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id5_3_cond_1_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      _ram_w4_l8192_id5_3_cond_2_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      ram_w4_l8192_id5_3_0_wdata <= 0;
      ram_w4_l8192_id5_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id5_4_1_addr <= 0;
      ram_w4_l8192_id5_4_1_wdata <= 0;
      ram_w4_l8192_id5_4_1_wenable <= 0;
      _ram_w4_l8192_id5_4_cond_0_1 <= 0;
      ram_w4_l8192_id5_4_0_addr <= 0;
      _ram_w4_l8192_id5_4_cond_1_1 <= 0;
      _tmp_660 <= 0;
      _ram_w4_l8192_id5_4_cond_2_1 <= 0;
      _ram_w4_l8192_id5_4_cond_2_2 <= 0;
      ram_w4_l8192_id5_4_0_wdata <= 0;
      ram_w4_l8192_id5_4_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id5_4_cond_2_2) begin
        _tmp_660 <= 0;
      end 
      if(_ram_w4_l8192_id5_4_cond_0_1) begin
        ram_w4_l8192_id5_4_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id5_4_cond_1_1) begin
        _tmp_660 <= 1;
      end 
      _ram_w4_l8192_id5_4_cond_2_2 <= _ram_w4_l8192_id5_4_cond_2_1;
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0)) begin
        ram_w4_l8192_id5_4_1_addr <= _tmp_188;
        ram_w4_l8192_id5_4_1_wdata <= _dataflow_slice_odata_41;
        ram_w4_l8192_id5_4_1_wenable <= _tmp_192 == 5;
      end 
      _ram_w4_l8192_id5_4_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17)) begin
        ram_w4_l8192_id5_4_0_addr <= _stream_conv2d_16_source_33_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id5_4_cond_1_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      _ram_w4_l8192_id5_4_cond_2_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      ram_w4_l8192_id5_4_0_wdata <= 0;
      ram_w4_l8192_id5_4_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id5_5_1_addr <= 0;
      ram_w4_l8192_id5_5_1_wdata <= 0;
      ram_w4_l8192_id5_5_1_wenable <= 0;
      _ram_w4_l8192_id5_5_cond_0_1 <= 0;
      ram_w4_l8192_id5_5_0_addr <= 0;
      _ram_w4_l8192_id5_5_cond_1_1 <= 0;
      _tmp_661 <= 0;
      _ram_w4_l8192_id5_5_cond_2_1 <= 0;
      _ram_w4_l8192_id5_5_cond_2_2 <= 0;
      ram_w4_l8192_id5_5_0_wdata <= 0;
      ram_w4_l8192_id5_5_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id5_5_cond_2_2) begin
        _tmp_661 <= 0;
      end 
      if(_ram_w4_l8192_id5_5_cond_0_1) begin
        ram_w4_l8192_id5_5_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id5_5_cond_1_1) begin
        _tmp_661 <= 1;
      end 
      _ram_w4_l8192_id5_5_cond_2_2 <= _ram_w4_l8192_id5_5_cond_2_1;
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0)) begin
        ram_w4_l8192_id5_5_1_addr <= _tmp_219;
        ram_w4_l8192_id5_5_1_wdata <= _dataflow_slice_odata_44;
        ram_w4_l8192_id5_5_1_wenable <= _tmp_223 == 5;
      end 
      _ram_w4_l8192_id5_5_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17)) begin
        ram_w4_l8192_id5_5_0_addr <= _stream_conv2d_16_source_33_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id5_5_cond_1_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      _ram_w4_l8192_id5_5_cond_2_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      ram_w4_l8192_id5_5_0_wdata <= 0;
      ram_w4_l8192_id5_5_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id5_6_1_addr <= 0;
      ram_w4_l8192_id5_6_1_wdata <= 0;
      ram_w4_l8192_id5_6_1_wenable <= 0;
      _ram_w4_l8192_id5_6_cond_0_1 <= 0;
      ram_w4_l8192_id5_6_0_addr <= 0;
      _ram_w4_l8192_id5_6_cond_1_1 <= 0;
      _tmp_662 <= 0;
      _ram_w4_l8192_id5_6_cond_2_1 <= 0;
      _ram_w4_l8192_id5_6_cond_2_2 <= 0;
      ram_w4_l8192_id5_6_0_wdata <= 0;
      ram_w4_l8192_id5_6_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id5_6_cond_2_2) begin
        _tmp_662 <= 0;
      end 
      if(_ram_w4_l8192_id5_6_cond_0_1) begin
        ram_w4_l8192_id5_6_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id5_6_cond_1_1) begin
        _tmp_662 <= 1;
      end 
      _ram_w4_l8192_id5_6_cond_2_2 <= _ram_w4_l8192_id5_6_cond_2_1;
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0)) begin
        ram_w4_l8192_id5_6_1_addr <= _tmp_250;
        ram_w4_l8192_id5_6_1_wdata <= _dataflow_slice_odata_47;
        ram_w4_l8192_id5_6_1_wenable <= _tmp_254 == 5;
      end 
      _ram_w4_l8192_id5_6_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17)) begin
        ram_w4_l8192_id5_6_0_addr <= _stream_conv2d_16_source_33_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id5_6_cond_1_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      _ram_w4_l8192_id5_6_cond_2_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      ram_w4_l8192_id5_6_0_wdata <= 0;
      ram_w4_l8192_id5_6_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id5_7_1_addr <= 0;
      ram_w4_l8192_id5_7_1_wdata <= 0;
      ram_w4_l8192_id5_7_1_wenable <= 0;
      _ram_w4_l8192_id5_7_cond_0_1 <= 0;
      ram_w4_l8192_id5_7_0_addr <= 0;
      _ram_w4_l8192_id5_7_cond_1_1 <= 0;
      _tmp_663 <= 0;
      _ram_w4_l8192_id5_7_cond_2_1 <= 0;
      _ram_w4_l8192_id5_7_cond_2_2 <= 0;
      ram_w4_l8192_id5_7_0_wdata <= 0;
      ram_w4_l8192_id5_7_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id5_7_cond_2_2) begin
        _tmp_663 <= 0;
      end 
      if(_ram_w4_l8192_id5_7_cond_0_1) begin
        ram_w4_l8192_id5_7_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id5_7_cond_1_1) begin
        _tmp_663 <= 1;
      end 
      _ram_w4_l8192_id5_7_cond_2_2 <= _ram_w4_l8192_id5_7_cond_2_1;
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0)) begin
        ram_w4_l8192_id5_7_1_addr <= _tmp_281;
        ram_w4_l8192_id5_7_1_wdata <= _dataflow_slice_odata_50;
        ram_w4_l8192_id5_7_1_wenable <= _tmp_285 == 5;
      end 
      _ram_w4_l8192_id5_7_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17)) begin
        ram_w4_l8192_id5_7_0_addr <= _stream_conv2d_16_source_33_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id5_7_cond_1_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      _ram_w4_l8192_id5_7_cond_2_1 <= _stream_conv2d_16_source_33_source_ram_renable && (_stream_conv2d_16_source_33_source_ram_sel == 17);
      ram_w4_l8192_id5_7_0_wdata <= 0;
      ram_w4_l8192_id5_7_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id6_0_1_addr <= 0;
      ram_w4_l8192_id6_0_1_wdata <= 0;
      ram_w4_l8192_id6_0_1_wenable <= 0;
      _ram_w4_l8192_id6_0_cond_0_1 <= 0;
      ram_w4_l8192_id6_0_0_addr <= 0;
      _ram_w4_l8192_id6_0_cond_1_1 <= 0;
      _tmp_670 <= 0;
      _ram_w4_l8192_id6_0_cond_2_1 <= 0;
      _ram_w4_l8192_id6_0_cond_2_2 <= 0;
      ram_w4_l8192_id6_0_0_wdata <= 0;
      ram_w4_l8192_id6_0_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id6_0_cond_2_2) begin
        _tmp_670 <= 0;
      end 
      if(_ram_w4_l8192_id6_0_cond_0_1) begin
        ram_w4_l8192_id6_0_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id6_0_cond_1_1) begin
        _tmp_670 <= 1;
      end 
      _ram_w4_l8192_id6_0_cond_2_2 <= _ram_w4_l8192_id6_0_cond_2_1;
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0)) begin
        ram_w4_l8192_id6_0_1_addr <= _tmp_65;
        ram_w4_l8192_id6_0_1_wdata <= _dataflow_slice_odata_29;
        ram_w4_l8192_id6_0_1_wenable <= _tmp_68 == 6;
      end 
      _ram_w4_l8192_id6_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18)) begin
        ram_w4_l8192_id6_0_0_addr <= _stream_conv2d_16_source_34_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id6_0_cond_1_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      _ram_w4_l8192_id6_0_cond_2_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      ram_w4_l8192_id6_0_0_wdata <= 0;
      ram_w4_l8192_id6_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id6_1_1_addr <= 0;
      ram_w4_l8192_id6_1_1_wdata <= 0;
      ram_w4_l8192_id6_1_1_wenable <= 0;
      _ram_w4_l8192_id6_1_cond_0_1 <= 0;
      ram_w4_l8192_id6_1_0_addr <= 0;
      _ram_w4_l8192_id6_1_cond_1_1 <= 0;
      _tmp_671 <= 0;
      _ram_w4_l8192_id6_1_cond_2_1 <= 0;
      _ram_w4_l8192_id6_1_cond_2_2 <= 0;
      ram_w4_l8192_id6_1_0_wdata <= 0;
      ram_w4_l8192_id6_1_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id6_1_cond_2_2) begin
        _tmp_671 <= 0;
      end 
      if(_ram_w4_l8192_id6_1_cond_0_1) begin
        ram_w4_l8192_id6_1_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id6_1_cond_1_1) begin
        _tmp_671 <= 1;
      end 
      _ram_w4_l8192_id6_1_cond_2_2 <= _ram_w4_l8192_id6_1_cond_2_1;
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0)) begin
        ram_w4_l8192_id6_1_1_addr <= _tmp_96;
        ram_w4_l8192_id6_1_1_wdata <= _dataflow_slice_odata_32;
        ram_w4_l8192_id6_1_1_wenable <= _tmp_99 == 6;
      end 
      _ram_w4_l8192_id6_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18)) begin
        ram_w4_l8192_id6_1_0_addr <= _stream_conv2d_16_source_34_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id6_1_cond_1_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      _ram_w4_l8192_id6_1_cond_2_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      ram_w4_l8192_id6_1_0_wdata <= 0;
      ram_w4_l8192_id6_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id6_2_1_addr <= 0;
      ram_w4_l8192_id6_2_1_wdata <= 0;
      ram_w4_l8192_id6_2_1_wenable <= 0;
      _ram_w4_l8192_id6_2_cond_0_1 <= 0;
      ram_w4_l8192_id6_2_0_addr <= 0;
      _ram_w4_l8192_id6_2_cond_1_1 <= 0;
      _tmp_672 <= 0;
      _ram_w4_l8192_id6_2_cond_2_1 <= 0;
      _ram_w4_l8192_id6_2_cond_2_2 <= 0;
      ram_w4_l8192_id6_2_0_wdata <= 0;
      ram_w4_l8192_id6_2_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id6_2_cond_2_2) begin
        _tmp_672 <= 0;
      end 
      if(_ram_w4_l8192_id6_2_cond_0_1) begin
        ram_w4_l8192_id6_2_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id6_2_cond_1_1) begin
        _tmp_672 <= 1;
      end 
      _ram_w4_l8192_id6_2_cond_2_2 <= _ram_w4_l8192_id6_2_cond_2_1;
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0)) begin
        ram_w4_l8192_id6_2_1_addr <= _tmp_127;
        ram_w4_l8192_id6_2_1_wdata <= _dataflow_slice_odata_35;
        ram_w4_l8192_id6_2_1_wenable <= _tmp_130 == 6;
      end 
      _ram_w4_l8192_id6_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18)) begin
        ram_w4_l8192_id6_2_0_addr <= _stream_conv2d_16_source_34_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id6_2_cond_1_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      _ram_w4_l8192_id6_2_cond_2_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      ram_w4_l8192_id6_2_0_wdata <= 0;
      ram_w4_l8192_id6_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id6_3_1_addr <= 0;
      ram_w4_l8192_id6_3_1_wdata <= 0;
      ram_w4_l8192_id6_3_1_wenable <= 0;
      _ram_w4_l8192_id6_3_cond_0_1 <= 0;
      ram_w4_l8192_id6_3_0_addr <= 0;
      _ram_w4_l8192_id6_3_cond_1_1 <= 0;
      _tmp_673 <= 0;
      _ram_w4_l8192_id6_3_cond_2_1 <= 0;
      _ram_w4_l8192_id6_3_cond_2_2 <= 0;
      ram_w4_l8192_id6_3_0_wdata <= 0;
      ram_w4_l8192_id6_3_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id6_3_cond_2_2) begin
        _tmp_673 <= 0;
      end 
      if(_ram_w4_l8192_id6_3_cond_0_1) begin
        ram_w4_l8192_id6_3_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id6_3_cond_1_1) begin
        _tmp_673 <= 1;
      end 
      _ram_w4_l8192_id6_3_cond_2_2 <= _ram_w4_l8192_id6_3_cond_2_1;
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0)) begin
        ram_w4_l8192_id6_3_1_addr <= _tmp_158;
        ram_w4_l8192_id6_3_1_wdata <= _dataflow_slice_odata_38;
        ram_w4_l8192_id6_3_1_wenable <= _tmp_161 == 6;
      end 
      _ram_w4_l8192_id6_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18)) begin
        ram_w4_l8192_id6_3_0_addr <= _stream_conv2d_16_source_34_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id6_3_cond_1_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      _ram_w4_l8192_id6_3_cond_2_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      ram_w4_l8192_id6_3_0_wdata <= 0;
      ram_w4_l8192_id6_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id6_4_1_addr <= 0;
      ram_w4_l8192_id6_4_1_wdata <= 0;
      ram_w4_l8192_id6_4_1_wenable <= 0;
      _ram_w4_l8192_id6_4_cond_0_1 <= 0;
      ram_w4_l8192_id6_4_0_addr <= 0;
      _ram_w4_l8192_id6_4_cond_1_1 <= 0;
      _tmp_674 <= 0;
      _ram_w4_l8192_id6_4_cond_2_1 <= 0;
      _ram_w4_l8192_id6_4_cond_2_2 <= 0;
      ram_w4_l8192_id6_4_0_wdata <= 0;
      ram_w4_l8192_id6_4_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id6_4_cond_2_2) begin
        _tmp_674 <= 0;
      end 
      if(_ram_w4_l8192_id6_4_cond_0_1) begin
        ram_w4_l8192_id6_4_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id6_4_cond_1_1) begin
        _tmp_674 <= 1;
      end 
      _ram_w4_l8192_id6_4_cond_2_2 <= _ram_w4_l8192_id6_4_cond_2_1;
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0)) begin
        ram_w4_l8192_id6_4_1_addr <= _tmp_189;
        ram_w4_l8192_id6_4_1_wdata <= _dataflow_slice_odata_41;
        ram_w4_l8192_id6_4_1_wenable <= _tmp_192 == 6;
      end 
      _ram_w4_l8192_id6_4_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18)) begin
        ram_w4_l8192_id6_4_0_addr <= _stream_conv2d_16_source_34_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id6_4_cond_1_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      _ram_w4_l8192_id6_4_cond_2_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      ram_w4_l8192_id6_4_0_wdata <= 0;
      ram_w4_l8192_id6_4_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id6_5_1_addr <= 0;
      ram_w4_l8192_id6_5_1_wdata <= 0;
      ram_w4_l8192_id6_5_1_wenable <= 0;
      _ram_w4_l8192_id6_5_cond_0_1 <= 0;
      ram_w4_l8192_id6_5_0_addr <= 0;
      _ram_w4_l8192_id6_5_cond_1_1 <= 0;
      _tmp_675 <= 0;
      _ram_w4_l8192_id6_5_cond_2_1 <= 0;
      _ram_w4_l8192_id6_5_cond_2_2 <= 0;
      ram_w4_l8192_id6_5_0_wdata <= 0;
      ram_w4_l8192_id6_5_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id6_5_cond_2_2) begin
        _tmp_675 <= 0;
      end 
      if(_ram_w4_l8192_id6_5_cond_0_1) begin
        ram_w4_l8192_id6_5_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id6_5_cond_1_1) begin
        _tmp_675 <= 1;
      end 
      _ram_w4_l8192_id6_5_cond_2_2 <= _ram_w4_l8192_id6_5_cond_2_1;
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0)) begin
        ram_w4_l8192_id6_5_1_addr <= _tmp_220;
        ram_w4_l8192_id6_5_1_wdata <= _dataflow_slice_odata_44;
        ram_w4_l8192_id6_5_1_wenable <= _tmp_223 == 6;
      end 
      _ram_w4_l8192_id6_5_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18)) begin
        ram_w4_l8192_id6_5_0_addr <= _stream_conv2d_16_source_34_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id6_5_cond_1_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      _ram_w4_l8192_id6_5_cond_2_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      ram_w4_l8192_id6_5_0_wdata <= 0;
      ram_w4_l8192_id6_5_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id6_6_1_addr <= 0;
      ram_w4_l8192_id6_6_1_wdata <= 0;
      ram_w4_l8192_id6_6_1_wenable <= 0;
      _ram_w4_l8192_id6_6_cond_0_1 <= 0;
      ram_w4_l8192_id6_6_0_addr <= 0;
      _ram_w4_l8192_id6_6_cond_1_1 <= 0;
      _tmp_676 <= 0;
      _ram_w4_l8192_id6_6_cond_2_1 <= 0;
      _ram_w4_l8192_id6_6_cond_2_2 <= 0;
      ram_w4_l8192_id6_6_0_wdata <= 0;
      ram_w4_l8192_id6_6_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id6_6_cond_2_2) begin
        _tmp_676 <= 0;
      end 
      if(_ram_w4_l8192_id6_6_cond_0_1) begin
        ram_w4_l8192_id6_6_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id6_6_cond_1_1) begin
        _tmp_676 <= 1;
      end 
      _ram_w4_l8192_id6_6_cond_2_2 <= _ram_w4_l8192_id6_6_cond_2_1;
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0)) begin
        ram_w4_l8192_id6_6_1_addr <= _tmp_251;
        ram_w4_l8192_id6_6_1_wdata <= _dataflow_slice_odata_47;
        ram_w4_l8192_id6_6_1_wenable <= _tmp_254 == 6;
      end 
      _ram_w4_l8192_id6_6_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18)) begin
        ram_w4_l8192_id6_6_0_addr <= _stream_conv2d_16_source_34_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id6_6_cond_1_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      _ram_w4_l8192_id6_6_cond_2_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      ram_w4_l8192_id6_6_0_wdata <= 0;
      ram_w4_l8192_id6_6_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id6_7_1_addr <= 0;
      ram_w4_l8192_id6_7_1_wdata <= 0;
      ram_w4_l8192_id6_7_1_wenable <= 0;
      _ram_w4_l8192_id6_7_cond_0_1 <= 0;
      ram_w4_l8192_id6_7_0_addr <= 0;
      _ram_w4_l8192_id6_7_cond_1_1 <= 0;
      _tmp_677 <= 0;
      _ram_w4_l8192_id6_7_cond_2_1 <= 0;
      _ram_w4_l8192_id6_7_cond_2_2 <= 0;
      ram_w4_l8192_id6_7_0_wdata <= 0;
      ram_w4_l8192_id6_7_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id6_7_cond_2_2) begin
        _tmp_677 <= 0;
      end 
      if(_ram_w4_l8192_id6_7_cond_0_1) begin
        ram_w4_l8192_id6_7_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id6_7_cond_1_1) begin
        _tmp_677 <= 1;
      end 
      _ram_w4_l8192_id6_7_cond_2_2 <= _ram_w4_l8192_id6_7_cond_2_1;
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0)) begin
        ram_w4_l8192_id6_7_1_addr <= _tmp_282;
        ram_w4_l8192_id6_7_1_wdata <= _dataflow_slice_odata_50;
        ram_w4_l8192_id6_7_1_wenable <= _tmp_285 == 6;
      end 
      _ram_w4_l8192_id6_7_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18)) begin
        ram_w4_l8192_id6_7_0_addr <= _stream_conv2d_16_source_34_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id6_7_cond_1_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      _ram_w4_l8192_id6_7_cond_2_1 <= _stream_conv2d_16_source_34_source_ram_renable && (_stream_conv2d_16_source_34_source_ram_sel == 18);
      ram_w4_l8192_id6_7_0_wdata <= 0;
      ram_w4_l8192_id6_7_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id7_0_1_addr <= 0;
      ram_w4_l8192_id7_0_1_wdata <= 0;
      ram_w4_l8192_id7_0_1_wenable <= 0;
      _ram_w4_l8192_id7_0_cond_0_1 <= 0;
      ram_w4_l8192_id7_0_0_addr <= 0;
      _ram_w4_l8192_id7_0_cond_1_1 <= 0;
      _tmp_684 <= 0;
      _ram_w4_l8192_id7_0_cond_2_1 <= 0;
      _ram_w4_l8192_id7_0_cond_2_2 <= 0;
      ram_w4_l8192_id7_0_0_wdata <= 0;
      ram_w4_l8192_id7_0_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id7_0_cond_2_2) begin
        _tmp_684 <= 0;
      end 
      if(_ram_w4_l8192_id7_0_cond_0_1) begin
        ram_w4_l8192_id7_0_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id7_0_cond_1_1) begin
        _tmp_684 <= 1;
      end 
      _ram_w4_l8192_id7_0_cond_2_2 <= _ram_w4_l8192_id7_0_cond_2_1;
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0)) begin
        ram_w4_l8192_id7_0_1_addr <= _tmp_66;
        ram_w4_l8192_id7_0_1_wdata <= _dataflow_slice_odata_29;
        ram_w4_l8192_id7_0_1_wenable <= _tmp_68 == 7;
      end 
      _ram_w4_l8192_id7_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19)) begin
        ram_w4_l8192_id7_0_0_addr <= _stream_conv2d_16_source_35_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id7_0_cond_1_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      _ram_w4_l8192_id7_0_cond_2_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      ram_w4_l8192_id7_0_0_wdata <= 0;
      ram_w4_l8192_id7_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id7_1_1_addr <= 0;
      ram_w4_l8192_id7_1_1_wdata <= 0;
      ram_w4_l8192_id7_1_1_wenable <= 0;
      _ram_w4_l8192_id7_1_cond_0_1 <= 0;
      ram_w4_l8192_id7_1_0_addr <= 0;
      _ram_w4_l8192_id7_1_cond_1_1 <= 0;
      _tmp_685 <= 0;
      _ram_w4_l8192_id7_1_cond_2_1 <= 0;
      _ram_w4_l8192_id7_1_cond_2_2 <= 0;
      ram_w4_l8192_id7_1_0_wdata <= 0;
      ram_w4_l8192_id7_1_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id7_1_cond_2_2) begin
        _tmp_685 <= 0;
      end 
      if(_ram_w4_l8192_id7_1_cond_0_1) begin
        ram_w4_l8192_id7_1_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id7_1_cond_1_1) begin
        _tmp_685 <= 1;
      end 
      _ram_w4_l8192_id7_1_cond_2_2 <= _ram_w4_l8192_id7_1_cond_2_1;
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0)) begin
        ram_w4_l8192_id7_1_1_addr <= _tmp_97;
        ram_w4_l8192_id7_1_1_wdata <= _dataflow_slice_odata_32;
        ram_w4_l8192_id7_1_1_wenable <= _tmp_99 == 7;
      end 
      _ram_w4_l8192_id7_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19)) begin
        ram_w4_l8192_id7_1_0_addr <= _stream_conv2d_16_source_35_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id7_1_cond_1_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      _ram_w4_l8192_id7_1_cond_2_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      ram_w4_l8192_id7_1_0_wdata <= 0;
      ram_w4_l8192_id7_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id7_2_1_addr <= 0;
      ram_w4_l8192_id7_2_1_wdata <= 0;
      ram_w4_l8192_id7_2_1_wenable <= 0;
      _ram_w4_l8192_id7_2_cond_0_1 <= 0;
      ram_w4_l8192_id7_2_0_addr <= 0;
      _ram_w4_l8192_id7_2_cond_1_1 <= 0;
      _tmp_686 <= 0;
      _ram_w4_l8192_id7_2_cond_2_1 <= 0;
      _ram_w4_l8192_id7_2_cond_2_2 <= 0;
      ram_w4_l8192_id7_2_0_wdata <= 0;
      ram_w4_l8192_id7_2_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id7_2_cond_2_2) begin
        _tmp_686 <= 0;
      end 
      if(_ram_w4_l8192_id7_2_cond_0_1) begin
        ram_w4_l8192_id7_2_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id7_2_cond_1_1) begin
        _tmp_686 <= 1;
      end 
      _ram_w4_l8192_id7_2_cond_2_2 <= _ram_w4_l8192_id7_2_cond_2_1;
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0)) begin
        ram_w4_l8192_id7_2_1_addr <= _tmp_128;
        ram_w4_l8192_id7_2_1_wdata <= _dataflow_slice_odata_35;
        ram_w4_l8192_id7_2_1_wenable <= _tmp_130 == 7;
      end 
      _ram_w4_l8192_id7_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19)) begin
        ram_w4_l8192_id7_2_0_addr <= _stream_conv2d_16_source_35_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id7_2_cond_1_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      _ram_w4_l8192_id7_2_cond_2_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      ram_w4_l8192_id7_2_0_wdata <= 0;
      ram_w4_l8192_id7_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id7_3_1_addr <= 0;
      ram_w4_l8192_id7_3_1_wdata <= 0;
      ram_w4_l8192_id7_3_1_wenable <= 0;
      _ram_w4_l8192_id7_3_cond_0_1 <= 0;
      ram_w4_l8192_id7_3_0_addr <= 0;
      _ram_w4_l8192_id7_3_cond_1_1 <= 0;
      _tmp_687 <= 0;
      _ram_w4_l8192_id7_3_cond_2_1 <= 0;
      _ram_w4_l8192_id7_3_cond_2_2 <= 0;
      ram_w4_l8192_id7_3_0_wdata <= 0;
      ram_w4_l8192_id7_3_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id7_3_cond_2_2) begin
        _tmp_687 <= 0;
      end 
      if(_ram_w4_l8192_id7_3_cond_0_1) begin
        ram_w4_l8192_id7_3_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id7_3_cond_1_1) begin
        _tmp_687 <= 1;
      end 
      _ram_w4_l8192_id7_3_cond_2_2 <= _ram_w4_l8192_id7_3_cond_2_1;
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0)) begin
        ram_w4_l8192_id7_3_1_addr <= _tmp_159;
        ram_w4_l8192_id7_3_1_wdata <= _dataflow_slice_odata_38;
        ram_w4_l8192_id7_3_1_wenable <= _tmp_161 == 7;
      end 
      _ram_w4_l8192_id7_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19)) begin
        ram_w4_l8192_id7_3_0_addr <= _stream_conv2d_16_source_35_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id7_3_cond_1_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      _ram_w4_l8192_id7_3_cond_2_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      ram_w4_l8192_id7_3_0_wdata <= 0;
      ram_w4_l8192_id7_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id7_4_1_addr <= 0;
      ram_w4_l8192_id7_4_1_wdata <= 0;
      ram_w4_l8192_id7_4_1_wenable <= 0;
      _ram_w4_l8192_id7_4_cond_0_1 <= 0;
      ram_w4_l8192_id7_4_0_addr <= 0;
      _ram_w4_l8192_id7_4_cond_1_1 <= 0;
      _tmp_688 <= 0;
      _ram_w4_l8192_id7_4_cond_2_1 <= 0;
      _ram_w4_l8192_id7_4_cond_2_2 <= 0;
      ram_w4_l8192_id7_4_0_wdata <= 0;
      ram_w4_l8192_id7_4_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id7_4_cond_2_2) begin
        _tmp_688 <= 0;
      end 
      if(_ram_w4_l8192_id7_4_cond_0_1) begin
        ram_w4_l8192_id7_4_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id7_4_cond_1_1) begin
        _tmp_688 <= 1;
      end 
      _ram_w4_l8192_id7_4_cond_2_2 <= _ram_w4_l8192_id7_4_cond_2_1;
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0)) begin
        ram_w4_l8192_id7_4_1_addr <= _tmp_190;
        ram_w4_l8192_id7_4_1_wdata <= _dataflow_slice_odata_41;
        ram_w4_l8192_id7_4_1_wenable <= _tmp_192 == 7;
      end 
      _ram_w4_l8192_id7_4_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19)) begin
        ram_w4_l8192_id7_4_0_addr <= _stream_conv2d_16_source_35_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id7_4_cond_1_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      _ram_w4_l8192_id7_4_cond_2_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      ram_w4_l8192_id7_4_0_wdata <= 0;
      ram_w4_l8192_id7_4_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id7_5_1_addr <= 0;
      ram_w4_l8192_id7_5_1_wdata <= 0;
      ram_w4_l8192_id7_5_1_wenable <= 0;
      _ram_w4_l8192_id7_5_cond_0_1 <= 0;
      ram_w4_l8192_id7_5_0_addr <= 0;
      _ram_w4_l8192_id7_5_cond_1_1 <= 0;
      _tmp_689 <= 0;
      _ram_w4_l8192_id7_5_cond_2_1 <= 0;
      _ram_w4_l8192_id7_5_cond_2_2 <= 0;
      ram_w4_l8192_id7_5_0_wdata <= 0;
      ram_w4_l8192_id7_5_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id7_5_cond_2_2) begin
        _tmp_689 <= 0;
      end 
      if(_ram_w4_l8192_id7_5_cond_0_1) begin
        ram_w4_l8192_id7_5_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id7_5_cond_1_1) begin
        _tmp_689 <= 1;
      end 
      _ram_w4_l8192_id7_5_cond_2_2 <= _ram_w4_l8192_id7_5_cond_2_1;
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0)) begin
        ram_w4_l8192_id7_5_1_addr <= _tmp_221;
        ram_w4_l8192_id7_5_1_wdata <= _dataflow_slice_odata_44;
        ram_w4_l8192_id7_5_1_wenable <= _tmp_223 == 7;
      end 
      _ram_w4_l8192_id7_5_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19)) begin
        ram_w4_l8192_id7_5_0_addr <= _stream_conv2d_16_source_35_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id7_5_cond_1_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      _ram_w4_l8192_id7_5_cond_2_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      ram_w4_l8192_id7_5_0_wdata <= 0;
      ram_w4_l8192_id7_5_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id7_6_1_addr <= 0;
      ram_w4_l8192_id7_6_1_wdata <= 0;
      ram_w4_l8192_id7_6_1_wenable <= 0;
      _ram_w4_l8192_id7_6_cond_0_1 <= 0;
      ram_w4_l8192_id7_6_0_addr <= 0;
      _ram_w4_l8192_id7_6_cond_1_1 <= 0;
      _tmp_690 <= 0;
      _ram_w4_l8192_id7_6_cond_2_1 <= 0;
      _ram_w4_l8192_id7_6_cond_2_2 <= 0;
      ram_w4_l8192_id7_6_0_wdata <= 0;
      ram_w4_l8192_id7_6_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id7_6_cond_2_2) begin
        _tmp_690 <= 0;
      end 
      if(_ram_w4_l8192_id7_6_cond_0_1) begin
        ram_w4_l8192_id7_6_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id7_6_cond_1_1) begin
        _tmp_690 <= 1;
      end 
      _ram_w4_l8192_id7_6_cond_2_2 <= _ram_w4_l8192_id7_6_cond_2_1;
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0)) begin
        ram_w4_l8192_id7_6_1_addr <= _tmp_252;
        ram_w4_l8192_id7_6_1_wdata <= _dataflow_slice_odata_47;
        ram_w4_l8192_id7_6_1_wenable <= _tmp_254 == 7;
      end 
      _ram_w4_l8192_id7_6_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19)) begin
        ram_w4_l8192_id7_6_0_addr <= _stream_conv2d_16_source_35_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id7_6_cond_1_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      _ram_w4_l8192_id7_6_cond_2_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      ram_w4_l8192_id7_6_0_wdata <= 0;
      ram_w4_l8192_id7_6_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id7_7_1_addr <= 0;
      ram_w4_l8192_id7_7_1_wdata <= 0;
      ram_w4_l8192_id7_7_1_wenable <= 0;
      _ram_w4_l8192_id7_7_cond_0_1 <= 0;
      ram_w4_l8192_id7_7_0_addr <= 0;
      _ram_w4_l8192_id7_7_cond_1_1 <= 0;
      _tmp_691 <= 0;
      _ram_w4_l8192_id7_7_cond_2_1 <= 0;
      _ram_w4_l8192_id7_7_cond_2_2 <= 0;
      ram_w4_l8192_id7_7_0_wdata <= 0;
      ram_w4_l8192_id7_7_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id7_7_cond_2_2) begin
        _tmp_691 <= 0;
      end 
      if(_ram_w4_l8192_id7_7_cond_0_1) begin
        ram_w4_l8192_id7_7_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id7_7_cond_1_1) begin
        _tmp_691 <= 1;
      end 
      _ram_w4_l8192_id7_7_cond_2_2 <= _ram_w4_l8192_id7_7_cond_2_1;
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0)) begin
        ram_w4_l8192_id7_7_1_addr <= _tmp_283;
        ram_w4_l8192_id7_7_1_wdata <= _dataflow_slice_odata_50;
        ram_w4_l8192_id7_7_1_wenable <= _tmp_285 == 7;
      end 
      _ram_w4_l8192_id7_7_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19)) begin
        ram_w4_l8192_id7_7_0_addr <= _stream_conv2d_16_source_35_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id7_7_cond_1_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      _ram_w4_l8192_id7_7_cond_2_1 <= _stream_conv2d_16_source_35_source_ram_renable && (_stream_conv2d_16_source_35_source_ram_sel == 19);
      ram_w4_l8192_id7_7_0_wdata <= 0;
      ram_w4_l8192_id7_7_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id8_0_1_addr <= 0;
      ram_w4_l8192_id8_0_1_wdata <= 0;
      ram_w4_l8192_id8_0_1_wenable <= 0;
      _ram_w4_l8192_id8_0_cond_0_1 <= 0;
      ram_w4_l8192_id8_0_0_addr <= 0;
      _ram_w4_l8192_id8_0_cond_1_1 <= 0;
      _tmp_698 <= 0;
      _ram_w4_l8192_id8_0_cond_2_1 <= 0;
      _ram_w4_l8192_id8_0_cond_2_2 <= 0;
      ram_w4_l8192_id8_0_0_wdata <= 0;
      ram_w4_l8192_id8_0_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id8_0_cond_2_2) begin
        _tmp_698 <= 0;
      end 
      if(_ram_w4_l8192_id8_0_cond_0_1) begin
        ram_w4_l8192_id8_0_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id8_0_cond_1_1) begin
        _tmp_698 <= 1;
      end 
      _ram_w4_l8192_id8_0_cond_2_2 <= _ram_w4_l8192_id8_0_cond_2_1;
      if(_dataflow_slice_ovalid_29 && ((_tmp_39 > 0) && !_tmp_40) && (_tmp_39 > 0)) begin
        ram_w4_l8192_id8_0_1_addr <= _tmp_67;
        ram_w4_l8192_id8_0_1_wdata <= _dataflow_slice_odata_29;
        ram_w4_l8192_id8_0_1_wenable <= _tmp_68 == 8;
      end 
      _ram_w4_l8192_id8_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20)) begin
        ram_w4_l8192_id8_0_0_addr <= _stream_conv2d_16_source_36_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id8_0_cond_1_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      _ram_w4_l8192_id8_0_cond_2_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      ram_w4_l8192_id8_0_0_wdata <= 0;
      ram_w4_l8192_id8_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id8_1_1_addr <= 0;
      ram_w4_l8192_id8_1_1_wdata <= 0;
      ram_w4_l8192_id8_1_1_wenable <= 0;
      _ram_w4_l8192_id8_1_cond_0_1 <= 0;
      ram_w4_l8192_id8_1_0_addr <= 0;
      _ram_w4_l8192_id8_1_cond_1_1 <= 0;
      _tmp_699 <= 0;
      _ram_w4_l8192_id8_1_cond_2_1 <= 0;
      _ram_w4_l8192_id8_1_cond_2_2 <= 0;
      ram_w4_l8192_id8_1_0_wdata <= 0;
      ram_w4_l8192_id8_1_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id8_1_cond_2_2) begin
        _tmp_699 <= 0;
      end 
      if(_ram_w4_l8192_id8_1_cond_0_1) begin
        ram_w4_l8192_id8_1_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id8_1_cond_1_1) begin
        _tmp_699 <= 1;
      end 
      _ram_w4_l8192_id8_1_cond_2_2 <= _ram_w4_l8192_id8_1_cond_2_1;
      if(_dataflow_slice_ovalid_32 && ((_tmp_70 > 0) && !_tmp_71) && (_tmp_70 > 0)) begin
        ram_w4_l8192_id8_1_1_addr <= _tmp_98;
        ram_w4_l8192_id8_1_1_wdata <= _dataflow_slice_odata_32;
        ram_w4_l8192_id8_1_1_wenable <= _tmp_99 == 8;
      end 
      _ram_w4_l8192_id8_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20)) begin
        ram_w4_l8192_id8_1_0_addr <= _stream_conv2d_16_source_36_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id8_1_cond_1_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      _ram_w4_l8192_id8_1_cond_2_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      ram_w4_l8192_id8_1_0_wdata <= 0;
      ram_w4_l8192_id8_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id8_2_1_addr <= 0;
      ram_w4_l8192_id8_2_1_wdata <= 0;
      ram_w4_l8192_id8_2_1_wenable <= 0;
      _ram_w4_l8192_id8_2_cond_0_1 <= 0;
      ram_w4_l8192_id8_2_0_addr <= 0;
      _ram_w4_l8192_id8_2_cond_1_1 <= 0;
      _tmp_700 <= 0;
      _ram_w4_l8192_id8_2_cond_2_1 <= 0;
      _ram_w4_l8192_id8_2_cond_2_2 <= 0;
      ram_w4_l8192_id8_2_0_wdata <= 0;
      ram_w4_l8192_id8_2_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id8_2_cond_2_2) begin
        _tmp_700 <= 0;
      end 
      if(_ram_w4_l8192_id8_2_cond_0_1) begin
        ram_w4_l8192_id8_2_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id8_2_cond_1_1) begin
        _tmp_700 <= 1;
      end 
      _ram_w4_l8192_id8_2_cond_2_2 <= _ram_w4_l8192_id8_2_cond_2_1;
      if(_dataflow_slice_ovalid_35 && ((_tmp_101 > 0) && !_tmp_102) && (_tmp_101 > 0)) begin
        ram_w4_l8192_id8_2_1_addr <= _tmp_129;
        ram_w4_l8192_id8_2_1_wdata <= _dataflow_slice_odata_35;
        ram_w4_l8192_id8_2_1_wenable <= _tmp_130 == 8;
      end 
      _ram_w4_l8192_id8_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20)) begin
        ram_w4_l8192_id8_2_0_addr <= _stream_conv2d_16_source_36_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id8_2_cond_1_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      _ram_w4_l8192_id8_2_cond_2_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      ram_w4_l8192_id8_2_0_wdata <= 0;
      ram_w4_l8192_id8_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id8_3_1_addr <= 0;
      ram_w4_l8192_id8_3_1_wdata <= 0;
      ram_w4_l8192_id8_3_1_wenable <= 0;
      _ram_w4_l8192_id8_3_cond_0_1 <= 0;
      ram_w4_l8192_id8_3_0_addr <= 0;
      _ram_w4_l8192_id8_3_cond_1_1 <= 0;
      _tmp_701 <= 0;
      _ram_w4_l8192_id8_3_cond_2_1 <= 0;
      _ram_w4_l8192_id8_3_cond_2_2 <= 0;
      ram_w4_l8192_id8_3_0_wdata <= 0;
      ram_w4_l8192_id8_3_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id8_3_cond_2_2) begin
        _tmp_701 <= 0;
      end 
      if(_ram_w4_l8192_id8_3_cond_0_1) begin
        ram_w4_l8192_id8_3_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id8_3_cond_1_1) begin
        _tmp_701 <= 1;
      end 
      _ram_w4_l8192_id8_3_cond_2_2 <= _ram_w4_l8192_id8_3_cond_2_1;
      if(_dataflow_slice_ovalid_38 && ((_tmp_132 > 0) && !_tmp_133) && (_tmp_132 > 0)) begin
        ram_w4_l8192_id8_3_1_addr <= _tmp_160;
        ram_w4_l8192_id8_3_1_wdata <= _dataflow_slice_odata_38;
        ram_w4_l8192_id8_3_1_wenable <= _tmp_161 == 8;
      end 
      _ram_w4_l8192_id8_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20)) begin
        ram_w4_l8192_id8_3_0_addr <= _stream_conv2d_16_source_36_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id8_3_cond_1_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      _ram_w4_l8192_id8_3_cond_2_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      ram_w4_l8192_id8_3_0_wdata <= 0;
      ram_w4_l8192_id8_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id8_4_1_addr <= 0;
      ram_w4_l8192_id8_4_1_wdata <= 0;
      ram_w4_l8192_id8_4_1_wenable <= 0;
      _ram_w4_l8192_id8_4_cond_0_1 <= 0;
      ram_w4_l8192_id8_4_0_addr <= 0;
      _ram_w4_l8192_id8_4_cond_1_1 <= 0;
      _tmp_702 <= 0;
      _ram_w4_l8192_id8_4_cond_2_1 <= 0;
      _ram_w4_l8192_id8_4_cond_2_2 <= 0;
      ram_w4_l8192_id8_4_0_wdata <= 0;
      ram_w4_l8192_id8_4_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id8_4_cond_2_2) begin
        _tmp_702 <= 0;
      end 
      if(_ram_w4_l8192_id8_4_cond_0_1) begin
        ram_w4_l8192_id8_4_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id8_4_cond_1_1) begin
        _tmp_702 <= 1;
      end 
      _ram_w4_l8192_id8_4_cond_2_2 <= _ram_w4_l8192_id8_4_cond_2_1;
      if(_dataflow_slice_ovalid_41 && ((_tmp_163 > 0) && !_tmp_164) && (_tmp_163 > 0)) begin
        ram_w4_l8192_id8_4_1_addr <= _tmp_191;
        ram_w4_l8192_id8_4_1_wdata <= _dataflow_slice_odata_41;
        ram_w4_l8192_id8_4_1_wenable <= _tmp_192 == 8;
      end 
      _ram_w4_l8192_id8_4_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20)) begin
        ram_w4_l8192_id8_4_0_addr <= _stream_conv2d_16_source_36_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id8_4_cond_1_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      _ram_w4_l8192_id8_4_cond_2_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      ram_w4_l8192_id8_4_0_wdata <= 0;
      ram_w4_l8192_id8_4_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id8_5_1_addr <= 0;
      ram_w4_l8192_id8_5_1_wdata <= 0;
      ram_w4_l8192_id8_5_1_wenable <= 0;
      _ram_w4_l8192_id8_5_cond_0_1 <= 0;
      ram_w4_l8192_id8_5_0_addr <= 0;
      _ram_w4_l8192_id8_5_cond_1_1 <= 0;
      _tmp_703 <= 0;
      _ram_w4_l8192_id8_5_cond_2_1 <= 0;
      _ram_w4_l8192_id8_5_cond_2_2 <= 0;
      ram_w4_l8192_id8_5_0_wdata <= 0;
      ram_w4_l8192_id8_5_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id8_5_cond_2_2) begin
        _tmp_703 <= 0;
      end 
      if(_ram_w4_l8192_id8_5_cond_0_1) begin
        ram_w4_l8192_id8_5_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id8_5_cond_1_1) begin
        _tmp_703 <= 1;
      end 
      _ram_w4_l8192_id8_5_cond_2_2 <= _ram_w4_l8192_id8_5_cond_2_1;
      if(_dataflow_slice_ovalid_44 && ((_tmp_194 > 0) && !_tmp_195) && (_tmp_194 > 0)) begin
        ram_w4_l8192_id8_5_1_addr <= _tmp_222;
        ram_w4_l8192_id8_5_1_wdata <= _dataflow_slice_odata_44;
        ram_w4_l8192_id8_5_1_wenable <= _tmp_223 == 8;
      end 
      _ram_w4_l8192_id8_5_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20)) begin
        ram_w4_l8192_id8_5_0_addr <= _stream_conv2d_16_source_36_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id8_5_cond_1_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      _ram_w4_l8192_id8_5_cond_2_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      ram_w4_l8192_id8_5_0_wdata <= 0;
      ram_w4_l8192_id8_5_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id8_6_1_addr <= 0;
      ram_w4_l8192_id8_6_1_wdata <= 0;
      ram_w4_l8192_id8_6_1_wenable <= 0;
      _ram_w4_l8192_id8_6_cond_0_1 <= 0;
      ram_w4_l8192_id8_6_0_addr <= 0;
      _ram_w4_l8192_id8_6_cond_1_1 <= 0;
      _tmp_704 <= 0;
      _ram_w4_l8192_id8_6_cond_2_1 <= 0;
      _ram_w4_l8192_id8_6_cond_2_2 <= 0;
      ram_w4_l8192_id8_6_0_wdata <= 0;
      ram_w4_l8192_id8_6_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id8_6_cond_2_2) begin
        _tmp_704 <= 0;
      end 
      if(_ram_w4_l8192_id8_6_cond_0_1) begin
        ram_w4_l8192_id8_6_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id8_6_cond_1_1) begin
        _tmp_704 <= 1;
      end 
      _ram_w4_l8192_id8_6_cond_2_2 <= _ram_w4_l8192_id8_6_cond_2_1;
      if(_dataflow_slice_ovalid_47 && ((_tmp_225 > 0) && !_tmp_226) && (_tmp_225 > 0)) begin
        ram_w4_l8192_id8_6_1_addr <= _tmp_253;
        ram_w4_l8192_id8_6_1_wdata <= _dataflow_slice_odata_47;
        ram_w4_l8192_id8_6_1_wenable <= _tmp_254 == 8;
      end 
      _ram_w4_l8192_id8_6_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20)) begin
        ram_w4_l8192_id8_6_0_addr <= _stream_conv2d_16_source_36_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id8_6_cond_1_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      _ram_w4_l8192_id8_6_cond_2_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      ram_w4_l8192_id8_6_0_wdata <= 0;
      ram_w4_l8192_id8_6_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w4_l8192_id8_7_1_addr <= 0;
      ram_w4_l8192_id8_7_1_wdata <= 0;
      ram_w4_l8192_id8_7_1_wenable <= 0;
      _ram_w4_l8192_id8_7_cond_0_1 <= 0;
      ram_w4_l8192_id8_7_0_addr <= 0;
      _ram_w4_l8192_id8_7_cond_1_1 <= 0;
      _tmp_705 <= 0;
      _ram_w4_l8192_id8_7_cond_2_1 <= 0;
      _ram_w4_l8192_id8_7_cond_2_2 <= 0;
      ram_w4_l8192_id8_7_0_wdata <= 0;
      ram_w4_l8192_id8_7_0_wenable <= 0;
    end else begin
      if(_ram_w4_l8192_id8_7_cond_2_2) begin
        _tmp_705 <= 0;
      end 
      if(_ram_w4_l8192_id8_7_cond_0_1) begin
        ram_w4_l8192_id8_7_1_wenable <= 0;
      end 
      if(_ram_w4_l8192_id8_7_cond_1_1) begin
        _tmp_705 <= 1;
      end 
      _ram_w4_l8192_id8_7_cond_2_2 <= _ram_w4_l8192_id8_7_cond_2_1;
      if(_dataflow_slice_ovalid_50 && ((_tmp_256 > 0) && !_tmp_257) && (_tmp_256 > 0)) begin
        ram_w4_l8192_id8_7_1_addr <= _tmp_284;
        ram_w4_l8192_id8_7_1_wdata <= _dataflow_slice_odata_50;
        ram_w4_l8192_id8_7_1_wenable <= _tmp_285 == 8;
      end 
      _ram_w4_l8192_id8_7_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20)) begin
        ram_w4_l8192_id8_7_0_addr <= _stream_conv2d_16_source_36_source_ram_raddr >> 3;
      end 
      _ram_w4_l8192_id8_7_cond_1_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      _ram_w4_l8192_id8_7_cond_2_1 <= _stream_conv2d_16_source_36_source_ram_renable && (_stream_conv2d_16_source_36_source_ram_sel == 20);
      ram_w4_l8192_id8_7_0_wdata <= 0;
      ram_w4_l8192_id8_7_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id0_0_1_addr <= 0;
      _tmp_25 <= 0;
      ram_w8_l2048_id0_0_1_wdata <= 0;
      ram_w8_l2048_id0_0_1_wenable <= 0;
      _tmp_26 <= 0;
      _ram_w8_l2048_id0_0_cond_0_1 <= 0;
      ram_w8_l2048_id0_0_0_addr <= 0;
      _ram_w8_l2048_id0_0_cond_1_1 <= 0;
      _tmp_476 <= 0;
      _ram_w8_l2048_id0_0_cond_2_1 <= 0;
      _ram_w8_l2048_id0_0_cond_2_2 <= 0;
      ram_w8_l2048_id0_0_0_wdata <= 0;
      ram_w8_l2048_id0_0_0_wenable <= 0;
      _ram_w8_l2048_id0_0_cond_3_1 <= 0;
      __tmp_1077_1 <= 0;
      __tmp_1078_1 <= 0;
      _tmp_1082 <= 0;
      _tmp_1072 <= 0;
      _tmp_1073 <= 0;
      _tmp_1080 <= 0;
      _tmp_1081 <= 0;
      _tmp_1079 <= 0;
      _tmp_1083 <= 0;
      _ram_w8_l2048_id0_0_cond_4_1 <= 0;
      _tmp_1182 <= 0;
      _ram_w8_l2048_id0_0_cond_5_1 <= 0;
      _ram_w8_l2048_id0_0_cond_5_2 <= 0;
    end else begin
      if(_ram_w8_l2048_id0_0_cond_2_2) begin
        _tmp_476 <= 0;
      end 
      if(_ram_w8_l2048_id0_0_cond_5_2) begin
        _tmp_1182 <= 0;
      end 
      if(_ram_w8_l2048_id0_0_cond_0_1) begin
        ram_w8_l2048_id0_0_1_wenable <= 0;
        _tmp_26 <= 0;
      end 
      if(_ram_w8_l2048_id0_0_cond_1_1) begin
        _tmp_476 <= 1;
      end 
      _ram_w8_l2048_id0_0_cond_2_2 <= _ram_w8_l2048_id0_0_cond_2_1;
      if(_ram_w8_l2048_id0_0_cond_3_1) begin
        ram_w8_l2048_id0_0_0_wenable <= 0;
      end 
      if(_ram_w8_l2048_id0_0_cond_4_1) begin
        _tmp_1182 <= 1;
      end 
      _ram_w8_l2048_id0_0_cond_5_2 <= _ram_w8_l2048_id0_0_cond_5_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 2) && (_tmp_25 == 0)) begin
        ram_w8_l2048_id0_0_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_25 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_16 && ((_tmp_25 > 0) && !_tmp_26) && (_tmp_25 > 0)) begin
        ram_w8_l2048_id0_0_1_addr <= ram_w8_l2048_id0_0_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id0_0_1_wdata <= _dataflow_slice_odata_16;
        ram_w8_l2048_id0_0_1_wenable <= 1;
        _tmp_25 <= _tmp_25 - 1;
      end 
      if(_dataflow_slice_ovalid_16 && ((_tmp_25 > 0) && !_tmp_26) && (_tmp_25 == 1)) begin
        _tmp_26 <= 1;
      end 
      _ram_w8_l2048_id0_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2)) begin
        ram_w8_l2048_id0_0_0_addr <= _stream_conv2d_16_source_8_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id0_0_cond_1_1 <= _stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2);
      _ram_w8_l2048_id0_0_cond_2_1 <= _stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2);
      if(_stream_max_pool_serial_18_sink_3_sink_wenable && (_stream_max_pool_serial_18_sink_3_sink_ram_sel == 2) && (_tmp_1037 == 0)) begin
        ram_w8_l2048_id0_0_0_addr <= _stream_max_pool_serial_18_sink_3_sink_waddr >> 2;
        ram_w8_l2048_id0_0_0_wdata <= _stream_max_pool_serial_18_sink_3_sink_wdata;
        ram_w8_l2048_id0_0_0_wenable <= 1;
      end 
      _ram_w8_l2048_id0_0_cond_3_1 <= _stream_max_pool_serial_18_sink_3_sink_wenable && (_stream_max_pool_serial_18_sink_3_sink_ram_sel == 2) && (_tmp_1037 == 0);
      __tmp_1077_1 <= _tmp_1077;
      __tmp_1078_1 <= _tmp_1078;
      if((_tmp_1074 || !_tmp_1072) && (_tmp_1075 || !_tmp_1073) && _tmp_1080) begin
        _tmp_1082 <= 0;
        _tmp_1072 <= 0;
        _tmp_1073 <= 0;
        _tmp_1080 <= 0;
      end 
      if((_tmp_1074 || !_tmp_1072) && (_tmp_1075 || !_tmp_1073) && _tmp_1079) begin
        _tmp_1072 <= 1;
        _tmp_1073 <= 1;
        _tmp_1082 <= _tmp_1081;
        _tmp_1081 <= 0;
        _tmp_1079 <= 0;
        _tmp_1080 <= 1;
      end 
      if(_maxi_write_start && (_maxi_write_op_sel == 2) && (_tmp_1083 == 0) && !_tmp_1081 && !_tmp_1082) begin
        ram_w8_l2048_id0_0_1_addr <= _maxi_write_local_addr;
        _tmp_1083 <= _maxi_write_size - 1;
        _tmp_1079 <= 1;
        _tmp_1081 <= _maxi_write_size == 1;
      end 
      if((_tmp_1074 || !_tmp_1072) && (_tmp_1075 || !_tmp_1073) && (_tmp_1083 > 0)) begin
        ram_w8_l2048_id0_0_1_addr <= ram_w8_l2048_id0_0_1_addr + _maxi_write_local_stride;
        _tmp_1083 <= _tmp_1083 - 1;
        _tmp_1079 <= 1;
        _tmp_1081 <= 0;
      end 
      if((_tmp_1074 || !_tmp_1072) && (_tmp_1075 || !_tmp_1073) && (_tmp_1083 == 1)) begin
        _tmp_1081 <= 1;
      end 
      if(_stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2)) begin
        ram_w8_l2048_id0_0_0_addr <= _stream_matmul_29_source_8_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id0_0_cond_4_1 <= _stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2);
      _ram_w8_l2048_id0_0_cond_5_1 <= _stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2);
    end
  end

  reg [32-1:0] _dataflow_cat_data_107;
  reg _dataflow_cat_valid_107;
  wire _dataflow_cat_ready_107;
  assign _tmp_1110 = 1 && ((_dataflow_cat_ready_107 || !_dataflow_cat_valid_107) && (_tmp_1108 && _tmp_1096 && _tmp_1084 && _tmp_1072));
  assign _tmp_1098 = 1 && ((_dataflow_cat_ready_107 || !_dataflow_cat_valid_107) && (_tmp_1108 && _tmp_1096 && _tmp_1084 && _tmp_1072));
  assign _tmp_1086 = 1 && ((_dataflow_cat_ready_107 || !_dataflow_cat_valid_107) && (_tmp_1108 && _tmp_1096 && _tmp_1084 && _tmp_1072));
  assign _tmp_1074 = 1 && ((_dataflow_cat_ready_107 || !_dataflow_cat_valid_107) && (_tmp_1108 && _tmp_1096 && _tmp_1084 && _tmp_1072));
  assign _dataflow_cat_odata_107 = _dataflow_cat_data_107;
  assign _dataflow_cat_ovalid_107 = _dataflow_cat_valid_107;
  assign _dataflow_cat_ready_107 = _dataflow_cat_oready_107;

  always @(posedge CLK) begin
    if(RST) begin
      _dataflow_cat_data_107 <= 0;
      _dataflow_cat_valid_107 <= 0;
    end else begin
      if((_dataflow_cat_ready_107 || !_dataflow_cat_valid_107) && (_tmp_1110 && _tmp_1098 && _tmp_1086 && _tmp_1074) && (_tmp_1108 && _tmp_1096 && _tmp_1084 && _tmp_1072)) begin
        _dataflow_cat_data_107 <= { _tmp_1114, _tmp_1102, _tmp_1090, _tmp_1078 };
      end 
      if(_dataflow_cat_valid_107 && _dataflow_cat_ready_107) begin
        _dataflow_cat_valid_107 <= 0;
      end 
      if((_dataflow_cat_ready_107 || !_dataflow_cat_valid_107) && (_tmp_1110 && _tmp_1098 && _tmp_1086 && _tmp_1074)) begin
        _dataflow_cat_valid_107 <= _tmp_1108 && _tmp_1096 && _tmp_1084 && _tmp_1072;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id0_1_1_addr <= 0;
      _tmp_27 <= 0;
      ram_w8_l2048_id0_1_1_wdata <= 0;
      ram_w8_l2048_id0_1_1_wenable <= 0;
      _tmp_28 <= 0;
      _ram_w8_l2048_id0_1_cond_0_1 <= 0;
      ram_w8_l2048_id0_1_0_addr <= 0;
      _ram_w8_l2048_id0_1_cond_1_1 <= 0;
      _tmp_477 <= 0;
      _ram_w8_l2048_id0_1_cond_2_1 <= 0;
      _ram_w8_l2048_id0_1_cond_2_2 <= 0;
      ram_w8_l2048_id0_1_0_wdata <= 0;
      ram_w8_l2048_id0_1_0_wenable <= 0;
      _ram_w8_l2048_id0_1_cond_3_1 <= 0;
      __tmp_1089_1 <= 0;
      __tmp_1090_1 <= 0;
      _tmp_1094 <= 0;
      _tmp_1084 <= 0;
      _tmp_1085 <= 0;
      _tmp_1092 <= 0;
      _tmp_1093 <= 0;
      _tmp_1091 <= 0;
      _tmp_1095 <= 0;
      _ram_w8_l2048_id0_1_cond_4_1 <= 0;
      _tmp_1183 <= 0;
      _ram_w8_l2048_id0_1_cond_5_1 <= 0;
      _ram_w8_l2048_id0_1_cond_5_2 <= 0;
    end else begin
      if(_ram_w8_l2048_id0_1_cond_2_2) begin
        _tmp_477 <= 0;
      end 
      if(_ram_w8_l2048_id0_1_cond_5_2) begin
        _tmp_1183 <= 0;
      end 
      if(_ram_w8_l2048_id0_1_cond_0_1) begin
        ram_w8_l2048_id0_1_1_wenable <= 0;
        _tmp_28 <= 0;
      end 
      if(_ram_w8_l2048_id0_1_cond_1_1) begin
        _tmp_477 <= 1;
      end 
      _ram_w8_l2048_id0_1_cond_2_2 <= _ram_w8_l2048_id0_1_cond_2_1;
      if(_ram_w8_l2048_id0_1_cond_3_1) begin
        ram_w8_l2048_id0_1_0_wenable <= 0;
      end 
      if(_ram_w8_l2048_id0_1_cond_4_1) begin
        _tmp_1183 <= 1;
      end 
      _ram_w8_l2048_id0_1_cond_5_2 <= _ram_w8_l2048_id0_1_cond_5_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 2) && (_tmp_27 == 0)) begin
        ram_w8_l2048_id0_1_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_27 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_19 && ((_tmp_27 > 0) && !_tmp_28) && (_tmp_27 > 0)) begin
        ram_w8_l2048_id0_1_1_addr <= ram_w8_l2048_id0_1_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id0_1_1_wdata <= _dataflow_slice_odata_19;
        ram_w8_l2048_id0_1_1_wenable <= 1;
        _tmp_27 <= _tmp_27 - 1;
      end 
      if(_dataflow_slice_ovalid_19 && ((_tmp_27 > 0) && !_tmp_28) && (_tmp_27 == 1)) begin
        _tmp_28 <= 1;
      end 
      _ram_w8_l2048_id0_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2)) begin
        ram_w8_l2048_id0_1_0_addr <= _stream_conv2d_16_source_8_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id0_1_cond_1_1 <= _stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2);
      _ram_w8_l2048_id0_1_cond_2_1 <= _stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2);
      if(_stream_max_pool_serial_18_sink_3_sink_wenable && (_stream_max_pool_serial_18_sink_3_sink_ram_sel == 2) && (_tmp_1037 == 1)) begin
        ram_w8_l2048_id0_1_0_addr <= _stream_max_pool_serial_18_sink_3_sink_waddr >> 2;
        ram_w8_l2048_id0_1_0_wdata <= _stream_max_pool_serial_18_sink_3_sink_wdata;
        ram_w8_l2048_id0_1_0_wenable <= 1;
      end 
      _ram_w8_l2048_id0_1_cond_3_1 <= _stream_max_pool_serial_18_sink_3_sink_wenable && (_stream_max_pool_serial_18_sink_3_sink_ram_sel == 2) && (_tmp_1037 == 1);
      __tmp_1089_1 <= _tmp_1089;
      __tmp_1090_1 <= _tmp_1090;
      if((_tmp_1086 || !_tmp_1084) && (_tmp_1087 || !_tmp_1085) && _tmp_1092) begin
        _tmp_1094 <= 0;
        _tmp_1084 <= 0;
        _tmp_1085 <= 0;
        _tmp_1092 <= 0;
      end 
      if((_tmp_1086 || !_tmp_1084) && (_tmp_1087 || !_tmp_1085) && _tmp_1091) begin
        _tmp_1084 <= 1;
        _tmp_1085 <= 1;
        _tmp_1094 <= _tmp_1093;
        _tmp_1093 <= 0;
        _tmp_1091 <= 0;
        _tmp_1092 <= 1;
      end 
      if(_maxi_write_start && (_maxi_write_op_sel == 2) && (_tmp_1095 == 0) && !_tmp_1093 && !_tmp_1094) begin
        ram_w8_l2048_id0_1_1_addr <= _maxi_write_local_addr;
        _tmp_1095 <= _maxi_write_size - 1;
        _tmp_1091 <= 1;
        _tmp_1093 <= _maxi_write_size == 1;
      end 
      if((_tmp_1086 || !_tmp_1084) && (_tmp_1087 || !_tmp_1085) && (_tmp_1095 > 0)) begin
        ram_w8_l2048_id0_1_1_addr <= ram_w8_l2048_id0_1_1_addr + _maxi_write_local_stride;
        _tmp_1095 <= _tmp_1095 - 1;
        _tmp_1091 <= 1;
        _tmp_1093 <= 0;
      end 
      if((_tmp_1086 || !_tmp_1084) && (_tmp_1087 || !_tmp_1085) && (_tmp_1095 == 1)) begin
        _tmp_1093 <= 1;
      end 
      if(_stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2)) begin
        ram_w8_l2048_id0_1_0_addr <= _stream_matmul_29_source_8_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id0_1_cond_4_1 <= _stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2);
      _ram_w8_l2048_id0_1_cond_5_1 <= _stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2);
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id0_2_1_addr <= 0;
      _tmp_29 <= 0;
      ram_w8_l2048_id0_2_1_wdata <= 0;
      ram_w8_l2048_id0_2_1_wenable <= 0;
      _tmp_30 <= 0;
      _ram_w8_l2048_id0_2_cond_0_1 <= 0;
      ram_w8_l2048_id0_2_0_addr <= 0;
      _ram_w8_l2048_id0_2_cond_1_1 <= 0;
      _tmp_478 <= 0;
      _ram_w8_l2048_id0_2_cond_2_1 <= 0;
      _ram_w8_l2048_id0_2_cond_2_2 <= 0;
      ram_w8_l2048_id0_2_0_wdata <= 0;
      ram_w8_l2048_id0_2_0_wenable <= 0;
      _ram_w8_l2048_id0_2_cond_3_1 <= 0;
      __tmp_1101_1 <= 0;
      __tmp_1102_1 <= 0;
      _tmp_1106 <= 0;
      _tmp_1096 <= 0;
      _tmp_1097 <= 0;
      _tmp_1104 <= 0;
      _tmp_1105 <= 0;
      _tmp_1103 <= 0;
      _tmp_1107 <= 0;
      _ram_w8_l2048_id0_2_cond_4_1 <= 0;
      _tmp_1184 <= 0;
      _ram_w8_l2048_id0_2_cond_5_1 <= 0;
      _ram_w8_l2048_id0_2_cond_5_2 <= 0;
    end else begin
      if(_ram_w8_l2048_id0_2_cond_2_2) begin
        _tmp_478 <= 0;
      end 
      if(_ram_w8_l2048_id0_2_cond_5_2) begin
        _tmp_1184 <= 0;
      end 
      if(_ram_w8_l2048_id0_2_cond_0_1) begin
        ram_w8_l2048_id0_2_1_wenable <= 0;
        _tmp_30 <= 0;
      end 
      if(_ram_w8_l2048_id0_2_cond_1_1) begin
        _tmp_478 <= 1;
      end 
      _ram_w8_l2048_id0_2_cond_2_2 <= _ram_w8_l2048_id0_2_cond_2_1;
      if(_ram_w8_l2048_id0_2_cond_3_1) begin
        ram_w8_l2048_id0_2_0_wenable <= 0;
      end 
      if(_ram_w8_l2048_id0_2_cond_4_1) begin
        _tmp_1184 <= 1;
      end 
      _ram_w8_l2048_id0_2_cond_5_2 <= _ram_w8_l2048_id0_2_cond_5_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 2) && (_tmp_29 == 0)) begin
        ram_w8_l2048_id0_2_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_29 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_22 && ((_tmp_29 > 0) && !_tmp_30) && (_tmp_29 > 0)) begin
        ram_w8_l2048_id0_2_1_addr <= ram_w8_l2048_id0_2_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id0_2_1_wdata <= _dataflow_slice_odata_22;
        ram_w8_l2048_id0_2_1_wenable <= 1;
        _tmp_29 <= _tmp_29 - 1;
      end 
      if(_dataflow_slice_ovalid_22 && ((_tmp_29 > 0) && !_tmp_30) && (_tmp_29 == 1)) begin
        _tmp_30 <= 1;
      end 
      _ram_w8_l2048_id0_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2)) begin
        ram_w8_l2048_id0_2_0_addr <= _stream_conv2d_16_source_8_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id0_2_cond_1_1 <= _stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2);
      _ram_w8_l2048_id0_2_cond_2_1 <= _stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2);
      if(_stream_max_pool_serial_18_sink_3_sink_wenable && (_stream_max_pool_serial_18_sink_3_sink_ram_sel == 2) && (_tmp_1037 == 2)) begin
        ram_w8_l2048_id0_2_0_addr <= _stream_max_pool_serial_18_sink_3_sink_waddr >> 2;
        ram_w8_l2048_id0_2_0_wdata <= _stream_max_pool_serial_18_sink_3_sink_wdata;
        ram_w8_l2048_id0_2_0_wenable <= 1;
      end 
      _ram_w8_l2048_id0_2_cond_3_1 <= _stream_max_pool_serial_18_sink_3_sink_wenable && (_stream_max_pool_serial_18_sink_3_sink_ram_sel == 2) && (_tmp_1037 == 2);
      __tmp_1101_1 <= _tmp_1101;
      __tmp_1102_1 <= _tmp_1102;
      if((_tmp_1098 || !_tmp_1096) && (_tmp_1099 || !_tmp_1097) && _tmp_1104) begin
        _tmp_1106 <= 0;
        _tmp_1096 <= 0;
        _tmp_1097 <= 0;
        _tmp_1104 <= 0;
      end 
      if((_tmp_1098 || !_tmp_1096) && (_tmp_1099 || !_tmp_1097) && _tmp_1103) begin
        _tmp_1096 <= 1;
        _tmp_1097 <= 1;
        _tmp_1106 <= _tmp_1105;
        _tmp_1105 <= 0;
        _tmp_1103 <= 0;
        _tmp_1104 <= 1;
      end 
      if(_maxi_write_start && (_maxi_write_op_sel == 2) && (_tmp_1107 == 0) && !_tmp_1105 && !_tmp_1106) begin
        ram_w8_l2048_id0_2_1_addr <= _maxi_write_local_addr;
        _tmp_1107 <= _maxi_write_size - 1;
        _tmp_1103 <= 1;
        _tmp_1105 <= _maxi_write_size == 1;
      end 
      if((_tmp_1098 || !_tmp_1096) && (_tmp_1099 || !_tmp_1097) && (_tmp_1107 > 0)) begin
        ram_w8_l2048_id0_2_1_addr <= ram_w8_l2048_id0_2_1_addr + _maxi_write_local_stride;
        _tmp_1107 <= _tmp_1107 - 1;
        _tmp_1103 <= 1;
        _tmp_1105 <= 0;
      end 
      if((_tmp_1098 || !_tmp_1096) && (_tmp_1099 || !_tmp_1097) && (_tmp_1107 == 1)) begin
        _tmp_1105 <= 1;
      end 
      if(_stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2)) begin
        ram_w8_l2048_id0_2_0_addr <= _stream_matmul_29_source_8_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id0_2_cond_4_1 <= _stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2);
      _ram_w8_l2048_id0_2_cond_5_1 <= _stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2);
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id0_3_1_addr <= 0;
      _tmp_31 <= 0;
      ram_w8_l2048_id0_3_1_wdata <= 0;
      ram_w8_l2048_id0_3_1_wenable <= 0;
      _tmp_32 <= 0;
      _ram_w8_l2048_id0_3_cond_0_1 <= 0;
      ram_w8_l2048_id0_3_0_addr <= 0;
      _ram_w8_l2048_id0_3_cond_1_1 <= 0;
      _tmp_479 <= 0;
      _ram_w8_l2048_id0_3_cond_2_1 <= 0;
      _ram_w8_l2048_id0_3_cond_2_2 <= 0;
      ram_w8_l2048_id0_3_0_wdata <= 0;
      ram_w8_l2048_id0_3_0_wenable <= 0;
      _ram_w8_l2048_id0_3_cond_3_1 <= 0;
      __tmp_1113_1 <= 0;
      __tmp_1114_1 <= 0;
      _tmp_1118 <= 0;
      _tmp_1108 <= 0;
      _tmp_1109 <= 0;
      _tmp_1116 <= 0;
      _tmp_1117 <= 0;
      _tmp_1115 <= 0;
      _tmp_1119 <= 0;
      _ram_w8_l2048_id0_3_cond_4_1 <= 0;
      _tmp_1185 <= 0;
      _ram_w8_l2048_id0_3_cond_5_1 <= 0;
      _ram_w8_l2048_id0_3_cond_5_2 <= 0;
    end else begin
      if(_ram_w8_l2048_id0_3_cond_2_2) begin
        _tmp_479 <= 0;
      end 
      if(_ram_w8_l2048_id0_3_cond_5_2) begin
        _tmp_1185 <= 0;
      end 
      if(_ram_w8_l2048_id0_3_cond_0_1) begin
        ram_w8_l2048_id0_3_1_wenable <= 0;
        _tmp_32 <= 0;
      end 
      if(_ram_w8_l2048_id0_3_cond_1_1) begin
        _tmp_479 <= 1;
      end 
      _ram_w8_l2048_id0_3_cond_2_2 <= _ram_w8_l2048_id0_3_cond_2_1;
      if(_ram_w8_l2048_id0_3_cond_3_1) begin
        ram_w8_l2048_id0_3_0_wenable <= 0;
      end 
      if(_ram_w8_l2048_id0_3_cond_4_1) begin
        _tmp_1185 <= 1;
      end 
      _ram_w8_l2048_id0_3_cond_5_2 <= _ram_w8_l2048_id0_3_cond_5_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 2) && (_tmp_31 == 0)) begin
        ram_w8_l2048_id0_3_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_31 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_25 && ((_tmp_31 > 0) && !_tmp_32) && (_tmp_31 > 0)) begin
        ram_w8_l2048_id0_3_1_addr <= ram_w8_l2048_id0_3_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id0_3_1_wdata <= _dataflow_slice_odata_25;
        ram_w8_l2048_id0_3_1_wenable <= 1;
        _tmp_31 <= _tmp_31 - 1;
      end 
      if(_dataflow_slice_ovalid_25 && ((_tmp_31 > 0) && !_tmp_32) && (_tmp_31 == 1)) begin
        _tmp_32 <= 1;
      end 
      _ram_w8_l2048_id0_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2)) begin
        ram_w8_l2048_id0_3_0_addr <= _stream_conv2d_16_source_8_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id0_3_cond_1_1 <= _stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2);
      _ram_w8_l2048_id0_3_cond_2_1 <= _stream_conv2d_16_source_8_source_ram_renable && (_stream_conv2d_16_source_8_source_ram_sel == 2);
      if(_stream_max_pool_serial_18_sink_3_sink_wenable && (_stream_max_pool_serial_18_sink_3_sink_ram_sel == 2) && (_tmp_1037 == 3)) begin
        ram_w8_l2048_id0_3_0_addr <= _stream_max_pool_serial_18_sink_3_sink_waddr >> 2;
        ram_w8_l2048_id0_3_0_wdata <= _stream_max_pool_serial_18_sink_3_sink_wdata;
        ram_w8_l2048_id0_3_0_wenable <= 1;
      end 
      _ram_w8_l2048_id0_3_cond_3_1 <= _stream_max_pool_serial_18_sink_3_sink_wenable && (_stream_max_pool_serial_18_sink_3_sink_ram_sel == 2) && (_tmp_1037 == 3);
      __tmp_1113_1 <= _tmp_1113;
      __tmp_1114_1 <= _tmp_1114;
      if((_tmp_1110 || !_tmp_1108) && (_tmp_1111 || !_tmp_1109) && _tmp_1116) begin
        _tmp_1118 <= 0;
        _tmp_1108 <= 0;
        _tmp_1109 <= 0;
        _tmp_1116 <= 0;
      end 
      if((_tmp_1110 || !_tmp_1108) && (_tmp_1111 || !_tmp_1109) && _tmp_1115) begin
        _tmp_1108 <= 1;
        _tmp_1109 <= 1;
        _tmp_1118 <= _tmp_1117;
        _tmp_1117 <= 0;
        _tmp_1115 <= 0;
        _tmp_1116 <= 1;
      end 
      if(_maxi_write_start && (_maxi_write_op_sel == 2) && (_tmp_1119 == 0) && !_tmp_1117 && !_tmp_1118) begin
        ram_w8_l2048_id0_3_1_addr <= _maxi_write_local_addr;
        _tmp_1119 <= _maxi_write_size - 1;
        _tmp_1115 <= 1;
        _tmp_1117 <= _maxi_write_size == 1;
      end 
      if((_tmp_1110 || !_tmp_1108) && (_tmp_1111 || !_tmp_1109) && (_tmp_1119 > 0)) begin
        ram_w8_l2048_id0_3_1_addr <= ram_w8_l2048_id0_3_1_addr + _maxi_write_local_stride;
        _tmp_1119 <= _tmp_1119 - 1;
        _tmp_1115 <= 1;
        _tmp_1117 <= 0;
      end 
      if((_tmp_1110 || !_tmp_1108) && (_tmp_1111 || !_tmp_1109) && (_tmp_1119 == 1)) begin
        _tmp_1117 <= 1;
      end 
      if(_stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2)) begin
        ram_w8_l2048_id0_3_0_addr <= _stream_matmul_29_source_8_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id0_3_cond_4_1 <= _stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2);
      _ram_w8_l2048_id0_3_cond_5_1 <= _stream_matmul_29_source_8_source_ram_renable && (_stream_matmul_29_source_8_source_ram_sel == 2);
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id1_0_1_addr <= 0;
      _tmp_12 <= 0;
      ram_w8_l2048_id1_0_1_wdata <= 0;
      ram_w8_l2048_id1_0_1_wenable <= 0;
      _tmp_13 <= 0;
      _ram_w8_l2048_id1_0_cond_0_1 <= 0;
      ram_w8_l2048_id1_0_0_addr <= 0;
      _ram_w8_l2048_id1_0_cond_1_1 <= 0;
      _tmp_465 <= 0;
      _ram_w8_l2048_id1_0_cond_2_1 <= 0;
      _ram_w8_l2048_id1_0_cond_2_2 <= 0;
      _ram_w8_l2048_id1_0_cond_3_1 <= 0;
      _tmp_1028 <= 0;
      _ram_w8_l2048_id1_0_cond_4_1 <= 0;
      _ram_w8_l2048_id1_0_cond_4_2 <= 0;
      ram_w8_l2048_id1_0_0_wdata <= 0;
      ram_w8_l2048_id1_0_0_wenable <= 0;
      _ram_w8_l2048_id1_0_cond_5_1 <= 0;
      __tmp_1314_1 <= 0;
      __tmp_1315_1 <= 0;
      _tmp_1319 <= 0;
      _tmp_1309 <= 0;
      _tmp_1310 <= 0;
      _tmp_1317 <= 0;
      _tmp_1318 <= 0;
      _tmp_1316 <= 0;
      _tmp_1320 <= 0;
    end else begin
      if(_ram_w8_l2048_id1_0_cond_2_2) begin
        _tmp_465 <= 0;
      end 
      if(_ram_w8_l2048_id1_0_cond_4_2) begin
        _tmp_1028 <= 0;
      end 
      if(_ram_w8_l2048_id1_0_cond_0_1) begin
        ram_w8_l2048_id1_0_1_wenable <= 0;
        _tmp_13 <= 0;
      end 
      if(_ram_w8_l2048_id1_0_cond_1_1) begin
        _tmp_465 <= 1;
      end 
      _ram_w8_l2048_id1_0_cond_2_2 <= _ram_w8_l2048_id1_0_cond_2_1;
      if(_ram_w8_l2048_id1_0_cond_3_1) begin
        _tmp_1028 <= 1;
      end 
      _ram_w8_l2048_id1_0_cond_4_2 <= _ram_w8_l2048_id1_0_cond_4_1;
      if(_ram_w8_l2048_id1_0_cond_5_1) begin
        ram_w8_l2048_id1_0_0_wenable <= 0;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 1) && (_tmp_12 == 0)) begin
        ram_w8_l2048_id1_0_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_12 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_3 && ((_tmp_12 > 0) && !_tmp_13) && (_tmp_12 > 0)) begin
        ram_w8_l2048_id1_0_1_addr <= ram_w8_l2048_id1_0_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id1_0_1_wdata <= _dataflow_slice_odata_3;
        ram_w8_l2048_id1_0_1_wenable <= 1;
        _tmp_12 <= _tmp_12 - 1;
      end 
      if(_dataflow_slice_ovalid_3 && ((_tmp_12 > 0) && !_tmp_13) && (_tmp_12 == 1)) begin
        _tmp_13 <= 1;
      end 
      _ram_w8_l2048_id1_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1)) begin
        ram_w8_l2048_id1_0_0_addr <= _stream_conv2d_16_source_6_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id1_0_cond_1_1 <= _stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1);
      _ram_w8_l2048_id1_0_cond_2_1 <= _stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1);
      if(_stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1)) begin
        ram_w8_l2048_id1_0_0_addr <= _stream_max_pool_serial_18_source_1_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id1_0_cond_3_1 <= _stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1);
      _ram_w8_l2048_id1_0_cond_4_1 <= _stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1);
      if(_stream_matmul_29_sink_21_sink_wenable && (_stream_matmul_29_sink_21_sink_ram_sel == 5) && (_tmp_1225 == 0)) begin
        ram_w8_l2048_id1_0_0_addr <= _stream_matmul_29_sink_21_sink_waddr >> 2;
        ram_w8_l2048_id1_0_0_wdata <= _stream_matmul_29_sink_21_sink_wdata;
        ram_w8_l2048_id1_0_0_wenable <= 1;
      end 
      _ram_w8_l2048_id1_0_cond_5_1 <= _stream_matmul_29_sink_21_sink_wenable && (_stream_matmul_29_sink_21_sink_ram_sel == 5) && (_tmp_1225 == 0);
      __tmp_1314_1 <= _tmp_1314;
      __tmp_1315_1 <= _tmp_1315;
      if((_tmp_1311 || !_tmp_1309) && (_tmp_1312 || !_tmp_1310) && _tmp_1317) begin
        _tmp_1319 <= 0;
        _tmp_1309 <= 0;
        _tmp_1310 <= 0;
        _tmp_1317 <= 0;
      end 
      if((_tmp_1311 || !_tmp_1309) && (_tmp_1312 || !_tmp_1310) && _tmp_1316) begin
        _tmp_1309 <= 1;
        _tmp_1310 <= 1;
        _tmp_1319 <= _tmp_1318;
        _tmp_1318 <= 0;
        _tmp_1316 <= 0;
        _tmp_1317 <= 1;
      end 
      if(_maxi_write_start && (_maxi_write_op_sel == 3) && (_tmp_1320 == 0) && !_tmp_1318 && !_tmp_1319) begin
        ram_w8_l2048_id1_0_1_addr <= _maxi_write_local_addr;
        _tmp_1320 <= _maxi_write_size - 1;
        _tmp_1316 <= 1;
        _tmp_1318 <= _maxi_write_size == 1;
      end 
      if((_tmp_1311 || !_tmp_1309) && (_tmp_1312 || !_tmp_1310) && (_tmp_1320 > 0)) begin
        ram_w8_l2048_id1_0_1_addr <= ram_w8_l2048_id1_0_1_addr + _maxi_write_local_stride;
        _tmp_1320 <= _tmp_1320 - 1;
        _tmp_1316 <= 1;
        _tmp_1318 <= 0;
      end 
      if((_tmp_1311 || !_tmp_1309) && (_tmp_1312 || !_tmp_1310) && (_tmp_1320 == 1)) begin
        _tmp_1318 <= 1;
      end 
    end
  end

  reg [32-1:0] _dataflow_cat_data_167;
  reg _dataflow_cat_valid_167;
  wire _dataflow_cat_ready_167;
  assign _tmp_1347 = 1 && ((_dataflow_cat_ready_167 || !_dataflow_cat_valid_167) && (_tmp_1345 && _tmp_1333 && _tmp_1321 && _tmp_1309));
  assign _tmp_1335 = 1 && ((_dataflow_cat_ready_167 || !_dataflow_cat_valid_167) && (_tmp_1345 && _tmp_1333 && _tmp_1321 && _tmp_1309));
  assign _tmp_1323 = 1 && ((_dataflow_cat_ready_167 || !_dataflow_cat_valid_167) && (_tmp_1345 && _tmp_1333 && _tmp_1321 && _tmp_1309));
  assign _tmp_1311 = 1 && ((_dataflow_cat_ready_167 || !_dataflow_cat_valid_167) && (_tmp_1345 && _tmp_1333 && _tmp_1321 && _tmp_1309));
  assign _dataflow_cat_odata_167 = _dataflow_cat_data_167;
  assign _dataflow_cat_ovalid_167 = _dataflow_cat_valid_167;
  assign _dataflow_cat_ready_167 = _dataflow_cat_oready_167;

  always @(posedge CLK) begin
    if(RST) begin
      _dataflow_cat_data_167 <= 0;
      _dataflow_cat_valid_167 <= 0;
    end else begin
      if((_dataflow_cat_ready_167 || !_dataflow_cat_valid_167) && (_tmp_1347 && _tmp_1335 && _tmp_1323 && _tmp_1311) && (_tmp_1345 && _tmp_1333 && _tmp_1321 && _tmp_1309)) begin
        _dataflow_cat_data_167 <= { _tmp_1351, _tmp_1339, _tmp_1327, _tmp_1315 };
      end 
      if(_dataflow_cat_valid_167 && _dataflow_cat_ready_167) begin
        _dataflow_cat_valid_167 <= 0;
      end 
      if((_dataflow_cat_ready_167 || !_dataflow_cat_valid_167) && (_tmp_1347 && _tmp_1335 && _tmp_1323 && _tmp_1311)) begin
        _dataflow_cat_valid_167 <= _tmp_1345 && _tmp_1333 && _tmp_1321 && _tmp_1309;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id1_1_1_addr <= 0;
      _tmp_14 <= 0;
      ram_w8_l2048_id1_1_1_wdata <= 0;
      ram_w8_l2048_id1_1_1_wenable <= 0;
      _tmp_15 <= 0;
      _ram_w8_l2048_id1_1_cond_0_1 <= 0;
      ram_w8_l2048_id1_1_0_addr <= 0;
      _ram_w8_l2048_id1_1_cond_1_1 <= 0;
      _tmp_466 <= 0;
      _ram_w8_l2048_id1_1_cond_2_1 <= 0;
      _ram_w8_l2048_id1_1_cond_2_2 <= 0;
      _ram_w8_l2048_id1_1_cond_3_1 <= 0;
      _tmp_1029 <= 0;
      _ram_w8_l2048_id1_1_cond_4_1 <= 0;
      _ram_w8_l2048_id1_1_cond_4_2 <= 0;
      ram_w8_l2048_id1_1_0_wdata <= 0;
      ram_w8_l2048_id1_1_0_wenable <= 0;
      _ram_w8_l2048_id1_1_cond_5_1 <= 0;
      __tmp_1326_1 <= 0;
      __tmp_1327_1 <= 0;
      _tmp_1331 <= 0;
      _tmp_1321 <= 0;
      _tmp_1322 <= 0;
      _tmp_1329 <= 0;
      _tmp_1330 <= 0;
      _tmp_1328 <= 0;
      _tmp_1332 <= 0;
    end else begin
      if(_ram_w8_l2048_id1_1_cond_2_2) begin
        _tmp_466 <= 0;
      end 
      if(_ram_w8_l2048_id1_1_cond_4_2) begin
        _tmp_1029 <= 0;
      end 
      if(_ram_w8_l2048_id1_1_cond_0_1) begin
        ram_w8_l2048_id1_1_1_wenable <= 0;
        _tmp_15 <= 0;
      end 
      if(_ram_w8_l2048_id1_1_cond_1_1) begin
        _tmp_466 <= 1;
      end 
      _ram_w8_l2048_id1_1_cond_2_2 <= _ram_w8_l2048_id1_1_cond_2_1;
      if(_ram_w8_l2048_id1_1_cond_3_1) begin
        _tmp_1029 <= 1;
      end 
      _ram_w8_l2048_id1_1_cond_4_2 <= _ram_w8_l2048_id1_1_cond_4_1;
      if(_ram_w8_l2048_id1_1_cond_5_1) begin
        ram_w8_l2048_id1_1_0_wenable <= 0;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 1) && (_tmp_14 == 0)) begin
        ram_w8_l2048_id1_1_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_14 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_6 && ((_tmp_14 > 0) && !_tmp_15) && (_tmp_14 > 0)) begin
        ram_w8_l2048_id1_1_1_addr <= ram_w8_l2048_id1_1_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id1_1_1_wdata <= _dataflow_slice_odata_6;
        ram_w8_l2048_id1_1_1_wenable <= 1;
        _tmp_14 <= _tmp_14 - 1;
      end 
      if(_dataflow_slice_ovalid_6 && ((_tmp_14 > 0) && !_tmp_15) && (_tmp_14 == 1)) begin
        _tmp_15 <= 1;
      end 
      _ram_w8_l2048_id1_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1)) begin
        ram_w8_l2048_id1_1_0_addr <= _stream_conv2d_16_source_6_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id1_1_cond_1_1 <= _stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1);
      _ram_w8_l2048_id1_1_cond_2_1 <= _stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1);
      if(_stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1)) begin
        ram_w8_l2048_id1_1_0_addr <= _stream_max_pool_serial_18_source_1_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id1_1_cond_3_1 <= _stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1);
      _ram_w8_l2048_id1_1_cond_4_1 <= _stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1);
      if(_stream_matmul_29_sink_21_sink_wenable && (_stream_matmul_29_sink_21_sink_ram_sel == 5) && (_tmp_1225 == 1)) begin
        ram_w8_l2048_id1_1_0_addr <= _stream_matmul_29_sink_21_sink_waddr >> 2;
        ram_w8_l2048_id1_1_0_wdata <= _stream_matmul_29_sink_21_sink_wdata;
        ram_w8_l2048_id1_1_0_wenable <= 1;
      end 
      _ram_w8_l2048_id1_1_cond_5_1 <= _stream_matmul_29_sink_21_sink_wenable && (_stream_matmul_29_sink_21_sink_ram_sel == 5) && (_tmp_1225 == 1);
      __tmp_1326_1 <= _tmp_1326;
      __tmp_1327_1 <= _tmp_1327;
      if((_tmp_1323 || !_tmp_1321) && (_tmp_1324 || !_tmp_1322) && _tmp_1329) begin
        _tmp_1331 <= 0;
        _tmp_1321 <= 0;
        _tmp_1322 <= 0;
        _tmp_1329 <= 0;
      end 
      if((_tmp_1323 || !_tmp_1321) && (_tmp_1324 || !_tmp_1322) && _tmp_1328) begin
        _tmp_1321 <= 1;
        _tmp_1322 <= 1;
        _tmp_1331 <= _tmp_1330;
        _tmp_1330 <= 0;
        _tmp_1328 <= 0;
        _tmp_1329 <= 1;
      end 
      if(_maxi_write_start && (_maxi_write_op_sel == 3) && (_tmp_1332 == 0) && !_tmp_1330 && !_tmp_1331) begin
        ram_w8_l2048_id1_1_1_addr <= _maxi_write_local_addr;
        _tmp_1332 <= _maxi_write_size - 1;
        _tmp_1328 <= 1;
        _tmp_1330 <= _maxi_write_size == 1;
      end 
      if((_tmp_1323 || !_tmp_1321) && (_tmp_1324 || !_tmp_1322) && (_tmp_1332 > 0)) begin
        ram_w8_l2048_id1_1_1_addr <= ram_w8_l2048_id1_1_1_addr + _maxi_write_local_stride;
        _tmp_1332 <= _tmp_1332 - 1;
        _tmp_1328 <= 1;
        _tmp_1330 <= 0;
      end 
      if((_tmp_1323 || !_tmp_1321) && (_tmp_1324 || !_tmp_1322) && (_tmp_1332 == 1)) begin
        _tmp_1330 <= 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id1_2_1_addr <= 0;
      _tmp_16 <= 0;
      ram_w8_l2048_id1_2_1_wdata <= 0;
      ram_w8_l2048_id1_2_1_wenable <= 0;
      _tmp_17 <= 0;
      _ram_w8_l2048_id1_2_cond_0_1 <= 0;
      ram_w8_l2048_id1_2_0_addr <= 0;
      _ram_w8_l2048_id1_2_cond_1_1 <= 0;
      _tmp_467 <= 0;
      _ram_w8_l2048_id1_2_cond_2_1 <= 0;
      _ram_w8_l2048_id1_2_cond_2_2 <= 0;
      _ram_w8_l2048_id1_2_cond_3_1 <= 0;
      _tmp_1030 <= 0;
      _ram_w8_l2048_id1_2_cond_4_1 <= 0;
      _ram_w8_l2048_id1_2_cond_4_2 <= 0;
      ram_w8_l2048_id1_2_0_wdata <= 0;
      ram_w8_l2048_id1_2_0_wenable <= 0;
      _ram_w8_l2048_id1_2_cond_5_1 <= 0;
      __tmp_1338_1 <= 0;
      __tmp_1339_1 <= 0;
      _tmp_1343 <= 0;
      _tmp_1333 <= 0;
      _tmp_1334 <= 0;
      _tmp_1341 <= 0;
      _tmp_1342 <= 0;
      _tmp_1340 <= 0;
      _tmp_1344 <= 0;
    end else begin
      if(_ram_w8_l2048_id1_2_cond_2_2) begin
        _tmp_467 <= 0;
      end 
      if(_ram_w8_l2048_id1_2_cond_4_2) begin
        _tmp_1030 <= 0;
      end 
      if(_ram_w8_l2048_id1_2_cond_0_1) begin
        ram_w8_l2048_id1_2_1_wenable <= 0;
        _tmp_17 <= 0;
      end 
      if(_ram_w8_l2048_id1_2_cond_1_1) begin
        _tmp_467 <= 1;
      end 
      _ram_w8_l2048_id1_2_cond_2_2 <= _ram_w8_l2048_id1_2_cond_2_1;
      if(_ram_w8_l2048_id1_2_cond_3_1) begin
        _tmp_1030 <= 1;
      end 
      _ram_w8_l2048_id1_2_cond_4_2 <= _ram_w8_l2048_id1_2_cond_4_1;
      if(_ram_w8_l2048_id1_2_cond_5_1) begin
        ram_w8_l2048_id1_2_0_wenable <= 0;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 1) && (_tmp_16 == 0)) begin
        ram_w8_l2048_id1_2_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_16 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_9 && ((_tmp_16 > 0) && !_tmp_17) && (_tmp_16 > 0)) begin
        ram_w8_l2048_id1_2_1_addr <= ram_w8_l2048_id1_2_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id1_2_1_wdata <= _dataflow_slice_odata_9;
        ram_w8_l2048_id1_2_1_wenable <= 1;
        _tmp_16 <= _tmp_16 - 1;
      end 
      if(_dataflow_slice_ovalid_9 && ((_tmp_16 > 0) && !_tmp_17) && (_tmp_16 == 1)) begin
        _tmp_17 <= 1;
      end 
      _ram_w8_l2048_id1_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1)) begin
        ram_w8_l2048_id1_2_0_addr <= _stream_conv2d_16_source_6_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id1_2_cond_1_1 <= _stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1);
      _ram_w8_l2048_id1_2_cond_2_1 <= _stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1);
      if(_stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1)) begin
        ram_w8_l2048_id1_2_0_addr <= _stream_max_pool_serial_18_source_1_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id1_2_cond_3_1 <= _stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1);
      _ram_w8_l2048_id1_2_cond_4_1 <= _stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1);
      if(_stream_matmul_29_sink_21_sink_wenable && (_stream_matmul_29_sink_21_sink_ram_sel == 5) && (_tmp_1225 == 2)) begin
        ram_w8_l2048_id1_2_0_addr <= _stream_matmul_29_sink_21_sink_waddr >> 2;
        ram_w8_l2048_id1_2_0_wdata <= _stream_matmul_29_sink_21_sink_wdata;
        ram_w8_l2048_id1_2_0_wenable <= 1;
      end 
      _ram_w8_l2048_id1_2_cond_5_1 <= _stream_matmul_29_sink_21_sink_wenable && (_stream_matmul_29_sink_21_sink_ram_sel == 5) && (_tmp_1225 == 2);
      __tmp_1338_1 <= _tmp_1338;
      __tmp_1339_1 <= _tmp_1339;
      if((_tmp_1335 || !_tmp_1333) && (_tmp_1336 || !_tmp_1334) && _tmp_1341) begin
        _tmp_1343 <= 0;
        _tmp_1333 <= 0;
        _tmp_1334 <= 0;
        _tmp_1341 <= 0;
      end 
      if((_tmp_1335 || !_tmp_1333) && (_tmp_1336 || !_tmp_1334) && _tmp_1340) begin
        _tmp_1333 <= 1;
        _tmp_1334 <= 1;
        _tmp_1343 <= _tmp_1342;
        _tmp_1342 <= 0;
        _tmp_1340 <= 0;
        _tmp_1341 <= 1;
      end 
      if(_maxi_write_start && (_maxi_write_op_sel == 3) && (_tmp_1344 == 0) && !_tmp_1342 && !_tmp_1343) begin
        ram_w8_l2048_id1_2_1_addr <= _maxi_write_local_addr;
        _tmp_1344 <= _maxi_write_size - 1;
        _tmp_1340 <= 1;
        _tmp_1342 <= _maxi_write_size == 1;
      end 
      if((_tmp_1335 || !_tmp_1333) && (_tmp_1336 || !_tmp_1334) && (_tmp_1344 > 0)) begin
        ram_w8_l2048_id1_2_1_addr <= ram_w8_l2048_id1_2_1_addr + _maxi_write_local_stride;
        _tmp_1344 <= _tmp_1344 - 1;
        _tmp_1340 <= 1;
        _tmp_1342 <= 0;
      end 
      if((_tmp_1335 || !_tmp_1333) && (_tmp_1336 || !_tmp_1334) && (_tmp_1344 == 1)) begin
        _tmp_1342 <= 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id1_3_1_addr <= 0;
      _tmp_18 <= 0;
      ram_w8_l2048_id1_3_1_wdata <= 0;
      ram_w8_l2048_id1_3_1_wenable <= 0;
      _tmp_19 <= 0;
      _ram_w8_l2048_id1_3_cond_0_1 <= 0;
      ram_w8_l2048_id1_3_0_addr <= 0;
      _ram_w8_l2048_id1_3_cond_1_1 <= 0;
      _tmp_468 <= 0;
      _ram_w8_l2048_id1_3_cond_2_1 <= 0;
      _ram_w8_l2048_id1_3_cond_2_2 <= 0;
      _ram_w8_l2048_id1_3_cond_3_1 <= 0;
      _tmp_1031 <= 0;
      _ram_w8_l2048_id1_3_cond_4_1 <= 0;
      _ram_w8_l2048_id1_3_cond_4_2 <= 0;
      ram_w8_l2048_id1_3_0_wdata <= 0;
      ram_w8_l2048_id1_3_0_wenable <= 0;
      _ram_w8_l2048_id1_3_cond_5_1 <= 0;
      __tmp_1350_1 <= 0;
      __tmp_1351_1 <= 0;
      _tmp_1355 <= 0;
      _tmp_1345 <= 0;
      _tmp_1346 <= 0;
      _tmp_1353 <= 0;
      _tmp_1354 <= 0;
      _tmp_1352 <= 0;
      _tmp_1356 <= 0;
    end else begin
      if(_ram_w8_l2048_id1_3_cond_2_2) begin
        _tmp_468 <= 0;
      end 
      if(_ram_w8_l2048_id1_3_cond_4_2) begin
        _tmp_1031 <= 0;
      end 
      if(_ram_w8_l2048_id1_3_cond_0_1) begin
        ram_w8_l2048_id1_3_1_wenable <= 0;
        _tmp_19 <= 0;
      end 
      if(_ram_w8_l2048_id1_3_cond_1_1) begin
        _tmp_468 <= 1;
      end 
      _ram_w8_l2048_id1_3_cond_2_2 <= _ram_w8_l2048_id1_3_cond_2_1;
      if(_ram_w8_l2048_id1_3_cond_3_1) begin
        _tmp_1031 <= 1;
      end 
      _ram_w8_l2048_id1_3_cond_4_2 <= _ram_w8_l2048_id1_3_cond_4_1;
      if(_ram_w8_l2048_id1_3_cond_5_1) begin
        ram_w8_l2048_id1_3_0_wenable <= 0;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 1) && (_tmp_18 == 0)) begin
        ram_w8_l2048_id1_3_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_18 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_12 && ((_tmp_18 > 0) && !_tmp_19) && (_tmp_18 > 0)) begin
        ram_w8_l2048_id1_3_1_addr <= ram_w8_l2048_id1_3_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id1_3_1_wdata <= _dataflow_slice_odata_12;
        ram_w8_l2048_id1_3_1_wenable <= 1;
        _tmp_18 <= _tmp_18 - 1;
      end 
      if(_dataflow_slice_ovalid_12 && ((_tmp_18 > 0) && !_tmp_19) && (_tmp_18 == 1)) begin
        _tmp_19 <= 1;
      end 
      _ram_w8_l2048_id1_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1)) begin
        ram_w8_l2048_id1_3_0_addr <= _stream_conv2d_16_source_6_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id1_3_cond_1_1 <= _stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1);
      _ram_w8_l2048_id1_3_cond_2_1 <= _stream_conv2d_16_source_6_source_ram_renable && (_stream_conv2d_16_source_6_source_ram_sel == 1);
      if(_stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1)) begin
        ram_w8_l2048_id1_3_0_addr <= _stream_max_pool_serial_18_source_1_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id1_3_cond_3_1 <= _stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1);
      _ram_w8_l2048_id1_3_cond_4_1 <= _stream_max_pool_serial_18_source_1_source_ram_renable && (_stream_max_pool_serial_18_source_1_source_ram_sel == 1);
      if(_stream_matmul_29_sink_21_sink_wenable && (_stream_matmul_29_sink_21_sink_ram_sel == 5) && (_tmp_1225 == 3)) begin
        ram_w8_l2048_id1_3_0_addr <= _stream_matmul_29_sink_21_sink_waddr >> 2;
        ram_w8_l2048_id1_3_0_wdata <= _stream_matmul_29_sink_21_sink_wdata;
        ram_w8_l2048_id1_3_0_wenable <= 1;
      end 
      _ram_w8_l2048_id1_3_cond_5_1 <= _stream_matmul_29_sink_21_sink_wenable && (_stream_matmul_29_sink_21_sink_ram_sel == 5) && (_tmp_1225 == 3);
      __tmp_1350_1 <= _tmp_1350;
      __tmp_1351_1 <= _tmp_1351;
      if((_tmp_1347 || !_tmp_1345) && (_tmp_1348 || !_tmp_1346) && _tmp_1353) begin
        _tmp_1355 <= 0;
        _tmp_1345 <= 0;
        _tmp_1346 <= 0;
        _tmp_1353 <= 0;
      end 
      if((_tmp_1347 || !_tmp_1345) && (_tmp_1348 || !_tmp_1346) && _tmp_1352) begin
        _tmp_1345 <= 1;
        _tmp_1346 <= 1;
        _tmp_1355 <= _tmp_1354;
        _tmp_1354 <= 0;
        _tmp_1352 <= 0;
        _tmp_1353 <= 1;
      end 
      if(_maxi_write_start && (_maxi_write_op_sel == 3) && (_tmp_1356 == 0) && !_tmp_1354 && !_tmp_1355) begin
        ram_w8_l2048_id1_3_1_addr <= _maxi_write_local_addr;
        _tmp_1356 <= _maxi_write_size - 1;
        _tmp_1352 <= 1;
        _tmp_1354 <= _maxi_write_size == 1;
      end 
      if((_tmp_1347 || !_tmp_1345) && (_tmp_1348 || !_tmp_1346) && (_tmp_1356 > 0)) begin
        ram_w8_l2048_id1_3_1_addr <= ram_w8_l2048_id1_3_1_addr + _maxi_write_local_stride;
        _tmp_1356 <= _tmp_1356 - 1;
        _tmp_1352 <= 1;
        _tmp_1354 <= 0;
      end 
      if((_tmp_1347 || !_tmp_1345) && (_tmp_1348 || !_tmp_1346) && (_tmp_1356 == 1)) begin
        _tmp_1354 <= 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_303 <= 0;
      _tmp_291 <= 0;
      _tmp_292 <= 0;
      _tmp_294 <= 0;
      _tmp_295 <= 0;
      _tmp_296 <= 0;
      ram_w8_l2048_id2_0_1_addr <= 0;
      ram_w8_l2048_id2_0_1_wdata <= 0;
      ram_w8_l2048_id2_0_1_wenable <= 0;
      _tmp_293 <= 0;
      _ram_w8_l2048_id2_0_cond_0_1 <= 0;
      _ram_w8_l2048_id2_0_cond_1_1 <= 0;
      ram_w8_l2048_id2_0_0_addr <= 0;
      _ram_w8_l2048_id2_0_cond_2_1 <= 0;
      _tmp_496 <= 0;
      _ram_w8_l2048_id2_0_cond_3_1 <= 0;
      _ram_w8_l2048_id2_0_cond_3_2 <= 0;
      _tmp_1124 <= 0;
      _tmp_1125 <= 0;
      _ram_w8_l2048_id2_0_cond_4_1 <= 0;
      _ram_w8_l2048_id2_0_cond_5_1 <= 0;
      _tmp_1171 <= 0;
      _ram_w8_l2048_id2_0_cond_6_1 <= 0;
      _ram_w8_l2048_id2_0_cond_6_2 <= 0;
      ram_w8_l2048_id2_0_0_wdata <= 0;
      ram_w8_l2048_id2_0_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id2_0_cond_3_2) begin
        _tmp_496 <= 0;
      end 
      if(_ram_w8_l2048_id2_0_cond_6_2) begin
        _tmp_1171 <= 0;
      end 
      if(_ram_w8_l2048_id2_0_cond_0_1) begin
        _tmp_293 <= 0;
      end 
      if(_ram_w8_l2048_id2_0_cond_1_1) begin
        ram_w8_l2048_id2_0_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id2_0_cond_2_1) begin
        _tmp_496 <= 1;
      end 
      _ram_w8_l2048_id2_0_cond_3_2 <= _ram_w8_l2048_id2_0_cond_3_1;
      if(_ram_w8_l2048_id2_0_cond_4_1) begin
        ram_w8_l2048_id2_0_1_wenable <= 0;
        _tmp_1125 <= 0;
      end 
      if(_ram_w8_l2048_id2_0_cond_5_1) begin
        _tmp_1171 <= 1;
      end 
      _ram_w8_l2048_id2_0_cond_6_2 <= _ram_w8_l2048_id2_0_cond_6_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_292 == 0)) begin
        _tmp_303 <= 0;
        _tmp_291 <= req_block_size_286 - 1;
        _tmp_292 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_292 == 0)) begin
        _tmp_294 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_292 == 0)) begin
        _tmp_295 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_292 == 0)) begin
        _tmp_296 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_54 && ((_tmp_292 > 0) && !_tmp_293) && (_tmp_292 > 0)) begin
        _tmp_291 <= _tmp_291 - 1;
        _tmp_292 <= _tmp_292 - 1;
      end 
      if(_dataflow_slice_ovalid_54 && ((_tmp_292 > 0) && !_tmp_293) && (_tmp_292 > 0) && (_tmp_291 == 0)) begin
        _tmp_291 <= req_block_size_286 - 1;
        _tmp_303 <= _tmp_303 + 1;
      end 
      if(_dataflow_slice_ovalid_54 && ((_tmp_292 > 0) && !_tmp_293) && (_tmp_292 > 0) && (_tmp_291 == 0) && (_tmp_303 == 2)) begin
        _tmp_303 <= 0;
      end 
      if(_dataflow_slice_ovalid_54 && ((_tmp_292 > 0) && !_tmp_293) && (_tmp_292 > 0) && (_tmp_303 == 0)) begin
        _tmp_294 <= _tmp_297;
      end 
      if(_dataflow_slice_ovalid_54 && ((_tmp_292 > 0) && !_tmp_293) && (_tmp_292 > 0) && (_tmp_303 == 1)) begin
        _tmp_295 <= _tmp_298;
      end 
      if(_dataflow_slice_ovalid_54 && ((_tmp_292 > 0) && !_tmp_293) && (_tmp_292 > 0) && (_tmp_303 == 2)) begin
        _tmp_296 <= _tmp_299;
      end 
      if(_dataflow_slice_ovalid_54 && ((_tmp_292 > 0) && !_tmp_293) && (_tmp_292 > 0)) begin
        ram_w8_l2048_id2_0_1_addr <= _tmp_300;
        ram_w8_l2048_id2_0_1_wdata <= _dataflow_slice_odata_54;
        ram_w8_l2048_id2_0_1_wenable <= _tmp_303 == 0;
      end 
      if(_dataflow_slice_ovalid_54 && ((_tmp_292 > 0) && !_tmp_293) && (_tmp_292 == 1)) begin
        _tmp_293 <= 1;
      end 
      _ram_w8_l2048_id2_0_cond_0_1 <= 1;
      _ram_w8_l2048_id2_0_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3)) begin
        ram_w8_l2048_id2_0_0_addr <= _stream_conv2d_16_source_19_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id2_0_cond_2_1 <= _stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3);
      _ram_w8_l2048_id2_0_cond_3_1 <= _stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3);
      if(_maxi_read_start && (_maxi_read_op_sel == 7) && (_tmp_1124 == 0)) begin
        ram_w8_l2048_id2_0_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1124 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_111 && ((_tmp_1124 > 0) && !_tmp_1125) && (_tmp_1124 > 0)) begin
        ram_w8_l2048_id2_0_1_addr <= ram_w8_l2048_id2_0_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id2_0_1_wdata <= _dataflow_slice_odata_111;
        ram_w8_l2048_id2_0_1_wenable <= 1;
        _tmp_1124 <= _tmp_1124 - 1;
      end 
      if(_dataflow_slice_ovalid_111 && ((_tmp_1124 > 0) && !_tmp_1125) && (_tmp_1124 == 1)) begin
        _tmp_1125 <= 1;
      end 
      _ram_w8_l2048_id2_0_cond_4_1 <= 1;
      if(_stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1)) begin
        ram_w8_l2048_id2_0_0_addr <= _stream_matmul_29_source_6_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id2_0_cond_5_1 <= _stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1);
      _ram_w8_l2048_id2_0_cond_6_1 <= _stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1);
      ram_w8_l2048_id2_0_0_wdata <= 0;
      ram_w8_l2048_id2_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_316 <= 0;
      _tmp_304 <= 0;
      _tmp_305 <= 0;
      _tmp_307 <= 0;
      _tmp_308 <= 0;
      _tmp_309 <= 0;
      ram_w8_l2048_id2_1_1_addr <= 0;
      ram_w8_l2048_id2_1_1_wdata <= 0;
      ram_w8_l2048_id2_1_1_wenable <= 0;
      _tmp_306 <= 0;
      _ram_w8_l2048_id2_1_cond_0_1 <= 0;
      _ram_w8_l2048_id2_1_cond_1_1 <= 0;
      ram_w8_l2048_id2_1_0_addr <= 0;
      _ram_w8_l2048_id2_1_cond_2_1 <= 0;
      _tmp_497 <= 0;
      _ram_w8_l2048_id2_1_cond_3_1 <= 0;
      _ram_w8_l2048_id2_1_cond_3_2 <= 0;
      _tmp_1126 <= 0;
      _tmp_1127 <= 0;
      _ram_w8_l2048_id2_1_cond_4_1 <= 0;
      _ram_w8_l2048_id2_1_cond_5_1 <= 0;
      _tmp_1172 <= 0;
      _ram_w8_l2048_id2_1_cond_6_1 <= 0;
      _ram_w8_l2048_id2_1_cond_6_2 <= 0;
      ram_w8_l2048_id2_1_0_wdata <= 0;
      ram_w8_l2048_id2_1_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id2_1_cond_3_2) begin
        _tmp_497 <= 0;
      end 
      if(_ram_w8_l2048_id2_1_cond_6_2) begin
        _tmp_1172 <= 0;
      end 
      if(_ram_w8_l2048_id2_1_cond_0_1) begin
        _tmp_306 <= 0;
      end 
      if(_ram_w8_l2048_id2_1_cond_1_1) begin
        ram_w8_l2048_id2_1_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id2_1_cond_2_1) begin
        _tmp_497 <= 1;
      end 
      _ram_w8_l2048_id2_1_cond_3_2 <= _ram_w8_l2048_id2_1_cond_3_1;
      if(_ram_w8_l2048_id2_1_cond_4_1) begin
        ram_w8_l2048_id2_1_1_wenable <= 0;
        _tmp_1127 <= 0;
      end 
      if(_ram_w8_l2048_id2_1_cond_5_1) begin
        _tmp_1172 <= 1;
      end 
      _ram_w8_l2048_id2_1_cond_6_2 <= _ram_w8_l2048_id2_1_cond_6_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_305 == 0)) begin
        _tmp_316 <= 0;
        _tmp_304 <= req_block_size_286 - 1;
        _tmp_305 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_305 == 0)) begin
        _tmp_307 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_305 == 0)) begin
        _tmp_308 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_305 == 0)) begin
        _tmp_309 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_57 && ((_tmp_305 > 0) && !_tmp_306) && (_tmp_305 > 0)) begin
        _tmp_304 <= _tmp_304 - 1;
        _tmp_305 <= _tmp_305 - 1;
      end 
      if(_dataflow_slice_ovalid_57 && ((_tmp_305 > 0) && !_tmp_306) && (_tmp_305 > 0) && (_tmp_304 == 0)) begin
        _tmp_304 <= req_block_size_286 - 1;
        _tmp_316 <= _tmp_316 + 1;
      end 
      if(_dataflow_slice_ovalid_57 && ((_tmp_305 > 0) && !_tmp_306) && (_tmp_305 > 0) && (_tmp_304 == 0) && (_tmp_316 == 2)) begin
        _tmp_316 <= 0;
      end 
      if(_dataflow_slice_ovalid_57 && ((_tmp_305 > 0) && !_tmp_306) && (_tmp_305 > 0) && (_tmp_316 == 0)) begin
        _tmp_307 <= _tmp_310;
      end 
      if(_dataflow_slice_ovalid_57 && ((_tmp_305 > 0) && !_tmp_306) && (_tmp_305 > 0) && (_tmp_316 == 1)) begin
        _tmp_308 <= _tmp_311;
      end 
      if(_dataflow_slice_ovalid_57 && ((_tmp_305 > 0) && !_tmp_306) && (_tmp_305 > 0) && (_tmp_316 == 2)) begin
        _tmp_309 <= _tmp_312;
      end 
      if(_dataflow_slice_ovalid_57 && ((_tmp_305 > 0) && !_tmp_306) && (_tmp_305 > 0)) begin
        ram_w8_l2048_id2_1_1_addr <= _tmp_313;
        ram_w8_l2048_id2_1_1_wdata <= _dataflow_slice_odata_57;
        ram_w8_l2048_id2_1_1_wenable <= _tmp_316 == 0;
      end 
      if(_dataflow_slice_ovalid_57 && ((_tmp_305 > 0) && !_tmp_306) && (_tmp_305 == 1)) begin
        _tmp_306 <= 1;
      end 
      _ram_w8_l2048_id2_1_cond_0_1 <= 1;
      _ram_w8_l2048_id2_1_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3)) begin
        ram_w8_l2048_id2_1_0_addr <= _stream_conv2d_16_source_19_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id2_1_cond_2_1 <= _stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3);
      _ram_w8_l2048_id2_1_cond_3_1 <= _stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3);
      if(_maxi_read_start && (_maxi_read_op_sel == 7) && (_tmp_1126 == 0)) begin
        ram_w8_l2048_id2_1_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1126 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_114 && ((_tmp_1126 > 0) && !_tmp_1127) && (_tmp_1126 > 0)) begin
        ram_w8_l2048_id2_1_1_addr <= ram_w8_l2048_id2_1_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id2_1_1_wdata <= _dataflow_slice_odata_114;
        ram_w8_l2048_id2_1_1_wenable <= 1;
        _tmp_1126 <= _tmp_1126 - 1;
      end 
      if(_dataflow_slice_ovalid_114 && ((_tmp_1126 > 0) && !_tmp_1127) && (_tmp_1126 == 1)) begin
        _tmp_1127 <= 1;
      end 
      _ram_w8_l2048_id2_1_cond_4_1 <= 1;
      if(_stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1)) begin
        ram_w8_l2048_id2_1_0_addr <= _stream_matmul_29_source_6_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id2_1_cond_5_1 <= _stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1);
      _ram_w8_l2048_id2_1_cond_6_1 <= _stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1);
      ram_w8_l2048_id2_1_0_wdata <= 0;
      ram_w8_l2048_id2_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_329 <= 0;
      _tmp_317 <= 0;
      _tmp_318 <= 0;
      _tmp_320 <= 0;
      _tmp_321 <= 0;
      _tmp_322 <= 0;
      ram_w8_l2048_id2_2_1_addr <= 0;
      ram_w8_l2048_id2_2_1_wdata <= 0;
      ram_w8_l2048_id2_2_1_wenable <= 0;
      _tmp_319 <= 0;
      _ram_w8_l2048_id2_2_cond_0_1 <= 0;
      _ram_w8_l2048_id2_2_cond_1_1 <= 0;
      ram_w8_l2048_id2_2_0_addr <= 0;
      _ram_w8_l2048_id2_2_cond_2_1 <= 0;
      _tmp_498 <= 0;
      _ram_w8_l2048_id2_2_cond_3_1 <= 0;
      _ram_w8_l2048_id2_2_cond_3_2 <= 0;
      _tmp_1128 <= 0;
      _tmp_1129 <= 0;
      _ram_w8_l2048_id2_2_cond_4_1 <= 0;
      _ram_w8_l2048_id2_2_cond_5_1 <= 0;
      _tmp_1173 <= 0;
      _ram_w8_l2048_id2_2_cond_6_1 <= 0;
      _ram_w8_l2048_id2_2_cond_6_2 <= 0;
      ram_w8_l2048_id2_2_0_wdata <= 0;
      ram_w8_l2048_id2_2_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id2_2_cond_3_2) begin
        _tmp_498 <= 0;
      end 
      if(_ram_w8_l2048_id2_2_cond_6_2) begin
        _tmp_1173 <= 0;
      end 
      if(_ram_w8_l2048_id2_2_cond_0_1) begin
        _tmp_319 <= 0;
      end 
      if(_ram_w8_l2048_id2_2_cond_1_1) begin
        ram_w8_l2048_id2_2_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id2_2_cond_2_1) begin
        _tmp_498 <= 1;
      end 
      _ram_w8_l2048_id2_2_cond_3_2 <= _ram_w8_l2048_id2_2_cond_3_1;
      if(_ram_w8_l2048_id2_2_cond_4_1) begin
        ram_w8_l2048_id2_2_1_wenable <= 0;
        _tmp_1129 <= 0;
      end 
      if(_ram_w8_l2048_id2_2_cond_5_1) begin
        _tmp_1173 <= 1;
      end 
      _ram_w8_l2048_id2_2_cond_6_2 <= _ram_w8_l2048_id2_2_cond_6_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_318 == 0)) begin
        _tmp_329 <= 0;
        _tmp_317 <= req_block_size_286 - 1;
        _tmp_318 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_318 == 0)) begin
        _tmp_320 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_318 == 0)) begin
        _tmp_321 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_318 == 0)) begin
        _tmp_322 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_60 && ((_tmp_318 > 0) && !_tmp_319) && (_tmp_318 > 0)) begin
        _tmp_317 <= _tmp_317 - 1;
        _tmp_318 <= _tmp_318 - 1;
      end 
      if(_dataflow_slice_ovalid_60 && ((_tmp_318 > 0) && !_tmp_319) && (_tmp_318 > 0) && (_tmp_317 == 0)) begin
        _tmp_317 <= req_block_size_286 - 1;
        _tmp_329 <= _tmp_329 + 1;
      end 
      if(_dataflow_slice_ovalid_60 && ((_tmp_318 > 0) && !_tmp_319) && (_tmp_318 > 0) && (_tmp_317 == 0) && (_tmp_329 == 2)) begin
        _tmp_329 <= 0;
      end 
      if(_dataflow_slice_ovalid_60 && ((_tmp_318 > 0) && !_tmp_319) && (_tmp_318 > 0) && (_tmp_329 == 0)) begin
        _tmp_320 <= _tmp_323;
      end 
      if(_dataflow_slice_ovalid_60 && ((_tmp_318 > 0) && !_tmp_319) && (_tmp_318 > 0) && (_tmp_329 == 1)) begin
        _tmp_321 <= _tmp_324;
      end 
      if(_dataflow_slice_ovalid_60 && ((_tmp_318 > 0) && !_tmp_319) && (_tmp_318 > 0) && (_tmp_329 == 2)) begin
        _tmp_322 <= _tmp_325;
      end 
      if(_dataflow_slice_ovalid_60 && ((_tmp_318 > 0) && !_tmp_319) && (_tmp_318 > 0)) begin
        ram_w8_l2048_id2_2_1_addr <= _tmp_326;
        ram_w8_l2048_id2_2_1_wdata <= _dataflow_slice_odata_60;
        ram_w8_l2048_id2_2_1_wenable <= _tmp_329 == 0;
      end 
      if(_dataflow_slice_ovalid_60 && ((_tmp_318 > 0) && !_tmp_319) && (_tmp_318 == 1)) begin
        _tmp_319 <= 1;
      end 
      _ram_w8_l2048_id2_2_cond_0_1 <= 1;
      _ram_w8_l2048_id2_2_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3)) begin
        ram_w8_l2048_id2_2_0_addr <= _stream_conv2d_16_source_19_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id2_2_cond_2_1 <= _stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3);
      _ram_w8_l2048_id2_2_cond_3_1 <= _stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3);
      if(_maxi_read_start && (_maxi_read_op_sel == 7) && (_tmp_1128 == 0)) begin
        ram_w8_l2048_id2_2_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1128 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_117 && ((_tmp_1128 > 0) && !_tmp_1129) && (_tmp_1128 > 0)) begin
        ram_w8_l2048_id2_2_1_addr <= ram_w8_l2048_id2_2_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id2_2_1_wdata <= _dataflow_slice_odata_117;
        ram_w8_l2048_id2_2_1_wenable <= 1;
        _tmp_1128 <= _tmp_1128 - 1;
      end 
      if(_dataflow_slice_ovalid_117 && ((_tmp_1128 > 0) && !_tmp_1129) && (_tmp_1128 == 1)) begin
        _tmp_1129 <= 1;
      end 
      _ram_w8_l2048_id2_2_cond_4_1 <= 1;
      if(_stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1)) begin
        ram_w8_l2048_id2_2_0_addr <= _stream_matmul_29_source_6_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id2_2_cond_5_1 <= _stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1);
      _ram_w8_l2048_id2_2_cond_6_1 <= _stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1);
      ram_w8_l2048_id2_2_0_wdata <= 0;
      ram_w8_l2048_id2_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_342 <= 0;
      _tmp_330 <= 0;
      _tmp_331 <= 0;
      _tmp_333 <= 0;
      _tmp_334 <= 0;
      _tmp_335 <= 0;
      ram_w8_l2048_id2_3_1_addr <= 0;
      ram_w8_l2048_id2_3_1_wdata <= 0;
      ram_w8_l2048_id2_3_1_wenable <= 0;
      _tmp_332 <= 0;
      _ram_w8_l2048_id2_3_cond_0_1 <= 0;
      _ram_w8_l2048_id2_3_cond_1_1 <= 0;
      ram_w8_l2048_id2_3_0_addr <= 0;
      _ram_w8_l2048_id2_3_cond_2_1 <= 0;
      _tmp_499 <= 0;
      _ram_w8_l2048_id2_3_cond_3_1 <= 0;
      _ram_w8_l2048_id2_3_cond_3_2 <= 0;
      _tmp_1130 <= 0;
      _tmp_1131 <= 0;
      _ram_w8_l2048_id2_3_cond_4_1 <= 0;
      _ram_w8_l2048_id2_3_cond_5_1 <= 0;
      _tmp_1174 <= 0;
      _ram_w8_l2048_id2_3_cond_6_1 <= 0;
      _ram_w8_l2048_id2_3_cond_6_2 <= 0;
      ram_w8_l2048_id2_3_0_wdata <= 0;
      ram_w8_l2048_id2_3_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id2_3_cond_3_2) begin
        _tmp_499 <= 0;
      end 
      if(_ram_w8_l2048_id2_3_cond_6_2) begin
        _tmp_1174 <= 0;
      end 
      if(_ram_w8_l2048_id2_3_cond_0_1) begin
        _tmp_332 <= 0;
      end 
      if(_ram_w8_l2048_id2_3_cond_1_1) begin
        ram_w8_l2048_id2_3_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id2_3_cond_2_1) begin
        _tmp_499 <= 1;
      end 
      _ram_w8_l2048_id2_3_cond_3_2 <= _ram_w8_l2048_id2_3_cond_3_1;
      if(_ram_w8_l2048_id2_3_cond_4_1) begin
        ram_w8_l2048_id2_3_1_wenable <= 0;
        _tmp_1131 <= 0;
      end 
      if(_ram_w8_l2048_id2_3_cond_5_1) begin
        _tmp_1174 <= 1;
      end 
      _ram_w8_l2048_id2_3_cond_6_2 <= _ram_w8_l2048_id2_3_cond_6_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_331 == 0)) begin
        _tmp_342 <= 0;
        _tmp_330 <= req_block_size_286 - 1;
        _tmp_331 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_331 == 0)) begin
        _tmp_333 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_331 == 0)) begin
        _tmp_334 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 4) && (_tmp_331 == 0)) begin
        _tmp_335 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_63 && ((_tmp_331 > 0) && !_tmp_332) && (_tmp_331 > 0)) begin
        _tmp_330 <= _tmp_330 - 1;
        _tmp_331 <= _tmp_331 - 1;
      end 
      if(_dataflow_slice_ovalid_63 && ((_tmp_331 > 0) && !_tmp_332) && (_tmp_331 > 0) && (_tmp_330 == 0)) begin
        _tmp_330 <= req_block_size_286 - 1;
        _tmp_342 <= _tmp_342 + 1;
      end 
      if(_dataflow_slice_ovalid_63 && ((_tmp_331 > 0) && !_tmp_332) && (_tmp_331 > 0) && (_tmp_330 == 0) && (_tmp_342 == 2)) begin
        _tmp_342 <= 0;
      end 
      if(_dataflow_slice_ovalid_63 && ((_tmp_331 > 0) && !_tmp_332) && (_tmp_331 > 0) && (_tmp_342 == 0)) begin
        _tmp_333 <= _tmp_336;
      end 
      if(_dataflow_slice_ovalid_63 && ((_tmp_331 > 0) && !_tmp_332) && (_tmp_331 > 0) && (_tmp_342 == 1)) begin
        _tmp_334 <= _tmp_337;
      end 
      if(_dataflow_slice_ovalid_63 && ((_tmp_331 > 0) && !_tmp_332) && (_tmp_331 > 0) && (_tmp_342 == 2)) begin
        _tmp_335 <= _tmp_338;
      end 
      if(_dataflow_slice_ovalid_63 && ((_tmp_331 > 0) && !_tmp_332) && (_tmp_331 > 0)) begin
        ram_w8_l2048_id2_3_1_addr <= _tmp_339;
        ram_w8_l2048_id2_3_1_wdata <= _dataflow_slice_odata_63;
        ram_w8_l2048_id2_3_1_wenable <= _tmp_342 == 0;
      end 
      if(_dataflow_slice_ovalid_63 && ((_tmp_331 > 0) && !_tmp_332) && (_tmp_331 == 1)) begin
        _tmp_332 <= 1;
      end 
      _ram_w8_l2048_id2_3_cond_0_1 <= 1;
      _ram_w8_l2048_id2_3_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3)) begin
        ram_w8_l2048_id2_3_0_addr <= _stream_conv2d_16_source_19_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id2_3_cond_2_1 <= _stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3);
      _ram_w8_l2048_id2_3_cond_3_1 <= _stream_conv2d_16_source_19_source_ram_renable && (_stream_conv2d_16_source_19_source_ram_sel == 3);
      if(_maxi_read_start && (_maxi_read_op_sel == 7) && (_tmp_1130 == 0)) begin
        ram_w8_l2048_id2_3_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1130 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_120 && ((_tmp_1130 > 0) && !_tmp_1131) && (_tmp_1130 > 0)) begin
        ram_w8_l2048_id2_3_1_addr <= ram_w8_l2048_id2_3_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id2_3_1_wdata <= _dataflow_slice_odata_120;
        ram_w8_l2048_id2_3_1_wenable <= 1;
        _tmp_1130 <= _tmp_1130 - 1;
      end 
      if(_dataflow_slice_ovalid_120 && ((_tmp_1130 > 0) && !_tmp_1131) && (_tmp_1130 == 1)) begin
        _tmp_1131 <= 1;
      end 
      _ram_w8_l2048_id2_3_cond_4_1 <= 1;
      if(_stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1)) begin
        ram_w8_l2048_id2_3_0_addr <= _stream_matmul_29_source_6_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id2_3_cond_5_1 <= _stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1);
      _ram_w8_l2048_id2_3_cond_6_1 <= _stream_matmul_29_source_6_source_ram_renable && (_stream_matmul_29_source_6_source_ram_sel == 1);
      ram_w8_l2048_id2_3_0_wdata <= 0;
      ram_w8_l2048_id2_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id3_0_1_addr <= 0;
      ram_w8_l2048_id3_0_1_wdata <= 0;
      ram_w8_l2048_id3_0_1_wenable <= 0;
      _ram_w8_l2048_id3_0_cond_0_1 <= 0;
      ram_w8_l2048_id3_0_0_addr <= 0;
      _ram_w8_l2048_id3_0_cond_1_1 <= 0;
      _tmp_506 <= 0;
      _ram_w8_l2048_id3_0_cond_2_1 <= 0;
      _ram_w8_l2048_id3_0_cond_2_2 <= 0;
      _tmp_1155 <= 0;
      _tmp_1156 <= 0;
      _ram_w8_l2048_id3_0_cond_3_1 <= 0;
      _ram_w8_l2048_id3_0_cond_4_1 <= 0;
      _tmp_1202 <= 0;
      _ram_w8_l2048_id3_0_cond_5_1 <= 0;
      _ram_w8_l2048_id3_0_cond_5_2 <= 0;
      ram_w8_l2048_id3_0_0_wdata <= 0;
      ram_w8_l2048_id3_0_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id3_0_cond_2_2) begin
        _tmp_506 <= 0;
      end 
      if(_ram_w8_l2048_id3_0_cond_5_2) begin
        _tmp_1202 <= 0;
      end 
      if(_ram_w8_l2048_id3_0_cond_0_1) begin
        ram_w8_l2048_id3_0_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id3_0_cond_1_1) begin
        _tmp_506 <= 1;
      end 
      _ram_w8_l2048_id3_0_cond_2_2 <= _ram_w8_l2048_id3_0_cond_2_1;
      if(_ram_w8_l2048_id3_0_cond_3_1) begin
        ram_w8_l2048_id3_0_1_wenable <= 0;
        _tmp_1156 <= 0;
      end 
      if(_ram_w8_l2048_id3_0_cond_4_1) begin
        _tmp_1202 <= 1;
      end 
      _ram_w8_l2048_id3_0_cond_5_2 <= _ram_w8_l2048_id3_0_cond_5_1;
      if(_dataflow_slice_ovalid_54 && ((_tmp_292 > 0) && !_tmp_293) && (_tmp_292 > 0)) begin
        ram_w8_l2048_id3_0_1_addr <= _tmp_301;
        ram_w8_l2048_id3_0_1_wdata <= _dataflow_slice_odata_54;
        ram_w8_l2048_id3_0_1_wenable <= _tmp_303 == 1;
      end 
      _ram_w8_l2048_id3_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4)) begin
        ram_w8_l2048_id3_0_0_addr <= _stream_conv2d_16_source_20_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id3_0_cond_1_1 <= _stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4);
      _ram_w8_l2048_id3_0_cond_2_1 <= _stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4);
      if(_maxi_read_start && (_maxi_read_op_sel == 9) && (_tmp_1155 == 0)) begin
        ram_w8_l2048_id3_0_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1155 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_149 && ((_tmp_1155 > 0) && !_tmp_1156) && (_tmp_1155 > 0)) begin
        ram_w8_l2048_id3_0_1_addr <= ram_w8_l2048_id3_0_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id3_0_1_wdata <= _dataflow_slice_odata_149;
        ram_w8_l2048_id3_0_1_wenable <= 1;
        _tmp_1155 <= _tmp_1155 - 1;
      end 
      if(_dataflow_slice_ovalid_149 && ((_tmp_1155 > 0) && !_tmp_1156) && (_tmp_1155 == 1)) begin
        _tmp_1156 <= 1;
      end 
      _ram_w8_l2048_id3_0_cond_3_1 <= 1;
      if(_stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3)) begin
        ram_w8_l2048_id3_0_0_addr <= _stream_matmul_29_source_19_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id3_0_cond_4_1 <= _stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3);
      _ram_w8_l2048_id3_0_cond_5_1 <= _stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3);
      ram_w8_l2048_id3_0_0_wdata <= 0;
      ram_w8_l2048_id3_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id3_1_1_addr <= 0;
      ram_w8_l2048_id3_1_1_wdata <= 0;
      ram_w8_l2048_id3_1_1_wenable <= 0;
      _ram_w8_l2048_id3_1_cond_0_1 <= 0;
      ram_w8_l2048_id3_1_0_addr <= 0;
      _ram_w8_l2048_id3_1_cond_1_1 <= 0;
      _tmp_507 <= 0;
      _ram_w8_l2048_id3_1_cond_2_1 <= 0;
      _ram_w8_l2048_id3_1_cond_2_2 <= 0;
      _tmp_1157 <= 0;
      _tmp_1158 <= 0;
      _ram_w8_l2048_id3_1_cond_3_1 <= 0;
      _ram_w8_l2048_id3_1_cond_4_1 <= 0;
      _tmp_1203 <= 0;
      _ram_w8_l2048_id3_1_cond_5_1 <= 0;
      _ram_w8_l2048_id3_1_cond_5_2 <= 0;
      ram_w8_l2048_id3_1_0_wdata <= 0;
      ram_w8_l2048_id3_1_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id3_1_cond_2_2) begin
        _tmp_507 <= 0;
      end 
      if(_ram_w8_l2048_id3_1_cond_5_2) begin
        _tmp_1203 <= 0;
      end 
      if(_ram_w8_l2048_id3_1_cond_0_1) begin
        ram_w8_l2048_id3_1_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id3_1_cond_1_1) begin
        _tmp_507 <= 1;
      end 
      _ram_w8_l2048_id3_1_cond_2_2 <= _ram_w8_l2048_id3_1_cond_2_1;
      if(_ram_w8_l2048_id3_1_cond_3_1) begin
        ram_w8_l2048_id3_1_1_wenable <= 0;
        _tmp_1158 <= 0;
      end 
      if(_ram_w8_l2048_id3_1_cond_4_1) begin
        _tmp_1203 <= 1;
      end 
      _ram_w8_l2048_id3_1_cond_5_2 <= _ram_w8_l2048_id3_1_cond_5_1;
      if(_dataflow_slice_ovalid_57 && ((_tmp_305 > 0) && !_tmp_306) && (_tmp_305 > 0)) begin
        ram_w8_l2048_id3_1_1_addr <= _tmp_314;
        ram_w8_l2048_id3_1_1_wdata <= _dataflow_slice_odata_57;
        ram_w8_l2048_id3_1_1_wenable <= _tmp_316 == 1;
      end 
      _ram_w8_l2048_id3_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4)) begin
        ram_w8_l2048_id3_1_0_addr <= _stream_conv2d_16_source_20_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id3_1_cond_1_1 <= _stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4);
      _ram_w8_l2048_id3_1_cond_2_1 <= _stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4);
      if(_maxi_read_start && (_maxi_read_op_sel == 9) && (_tmp_1157 == 0)) begin
        ram_w8_l2048_id3_1_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1157 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_152 && ((_tmp_1157 > 0) && !_tmp_1158) && (_tmp_1157 > 0)) begin
        ram_w8_l2048_id3_1_1_addr <= ram_w8_l2048_id3_1_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id3_1_1_wdata <= _dataflow_slice_odata_152;
        ram_w8_l2048_id3_1_1_wenable <= 1;
        _tmp_1157 <= _tmp_1157 - 1;
      end 
      if(_dataflow_slice_ovalid_152 && ((_tmp_1157 > 0) && !_tmp_1158) && (_tmp_1157 == 1)) begin
        _tmp_1158 <= 1;
      end 
      _ram_w8_l2048_id3_1_cond_3_1 <= 1;
      if(_stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3)) begin
        ram_w8_l2048_id3_1_0_addr <= _stream_matmul_29_source_19_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id3_1_cond_4_1 <= _stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3);
      _ram_w8_l2048_id3_1_cond_5_1 <= _stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3);
      ram_w8_l2048_id3_1_0_wdata <= 0;
      ram_w8_l2048_id3_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id3_2_1_addr <= 0;
      ram_w8_l2048_id3_2_1_wdata <= 0;
      ram_w8_l2048_id3_2_1_wenable <= 0;
      _ram_w8_l2048_id3_2_cond_0_1 <= 0;
      ram_w8_l2048_id3_2_0_addr <= 0;
      _ram_w8_l2048_id3_2_cond_1_1 <= 0;
      _tmp_508 <= 0;
      _ram_w8_l2048_id3_2_cond_2_1 <= 0;
      _ram_w8_l2048_id3_2_cond_2_2 <= 0;
      _tmp_1159 <= 0;
      _tmp_1160 <= 0;
      _ram_w8_l2048_id3_2_cond_3_1 <= 0;
      _ram_w8_l2048_id3_2_cond_4_1 <= 0;
      _tmp_1204 <= 0;
      _ram_w8_l2048_id3_2_cond_5_1 <= 0;
      _ram_w8_l2048_id3_2_cond_5_2 <= 0;
      ram_w8_l2048_id3_2_0_wdata <= 0;
      ram_w8_l2048_id3_2_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id3_2_cond_2_2) begin
        _tmp_508 <= 0;
      end 
      if(_ram_w8_l2048_id3_2_cond_5_2) begin
        _tmp_1204 <= 0;
      end 
      if(_ram_w8_l2048_id3_2_cond_0_1) begin
        ram_w8_l2048_id3_2_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id3_2_cond_1_1) begin
        _tmp_508 <= 1;
      end 
      _ram_w8_l2048_id3_2_cond_2_2 <= _ram_w8_l2048_id3_2_cond_2_1;
      if(_ram_w8_l2048_id3_2_cond_3_1) begin
        ram_w8_l2048_id3_2_1_wenable <= 0;
        _tmp_1160 <= 0;
      end 
      if(_ram_w8_l2048_id3_2_cond_4_1) begin
        _tmp_1204 <= 1;
      end 
      _ram_w8_l2048_id3_2_cond_5_2 <= _ram_w8_l2048_id3_2_cond_5_1;
      if(_dataflow_slice_ovalid_60 && ((_tmp_318 > 0) && !_tmp_319) && (_tmp_318 > 0)) begin
        ram_w8_l2048_id3_2_1_addr <= _tmp_327;
        ram_w8_l2048_id3_2_1_wdata <= _dataflow_slice_odata_60;
        ram_w8_l2048_id3_2_1_wenable <= _tmp_329 == 1;
      end 
      _ram_w8_l2048_id3_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4)) begin
        ram_w8_l2048_id3_2_0_addr <= _stream_conv2d_16_source_20_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id3_2_cond_1_1 <= _stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4);
      _ram_w8_l2048_id3_2_cond_2_1 <= _stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4);
      if(_maxi_read_start && (_maxi_read_op_sel == 9) && (_tmp_1159 == 0)) begin
        ram_w8_l2048_id3_2_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1159 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_155 && ((_tmp_1159 > 0) && !_tmp_1160) && (_tmp_1159 > 0)) begin
        ram_w8_l2048_id3_2_1_addr <= ram_w8_l2048_id3_2_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id3_2_1_wdata <= _dataflow_slice_odata_155;
        ram_w8_l2048_id3_2_1_wenable <= 1;
        _tmp_1159 <= _tmp_1159 - 1;
      end 
      if(_dataflow_slice_ovalid_155 && ((_tmp_1159 > 0) && !_tmp_1160) && (_tmp_1159 == 1)) begin
        _tmp_1160 <= 1;
      end 
      _ram_w8_l2048_id3_2_cond_3_1 <= 1;
      if(_stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3)) begin
        ram_w8_l2048_id3_2_0_addr <= _stream_matmul_29_source_19_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id3_2_cond_4_1 <= _stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3);
      _ram_w8_l2048_id3_2_cond_5_1 <= _stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3);
      ram_w8_l2048_id3_2_0_wdata <= 0;
      ram_w8_l2048_id3_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id3_3_1_addr <= 0;
      ram_w8_l2048_id3_3_1_wdata <= 0;
      ram_w8_l2048_id3_3_1_wenable <= 0;
      _ram_w8_l2048_id3_3_cond_0_1 <= 0;
      ram_w8_l2048_id3_3_0_addr <= 0;
      _ram_w8_l2048_id3_3_cond_1_1 <= 0;
      _tmp_509 <= 0;
      _ram_w8_l2048_id3_3_cond_2_1 <= 0;
      _ram_w8_l2048_id3_3_cond_2_2 <= 0;
      _tmp_1161 <= 0;
      _tmp_1162 <= 0;
      _ram_w8_l2048_id3_3_cond_3_1 <= 0;
      _ram_w8_l2048_id3_3_cond_4_1 <= 0;
      _tmp_1205 <= 0;
      _ram_w8_l2048_id3_3_cond_5_1 <= 0;
      _ram_w8_l2048_id3_3_cond_5_2 <= 0;
      ram_w8_l2048_id3_3_0_wdata <= 0;
      ram_w8_l2048_id3_3_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id3_3_cond_2_2) begin
        _tmp_509 <= 0;
      end 
      if(_ram_w8_l2048_id3_3_cond_5_2) begin
        _tmp_1205 <= 0;
      end 
      if(_ram_w8_l2048_id3_3_cond_0_1) begin
        ram_w8_l2048_id3_3_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id3_3_cond_1_1) begin
        _tmp_509 <= 1;
      end 
      _ram_w8_l2048_id3_3_cond_2_2 <= _ram_w8_l2048_id3_3_cond_2_1;
      if(_ram_w8_l2048_id3_3_cond_3_1) begin
        ram_w8_l2048_id3_3_1_wenable <= 0;
        _tmp_1162 <= 0;
      end 
      if(_ram_w8_l2048_id3_3_cond_4_1) begin
        _tmp_1205 <= 1;
      end 
      _ram_w8_l2048_id3_3_cond_5_2 <= _ram_w8_l2048_id3_3_cond_5_1;
      if(_dataflow_slice_ovalid_63 && ((_tmp_331 > 0) && !_tmp_332) && (_tmp_331 > 0)) begin
        ram_w8_l2048_id3_3_1_addr <= _tmp_340;
        ram_w8_l2048_id3_3_1_wdata <= _dataflow_slice_odata_63;
        ram_w8_l2048_id3_3_1_wenable <= _tmp_342 == 1;
      end 
      _ram_w8_l2048_id3_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4)) begin
        ram_w8_l2048_id3_3_0_addr <= _stream_conv2d_16_source_20_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id3_3_cond_1_1 <= _stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4);
      _ram_w8_l2048_id3_3_cond_2_1 <= _stream_conv2d_16_source_20_source_ram_renable && (_stream_conv2d_16_source_20_source_ram_sel == 4);
      if(_maxi_read_start && (_maxi_read_op_sel == 9) && (_tmp_1161 == 0)) begin
        ram_w8_l2048_id3_3_1_addr <= _maxi_read_local_addr - _maxi_read_local_stride;
        _tmp_1161 <= _maxi_read_size;
      end 
      if(_dataflow_slice_ovalid_158 && ((_tmp_1161 > 0) && !_tmp_1162) && (_tmp_1161 > 0)) begin
        ram_w8_l2048_id3_3_1_addr <= ram_w8_l2048_id3_3_1_addr + _maxi_read_local_stride;
        ram_w8_l2048_id3_3_1_wdata <= _dataflow_slice_odata_158;
        ram_w8_l2048_id3_3_1_wenable <= 1;
        _tmp_1161 <= _tmp_1161 - 1;
      end 
      if(_dataflow_slice_ovalid_158 && ((_tmp_1161 > 0) && !_tmp_1162) && (_tmp_1161 == 1)) begin
        _tmp_1162 <= 1;
      end 
      _ram_w8_l2048_id3_3_cond_3_1 <= 1;
      if(_stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3)) begin
        ram_w8_l2048_id3_3_0_addr <= _stream_matmul_29_source_19_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id3_3_cond_4_1 <= _stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3);
      _ram_w8_l2048_id3_3_cond_5_1 <= _stream_matmul_29_source_19_source_ram_renable && (_stream_matmul_29_source_19_source_ram_sel == 3);
      ram_w8_l2048_id3_3_0_wdata <= 0;
      ram_w8_l2048_id3_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id4_0_1_addr <= 0;
      ram_w8_l2048_id4_0_1_wdata <= 0;
      ram_w8_l2048_id4_0_1_wenable <= 0;
      _ram_w8_l2048_id4_0_cond_0_1 <= 0;
      ram_w8_l2048_id4_0_0_addr <= 0;
      _ram_w8_l2048_id4_0_cond_1_1 <= 0;
      _tmp_516 <= 0;
      _ram_w8_l2048_id4_0_cond_2_1 <= 0;
      _ram_w8_l2048_id4_0_cond_2_2 <= 0;
      ram_w8_l2048_id4_0_0_wdata <= 0;
      ram_w8_l2048_id4_0_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id4_0_cond_2_2) begin
        _tmp_516 <= 0;
      end 
      if(_ram_w8_l2048_id4_0_cond_0_1) begin
        ram_w8_l2048_id4_0_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id4_0_cond_1_1) begin
        _tmp_516 <= 1;
      end 
      _ram_w8_l2048_id4_0_cond_2_2 <= _ram_w8_l2048_id4_0_cond_2_1;
      if(_dataflow_slice_ovalid_54 && ((_tmp_292 > 0) && !_tmp_293) && (_tmp_292 > 0)) begin
        ram_w8_l2048_id4_0_1_addr <= _tmp_302;
        ram_w8_l2048_id4_0_1_wdata <= _dataflow_slice_odata_54;
        ram_w8_l2048_id4_0_1_wenable <= _tmp_303 == 2;
      end 
      _ram_w8_l2048_id4_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5)) begin
        ram_w8_l2048_id4_0_0_addr <= _stream_conv2d_16_source_21_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id4_0_cond_1_1 <= _stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5);
      _ram_w8_l2048_id4_0_cond_2_1 <= _stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5);
      ram_w8_l2048_id4_0_0_wdata <= 0;
      ram_w8_l2048_id4_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id4_1_1_addr <= 0;
      ram_w8_l2048_id4_1_1_wdata <= 0;
      ram_w8_l2048_id4_1_1_wenable <= 0;
      _ram_w8_l2048_id4_1_cond_0_1 <= 0;
      ram_w8_l2048_id4_1_0_addr <= 0;
      _ram_w8_l2048_id4_1_cond_1_1 <= 0;
      _tmp_517 <= 0;
      _ram_w8_l2048_id4_1_cond_2_1 <= 0;
      _ram_w8_l2048_id4_1_cond_2_2 <= 0;
      ram_w8_l2048_id4_1_0_wdata <= 0;
      ram_w8_l2048_id4_1_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id4_1_cond_2_2) begin
        _tmp_517 <= 0;
      end 
      if(_ram_w8_l2048_id4_1_cond_0_1) begin
        ram_w8_l2048_id4_1_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id4_1_cond_1_1) begin
        _tmp_517 <= 1;
      end 
      _ram_w8_l2048_id4_1_cond_2_2 <= _ram_w8_l2048_id4_1_cond_2_1;
      if(_dataflow_slice_ovalid_57 && ((_tmp_305 > 0) && !_tmp_306) && (_tmp_305 > 0)) begin
        ram_w8_l2048_id4_1_1_addr <= _tmp_315;
        ram_w8_l2048_id4_1_1_wdata <= _dataflow_slice_odata_57;
        ram_w8_l2048_id4_1_1_wenable <= _tmp_316 == 2;
      end 
      _ram_w8_l2048_id4_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5)) begin
        ram_w8_l2048_id4_1_0_addr <= _stream_conv2d_16_source_21_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id4_1_cond_1_1 <= _stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5);
      _ram_w8_l2048_id4_1_cond_2_1 <= _stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5);
      ram_w8_l2048_id4_1_0_wdata <= 0;
      ram_w8_l2048_id4_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id4_2_1_addr <= 0;
      ram_w8_l2048_id4_2_1_wdata <= 0;
      ram_w8_l2048_id4_2_1_wenable <= 0;
      _ram_w8_l2048_id4_2_cond_0_1 <= 0;
      ram_w8_l2048_id4_2_0_addr <= 0;
      _ram_w8_l2048_id4_2_cond_1_1 <= 0;
      _tmp_518 <= 0;
      _ram_w8_l2048_id4_2_cond_2_1 <= 0;
      _ram_w8_l2048_id4_2_cond_2_2 <= 0;
      ram_w8_l2048_id4_2_0_wdata <= 0;
      ram_w8_l2048_id4_2_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id4_2_cond_2_2) begin
        _tmp_518 <= 0;
      end 
      if(_ram_w8_l2048_id4_2_cond_0_1) begin
        ram_w8_l2048_id4_2_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id4_2_cond_1_1) begin
        _tmp_518 <= 1;
      end 
      _ram_w8_l2048_id4_2_cond_2_2 <= _ram_w8_l2048_id4_2_cond_2_1;
      if(_dataflow_slice_ovalid_60 && ((_tmp_318 > 0) && !_tmp_319) && (_tmp_318 > 0)) begin
        ram_w8_l2048_id4_2_1_addr <= _tmp_328;
        ram_w8_l2048_id4_2_1_wdata <= _dataflow_slice_odata_60;
        ram_w8_l2048_id4_2_1_wenable <= _tmp_329 == 2;
      end 
      _ram_w8_l2048_id4_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5)) begin
        ram_w8_l2048_id4_2_0_addr <= _stream_conv2d_16_source_21_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id4_2_cond_1_1 <= _stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5);
      _ram_w8_l2048_id4_2_cond_2_1 <= _stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5);
      ram_w8_l2048_id4_2_0_wdata <= 0;
      ram_w8_l2048_id4_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id4_3_1_addr <= 0;
      ram_w8_l2048_id4_3_1_wdata <= 0;
      ram_w8_l2048_id4_3_1_wenable <= 0;
      _ram_w8_l2048_id4_3_cond_0_1 <= 0;
      ram_w8_l2048_id4_3_0_addr <= 0;
      _ram_w8_l2048_id4_3_cond_1_1 <= 0;
      _tmp_519 <= 0;
      _ram_w8_l2048_id4_3_cond_2_1 <= 0;
      _ram_w8_l2048_id4_3_cond_2_2 <= 0;
      ram_w8_l2048_id4_3_0_wdata <= 0;
      ram_w8_l2048_id4_3_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id4_3_cond_2_2) begin
        _tmp_519 <= 0;
      end 
      if(_ram_w8_l2048_id4_3_cond_0_1) begin
        ram_w8_l2048_id4_3_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id4_3_cond_1_1) begin
        _tmp_519 <= 1;
      end 
      _ram_w8_l2048_id4_3_cond_2_2 <= _ram_w8_l2048_id4_3_cond_2_1;
      if(_dataflow_slice_ovalid_63 && ((_tmp_331 > 0) && !_tmp_332) && (_tmp_331 > 0)) begin
        ram_w8_l2048_id4_3_1_addr <= _tmp_341;
        ram_w8_l2048_id4_3_1_wdata <= _dataflow_slice_odata_63;
        ram_w8_l2048_id4_3_1_wenable <= _tmp_342 == 2;
      end 
      _ram_w8_l2048_id4_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5)) begin
        ram_w8_l2048_id4_3_0_addr <= _stream_conv2d_16_source_21_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id4_3_cond_1_1 <= _stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5);
      _ram_w8_l2048_id4_3_cond_2_1 <= _stream_conv2d_16_source_21_source_ram_renable && (_stream_conv2d_16_source_21_source_ram_sel == 5);
      ram_w8_l2048_id4_3_0_wdata <= 0;
      ram_w8_l2048_id4_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_360 <= 0;
      _tmp_348 <= 0;
      _tmp_349 <= 0;
      _tmp_351 <= 0;
      _tmp_352 <= 0;
      _tmp_353 <= 0;
      ram_w8_l2048_id5_0_1_addr <= 0;
      ram_w8_l2048_id5_0_1_wdata <= 0;
      ram_w8_l2048_id5_0_1_wenable <= 0;
      _tmp_350 <= 0;
      _ram_w8_l2048_id5_0_cond_0_1 <= 0;
      _ram_w8_l2048_id5_0_cond_1_1 <= 0;
      ram_w8_l2048_id5_0_0_addr <= 0;
      _ram_w8_l2048_id5_0_cond_2_1 <= 0;
      _tmp_526 <= 0;
      _ram_w8_l2048_id5_0_cond_3_1 <= 0;
      _ram_w8_l2048_id5_0_cond_3_2 <= 0;
      ram_w8_l2048_id5_0_0_wdata <= 0;
      ram_w8_l2048_id5_0_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id5_0_cond_3_2) begin
        _tmp_526 <= 0;
      end 
      if(_ram_w8_l2048_id5_0_cond_0_1) begin
        _tmp_350 <= 0;
      end 
      if(_ram_w8_l2048_id5_0_cond_1_1) begin
        ram_w8_l2048_id5_0_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id5_0_cond_2_1) begin
        _tmp_526 <= 1;
      end 
      _ram_w8_l2048_id5_0_cond_3_2 <= _ram_w8_l2048_id5_0_cond_3_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_349 == 0)) begin
        _tmp_360 <= 0;
        _tmp_348 <= req_block_size_343 - 1;
        _tmp_349 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_349 == 0)) begin
        _tmp_351 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_349 == 0)) begin
        _tmp_352 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_349 == 0)) begin
        _tmp_353 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_67 && ((_tmp_349 > 0) && !_tmp_350) && (_tmp_349 > 0)) begin
        _tmp_348 <= _tmp_348 - 1;
        _tmp_349 <= _tmp_349 - 1;
      end 
      if(_dataflow_slice_ovalid_67 && ((_tmp_349 > 0) && !_tmp_350) && (_tmp_349 > 0) && (_tmp_348 == 0)) begin
        _tmp_348 <= req_block_size_343 - 1;
        _tmp_360 <= _tmp_360 + 1;
      end 
      if(_dataflow_slice_ovalid_67 && ((_tmp_349 > 0) && !_tmp_350) && (_tmp_349 > 0) && (_tmp_348 == 0) && (_tmp_360 == 2)) begin
        _tmp_360 <= 0;
      end 
      if(_dataflow_slice_ovalid_67 && ((_tmp_349 > 0) && !_tmp_350) && (_tmp_349 > 0) && (_tmp_360 == 0)) begin
        _tmp_351 <= _tmp_354;
      end 
      if(_dataflow_slice_ovalid_67 && ((_tmp_349 > 0) && !_tmp_350) && (_tmp_349 > 0) && (_tmp_360 == 1)) begin
        _tmp_352 <= _tmp_355;
      end 
      if(_dataflow_slice_ovalid_67 && ((_tmp_349 > 0) && !_tmp_350) && (_tmp_349 > 0) && (_tmp_360 == 2)) begin
        _tmp_353 <= _tmp_356;
      end 
      if(_dataflow_slice_ovalid_67 && ((_tmp_349 > 0) && !_tmp_350) && (_tmp_349 > 0)) begin
        ram_w8_l2048_id5_0_1_addr <= _tmp_357;
        ram_w8_l2048_id5_0_1_wdata <= _dataflow_slice_odata_67;
        ram_w8_l2048_id5_0_1_wenable <= _tmp_360 == 0;
      end 
      if(_dataflow_slice_ovalid_67 && ((_tmp_349 > 0) && !_tmp_350) && (_tmp_349 == 1)) begin
        _tmp_350 <= 1;
      end 
      _ram_w8_l2048_id5_0_cond_0_1 <= 1;
      _ram_w8_l2048_id5_0_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6)) begin
        ram_w8_l2048_id5_0_0_addr <= _stream_conv2d_16_source_22_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id5_0_cond_2_1 <= _stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6);
      _ram_w8_l2048_id5_0_cond_3_1 <= _stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6);
      ram_w8_l2048_id5_0_0_wdata <= 0;
      ram_w8_l2048_id5_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_373 <= 0;
      _tmp_361 <= 0;
      _tmp_362 <= 0;
      _tmp_364 <= 0;
      _tmp_365 <= 0;
      _tmp_366 <= 0;
      ram_w8_l2048_id5_1_1_addr <= 0;
      ram_w8_l2048_id5_1_1_wdata <= 0;
      ram_w8_l2048_id5_1_1_wenable <= 0;
      _tmp_363 <= 0;
      _ram_w8_l2048_id5_1_cond_0_1 <= 0;
      _ram_w8_l2048_id5_1_cond_1_1 <= 0;
      ram_w8_l2048_id5_1_0_addr <= 0;
      _ram_w8_l2048_id5_1_cond_2_1 <= 0;
      _tmp_527 <= 0;
      _ram_w8_l2048_id5_1_cond_3_1 <= 0;
      _ram_w8_l2048_id5_1_cond_3_2 <= 0;
      ram_w8_l2048_id5_1_0_wdata <= 0;
      ram_w8_l2048_id5_1_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id5_1_cond_3_2) begin
        _tmp_527 <= 0;
      end 
      if(_ram_w8_l2048_id5_1_cond_0_1) begin
        _tmp_363 <= 0;
      end 
      if(_ram_w8_l2048_id5_1_cond_1_1) begin
        ram_w8_l2048_id5_1_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id5_1_cond_2_1) begin
        _tmp_527 <= 1;
      end 
      _ram_w8_l2048_id5_1_cond_3_2 <= _ram_w8_l2048_id5_1_cond_3_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_362 == 0)) begin
        _tmp_373 <= 0;
        _tmp_361 <= req_block_size_343 - 1;
        _tmp_362 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_362 == 0)) begin
        _tmp_364 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_362 == 0)) begin
        _tmp_365 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_362 == 0)) begin
        _tmp_366 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_70 && ((_tmp_362 > 0) && !_tmp_363) && (_tmp_362 > 0)) begin
        _tmp_361 <= _tmp_361 - 1;
        _tmp_362 <= _tmp_362 - 1;
      end 
      if(_dataflow_slice_ovalid_70 && ((_tmp_362 > 0) && !_tmp_363) && (_tmp_362 > 0) && (_tmp_361 == 0)) begin
        _tmp_361 <= req_block_size_343 - 1;
        _tmp_373 <= _tmp_373 + 1;
      end 
      if(_dataflow_slice_ovalid_70 && ((_tmp_362 > 0) && !_tmp_363) && (_tmp_362 > 0) && (_tmp_361 == 0) && (_tmp_373 == 2)) begin
        _tmp_373 <= 0;
      end 
      if(_dataflow_slice_ovalid_70 && ((_tmp_362 > 0) && !_tmp_363) && (_tmp_362 > 0) && (_tmp_373 == 0)) begin
        _tmp_364 <= _tmp_367;
      end 
      if(_dataflow_slice_ovalid_70 && ((_tmp_362 > 0) && !_tmp_363) && (_tmp_362 > 0) && (_tmp_373 == 1)) begin
        _tmp_365 <= _tmp_368;
      end 
      if(_dataflow_slice_ovalid_70 && ((_tmp_362 > 0) && !_tmp_363) && (_tmp_362 > 0) && (_tmp_373 == 2)) begin
        _tmp_366 <= _tmp_369;
      end 
      if(_dataflow_slice_ovalid_70 && ((_tmp_362 > 0) && !_tmp_363) && (_tmp_362 > 0)) begin
        ram_w8_l2048_id5_1_1_addr <= _tmp_370;
        ram_w8_l2048_id5_1_1_wdata <= _dataflow_slice_odata_70;
        ram_w8_l2048_id5_1_1_wenable <= _tmp_373 == 0;
      end 
      if(_dataflow_slice_ovalid_70 && ((_tmp_362 > 0) && !_tmp_363) && (_tmp_362 == 1)) begin
        _tmp_363 <= 1;
      end 
      _ram_w8_l2048_id5_1_cond_0_1 <= 1;
      _ram_w8_l2048_id5_1_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6)) begin
        ram_w8_l2048_id5_1_0_addr <= _stream_conv2d_16_source_22_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id5_1_cond_2_1 <= _stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6);
      _ram_w8_l2048_id5_1_cond_3_1 <= _stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6);
      ram_w8_l2048_id5_1_0_wdata <= 0;
      ram_w8_l2048_id5_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_386 <= 0;
      _tmp_374 <= 0;
      _tmp_375 <= 0;
      _tmp_377 <= 0;
      _tmp_378 <= 0;
      _tmp_379 <= 0;
      ram_w8_l2048_id5_2_1_addr <= 0;
      ram_w8_l2048_id5_2_1_wdata <= 0;
      ram_w8_l2048_id5_2_1_wenable <= 0;
      _tmp_376 <= 0;
      _ram_w8_l2048_id5_2_cond_0_1 <= 0;
      _ram_w8_l2048_id5_2_cond_1_1 <= 0;
      ram_w8_l2048_id5_2_0_addr <= 0;
      _ram_w8_l2048_id5_2_cond_2_1 <= 0;
      _tmp_528 <= 0;
      _ram_w8_l2048_id5_2_cond_3_1 <= 0;
      _ram_w8_l2048_id5_2_cond_3_2 <= 0;
      ram_w8_l2048_id5_2_0_wdata <= 0;
      ram_w8_l2048_id5_2_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id5_2_cond_3_2) begin
        _tmp_528 <= 0;
      end 
      if(_ram_w8_l2048_id5_2_cond_0_1) begin
        _tmp_376 <= 0;
      end 
      if(_ram_w8_l2048_id5_2_cond_1_1) begin
        ram_w8_l2048_id5_2_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id5_2_cond_2_1) begin
        _tmp_528 <= 1;
      end 
      _ram_w8_l2048_id5_2_cond_3_2 <= _ram_w8_l2048_id5_2_cond_3_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_375 == 0)) begin
        _tmp_386 <= 0;
        _tmp_374 <= req_block_size_343 - 1;
        _tmp_375 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_375 == 0)) begin
        _tmp_377 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_375 == 0)) begin
        _tmp_378 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_375 == 0)) begin
        _tmp_379 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_73 && ((_tmp_375 > 0) && !_tmp_376) && (_tmp_375 > 0)) begin
        _tmp_374 <= _tmp_374 - 1;
        _tmp_375 <= _tmp_375 - 1;
      end 
      if(_dataflow_slice_ovalid_73 && ((_tmp_375 > 0) && !_tmp_376) && (_tmp_375 > 0) && (_tmp_374 == 0)) begin
        _tmp_374 <= req_block_size_343 - 1;
        _tmp_386 <= _tmp_386 + 1;
      end 
      if(_dataflow_slice_ovalid_73 && ((_tmp_375 > 0) && !_tmp_376) && (_tmp_375 > 0) && (_tmp_374 == 0) && (_tmp_386 == 2)) begin
        _tmp_386 <= 0;
      end 
      if(_dataflow_slice_ovalid_73 && ((_tmp_375 > 0) && !_tmp_376) && (_tmp_375 > 0) && (_tmp_386 == 0)) begin
        _tmp_377 <= _tmp_380;
      end 
      if(_dataflow_slice_ovalid_73 && ((_tmp_375 > 0) && !_tmp_376) && (_tmp_375 > 0) && (_tmp_386 == 1)) begin
        _tmp_378 <= _tmp_381;
      end 
      if(_dataflow_slice_ovalid_73 && ((_tmp_375 > 0) && !_tmp_376) && (_tmp_375 > 0) && (_tmp_386 == 2)) begin
        _tmp_379 <= _tmp_382;
      end 
      if(_dataflow_slice_ovalid_73 && ((_tmp_375 > 0) && !_tmp_376) && (_tmp_375 > 0)) begin
        ram_w8_l2048_id5_2_1_addr <= _tmp_383;
        ram_w8_l2048_id5_2_1_wdata <= _dataflow_slice_odata_73;
        ram_w8_l2048_id5_2_1_wenable <= _tmp_386 == 0;
      end 
      if(_dataflow_slice_ovalid_73 && ((_tmp_375 > 0) && !_tmp_376) && (_tmp_375 == 1)) begin
        _tmp_376 <= 1;
      end 
      _ram_w8_l2048_id5_2_cond_0_1 <= 1;
      _ram_w8_l2048_id5_2_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6)) begin
        ram_w8_l2048_id5_2_0_addr <= _stream_conv2d_16_source_22_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id5_2_cond_2_1 <= _stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6);
      _ram_w8_l2048_id5_2_cond_3_1 <= _stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6);
      ram_w8_l2048_id5_2_0_wdata <= 0;
      ram_w8_l2048_id5_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_399 <= 0;
      _tmp_387 <= 0;
      _tmp_388 <= 0;
      _tmp_390 <= 0;
      _tmp_391 <= 0;
      _tmp_392 <= 0;
      ram_w8_l2048_id5_3_1_addr <= 0;
      ram_w8_l2048_id5_3_1_wdata <= 0;
      ram_w8_l2048_id5_3_1_wenable <= 0;
      _tmp_389 <= 0;
      _ram_w8_l2048_id5_3_cond_0_1 <= 0;
      _ram_w8_l2048_id5_3_cond_1_1 <= 0;
      ram_w8_l2048_id5_3_0_addr <= 0;
      _ram_w8_l2048_id5_3_cond_2_1 <= 0;
      _tmp_529 <= 0;
      _ram_w8_l2048_id5_3_cond_3_1 <= 0;
      _ram_w8_l2048_id5_3_cond_3_2 <= 0;
      ram_w8_l2048_id5_3_0_wdata <= 0;
      ram_w8_l2048_id5_3_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id5_3_cond_3_2) begin
        _tmp_529 <= 0;
      end 
      if(_ram_w8_l2048_id5_3_cond_0_1) begin
        _tmp_389 <= 0;
      end 
      if(_ram_w8_l2048_id5_3_cond_1_1) begin
        ram_w8_l2048_id5_3_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id5_3_cond_2_1) begin
        _tmp_529 <= 1;
      end 
      _ram_w8_l2048_id5_3_cond_3_2 <= _ram_w8_l2048_id5_3_cond_3_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_388 == 0)) begin
        _tmp_399 <= 0;
        _tmp_387 <= req_block_size_343 - 1;
        _tmp_388 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_388 == 0)) begin
        _tmp_390 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_388 == 0)) begin
        _tmp_391 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 5) && (_tmp_388 == 0)) begin
        _tmp_392 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_76 && ((_tmp_388 > 0) && !_tmp_389) && (_tmp_388 > 0)) begin
        _tmp_387 <= _tmp_387 - 1;
        _tmp_388 <= _tmp_388 - 1;
      end 
      if(_dataflow_slice_ovalid_76 && ((_tmp_388 > 0) && !_tmp_389) && (_tmp_388 > 0) && (_tmp_387 == 0)) begin
        _tmp_387 <= req_block_size_343 - 1;
        _tmp_399 <= _tmp_399 + 1;
      end 
      if(_dataflow_slice_ovalid_76 && ((_tmp_388 > 0) && !_tmp_389) && (_tmp_388 > 0) && (_tmp_387 == 0) && (_tmp_399 == 2)) begin
        _tmp_399 <= 0;
      end 
      if(_dataflow_slice_ovalid_76 && ((_tmp_388 > 0) && !_tmp_389) && (_tmp_388 > 0) && (_tmp_399 == 0)) begin
        _tmp_390 <= _tmp_393;
      end 
      if(_dataflow_slice_ovalid_76 && ((_tmp_388 > 0) && !_tmp_389) && (_tmp_388 > 0) && (_tmp_399 == 1)) begin
        _tmp_391 <= _tmp_394;
      end 
      if(_dataflow_slice_ovalid_76 && ((_tmp_388 > 0) && !_tmp_389) && (_tmp_388 > 0) && (_tmp_399 == 2)) begin
        _tmp_392 <= _tmp_395;
      end 
      if(_dataflow_slice_ovalid_76 && ((_tmp_388 > 0) && !_tmp_389) && (_tmp_388 > 0)) begin
        ram_w8_l2048_id5_3_1_addr <= _tmp_396;
        ram_w8_l2048_id5_3_1_wdata <= _dataflow_slice_odata_76;
        ram_w8_l2048_id5_3_1_wenable <= _tmp_399 == 0;
      end 
      if(_dataflow_slice_ovalid_76 && ((_tmp_388 > 0) && !_tmp_389) && (_tmp_388 == 1)) begin
        _tmp_389 <= 1;
      end 
      _ram_w8_l2048_id5_3_cond_0_1 <= 1;
      _ram_w8_l2048_id5_3_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6)) begin
        ram_w8_l2048_id5_3_0_addr <= _stream_conv2d_16_source_22_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id5_3_cond_2_1 <= _stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6);
      _ram_w8_l2048_id5_3_cond_3_1 <= _stream_conv2d_16_source_22_source_ram_renable && (_stream_conv2d_16_source_22_source_ram_sel == 6);
      ram_w8_l2048_id5_3_0_wdata <= 0;
      ram_w8_l2048_id5_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id6_0_1_addr <= 0;
      ram_w8_l2048_id6_0_1_wdata <= 0;
      ram_w8_l2048_id6_0_1_wenable <= 0;
      _ram_w8_l2048_id6_0_cond_0_1 <= 0;
      ram_w8_l2048_id6_0_0_addr <= 0;
      _ram_w8_l2048_id6_0_cond_1_1 <= 0;
      _tmp_536 <= 0;
      _ram_w8_l2048_id6_0_cond_2_1 <= 0;
      _ram_w8_l2048_id6_0_cond_2_2 <= 0;
      ram_w8_l2048_id6_0_0_wdata <= 0;
      ram_w8_l2048_id6_0_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id6_0_cond_2_2) begin
        _tmp_536 <= 0;
      end 
      if(_ram_w8_l2048_id6_0_cond_0_1) begin
        ram_w8_l2048_id6_0_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id6_0_cond_1_1) begin
        _tmp_536 <= 1;
      end 
      _ram_w8_l2048_id6_0_cond_2_2 <= _ram_w8_l2048_id6_0_cond_2_1;
      if(_dataflow_slice_ovalid_67 && ((_tmp_349 > 0) && !_tmp_350) && (_tmp_349 > 0)) begin
        ram_w8_l2048_id6_0_1_addr <= _tmp_358;
        ram_w8_l2048_id6_0_1_wdata <= _dataflow_slice_odata_67;
        ram_w8_l2048_id6_0_1_wenable <= _tmp_360 == 1;
      end 
      _ram_w8_l2048_id6_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7)) begin
        ram_w8_l2048_id6_0_0_addr <= _stream_conv2d_16_source_23_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id6_0_cond_1_1 <= _stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7);
      _ram_w8_l2048_id6_0_cond_2_1 <= _stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7);
      ram_w8_l2048_id6_0_0_wdata <= 0;
      ram_w8_l2048_id6_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id6_1_1_addr <= 0;
      ram_w8_l2048_id6_1_1_wdata <= 0;
      ram_w8_l2048_id6_1_1_wenable <= 0;
      _ram_w8_l2048_id6_1_cond_0_1 <= 0;
      ram_w8_l2048_id6_1_0_addr <= 0;
      _ram_w8_l2048_id6_1_cond_1_1 <= 0;
      _tmp_537 <= 0;
      _ram_w8_l2048_id6_1_cond_2_1 <= 0;
      _ram_w8_l2048_id6_1_cond_2_2 <= 0;
      ram_w8_l2048_id6_1_0_wdata <= 0;
      ram_w8_l2048_id6_1_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id6_1_cond_2_2) begin
        _tmp_537 <= 0;
      end 
      if(_ram_w8_l2048_id6_1_cond_0_1) begin
        ram_w8_l2048_id6_1_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id6_1_cond_1_1) begin
        _tmp_537 <= 1;
      end 
      _ram_w8_l2048_id6_1_cond_2_2 <= _ram_w8_l2048_id6_1_cond_2_1;
      if(_dataflow_slice_ovalid_70 && ((_tmp_362 > 0) && !_tmp_363) && (_tmp_362 > 0)) begin
        ram_w8_l2048_id6_1_1_addr <= _tmp_371;
        ram_w8_l2048_id6_1_1_wdata <= _dataflow_slice_odata_70;
        ram_w8_l2048_id6_1_1_wenable <= _tmp_373 == 1;
      end 
      _ram_w8_l2048_id6_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7)) begin
        ram_w8_l2048_id6_1_0_addr <= _stream_conv2d_16_source_23_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id6_1_cond_1_1 <= _stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7);
      _ram_w8_l2048_id6_1_cond_2_1 <= _stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7);
      ram_w8_l2048_id6_1_0_wdata <= 0;
      ram_w8_l2048_id6_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id6_2_1_addr <= 0;
      ram_w8_l2048_id6_2_1_wdata <= 0;
      ram_w8_l2048_id6_2_1_wenable <= 0;
      _ram_w8_l2048_id6_2_cond_0_1 <= 0;
      ram_w8_l2048_id6_2_0_addr <= 0;
      _ram_w8_l2048_id6_2_cond_1_1 <= 0;
      _tmp_538 <= 0;
      _ram_w8_l2048_id6_2_cond_2_1 <= 0;
      _ram_w8_l2048_id6_2_cond_2_2 <= 0;
      ram_w8_l2048_id6_2_0_wdata <= 0;
      ram_w8_l2048_id6_2_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id6_2_cond_2_2) begin
        _tmp_538 <= 0;
      end 
      if(_ram_w8_l2048_id6_2_cond_0_1) begin
        ram_w8_l2048_id6_2_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id6_2_cond_1_1) begin
        _tmp_538 <= 1;
      end 
      _ram_w8_l2048_id6_2_cond_2_2 <= _ram_w8_l2048_id6_2_cond_2_1;
      if(_dataflow_slice_ovalid_73 && ((_tmp_375 > 0) && !_tmp_376) && (_tmp_375 > 0)) begin
        ram_w8_l2048_id6_2_1_addr <= _tmp_384;
        ram_w8_l2048_id6_2_1_wdata <= _dataflow_slice_odata_73;
        ram_w8_l2048_id6_2_1_wenable <= _tmp_386 == 1;
      end 
      _ram_w8_l2048_id6_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7)) begin
        ram_w8_l2048_id6_2_0_addr <= _stream_conv2d_16_source_23_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id6_2_cond_1_1 <= _stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7);
      _ram_w8_l2048_id6_2_cond_2_1 <= _stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7);
      ram_w8_l2048_id6_2_0_wdata <= 0;
      ram_w8_l2048_id6_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id6_3_1_addr <= 0;
      ram_w8_l2048_id6_3_1_wdata <= 0;
      ram_w8_l2048_id6_3_1_wenable <= 0;
      _ram_w8_l2048_id6_3_cond_0_1 <= 0;
      ram_w8_l2048_id6_3_0_addr <= 0;
      _ram_w8_l2048_id6_3_cond_1_1 <= 0;
      _tmp_539 <= 0;
      _ram_w8_l2048_id6_3_cond_2_1 <= 0;
      _ram_w8_l2048_id6_3_cond_2_2 <= 0;
      ram_w8_l2048_id6_3_0_wdata <= 0;
      ram_w8_l2048_id6_3_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id6_3_cond_2_2) begin
        _tmp_539 <= 0;
      end 
      if(_ram_w8_l2048_id6_3_cond_0_1) begin
        ram_w8_l2048_id6_3_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id6_3_cond_1_1) begin
        _tmp_539 <= 1;
      end 
      _ram_w8_l2048_id6_3_cond_2_2 <= _ram_w8_l2048_id6_3_cond_2_1;
      if(_dataflow_slice_ovalid_76 && ((_tmp_388 > 0) && !_tmp_389) && (_tmp_388 > 0)) begin
        ram_w8_l2048_id6_3_1_addr <= _tmp_397;
        ram_w8_l2048_id6_3_1_wdata <= _dataflow_slice_odata_76;
        ram_w8_l2048_id6_3_1_wenable <= _tmp_399 == 1;
      end 
      _ram_w8_l2048_id6_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7)) begin
        ram_w8_l2048_id6_3_0_addr <= _stream_conv2d_16_source_23_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id6_3_cond_1_1 <= _stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7);
      _ram_w8_l2048_id6_3_cond_2_1 <= _stream_conv2d_16_source_23_source_ram_renable && (_stream_conv2d_16_source_23_source_ram_sel == 7);
      ram_w8_l2048_id6_3_0_wdata <= 0;
      ram_w8_l2048_id6_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id7_0_1_addr <= 0;
      ram_w8_l2048_id7_0_1_wdata <= 0;
      ram_w8_l2048_id7_0_1_wenable <= 0;
      _ram_w8_l2048_id7_0_cond_0_1 <= 0;
      ram_w8_l2048_id7_0_0_addr <= 0;
      _ram_w8_l2048_id7_0_cond_1_1 <= 0;
      _tmp_546 <= 0;
      _ram_w8_l2048_id7_0_cond_2_1 <= 0;
      _ram_w8_l2048_id7_0_cond_2_2 <= 0;
      ram_w8_l2048_id7_0_0_wdata <= 0;
      ram_w8_l2048_id7_0_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id7_0_cond_2_2) begin
        _tmp_546 <= 0;
      end 
      if(_ram_w8_l2048_id7_0_cond_0_1) begin
        ram_w8_l2048_id7_0_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id7_0_cond_1_1) begin
        _tmp_546 <= 1;
      end 
      _ram_w8_l2048_id7_0_cond_2_2 <= _ram_w8_l2048_id7_0_cond_2_1;
      if(_dataflow_slice_ovalid_67 && ((_tmp_349 > 0) && !_tmp_350) && (_tmp_349 > 0)) begin
        ram_w8_l2048_id7_0_1_addr <= _tmp_359;
        ram_w8_l2048_id7_0_1_wdata <= _dataflow_slice_odata_67;
        ram_w8_l2048_id7_0_1_wenable <= _tmp_360 == 2;
      end 
      _ram_w8_l2048_id7_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8)) begin
        ram_w8_l2048_id7_0_0_addr <= _stream_conv2d_16_source_24_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id7_0_cond_1_1 <= _stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8);
      _ram_w8_l2048_id7_0_cond_2_1 <= _stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8);
      ram_w8_l2048_id7_0_0_wdata <= 0;
      ram_w8_l2048_id7_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id7_1_1_addr <= 0;
      ram_w8_l2048_id7_1_1_wdata <= 0;
      ram_w8_l2048_id7_1_1_wenable <= 0;
      _ram_w8_l2048_id7_1_cond_0_1 <= 0;
      ram_w8_l2048_id7_1_0_addr <= 0;
      _ram_w8_l2048_id7_1_cond_1_1 <= 0;
      _tmp_547 <= 0;
      _ram_w8_l2048_id7_1_cond_2_1 <= 0;
      _ram_w8_l2048_id7_1_cond_2_2 <= 0;
      ram_w8_l2048_id7_1_0_wdata <= 0;
      ram_w8_l2048_id7_1_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id7_1_cond_2_2) begin
        _tmp_547 <= 0;
      end 
      if(_ram_w8_l2048_id7_1_cond_0_1) begin
        ram_w8_l2048_id7_1_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id7_1_cond_1_1) begin
        _tmp_547 <= 1;
      end 
      _ram_w8_l2048_id7_1_cond_2_2 <= _ram_w8_l2048_id7_1_cond_2_1;
      if(_dataflow_slice_ovalid_70 && ((_tmp_362 > 0) && !_tmp_363) && (_tmp_362 > 0)) begin
        ram_w8_l2048_id7_1_1_addr <= _tmp_372;
        ram_w8_l2048_id7_1_1_wdata <= _dataflow_slice_odata_70;
        ram_w8_l2048_id7_1_1_wenable <= _tmp_373 == 2;
      end 
      _ram_w8_l2048_id7_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8)) begin
        ram_w8_l2048_id7_1_0_addr <= _stream_conv2d_16_source_24_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id7_1_cond_1_1 <= _stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8);
      _ram_w8_l2048_id7_1_cond_2_1 <= _stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8);
      ram_w8_l2048_id7_1_0_wdata <= 0;
      ram_w8_l2048_id7_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id7_2_1_addr <= 0;
      ram_w8_l2048_id7_2_1_wdata <= 0;
      ram_w8_l2048_id7_2_1_wenable <= 0;
      _ram_w8_l2048_id7_2_cond_0_1 <= 0;
      ram_w8_l2048_id7_2_0_addr <= 0;
      _ram_w8_l2048_id7_2_cond_1_1 <= 0;
      _tmp_548 <= 0;
      _ram_w8_l2048_id7_2_cond_2_1 <= 0;
      _ram_w8_l2048_id7_2_cond_2_2 <= 0;
      ram_w8_l2048_id7_2_0_wdata <= 0;
      ram_w8_l2048_id7_2_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id7_2_cond_2_2) begin
        _tmp_548 <= 0;
      end 
      if(_ram_w8_l2048_id7_2_cond_0_1) begin
        ram_w8_l2048_id7_2_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id7_2_cond_1_1) begin
        _tmp_548 <= 1;
      end 
      _ram_w8_l2048_id7_2_cond_2_2 <= _ram_w8_l2048_id7_2_cond_2_1;
      if(_dataflow_slice_ovalid_73 && ((_tmp_375 > 0) && !_tmp_376) && (_tmp_375 > 0)) begin
        ram_w8_l2048_id7_2_1_addr <= _tmp_385;
        ram_w8_l2048_id7_2_1_wdata <= _dataflow_slice_odata_73;
        ram_w8_l2048_id7_2_1_wenable <= _tmp_386 == 2;
      end 
      _ram_w8_l2048_id7_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8)) begin
        ram_w8_l2048_id7_2_0_addr <= _stream_conv2d_16_source_24_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id7_2_cond_1_1 <= _stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8);
      _ram_w8_l2048_id7_2_cond_2_1 <= _stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8);
      ram_w8_l2048_id7_2_0_wdata <= 0;
      ram_w8_l2048_id7_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id7_3_1_addr <= 0;
      ram_w8_l2048_id7_3_1_wdata <= 0;
      ram_w8_l2048_id7_3_1_wenable <= 0;
      _ram_w8_l2048_id7_3_cond_0_1 <= 0;
      ram_w8_l2048_id7_3_0_addr <= 0;
      _ram_w8_l2048_id7_3_cond_1_1 <= 0;
      _tmp_549 <= 0;
      _ram_w8_l2048_id7_3_cond_2_1 <= 0;
      _ram_w8_l2048_id7_3_cond_2_2 <= 0;
      ram_w8_l2048_id7_3_0_wdata <= 0;
      ram_w8_l2048_id7_3_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id7_3_cond_2_2) begin
        _tmp_549 <= 0;
      end 
      if(_ram_w8_l2048_id7_3_cond_0_1) begin
        ram_w8_l2048_id7_3_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id7_3_cond_1_1) begin
        _tmp_549 <= 1;
      end 
      _ram_w8_l2048_id7_3_cond_2_2 <= _ram_w8_l2048_id7_3_cond_2_1;
      if(_dataflow_slice_ovalid_76 && ((_tmp_388 > 0) && !_tmp_389) && (_tmp_388 > 0)) begin
        ram_w8_l2048_id7_3_1_addr <= _tmp_398;
        ram_w8_l2048_id7_3_1_wdata <= _dataflow_slice_odata_76;
        ram_w8_l2048_id7_3_1_wenable <= _tmp_399 == 2;
      end 
      _ram_w8_l2048_id7_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8)) begin
        ram_w8_l2048_id7_3_0_addr <= _stream_conv2d_16_source_24_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id7_3_cond_1_1 <= _stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8);
      _ram_w8_l2048_id7_3_cond_2_1 <= _stream_conv2d_16_source_24_source_ram_renable && (_stream_conv2d_16_source_24_source_ram_sel == 8);
      ram_w8_l2048_id7_3_0_wdata <= 0;
      ram_w8_l2048_id7_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_417 <= 0;
      _tmp_405 <= 0;
      _tmp_406 <= 0;
      _tmp_408 <= 0;
      _tmp_409 <= 0;
      _tmp_410 <= 0;
      ram_w8_l2048_id8_0_1_addr <= 0;
      ram_w8_l2048_id8_0_1_wdata <= 0;
      ram_w8_l2048_id8_0_1_wenable <= 0;
      _tmp_407 <= 0;
      _ram_w8_l2048_id8_0_cond_0_1 <= 0;
      _ram_w8_l2048_id8_0_cond_1_1 <= 0;
      ram_w8_l2048_id8_0_0_addr <= 0;
      _ram_w8_l2048_id8_0_cond_2_1 <= 0;
      _tmp_556 <= 0;
      _ram_w8_l2048_id8_0_cond_3_1 <= 0;
      _ram_w8_l2048_id8_0_cond_3_2 <= 0;
      ram_w8_l2048_id8_0_0_wdata <= 0;
      ram_w8_l2048_id8_0_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id8_0_cond_3_2) begin
        _tmp_556 <= 0;
      end 
      if(_ram_w8_l2048_id8_0_cond_0_1) begin
        _tmp_407 <= 0;
      end 
      if(_ram_w8_l2048_id8_0_cond_1_1) begin
        ram_w8_l2048_id8_0_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id8_0_cond_2_1) begin
        _tmp_556 <= 1;
      end 
      _ram_w8_l2048_id8_0_cond_3_2 <= _ram_w8_l2048_id8_0_cond_3_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_406 == 0)) begin
        _tmp_417 <= 0;
        _tmp_405 <= req_block_size_400 - 1;
        _tmp_406 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_406 == 0)) begin
        _tmp_408 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_406 == 0)) begin
        _tmp_409 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_406 == 0)) begin
        _tmp_410 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_80 && ((_tmp_406 > 0) && !_tmp_407) && (_tmp_406 > 0)) begin
        _tmp_405 <= _tmp_405 - 1;
        _tmp_406 <= _tmp_406 - 1;
      end 
      if(_dataflow_slice_ovalid_80 && ((_tmp_406 > 0) && !_tmp_407) && (_tmp_406 > 0) && (_tmp_405 == 0)) begin
        _tmp_405 <= req_block_size_400 - 1;
        _tmp_417 <= _tmp_417 + 1;
      end 
      if(_dataflow_slice_ovalid_80 && ((_tmp_406 > 0) && !_tmp_407) && (_tmp_406 > 0) && (_tmp_405 == 0) && (_tmp_417 == 2)) begin
        _tmp_417 <= 0;
      end 
      if(_dataflow_slice_ovalid_80 && ((_tmp_406 > 0) && !_tmp_407) && (_tmp_406 > 0) && (_tmp_417 == 0)) begin
        _tmp_408 <= _tmp_411;
      end 
      if(_dataflow_slice_ovalid_80 && ((_tmp_406 > 0) && !_tmp_407) && (_tmp_406 > 0) && (_tmp_417 == 1)) begin
        _tmp_409 <= _tmp_412;
      end 
      if(_dataflow_slice_ovalid_80 && ((_tmp_406 > 0) && !_tmp_407) && (_tmp_406 > 0) && (_tmp_417 == 2)) begin
        _tmp_410 <= _tmp_413;
      end 
      if(_dataflow_slice_ovalid_80 && ((_tmp_406 > 0) && !_tmp_407) && (_tmp_406 > 0)) begin
        ram_w8_l2048_id8_0_1_addr <= _tmp_414;
        ram_w8_l2048_id8_0_1_wdata <= _dataflow_slice_odata_80;
        ram_w8_l2048_id8_0_1_wenable <= _tmp_417 == 0;
      end 
      if(_dataflow_slice_ovalid_80 && ((_tmp_406 > 0) && !_tmp_407) && (_tmp_406 == 1)) begin
        _tmp_407 <= 1;
      end 
      _ram_w8_l2048_id8_0_cond_0_1 <= 1;
      _ram_w8_l2048_id8_0_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9)) begin
        ram_w8_l2048_id8_0_0_addr <= _stream_conv2d_16_source_25_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id8_0_cond_2_1 <= _stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9);
      _ram_w8_l2048_id8_0_cond_3_1 <= _stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9);
      ram_w8_l2048_id8_0_0_wdata <= 0;
      ram_w8_l2048_id8_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_430 <= 0;
      _tmp_418 <= 0;
      _tmp_419 <= 0;
      _tmp_421 <= 0;
      _tmp_422 <= 0;
      _tmp_423 <= 0;
      ram_w8_l2048_id8_1_1_addr <= 0;
      ram_w8_l2048_id8_1_1_wdata <= 0;
      ram_w8_l2048_id8_1_1_wenable <= 0;
      _tmp_420 <= 0;
      _ram_w8_l2048_id8_1_cond_0_1 <= 0;
      _ram_w8_l2048_id8_1_cond_1_1 <= 0;
      ram_w8_l2048_id8_1_0_addr <= 0;
      _ram_w8_l2048_id8_1_cond_2_1 <= 0;
      _tmp_557 <= 0;
      _ram_w8_l2048_id8_1_cond_3_1 <= 0;
      _ram_w8_l2048_id8_1_cond_3_2 <= 0;
      ram_w8_l2048_id8_1_0_wdata <= 0;
      ram_w8_l2048_id8_1_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id8_1_cond_3_2) begin
        _tmp_557 <= 0;
      end 
      if(_ram_w8_l2048_id8_1_cond_0_1) begin
        _tmp_420 <= 0;
      end 
      if(_ram_w8_l2048_id8_1_cond_1_1) begin
        ram_w8_l2048_id8_1_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id8_1_cond_2_1) begin
        _tmp_557 <= 1;
      end 
      _ram_w8_l2048_id8_1_cond_3_2 <= _ram_w8_l2048_id8_1_cond_3_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_419 == 0)) begin
        _tmp_430 <= 0;
        _tmp_418 <= req_block_size_400 - 1;
        _tmp_419 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_419 == 0)) begin
        _tmp_421 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_419 == 0)) begin
        _tmp_422 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_419 == 0)) begin
        _tmp_423 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_83 && ((_tmp_419 > 0) && !_tmp_420) && (_tmp_419 > 0)) begin
        _tmp_418 <= _tmp_418 - 1;
        _tmp_419 <= _tmp_419 - 1;
      end 
      if(_dataflow_slice_ovalid_83 && ((_tmp_419 > 0) && !_tmp_420) && (_tmp_419 > 0) && (_tmp_418 == 0)) begin
        _tmp_418 <= req_block_size_400 - 1;
        _tmp_430 <= _tmp_430 + 1;
      end 
      if(_dataflow_slice_ovalid_83 && ((_tmp_419 > 0) && !_tmp_420) && (_tmp_419 > 0) && (_tmp_418 == 0) && (_tmp_430 == 2)) begin
        _tmp_430 <= 0;
      end 
      if(_dataflow_slice_ovalid_83 && ((_tmp_419 > 0) && !_tmp_420) && (_tmp_419 > 0) && (_tmp_430 == 0)) begin
        _tmp_421 <= _tmp_424;
      end 
      if(_dataflow_slice_ovalid_83 && ((_tmp_419 > 0) && !_tmp_420) && (_tmp_419 > 0) && (_tmp_430 == 1)) begin
        _tmp_422 <= _tmp_425;
      end 
      if(_dataflow_slice_ovalid_83 && ((_tmp_419 > 0) && !_tmp_420) && (_tmp_419 > 0) && (_tmp_430 == 2)) begin
        _tmp_423 <= _tmp_426;
      end 
      if(_dataflow_slice_ovalid_83 && ((_tmp_419 > 0) && !_tmp_420) && (_tmp_419 > 0)) begin
        ram_w8_l2048_id8_1_1_addr <= _tmp_427;
        ram_w8_l2048_id8_1_1_wdata <= _dataflow_slice_odata_83;
        ram_w8_l2048_id8_1_1_wenable <= _tmp_430 == 0;
      end 
      if(_dataflow_slice_ovalid_83 && ((_tmp_419 > 0) && !_tmp_420) && (_tmp_419 == 1)) begin
        _tmp_420 <= 1;
      end 
      _ram_w8_l2048_id8_1_cond_0_1 <= 1;
      _ram_w8_l2048_id8_1_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9)) begin
        ram_w8_l2048_id8_1_0_addr <= _stream_conv2d_16_source_25_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id8_1_cond_2_1 <= _stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9);
      _ram_w8_l2048_id8_1_cond_3_1 <= _stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9);
      ram_w8_l2048_id8_1_0_wdata <= 0;
      ram_w8_l2048_id8_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_443 <= 0;
      _tmp_431 <= 0;
      _tmp_432 <= 0;
      _tmp_434 <= 0;
      _tmp_435 <= 0;
      _tmp_436 <= 0;
      ram_w8_l2048_id8_2_1_addr <= 0;
      ram_w8_l2048_id8_2_1_wdata <= 0;
      ram_w8_l2048_id8_2_1_wenable <= 0;
      _tmp_433 <= 0;
      _ram_w8_l2048_id8_2_cond_0_1 <= 0;
      _ram_w8_l2048_id8_2_cond_1_1 <= 0;
      ram_w8_l2048_id8_2_0_addr <= 0;
      _ram_w8_l2048_id8_2_cond_2_1 <= 0;
      _tmp_558 <= 0;
      _ram_w8_l2048_id8_2_cond_3_1 <= 0;
      _ram_w8_l2048_id8_2_cond_3_2 <= 0;
      ram_w8_l2048_id8_2_0_wdata <= 0;
      ram_w8_l2048_id8_2_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id8_2_cond_3_2) begin
        _tmp_558 <= 0;
      end 
      if(_ram_w8_l2048_id8_2_cond_0_1) begin
        _tmp_433 <= 0;
      end 
      if(_ram_w8_l2048_id8_2_cond_1_1) begin
        ram_w8_l2048_id8_2_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id8_2_cond_2_1) begin
        _tmp_558 <= 1;
      end 
      _ram_w8_l2048_id8_2_cond_3_2 <= _ram_w8_l2048_id8_2_cond_3_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_432 == 0)) begin
        _tmp_443 <= 0;
        _tmp_431 <= req_block_size_400 - 1;
        _tmp_432 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_432 == 0)) begin
        _tmp_434 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_432 == 0)) begin
        _tmp_435 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_432 == 0)) begin
        _tmp_436 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_86 && ((_tmp_432 > 0) && !_tmp_433) && (_tmp_432 > 0)) begin
        _tmp_431 <= _tmp_431 - 1;
        _tmp_432 <= _tmp_432 - 1;
      end 
      if(_dataflow_slice_ovalid_86 && ((_tmp_432 > 0) && !_tmp_433) && (_tmp_432 > 0) && (_tmp_431 == 0)) begin
        _tmp_431 <= req_block_size_400 - 1;
        _tmp_443 <= _tmp_443 + 1;
      end 
      if(_dataflow_slice_ovalid_86 && ((_tmp_432 > 0) && !_tmp_433) && (_tmp_432 > 0) && (_tmp_431 == 0) && (_tmp_443 == 2)) begin
        _tmp_443 <= 0;
      end 
      if(_dataflow_slice_ovalid_86 && ((_tmp_432 > 0) && !_tmp_433) && (_tmp_432 > 0) && (_tmp_443 == 0)) begin
        _tmp_434 <= _tmp_437;
      end 
      if(_dataflow_slice_ovalid_86 && ((_tmp_432 > 0) && !_tmp_433) && (_tmp_432 > 0) && (_tmp_443 == 1)) begin
        _tmp_435 <= _tmp_438;
      end 
      if(_dataflow_slice_ovalid_86 && ((_tmp_432 > 0) && !_tmp_433) && (_tmp_432 > 0) && (_tmp_443 == 2)) begin
        _tmp_436 <= _tmp_439;
      end 
      if(_dataflow_slice_ovalid_86 && ((_tmp_432 > 0) && !_tmp_433) && (_tmp_432 > 0)) begin
        ram_w8_l2048_id8_2_1_addr <= _tmp_440;
        ram_w8_l2048_id8_2_1_wdata <= _dataflow_slice_odata_86;
        ram_w8_l2048_id8_2_1_wenable <= _tmp_443 == 0;
      end 
      if(_dataflow_slice_ovalid_86 && ((_tmp_432 > 0) && !_tmp_433) && (_tmp_432 == 1)) begin
        _tmp_433 <= 1;
      end 
      _ram_w8_l2048_id8_2_cond_0_1 <= 1;
      _ram_w8_l2048_id8_2_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9)) begin
        ram_w8_l2048_id8_2_0_addr <= _stream_conv2d_16_source_25_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id8_2_cond_2_1 <= _stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9);
      _ram_w8_l2048_id8_2_cond_3_1 <= _stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9);
      ram_w8_l2048_id8_2_0_wdata <= 0;
      ram_w8_l2048_id8_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_456 <= 0;
      _tmp_444 <= 0;
      _tmp_445 <= 0;
      _tmp_447 <= 0;
      _tmp_448 <= 0;
      _tmp_449 <= 0;
      ram_w8_l2048_id8_3_1_addr <= 0;
      ram_w8_l2048_id8_3_1_wdata <= 0;
      ram_w8_l2048_id8_3_1_wenable <= 0;
      _tmp_446 <= 0;
      _ram_w8_l2048_id8_3_cond_0_1 <= 0;
      _ram_w8_l2048_id8_3_cond_1_1 <= 0;
      ram_w8_l2048_id8_3_0_addr <= 0;
      _ram_w8_l2048_id8_3_cond_2_1 <= 0;
      _tmp_559 <= 0;
      _ram_w8_l2048_id8_3_cond_3_1 <= 0;
      _ram_w8_l2048_id8_3_cond_3_2 <= 0;
      ram_w8_l2048_id8_3_0_wdata <= 0;
      ram_w8_l2048_id8_3_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id8_3_cond_3_2) begin
        _tmp_559 <= 0;
      end 
      if(_ram_w8_l2048_id8_3_cond_0_1) begin
        _tmp_446 <= 0;
      end 
      if(_ram_w8_l2048_id8_3_cond_1_1) begin
        ram_w8_l2048_id8_3_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id8_3_cond_2_1) begin
        _tmp_559 <= 1;
      end 
      _ram_w8_l2048_id8_3_cond_3_2 <= _ram_w8_l2048_id8_3_cond_3_1;
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_445 == 0)) begin
        _tmp_456 <= 0;
        _tmp_444 <= req_block_size_400 - 1;
        _tmp_445 <= _maxi_read_size;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_445 == 0)) begin
        _tmp_447 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_445 == 0)) begin
        _tmp_448 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_maxi_read_start && (_maxi_read_op_sel == 6) && (_tmp_445 == 0)) begin
        _tmp_449 <= _maxi_read_local_addr - _maxi_read_local_stride;
      end 
      if(_dataflow_slice_ovalid_89 && ((_tmp_445 > 0) && !_tmp_446) && (_tmp_445 > 0)) begin
        _tmp_444 <= _tmp_444 - 1;
        _tmp_445 <= _tmp_445 - 1;
      end 
      if(_dataflow_slice_ovalid_89 && ((_tmp_445 > 0) && !_tmp_446) && (_tmp_445 > 0) && (_tmp_444 == 0)) begin
        _tmp_444 <= req_block_size_400 - 1;
        _tmp_456 <= _tmp_456 + 1;
      end 
      if(_dataflow_slice_ovalid_89 && ((_tmp_445 > 0) && !_tmp_446) && (_tmp_445 > 0) && (_tmp_444 == 0) && (_tmp_456 == 2)) begin
        _tmp_456 <= 0;
      end 
      if(_dataflow_slice_ovalid_89 && ((_tmp_445 > 0) && !_tmp_446) && (_tmp_445 > 0) && (_tmp_456 == 0)) begin
        _tmp_447 <= _tmp_450;
      end 
      if(_dataflow_slice_ovalid_89 && ((_tmp_445 > 0) && !_tmp_446) && (_tmp_445 > 0) && (_tmp_456 == 1)) begin
        _tmp_448 <= _tmp_451;
      end 
      if(_dataflow_slice_ovalid_89 && ((_tmp_445 > 0) && !_tmp_446) && (_tmp_445 > 0) && (_tmp_456 == 2)) begin
        _tmp_449 <= _tmp_452;
      end 
      if(_dataflow_slice_ovalid_89 && ((_tmp_445 > 0) && !_tmp_446) && (_tmp_445 > 0)) begin
        ram_w8_l2048_id8_3_1_addr <= _tmp_453;
        ram_w8_l2048_id8_3_1_wdata <= _dataflow_slice_odata_89;
        ram_w8_l2048_id8_3_1_wenable <= _tmp_456 == 0;
      end 
      if(_dataflow_slice_ovalid_89 && ((_tmp_445 > 0) && !_tmp_446) && (_tmp_445 == 1)) begin
        _tmp_446 <= 1;
      end 
      _ram_w8_l2048_id8_3_cond_0_1 <= 1;
      _ram_w8_l2048_id8_3_cond_1_1 <= 1;
      if(_stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9)) begin
        ram_w8_l2048_id8_3_0_addr <= _stream_conv2d_16_source_25_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id8_3_cond_2_1 <= _stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9);
      _ram_w8_l2048_id8_3_cond_3_1 <= _stream_conv2d_16_source_25_source_ram_renable && (_stream_conv2d_16_source_25_source_ram_sel == 9);
      ram_w8_l2048_id8_3_0_wdata <= 0;
      ram_w8_l2048_id8_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id9_0_1_addr <= 0;
      ram_w8_l2048_id9_0_1_wdata <= 0;
      ram_w8_l2048_id9_0_1_wenable <= 0;
      _ram_w8_l2048_id9_0_cond_0_1 <= 0;
      ram_w8_l2048_id9_0_0_addr <= 0;
      _ram_w8_l2048_id9_0_cond_1_1 <= 0;
      _tmp_566 <= 0;
      _ram_w8_l2048_id9_0_cond_2_1 <= 0;
      _ram_w8_l2048_id9_0_cond_2_2 <= 0;
      ram_w8_l2048_id9_0_0_wdata <= 0;
      ram_w8_l2048_id9_0_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id9_0_cond_2_2) begin
        _tmp_566 <= 0;
      end 
      if(_ram_w8_l2048_id9_0_cond_0_1) begin
        ram_w8_l2048_id9_0_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id9_0_cond_1_1) begin
        _tmp_566 <= 1;
      end 
      _ram_w8_l2048_id9_0_cond_2_2 <= _ram_w8_l2048_id9_0_cond_2_1;
      if(_dataflow_slice_ovalid_80 && ((_tmp_406 > 0) && !_tmp_407) && (_tmp_406 > 0)) begin
        ram_w8_l2048_id9_0_1_addr <= _tmp_415;
        ram_w8_l2048_id9_0_1_wdata <= _dataflow_slice_odata_80;
        ram_w8_l2048_id9_0_1_wenable <= _tmp_417 == 1;
      end 
      _ram_w8_l2048_id9_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10)) begin
        ram_w8_l2048_id9_0_0_addr <= _stream_conv2d_16_source_26_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id9_0_cond_1_1 <= _stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10);
      _ram_w8_l2048_id9_0_cond_2_1 <= _stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10);
      ram_w8_l2048_id9_0_0_wdata <= 0;
      ram_w8_l2048_id9_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id9_1_1_addr <= 0;
      ram_w8_l2048_id9_1_1_wdata <= 0;
      ram_w8_l2048_id9_1_1_wenable <= 0;
      _ram_w8_l2048_id9_1_cond_0_1 <= 0;
      ram_w8_l2048_id9_1_0_addr <= 0;
      _ram_w8_l2048_id9_1_cond_1_1 <= 0;
      _tmp_567 <= 0;
      _ram_w8_l2048_id9_1_cond_2_1 <= 0;
      _ram_w8_l2048_id9_1_cond_2_2 <= 0;
      ram_w8_l2048_id9_1_0_wdata <= 0;
      ram_w8_l2048_id9_1_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id9_1_cond_2_2) begin
        _tmp_567 <= 0;
      end 
      if(_ram_w8_l2048_id9_1_cond_0_1) begin
        ram_w8_l2048_id9_1_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id9_1_cond_1_1) begin
        _tmp_567 <= 1;
      end 
      _ram_w8_l2048_id9_1_cond_2_2 <= _ram_w8_l2048_id9_1_cond_2_1;
      if(_dataflow_slice_ovalid_83 && ((_tmp_419 > 0) && !_tmp_420) && (_tmp_419 > 0)) begin
        ram_w8_l2048_id9_1_1_addr <= _tmp_428;
        ram_w8_l2048_id9_1_1_wdata <= _dataflow_slice_odata_83;
        ram_w8_l2048_id9_1_1_wenable <= _tmp_430 == 1;
      end 
      _ram_w8_l2048_id9_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10)) begin
        ram_w8_l2048_id9_1_0_addr <= _stream_conv2d_16_source_26_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id9_1_cond_1_1 <= _stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10);
      _ram_w8_l2048_id9_1_cond_2_1 <= _stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10);
      ram_w8_l2048_id9_1_0_wdata <= 0;
      ram_w8_l2048_id9_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id9_2_1_addr <= 0;
      ram_w8_l2048_id9_2_1_wdata <= 0;
      ram_w8_l2048_id9_2_1_wenable <= 0;
      _ram_w8_l2048_id9_2_cond_0_1 <= 0;
      ram_w8_l2048_id9_2_0_addr <= 0;
      _ram_w8_l2048_id9_2_cond_1_1 <= 0;
      _tmp_568 <= 0;
      _ram_w8_l2048_id9_2_cond_2_1 <= 0;
      _ram_w8_l2048_id9_2_cond_2_2 <= 0;
      ram_w8_l2048_id9_2_0_wdata <= 0;
      ram_w8_l2048_id9_2_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id9_2_cond_2_2) begin
        _tmp_568 <= 0;
      end 
      if(_ram_w8_l2048_id9_2_cond_0_1) begin
        ram_w8_l2048_id9_2_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id9_2_cond_1_1) begin
        _tmp_568 <= 1;
      end 
      _ram_w8_l2048_id9_2_cond_2_2 <= _ram_w8_l2048_id9_2_cond_2_1;
      if(_dataflow_slice_ovalid_86 && ((_tmp_432 > 0) && !_tmp_433) && (_tmp_432 > 0)) begin
        ram_w8_l2048_id9_2_1_addr <= _tmp_441;
        ram_w8_l2048_id9_2_1_wdata <= _dataflow_slice_odata_86;
        ram_w8_l2048_id9_2_1_wenable <= _tmp_443 == 1;
      end 
      _ram_w8_l2048_id9_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10)) begin
        ram_w8_l2048_id9_2_0_addr <= _stream_conv2d_16_source_26_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id9_2_cond_1_1 <= _stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10);
      _ram_w8_l2048_id9_2_cond_2_1 <= _stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10);
      ram_w8_l2048_id9_2_0_wdata <= 0;
      ram_w8_l2048_id9_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id9_3_1_addr <= 0;
      ram_w8_l2048_id9_3_1_wdata <= 0;
      ram_w8_l2048_id9_3_1_wenable <= 0;
      _ram_w8_l2048_id9_3_cond_0_1 <= 0;
      ram_w8_l2048_id9_3_0_addr <= 0;
      _ram_w8_l2048_id9_3_cond_1_1 <= 0;
      _tmp_569 <= 0;
      _ram_w8_l2048_id9_3_cond_2_1 <= 0;
      _ram_w8_l2048_id9_3_cond_2_2 <= 0;
      ram_w8_l2048_id9_3_0_wdata <= 0;
      ram_w8_l2048_id9_3_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id9_3_cond_2_2) begin
        _tmp_569 <= 0;
      end 
      if(_ram_w8_l2048_id9_3_cond_0_1) begin
        ram_w8_l2048_id9_3_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id9_3_cond_1_1) begin
        _tmp_569 <= 1;
      end 
      _ram_w8_l2048_id9_3_cond_2_2 <= _ram_w8_l2048_id9_3_cond_2_1;
      if(_dataflow_slice_ovalid_89 && ((_tmp_445 > 0) && !_tmp_446) && (_tmp_445 > 0)) begin
        ram_w8_l2048_id9_3_1_addr <= _tmp_454;
        ram_w8_l2048_id9_3_1_wdata <= _dataflow_slice_odata_89;
        ram_w8_l2048_id9_3_1_wenable <= _tmp_456 == 1;
      end 
      _ram_w8_l2048_id9_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10)) begin
        ram_w8_l2048_id9_3_0_addr <= _stream_conv2d_16_source_26_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id9_3_cond_1_1 <= _stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10);
      _ram_w8_l2048_id9_3_cond_2_1 <= _stream_conv2d_16_source_26_source_ram_renable && (_stream_conv2d_16_source_26_source_ram_sel == 10);
      ram_w8_l2048_id9_3_0_wdata <= 0;
      ram_w8_l2048_id9_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id10_0_1_addr <= 0;
      ram_w8_l2048_id10_0_1_wdata <= 0;
      ram_w8_l2048_id10_0_1_wenable <= 0;
      _ram_w8_l2048_id10_0_cond_0_1 <= 0;
      ram_w8_l2048_id10_0_0_addr <= 0;
      _ram_w8_l2048_id10_0_cond_1_1 <= 0;
      _tmp_576 <= 0;
      _ram_w8_l2048_id10_0_cond_2_1 <= 0;
      _ram_w8_l2048_id10_0_cond_2_2 <= 0;
      ram_w8_l2048_id10_0_0_wdata <= 0;
      ram_w8_l2048_id10_0_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id10_0_cond_2_2) begin
        _tmp_576 <= 0;
      end 
      if(_ram_w8_l2048_id10_0_cond_0_1) begin
        ram_w8_l2048_id10_0_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id10_0_cond_1_1) begin
        _tmp_576 <= 1;
      end 
      _ram_w8_l2048_id10_0_cond_2_2 <= _ram_w8_l2048_id10_0_cond_2_1;
      if(_dataflow_slice_ovalid_80 && ((_tmp_406 > 0) && !_tmp_407) && (_tmp_406 > 0)) begin
        ram_w8_l2048_id10_0_1_addr <= _tmp_416;
        ram_w8_l2048_id10_0_1_wdata <= _dataflow_slice_odata_80;
        ram_w8_l2048_id10_0_1_wenable <= _tmp_417 == 2;
      end 
      _ram_w8_l2048_id10_0_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11)) begin
        ram_w8_l2048_id10_0_0_addr <= _stream_conv2d_16_source_27_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id10_0_cond_1_1 <= _stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11);
      _ram_w8_l2048_id10_0_cond_2_1 <= _stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11);
      ram_w8_l2048_id10_0_0_wdata <= 0;
      ram_w8_l2048_id10_0_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id10_1_1_addr <= 0;
      ram_w8_l2048_id10_1_1_wdata <= 0;
      ram_w8_l2048_id10_1_1_wenable <= 0;
      _ram_w8_l2048_id10_1_cond_0_1 <= 0;
      ram_w8_l2048_id10_1_0_addr <= 0;
      _ram_w8_l2048_id10_1_cond_1_1 <= 0;
      _tmp_577 <= 0;
      _ram_w8_l2048_id10_1_cond_2_1 <= 0;
      _ram_w8_l2048_id10_1_cond_2_2 <= 0;
      ram_w8_l2048_id10_1_0_wdata <= 0;
      ram_w8_l2048_id10_1_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id10_1_cond_2_2) begin
        _tmp_577 <= 0;
      end 
      if(_ram_w8_l2048_id10_1_cond_0_1) begin
        ram_w8_l2048_id10_1_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id10_1_cond_1_1) begin
        _tmp_577 <= 1;
      end 
      _ram_w8_l2048_id10_1_cond_2_2 <= _ram_w8_l2048_id10_1_cond_2_1;
      if(_dataflow_slice_ovalid_83 && ((_tmp_419 > 0) && !_tmp_420) && (_tmp_419 > 0)) begin
        ram_w8_l2048_id10_1_1_addr <= _tmp_429;
        ram_w8_l2048_id10_1_1_wdata <= _dataflow_slice_odata_83;
        ram_w8_l2048_id10_1_1_wenable <= _tmp_430 == 2;
      end 
      _ram_w8_l2048_id10_1_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11)) begin
        ram_w8_l2048_id10_1_0_addr <= _stream_conv2d_16_source_27_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id10_1_cond_1_1 <= _stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11);
      _ram_w8_l2048_id10_1_cond_2_1 <= _stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11);
      ram_w8_l2048_id10_1_0_wdata <= 0;
      ram_w8_l2048_id10_1_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id10_2_1_addr <= 0;
      ram_w8_l2048_id10_2_1_wdata <= 0;
      ram_w8_l2048_id10_2_1_wenable <= 0;
      _ram_w8_l2048_id10_2_cond_0_1 <= 0;
      ram_w8_l2048_id10_2_0_addr <= 0;
      _ram_w8_l2048_id10_2_cond_1_1 <= 0;
      _tmp_578 <= 0;
      _ram_w8_l2048_id10_2_cond_2_1 <= 0;
      _ram_w8_l2048_id10_2_cond_2_2 <= 0;
      ram_w8_l2048_id10_2_0_wdata <= 0;
      ram_w8_l2048_id10_2_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id10_2_cond_2_2) begin
        _tmp_578 <= 0;
      end 
      if(_ram_w8_l2048_id10_2_cond_0_1) begin
        ram_w8_l2048_id10_2_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id10_2_cond_1_1) begin
        _tmp_578 <= 1;
      end 
      _ram_w8_l2048_id10_2_cond_2_2 <= _ram_w8_l2048_id10_2_cond_2_1;
      if(_dataflow_slice_ovalid_86 && ((_tmp_432 > 0) && !_tmp_433) && (_tmp_432 > 0)) begin
        ram_w8_l2048_id10_2_1_addr <= _tmp_442;
        ram_w8_l2048_id10_2_1_wdata <= _dataflow_slice_odata_86;
        ram_w8_l2048_id10_2_1_wenable <= _tmp_443 == 2;
      end 
      _ram_w8_l2048_id10_2_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11)) begin
        ram_w8_l2048_id10_2_0_addr <= _stream_conv2d_16_source_27_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id10_2_cond_1_1 <= _stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11);
      _ram_w8_l2048_id10_2_cond_2_1 <= _stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11);
      ram_w8_l2048_id10_2_0_wdata <= 0;
      ram_w8_l2048_id10_2_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id10_3_1_addr <= 0;
      ram_w8_l2048_id10_3_1_wdata <= 0;
      ram_w8_l2048_id10_3_1_wenable <= 0;
      _ram_w8_l2048_id10_3_cond_0_1 <= 0;
      ram_w8_l2048_id10_3_0_addr <= 0;
      _ram_w8_l2048_id10_3_cond_1_1 <= 0;
      _tmp_579 <= 0;
      _ram_w8_l2048_id10_3_cond_2_1 <= 0;
      _ram_w8_l2048_id10_3_cond_2_2 <= 0;
      ram_w8_l2048_id10_3_0_wdata <= 0;
      ram_w8_l2048_id10_3_0_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id10_3_cond_2_2) begin
        _tmp_579 <= 0;
      end 
      if(_ram_w8_l2048_id10_3_cond_0_1) begin
        ram_w8_l2048_id10_3_1_wenable <= 0;
      end 
      if(_ram_w8_l2048_id10_3_cond_1_1) begin
        _tmp_579 <= 1;
      end 
      _ram_w8_l2048_id10_3_cond_2_2 <= _ram_w8_l2048_id10_3_cond_2_1;
      if(_dataflow_slice_ovalid_89 && ((_tmp_445 > 0) && !_tmp_446) && (_tmp_445 > 0)) begin
        ram_w8_l2048_id10_3_1_addr <= _tmp_455;
        ram_w8_l2048_id10_3_1_wdata <= _dataflow_slice_odata_89;
        ram_w8_l2048_id10_3_1_wenable <= _tmp_456 == 2;
      end 
      _ram_w8_l2048_id10_3_cond_0_1 <= 1;
      if(_stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11)) begin
        ram_w8_l2048_id10_3_0_addr <= _stream_conv2d_16_source_27_source_ram_raddr >> 2;
      end 
      _ram_w8_l2048_id10_3_cond_1_1 <= _stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11);
      _ram_w8_l2048_id10_3_cond_2_1 <= _stream_conv2d_16_source_27_source_ram_renable && (_stream_conv2d_16_source_27_source_ram_sel == 11);
      ram_w8_l2048_id10_3_0_wdata <= 0;
      ram_w8_l2048_id10_3_0_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id11_0_0_addr <= 0;
      ram_w8_l2048_id11_0_0_wdata <= 0;
      ram_w8_l2048_id11_0_0_wenable <= 0;
      _ram_w8_l2048_id11_0_cond_0_1 <= 0;
      __tmp_976_1 <= 0;
      __tmp_977_1 <= 0;
      _tmp_981 <= 0;
      _tmp_971 <= 0;
      _tmp_972 <= 0;
      _tmp_979 <= 0;
      _tmp_980 <= 0;
      _tmp_978 <= 0;
      ram_w8_l2048_id11_0_1_addr <= 0;
      _tmp_982 <= 0;
      ram_w8_l2048_id11_0_1_wdata <= 0;
      ram_w8_l2048_id11_0_1_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id11_0_cond_0_1) begin
        ram_w8_l2048_id11_0_0_wenable <= 0;
      end 
      if(_stream_conv2d_16_sink_37_sink_wenable && (_stream_conv2d_16_sink_37_sink_ram_sel == 21) && (_tmp_711 == 0)) begin
        ram_w8_l2048_id11_0_0_addr <= _stream_conv2d_16_sink_37_sink_waddr >> 2;
        ram_w8_l2048_id11_0_0_wdata <= _stream_conv2d_16_sink_37_sink_wdata;
        ram_w8_l2048_id11_0_0_wenable <= 1;
      end 
      _ram_w8_l2048_id11_0_cond_0_1 <= _stream_conv2d_16_sink_37_sink_wenable && (_stream_conv2d_16_sink_37_sink_ram_sel == 21) && (_tmp_711 == 0);
      __tmp_976_1 <= _tmp_976;
      __tmp_977_1 <= _tmp_977;
      if((_tmp_973 || !_tmp_971) && (_tmp_974 || !_tmp_972) && _tmp_979) begin
        _tmp_981 <= 0;
        _tmp_971 <= 0;
        _tmp_972 <= 0;
        _tmp_979 <= 0;
      end 
      if((_tmp_973 || !_tmp_971) && (_tmp_974 || !_tmp_972) && _tmp_978) begin
        _tmp_971 <= 1;
        _tmp_972 <= 1;
        _tmp_981 <= _tmp_980;
        _tmp_980 <= 0;
        _tmp_978 <= 0;
        _tmp_979 <= 1;
      end 
      if(_maxi_write_start && (_maxi_write_op_sel == 1) && (_tmp_982 == 0) && !_tmp_980 && !_tmp_981) begin
        ram_w8_l2048_id11_0_1_addr <= _maxi_write_local_addr;
        _tmp_982 <= _maxi_write_size - 1;
        _tmp_978 <= 1;
        _tmp_980 <= _maxi_write_size == 1;
      end 
      if((_tmp_973 || !_tmp_971) && (_tmp_974 || !_tmp_972) && (_tmp_982 > 0)) begin
        ram_w8_l2048_id11_0_1_addr <= ram_w8_l2048_id11_0_1_addr + _maxi_write_local_stride;
        _tmp_982 <= _tmp_982 - 1;
        _tmp_978 <= 1;
        _tmp_980 <= 0;
      end 
      if((_tmp_973 || !_tmp_971) && (_tmp_974 || !_tmp_972) && (_tmp_982 == 1)) begin
        _tmp_980 <= 1;
      end 
      ram_w8_l2048_id11_0_1_wdata <= 0;
      ram_w8_l2048_id11_0_1_wenable <= 0;
    end
  end

  reg [32-1:0] _dataflow_cat_data_98;
  reg _dataflow_cat_valid_98;
  wire _dataflow_cat_ready_98;
  assign _tmp_1009 = 1 && ((_dataflow_cat_ready_98 || !_dataflow_cat_valid_98) && (_tmp_1007 && _tmp_995 && _tmp_983 && _tmp_971));
  assign _tmp_997 = 1 && ((_dataflow_cat_ready_98 || !_dataflow_cat_valid_98) && (_tmp_1007 && _tmp_995 && _tmp_983 && _tmp_971));
  assign _tmp_985 = 1 && ((_dataflow_cat_ready_98 || !_dataflow_cat_valid_98) && (_tmp_1007 && _tmp_995 && _tmp_983 && _tmp_971));
  assign _tmp_973 = 1 && ((_dataflow_cat_ready_98 || !_dataflow_cat_valid_98) && (_tmp_1007 && _tmp_995 && _tmp_983 && _tmp_971));
  assign _dataflow_cat_odata_98 = _dataflow_cat_data_98;
  assign _dataflow_cat_ovalid_98 = _dataflow_cat_valid_98;
  assign _dataflow_cat_ready_98 = _dataflow_cat_oready_98;

  always @(posedge CLK) begin
    if(RST) begin
      _dataflow_cat_data_98 <= 0;
      _dataflow_cat_valid_98 <= 0;
    end else begin
      if((_dataflow_cat_ready_98 || !_dataflow_cat_valid_98) && (_tmp_1009 && _tmp_997 && _tmp_985 && _tmp_973) && (_tmp_1007 && _tmp_995 && _tmp_983 && _tmp_971)) begin
        _dataflow_cat_data_98 <= { _tmp_1013, _tmp_1001, _tmp_989, _tmp_977 };
      end 
      if(_dataflow_cat_valid_98 && _dataflow_cat_ready_98) begin
        _dataflow_cat_valid_98 <= 0;
      end 
      if((_dataflow_cat_ready_98 || !_dataflow_cat_valid_98) && (_tmp_1009 && _tmp_997 && _tmp_985 && _tmp_973)) begin
        _dataflow_cat_valid_98 <= _tmp_1007 && _tmp_995 && _tmp_983 && _tmp_971;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id11_1_0_addr <= 0;
      ram_w8_l2048_id11_1_0_wdata <= 0;
      ram_w8_l2048_id11_1_0_wenable <= 0;
      _ram_w8_l2048_id11_1_cond_0_1 <= 0;
      __tmp_988_1 <= 0;
      __tmp_989_1 <= 0;
      _tmp_993 <= 0;
      _tmp_983 <= 0;
      _tmp_984 <= 0;
      _tmp_991 <= 0;
      _tmp_992 <= 0;
      _tmp_990 <= 0;
      ram_w8_l2048_id11_1_1_addr <= 0;
      _tmp_994 <= 0;
      ram_w8_l2048_id11_1_1_wdata <= 0;
      ram_w8_l2048_id11_1_1_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id11_1_cond_0_1) begin
        ram_w8_l2048_id11_1_0_wenable <= 0;
      end 
      if(_stream_conv2d_16_sink_37_sink_wenable && (_stream_conv2d_16_sink_37_sink_ram_sel == 21) && (_tmp_711 == 1)) begin
        ram_w8_l2048_id11_1_0_addr <= _stream_conv2d_16_sink_37_sink_waddr >> 2;
        ram_w8_l2048_id11_1_0_wdata <= _stream_conv2d_16_sink_37_sink_wdata;
        ram_w8_l2048_id11_1_0_wenable <= 1;
      end 
      _ram_w8_l2048_id11_1_cond_0_1 <= _stream_conv2d_16_sink_37_sink_wenable && (_stream_conv2d_16_sink_37_sink_ram_sel == 21) && (_tmp_711 == 1);
      __tmp_988_1 <= _tmp_988;
      __tmp_989_1 <= _tmp_989;
      if((_tmp_985 || !_tmp_983) && (_tmp_986 || !_tmp_984) && _tmp_991) begin
        _tmp_993 <= 0;
        _tmp_983 <= 0;
        _tmp_984 <= 0;
        _tmp_991 <= 0;
      end 
      if((_tmp_985 || !_tmp_983) && (_tmp_986 || !_tmp_984) && _tmp_990) begin
        _tmp_983 <= 1;
        _tmp_984 <= 1;
        _tmp_993 <= _tmp_992;
        _tmp_992 <= 0;
        _tmp_990 <= 0;
        _tmp_991 <= 1;
      end 
      if(_maxi_write_start && (_maxi_write_op_sel == 1) && (_tmp_994 == 0) && !_tmp_992 && !_tmp_993) begin
        ram_w8_l2048_id11_1_1_addr <= _maxi_write_local_addr;
        _tmp_994 <= _maxi_write_size - 1;
        _tmp_990 <= 1;
        _tmp_992 <= _maxi_write_size == 1;
      end 
      if((_tmp_985 || !_tmp_983) && (_tmp_986 || !_tmp_984) && (_tmp_994 > 0)) begin
        ram_w8_l2048_id11_1_1_addr <= ram_w8_l2048_id11_1_1_addr + _maxi_write_local_stride;
        _tmp_994 <= _tmp_994 - 1;
        _tmp_990 <= 1;
        _tmp_992 <= 0;
      end 
      if((_tmp_985 || !_tmp_983) && (_tmp_986 || !_tmp_984) && (_tmp_994 == 1)) begin
        _tmp_992 <= 1;
      end 
      ram_w8_l2048_id11_1_1_wdata <= 0;
      ram_w8_l2048_id11_1_1_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id11_2_0_addr <= 0;
      ram_w8_l2048_id11_2_0_wdata <= 0;
      ram_w8_l2048_id11_2_0_wenable <= 0;
      _ram_w8_l2048_id11_2_cond_0_1 <= 0;
      __tmp_1000_1 <= 0;
      __tmp_1001_1 <= 0;
      _tmp_1005 <= 0;
      _tmp_995 <= 0;
      _tmp_996 <= 0;
      _tmp_1003 <= 0;
      _tmp_1004 <= 0;
      _tmp_1002 <= 0;
      ram_w8_l2048_id11_2_1_addr <= 0;
      _tmp_1006 <= 0;
      ram_w8_l2048_id11_2_1_wdata <= 0;
      ram_w8_l2048_id11_2_1_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id11_2_cond_0_1) begin
        ram_w8_l2048_id11_2_0_wenable <= 0;
      end 
      if(_stream_conv2d_16_sink_37_sink_wenable && (_stream_conv2d_16_sink_37_sink_ram_sel == 21) && (_tmp_711 == 2)) begin
        ram_w8_l2048_id11_2_0_addr <= _stream_conv2d_16_sink_37_sink_waddr >> 2;
        ram_w8_l2048_id11_2_0_wdata <= _stream_conv2d_16_sink_37_sink_wdata;
        ram_w8_l2048_id11_2_0_wenable <= 1;
      end 
      _ram_w8_l2048_id11_2_cond_0_1 <= _stream_conv2d_16_sink_37_sink_wenable && (_stream_conv2d_16_sink_37_sink_ram_sel == 21) && (_tmp_711 == 2);
      __tmp_1000_1 <= _tmp_1000;
      __tmp_1001_1 <= _tmp_1001;
      if((_tmp_997 || !_tmp_995) && (_tmp_998 || !_tmp_996) && _tmp_1003) begin
        _tmp_1005 <= 0;
        _tmp_995 <= 0;
        _tmp_996 <= 0;
        _tmp_1003 <= 0;
      end 
      if((_tmp_997 || !_tmp_995) && (_tmp_998 || !_tmp_996) && _tmp_1002) begin
        _tmp_995 <= 1;
        _tmp_996 <= 1;
        _tmp_1005 <= _tmp_1004;
        _tmp_1004 <= 0;
        _tmp_1002 <= 0;
        _tmp_1003 <= 1;
      end 
      if(_maxi_write_start && (_maxi_write_op_sel == 1) && (_tmp_1006 == 0) && !_tmp_1004 && !_tmp_1005) begin
        ram_w8_l2048_id11_2_1_addr <= _maxi_write_local_addr;
        _tmp_1006 <= _maxi_write_size - 1;
        _tmp_1002 <= 1;
        _tmp_1004 <= _maxi_write_size == 1;
      end 
      if((_tmp_997 || !_tmp_995) && (_tmp_998 || !_tmp_996) && (_tmp_1006 > 0)) begin
        ram_w8_l2048_id11_2_1_addr <= ram_w8_l2048_id11_2_1_addr + _maxi_write_local_stride;
        _tmp_1006 <= _tmp_1006 - 1;
        _tmp_1002 <= 1;
        _tmp_1004 <= 0;
      end 
      if((_tmp_997 || !_tmp_995) && (_tmp_998 || !_tmp_996) && (_tmp_1006 == 1)) begin
        _tmp_1004 <= 1;
      end 
      ram_w8_l2048_id11_2_1_wdata <= 0;
      ram_w8_l2048_id11_2_1_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      ram_w8_l2048_id11_3_0_addr <= 0;
      ram_w8_l2048_id11_3_0_wdata <= 0;
      ram_w8_l2048_id11_3_0_wenable <= 0;
      _ram_w8_l2048_id11_3_cond_0_1 <= 0;
      __tmp_1012_1 <= 0;
      __tmp_1013_1 <= 0;
      _tmp_1017 <= 0;
      _tmp_1007 <= 0;
      _tmp_1008 <= 0;
      _tmp_1015 <= 0;
      _tmp_1016 <= 0;
      _tmp_1014 <= 0;
      ram_w8_l2048_id11_3_1_addr <= 0;
      _tmp_1018 <= 0;
      ram_w8_l2048_id11_3_1_wdata <= 0;
      ram_w8_l2048_id11_3_1_wenable <= 0;
    end else begin
      if(_ram_w8_l2048_id11_3_cond_0_1) begin
        ram_w8_l2048_id11_3_0_wenable <= 0;
      end 
      if(_stream_conv2d_16_sink_37_sink_wenable && (_stream_conv2d_16_sink_37_sink_ram_sel == 21) && (_tmp_711 == 3)) begin
        ram_w8_l2048_id11_3_0_addr <= _stream_conv2d_16_sink_37_sink_waddr >> 2;
        ram_w8_l2048_id11_3_0_wdata <= _stream_conv2d_16_sink_37_sink_wdata;
        ram_w8_l2048_id11_3_0_wenable <= 1;
      end 
      _ram_w8_l2048_id11_3_cond_0_1 <= _stream_conv2d_16_sink_37_sink_wenable && (_stream_conv2d_16_sink_37_sink_ram_sel == 21) && (_tmp_711 == 3);
      __tmp_1012_1 <= _tmp_1012;
      __tmp_1013_1 <= _tmp_1013;
      if((_tmp_1009 || !_tmp_1007) && (_tmp_1010 || !_tmp_1008) && _tmp_1015) begin
        _tmp_1017 <= 0;
        _tmp_1007 <= 0;
        _tmp_1008 <= 0;
        _tmp_1015 <= 0;
      end 
      if((_tmp_1009 || !_tmp_1007) && (_tmp_1010 || !_tmp_1008) && _tmp_1014) begin
        _tmp_1007 <= 1;
        _tmp_1008 <= 1;
        _tmp_1017 <= _tmp_1016;
        _tmp_1016 <= 0;
        _tmp_1014 <= 0;
        _tmp_1015 <= 1;
      end 
      if(_maxi_write_start && (_maxi_write_op_sel == 1) && (_tmp_1018 == 0) && !_tmp_1016 && !_tmp_1017) begin
        ram_w8_l2048_id11_3_1_addr <= _maxi_write_local_addr;
        _tmp_1018 <= _maxi_write_size - 1;
        _tmp_1014 <= 1;
        _tmp_1016 <= _maxi_write_size == 1;
      end 
      if((_tmp_1009 || !_tmp_1007) && (_tmp_1010 || !_tmp_1008) && (_tmp_1018 > 0)) begin
        ram_w8_l2048_id11_3_1_addr <= ram_w8_l2048_id11_3_1_addr + _maxi_write_local_stride;
        _tmp_1018 <= _tmp_1018 - 1;
        _tmp_1014 <= 1;
        _tmp_1016 <= 0;
      end 
      if((_tmp_1009 || !_tmp_1007) && (_tmp_1010 || !_tmp_1008) && (_tmp_1018 == 1)) begin
        _tmp_1016 <= 1;
      end 
      ram_w8_l2048_id11_3_1_wdata <= 0;
      ram_w8_l2048_id11_3_1_wenable <= 0;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _acc_0_x_idle <= 1;
      _acc_0_x_source_ram_rvalid <= 0;
      _acc_0_rshift_idle <= 1;
      _acc_0_rshift_source_ram_rvalid <= 0;
      _acc_0_sum_sink_wenable <= 0;
      _acc_0_valid_sink_wenable <= 0;
      _greaterthan_data_3 <= 0;
      _minus_data_5 <= 0;
      _reduceadd_data_17 <= 1'sd0;
      _reduceadd_count_17 <= 0;
      _pulse_data_19 <= 1'sd0;
      _pulse_count_19 <= 0;
      __delay_data_751 <= 0;
      _sll_data_7 <= 0;
      __delay_data_748 <= 0;
      __delay_data_749 <= 0;
      __delay_data_752 <= 0;
      __delay_data_755 <= 0;
      _cond_data_13 <= 0;
      __delay_data_750 <= 0;
      __delay_data_753 <= 0;
      __delay_data_756 <= 0;
      _plus_data_20 <= 0;
      __delay_data_754 <= 0;
      __delay_data_757 <= 0;
      _sra_data_21 <= 0;
      __delay_data_758 <= 0;
      __variable_wdata_0 <= 0;
      __variable_wdata_1 <= 0;
      __variable_wdata_2 <= 0;
      __tmp_943_1 <= 0;
      __tmp_943_2 <= 0;
      __tmp_943_3 <= 0;
      __tmp_943_4 <= 0;
      __tmp_943_5 <= 0;
      __tmp_943_6 <= 0;
      __tmp_943_7 <= 0;
      __tmp_943_8 <= 0;
      __tmp_943_9 <= 0;
      __tmp_945_1 <= 0;
      __tmp_945_2 <= 0;
      __tmp_945_3 <= 0;
      __tmp_945_4 <= 0;
      __tmp_945_5 <= 0;
      __tmp_945_6 <= 0;
      __tmp_945_7 <= 0;
      __tmp_945_8 <= 0;
      __tmp_945_9 <= 0;
      __tmp_947_1 <= 0;
      __tmp_947_2 <= 0;
      __tmp_947_3 <= 0;
      __tmp_947_4 <= 0;
      __tmp_947_5 <= 0;
      __tmp_947_6 <= 0;
      __tmp_947_7 <= 0;
      __tmp_947_8 <= 0;
      __tmp_947_9 <= 0;
      __tmp_1281_1 <= 0;
      __tmp_1281_2 <= 0;
      __tmp_1281_3 <= 0;
      __tmp_1281_4 <= 0;
      __tmp_1281_5 <= 0;
      __tmp_1281_6 <= 0;
      __tmp_1281_7 <= 0;
      __tmp_1281_8 <= 0;
      __tmp_1281_9 <= 0;
      __tmp_1283_1 <= 0;
      __tmp_1283_2 <= 0;
      __tmp_1283_3 <= 0;
      __tmp_1283_4 <= 0;
      __tmp_1283_5 <= 0;
      __tmp_1283_6 <= 0;
      __tmp_1283_7 <= 0;
      __tmp_1283_8 <= 0;
      __tmp_1283_9 <= 0;
      __tmp_1285_1 <= 0;
      __tmp_1285_2 <= 0;
      __tmp_1285_3 <= 0;
      __tmp_1285_4 <= 0;
      __tmp_1285_5 <= 0;
      __tmp_1285_6 <= 0;
      __tmp_1285_7 <= 0;
      __tmp_1285_8 <= 0;
      __tmp_1285_9 <= 0;
    end else begin
      _acc_0_x_idle <= _acc_0_x_idle;
      _acc_0_x_source_ram_rvalid <= 0;
      _acc_0_rshift_idle <= _acc_0_rshift_idle;
      _acc_0_rshift_source_ram_rvalid <= 0;
      _acc_0_sum_sink_wenable <= 0;
      _acc_0_valid_sink_wenable <= 0;
      _greaterthan_data_3 <= acc_0_rshift_data > 1'sd0;
      _minus_data_5 <= acc_0_rshift_data - 2'sd1;
      _reduceadd_data_17 <= _reduceadd_data_17 + acc_0_x_data;
      _reduceadd_count_17 <= (_reduceadd_count_17 >= acc_0_size_data - 1)? 0 : _reduceadd_count_17 + 1;
      if(_acc_0_reduce_reset) begin
        _reduceadd_data_17 <= 1'sd0 + acc_0_x_data;
      end 
      if(_acc_0_reduce_reset) begin
        _reduceadd_count_17 <= 0;
      end 
      if(_reduceadd_count_17 == 0) begin
        _reduceadd_data_17 <= 1'sd0 + acc_0_x_data;
      end 
      _pulse_data_19 <= _pulse_count_19 >= acc_0_size_data - 1;
      _pulse_count_19 <= (_pulse_count_19 >= acc_0_size_data - 1)? 0 : _pulse_count_19 + 1;
      if(_acc_0_reduce_reset) begin
        _pulse_data_19 <= _pulse_count_19 >= acc_0_size_data - 1;
      end 
      if(_acc_0_reduce_reset) begin
        _pulse_count_19 <= 0;
      end 
      if(_pulse_count_19 == 0) begin
        _pulse_data_19 <= _pulse_count_19 >= acc_0_size_data - 1;
      end 
      __delay_data_751 <= acc_0_rshift_data;
      _sll_data_7 <= 2'sd1 << _minus_data_5;
      __delay_data_748 <= _greaterthan_data_3;
      __delay_data_749 <= _reduceadd_data_17;
      __delay_data_752 <= __delay_data_751;
      __delay_data_755 <= _pulse_data_19;
      _cond_data_13 <= (__delay_data_748)? _sll_data_7 : 1'sd0;
      __delay_data_750 <= __delay_data_749;
      __delay_data_753 <= __delay_data_752;
      __delay_data_756 <= __delay_data_755;
      _plus_data_20 <= __delay_data_750 + _cond_data_13;
      __delay_data_754 <= __delay_data_753;
      __delay_data_757 <= __delay_data_756;
      _sra_data_21 <= _plus_data_20 >>> __delay_data_754;
      __delay_data_758 <= __delay_data_757;
      if(_substream_acc_0_x_data_cond_747_36) begin
        __variable_wdata_0 <= __substreamoutput_data_746;
      end 
      if(_substream_acc_0_rshift_data_cond_747_37) begin
        __variable_wdata_1 <= __delay_data_1288;
      end 
      if(_substream_acc_0_size_data_cond_747_38) begin
        __variable_wdata_2 <= __delay_data_1310;
      end 
      __tmp_943_1 <= _tmp_943;
      __tmp_943_2 <= __tmp_943_1;
      __tmp_943_3 <= __tmp_943_2;
      __tmp_943_4 <= __tmp_943_3;
      __tmp_943_5 <= __tmp_943_4;
      __tmp_943_6 <= __tmp_943_5;
      __tmp_943_7 <= __tmp_943_6;
      __tmp_943_8 <= __tmp_943_7;
      __tmp_943_9 <= __tmp_943_8;
      __tmp_945_1 <= _tmp_945;
      __tmp_945_2 <= __tmp_945_1;
      __tmp_945_3 <= __tmp_945_2;
      __tmp_945_4 <= __tmp_945_3;
      __tmp_945_5 <= __tmp_945_4;
      __tmp_945_6 <= __tmp_945_5;
      __tmp_945_7 <= __tmp_945_6;
      __tmp_945_8 <= __tmp_945_7;
      __tmp_945_9 <= __tmp_945_8;
      __tmp_947_1 <= _tmp_947;
      __tmp_947_2 <= __tmp_947_1;
      __tmp_947_3 <= __tmp_947_2;
      __tmp_947_4 <= __tmp_947_3;
      __tmp_947_5 <= __tmp_947_4;
      __tmp_947_6 <= __tmp_947_5;
      __tmp_947_7 <= __tmp_947_6;
      __tmp_947_8 <= __tmp_947_7;
      __tmp_947_9 <= __tmp_947_8;
      if(_substream_acc_0_x_data_cond_879_48) begin
        __variable_wdata_0 <= __substreamoutput_data_878;
      end 
      if(_substream_acc_0_rshift_data_cond_879_49) begin
        __variable_wdata_1 <= __delay_data_1443;
      end 
      if(_substream_acc_0_size_data_cond_879_50) begin
        __variable_wdata_2 <= __delay_data_1459;
      end 
      __tmp_1281_1 <= _tmp_1281;
      __tmp_1281_2 <= __tmp_1281_1;
      __tmp_1281_3 <= __tmp_1281_2;
      __tmp_1281_4 <= __tmp_1281_3;
      __tmp_1281_5 <= __tmp_1281_4;
      __tmp_1281_6 <= __tmp_1281_5;
      __tmp_1281_7 <= __tmp_1281_6;
      __tmp_1281_8 <= __tmp_1281_7;
      __tmp_1281_9 <= __tmp_1281_8;
      __tmp_1283_1 <= _tmp_1283;
      __tmp_1283_2 <= __tmp_1283_1;
      __tmp_1283_3 <= __tmp_1283_2;
      __tmp_1283_4 <= __tmp_1283_3;
      __tmp_1283_5 <= __tmp_1283_4;
      __tmp_1283_6 <= __tmp_1283_5;
      __tmp_1283_7 <= __tmp_1283_6;
      __tmp_1283_8 <= __tmp_1283_7;
      __tmp_1283_9 <= __tmp_1283_8;
      __tmp_1285_1 <= _tmp_1285;
      __tmp_1285_2 <= __tmp_1285_1;
      __tmp_1285_3 <= __tmp_1285_2;
      __tmp_1285_4 <= __tmp_1285_3;
      __tmp_1285_5 <= __tmp_1285_4;
      __tmp_1285_6 <= __tmp_1285_5;
      __tmp_1285_7 <= __tmp_1285_6;
      __tmp_1285_8 <= __tmp_1285_7;
      __tmp_1285_9 <= __tmp_1285_8;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _acc_0_fsm <= _acc_0_fsm_init;
      _acc_0_source_busy <= 0;
      _acc_0_reduce_reset <= 1;
      _substream_acc_0_x_data_cond_747_36 <= 0;
      _substream_acc_0_rshift_data_cond_747_37 <= 0;
      _substream_acc_0_size_data_cond_747_38 <= 0;
      _acc_0_sink_busy <= 0;
      _acc_0_sink_wait_count <= 0;
      _substream_acc_0_x_data_cond_879_48 <= 0;
      _substream_acc_0_rshift_data_cond_879_49 <= 0;
      _substream_acc_0_size_data_cond_879_50 <= 0;
    end else begin
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _acc_0_source_busy <= 1;
      end 
      if(__tmp_787_28) begin
        _acc_0_reduce_reset <= 0;
      end 
      if(__tmp_789_26) begin
        _substream_acc_0_x_data_cond_747_36 <= 1;
      end 
      if(__tmp_791_26) begin
        _substream_acc_0_rshift_data_cond_747_37 <= 1;
      end 
      if(__tmp_793_26) begin
        _substream_acc_0_size_data_cond_747_38 <= 1;
      end 
      if(_stream_conv2d_16_fsm == 3) begin
        _acc_0_source_busy <= 0;
      end 
      if(__tmp_935_24) begin
        _acc_0_reduce_reset <= 1;
      end 
      if(__tmp_937_23) begin
        _substream_acc_0_x_data_cond_747_36 <= 0;
      end 
      if(__tmp_939_23) begin
        _substream_acc_0_rshift_data_cond_747_37 <= 0;
      end 
      if(__tmp_941_23) begin
        _substream_acc_0_size_data_cond_747_38 <= 0;
      end 
      if((_acc_0_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_943_9) begin
        _acc_0_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _acc_0_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_945_9) begin
        _acc_0_sink_wait_count <= _acc_0_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_947_9) begin
        _acc_0_sink_wait_count <= _acc_0_sink_wait_count + 1;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) begin
        _acc_0_source_busy <= 1;
      end 
      if(__tmp_1237_22) begin
        _acc_0_reduce_reset <= 0;
      end 
      if(__tmp_1239_20) begin
        _substream_acc_0_x_data_cond_879_48 <= 1;
      end 
      if(__tmp_1241_20) begin
        _substream_acc_0_rshift_data_cond_879_49 <= 1;
      end 
      if(__tmp_1243_20) begin
        _substream_acc_0_size_data_cond_879_50 <= 1;
      end 
      if(_stream_matmul_29_fsm == 3) begin
        _acc_0_source_busy <= 0;
      end 
      if(__tmp_1273_18) begin
        _acc_0_reduce_reset <= 1;
      end 
      if(__tmp_1275_17) begin
        _substream_acc_0_x_data_cond_879_48 <= 0;
      end 
      if(__tmp_1277_17) begin
        _substream_acc_0_rshift_data_cond_879_49 <= 0;
      end 
      if(__tmp_1279_17) begin
        _substream_acc_0_size_data_cond_879_50 <= 0;
      end 
      if((_acc_0_sink_wait_count == 1) && !((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) && __tmp_1281_9) begin
        _acc_0_sink_busy <= 0;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) begin
        _acc_0_sink_busy <= 1;
      end 
      if(!((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) && __tmp_1283_9) begin
        _acc_0_sink_wait_count <= _acc_0_sink_wait_count - 1;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag && !__tmp_1285_9) begin
        _acc_0_sink_wait_count <= _acc_0_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_1_var0_idle <= 1;
      _add_tree_1_var0_source_ram_rvalid <= 0;
      _add_tree_1_sum_sink_wenable <= 0;
      __variable_wdata_22 <= 0;
      __tmp_1267_1 <= 0;
      __tmp_1267_2 <= 0;
      __tmp_1267_3 <= 0;
      __tmp_1267_4 <= 0;
      __tmp_1269_1 <= 0;
      __tmp_1269_2 <= 0;
      __tmp_1269_3 <= 0;
      __tmp_1269_4 <= 0;
      __tmp_1271_1 <= 0;
      __tmp_1271_2 <= 0;
      __tmp_1271_3 <= 0;
      __tmp_1271_4 <= 0;
    end else begin
      _add_tree_1_var0_idle <= _add_tree_1_var0_idle;
      _add_tree_1_var0_source_ram_rvalid <= 0;
      _add_tree_1_sum_sink_wenable <= 0;
      if(_substream_add_tree_1_var0_data_cond_877_47) begin
        __variable_wdata_22 <= __substreamoutput_data_876;
      end 
      __tmp_1267_1 <= _tmp_1267;
      __tmp_1267_2 <= __tmp_1267_1;
      __tmp_1267_3 <= __tmp_1267_2;
      __tmp_1267_4 <= __tmp_1267_3;
      __tmp_1269_1 <= _tmp_1269;
      __tmp_1269_2 <= __tmp_1269_1;
      __tmp_1269_3 <= __tmp_1269_2;
      __tmp_1269_4 <= __tmp_1269_3;
      __tmp_1271_1 <= _tmp_1271;
      __tmp_1271_2 <= __tmp_1271_1;
      __tmp_1271_3 <= __tmp_1271_2;
      __tmp_1271_4 <= __tmp_1271_3;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_1_fsm <= _add_tree_1_fsm_init;
      _add_tree_1_source_busy <= 0;
      _substream_add_tree_1_var0_data_cond_877_47 <= 0;
      _add_tree_1_sink_busy <= 0;
      _add_tree_1_sink_wait_count <= 0;
    end else begin
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) begin
        _add_tree_1_source_busy <= 1;
      end 
      if(__tmp_1235_18) begin
        _substream_add_tree_1_var0_data_cond_877_47 <= 1;
      end 
      if(_stream_matmul_29_fsm == 3) begin
        _add_tree_1_source_busy <= 0;
      end 
      if(__tmp_1265_15) begin
        _substream_add_tree_1_var0_data_cond_877_47 <= 0;
      end 
      if((_add_tree_1_sink_wait_count == 1) && !((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) && __tmp_1267_4) begin
        _add_tree_1_sink_busy <= 0;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) begin
        _add_tree_1_sink_busy <= 1;
      end 
      if(!((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) && __tmp_1269_4) begin
        _add_tree_1_sink_wait_count <= _add_tree_1_sink_wait_count - 1;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag && !__tmp_1271_4) begin
        _add_tree_1_sink_wait_count <= _add_tree_1_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_2_var0_idle <= 1;
      _add_tree_2_var0_source_ram_rvalid <= 0;
      _add_tree_2_var1_idle <= 1;
      _add_tree_2_var1_source_ram_rvalid <= 0;
      _add_tree_2_var2_idle <= 1;
      _add_tree_2_var2_source_ram_rvalid <= 0;
      _add_tree_2_var3_idle <= 1;
      _add_tree_2_var3_source_ram_rvalid <= 0;
      _add_tree_2_var4_idle <= 1;
      _add_tree_2_var4_source_ram_rvalid <= 0;
      _add_tree_2_var5_idle <= 1;
      _add_tree_2_var5_source_ram_rvalid <= 0;
      _add_tree_2_var6_idle <= 1;
      _add_tree_2_var6_source_ram_rvalid <= 0;
      _add_tree_2_var7_idle <= 1;
      _add_tree_2_var7_source_ram_rvalid <= 0;
      _add_tree_2_var8_idle <= 1;
      _add_tree_2_var8_source_ram_rvalid <= 0;
      _add_tree_2_sum_sink_wenable <= 0;
      __plusn_data_34 <= 0;
      __plusn_data_35 <= 0;
      __plusn_data_36 <= 0;
      __plusn_data_37 <= 0;
      __variable_wdata_24 <= 0;
      __variable_wdata_25 <= 0;
      __variable_wdata_26 <= 0;
      __variable_wdata_27 <= 0;
      __variable_wdata_28 <= 0;
      __variable_wdata_29 <= 0;
      __variable_wdata_30 <= 0;
      __variable_wdata_31 <= 0;
      __variable_wdata_32 <= 0;
      __tmp_929_1 <= 0;
      __tmp_929_2 <= 0;
      __tmp_929_3 <= 0;
      __tmp_929_4 <= 0;
      __tmp_929_5 <= 0;
      __tmp_929_6 <= 0;
      __tmp_931_1 <= 0;
      __tmp_931_2 <= 0;
      __tmp_931_3 <= 0;
      __tmp_931_4 <= 0;
      __tmp_931_5 <= 0;
      __tmp_931_6 <= 0;
      __tmp_933_1 <= 0;
      __tmp_933_2 <= 0;
      __tmp_933_3 <= 0;
      __tmp_933_4 <= 0;
      __tmp_933_5 <= 0;
      __tmp_933_6 <= 0;
    end else begin
      _add_tree_2_var0_idle <= _add_tree_2_var0_idle;
      _add_tree_2_var0_source_ram_rvalid <= 0;
      _add_tree_2_var1_idle <= _add_tree_2_var1_idle;
      _add_tree_2_var1_source_ram_rvalid <= 0;
      _add_tree_2_var2_idle <= _add_tree_2_var2_idle;
      _add_tree_2_var2_source_ram_rvalid <= 0;
      _add_tree_2_var3_idle <= _add_tree_2_var3_idle;
      _add_tree_2_var3_source_ram_rvalid <= 0;
      _add_tree_2_var4_idle <= _add_tree_2_var4_idle;
      _add_tree_2_var4_source_ram_rvalid <= 0;
      _add_tree_2_var5_idle <= _add_tree_2_var5_idle;
      _add_tree_2_var5_source_ram_rvalid <= 0;
      _add_tree_2_var6_idle <= _add_tree_2_var6_idle;
      _add_tree_2_var6_source_ram_rvalid <= 0;
      _add_tree_2_var7_idle <= _add_tree_2_var7_idle;
      _add_tree_2_var7_source_ram_rvalid <= 0;
      _add_tree_2_var8_idle <= _add_tree_2_var8_idle;
      _add_tree_2_var8_source_ram_rvalid <= 0;
      _add_tree_2_sum_sink_wenable <= 0;
      __plusn_data_34 <= add_tree_2_var0_data + add_tree_2_var1_data + add_tree_2_var2_data;
      __plusn_data_35 <= add_tree_2_var3_data + add_tree_2_var4_data + add_tree_2_var5_data;
      __plusn_data_36 <= add_tree_2_var6_data + add_tree_2_var7_data + add_tree_2_var8_data;
      __plusn_data_37 <= __plusn_data_34 + __plusn_data_35 + __plusn_data_36;
      if(_substream_add_tree_2_var0_data_cond_745_27) begin
        __variable_wdata_24 <= __substreamoutput_data_608;
      end 
      if(_substream_add_tree_2_var1_data_cond_745_28) begin
        __variable_wdata_25 <= __substreamoutput_data_625;
      end 
      if(_substream_add_tree_2_var2_data_cond_745_29) begin
        __variable_wdata_26 <= __substreamoutput_data_642;
      end 
      if(_substream_add_tree_2_var3_data_cond_745_30) begin
        __variable_wdata_27 <= __substreamoutput_data_659;
      end 
      if(_substream_add_tree_2_var4_data_cond_745_31) begin
        __variable_wdata_28 <= __substreamoutput_data_676;
      end 
      if(_substream_add_tree_2_var5_data_cond_745_32) begin
        __variable_wdata_29 <= __substreamoutput_data_693;
      end 
      if(_substream_add_tree_2_var6_data_cond_745_33) begin
        __variable_wdata_30 <= __substreamoutput_data_710;
      end 
      if(_substream_add_tree_2_var7_data_cond_745_34) begin
        __variable_wdata_31 <= __substreamoutput_data_727;
      end 
      if(_substream_add_tree_2_var8_data_cond_745_35) begin
        __variable_wdata_32 <= __substreamoutput_data_744;
      end 
      __tmp_929_1 <= _tmp_929;
      __tmp_929_2 <= __tmp_929_1;
      __tmp_929_3 <= __tmp_929_2;
      __tmp_929_4 <= __tmp_929_3;
      __tmp_929_5 <= __tmp_929_4;
      __tmp_929_6 <= __tmp_929_5;
      __tmp_931_1 <= _tmp_931;
      __tmp_931_2 <= __tmp_931_1;
      __tmp_931_3 <= __tmp_931_2;
      __tmp_931_4 <= __tmp_931_3;
      __tmp_931_5 <= __tmp_931_4;
      __tmp_931_6 <= __tmp_931_5;
      __tmp_933_1 <= _tmp_933;
      __tmp_933_2 <= __tmp_933_1;
      __tmp_933_3 <= __tmp_933_2;
      __tmp_933_4 <= __tmp_933_3;
      __tmp_933_5 <= __tmp_933_4;
      __tmp_933_6 <= __tmp_933_5;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_2_fsm <= _add_tree_2_fsm_init;
      _add_tree_2_source_busy <= 0;
      _substream_add_tree_2_var0_data_cond_745_27 <= 0;
      _substream_add_tree_2_var1_data_cond_745_28 <= 0;
      _substream_add_tree_2_var2_data_cond_745_29 <= 0;
      _substream_add_tree_2_var3_data_cond_745_30 <= 0;
      _substream_add_tree_2_var4_data_cond_745_31 <= 0;
      _substream_add_tree_2_var5_data_cond_745_32 <= 0;
      _substream_add_tree_2_var6_data_cond_745_33 <= 0;
      _substream_add_tree_2_var7_data_cond_745_34 <= 0;
      _substream_add_tree_2_var8_data_cond_745_35 <= 0;
      _add_tree_2_sink_busy <= 0;
      _add_tree_2_sink_wait_count <= 0;
    end else begin
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _add_tree_2_source_busy <= 1;
      end 
      if(__tmp_769_22) begin
        _substream_add_tree_2_var0_data_cond_745_27 <= 1;
      end 
      if(__tmp_771_22) begin
        _substream_add_tree_2_var1_data_cond_745_28 <= 1;
      end 
      if(__tmp_773_22) begin
        _substream_add_tree_2_var2_data_cond_745_29 <= 1;
      end 
      if(__tmp_775_22) begin
        _substream_add_tree_2_var3_data_cond_745_30 <= 1;
      end 
      if(__tmp_777_22) begin
        _substream_add_tree_2_var4_data_cond_745_31 <= 1;
      end 
      if(__tmp_779_22) begin
        _substream_add_tree_2_var5_data_cond_745_32 <= 1;
      end 
      if(__tmp_781_22) begin
        _substream_add_tree_2_var6_data_cond_745_33 <= 1;
      end 
      if(__tmp_783_22) begin
        _substream_add_tree_2_var7_data_cond_745_34 <= 1;
      end 
      if(__tmp_785_22) begin
        _substream_add_tree_2_var8_data_cond_745_35 <= 1;
      end 
      if(_stream_conv2d_16_fsm == 3) begin
        _add_tree_2_source_busy <= 0;
      end 
      if(__tmp_911_19) begin
        _substream_add_tree_2_var0_data_cond_745_27 <= 0;
      end 
      if(__tmp_913_19) begin
        _substream_add_tree_2_var1_data_cond_745_28 <= 0;
      end 
      if(__tmp_915_19) begin
        _substream_add_tree_2_var2_data_cond_745_29 <= 0;
      end 
      if(__tmp_917_19) begin
        _substream_add_tree_2_var3_data_cond_745_30 <= 0;
      end 
      if(__tmp_919_19) begin
        _substream_add_tree_2_var4_data_cond_745_31 <= 0;
      end 
      if(__tmp_921_19) begin
        _substream_add_tree_2_var5_data_cond_745_32 <= 0;
      end 
      if(__tmp_923_19) begin
        _substream_add_tree_2_var6_data_cond_745_33 <= 0;
      end 
      if(__tmp_925_19) begin
        _substream_add_tree_2_var7_data_cond_745_34 <= 0;
      end 
      if(__tmp_927_19) begin
        _substream_add_tree_2_var8_data_cond_745_35 <= 0;
      end 
      if((_add_tree_2_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_929_6) begin
        _add_tree_2_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _add_tree_2_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_931_6) begin
        _add_tree_2_sink_wait_count <= _add_tree_2_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_933_6) begin
        _add_tree_2_sink_wait_count <= _add_tree_2_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_clip_3_x_idle <= 1;
      _mul_rshift_clip_3_x_source_ram_rvalid <= 0;
      _mul_rshift_clip_3_y_idle <= 1;
      _mul_rshift_clip_3_y_source_ram_rvalid <= 0;
      _mul_rshift_clip_3_rshift_idle <= 1;
      _mul_rshift_clip_3_rshift_source_ram_rvalid <= 0;
      _mul_rshift_clip_3_z_sink_wenable <= 0;
      _times_mul_odata_reg_41 <= 0;
      __delay_data_764 <= 0;
      __delay_data_765 <= 0;
      __delay_data_766 <= 0;
      __delay_data_767 <= 0;
      _sra_data_42 <= 0;
      _greaterthan_data_43 <= 0;
      _lessthan_data_47 <= 0;
      _greatereq_data_51 <= 0;
      __delay_data_768 <= 0;
      _cond_data_45 <= 0;
      _cond_data_49 <= 0;
      __delay_data_769 <= 0;
      _cond_data_53 <= 0;
      __variable_wdata_38 <= 0;
      __variable_wdata_39 <= 0;
      __variable_wdata_40 <= 0;
      __tmp_955_1 <= 0;
      __tmp_955_2 <= 0;
      __tmp_955_3 <= 0;
      __tmp_955_4 <= 0;
      __tmp_955_5 <= 0;
      __tmp_955_6 <= 0;
      __tmp_955_7 <= 0;
      __tmp_955_8 <= 0;
      __tmp_955_9 <= 0;
      __tmp_955_10 <= 0;
      __tmp_955_11 <= 0;
      __tmp_955_12 <= 0;
      __tmp_957_1 <= 0;
      __tmp_957_2 <= 0;
      __tmp_957_3 <= 0;
      __tmp_957_4 <= 0;
      __tmp_957_5 <= 0;
      __tmp_957_6 <= 0;
      __tmp_957_7 <= 0;
      __tmp_957_8 <= 0;
      __tmp_957_9 <= 0;
      __tmp_957_10 <= 0;
      __tmp_957_11 <= 0;
      __tmp_957_12 <= 0;
      __tmp_959_1 <= 0;
      __tmp_959_2 <= 0;
      __tmp_959_3 <= 0;
      __tmp_959_4 <= 0;
      __tmp_959_5 <= 0;
      __tmp_959_6 <= 0;
      __tmp_959_7 <= 0;
      __tmp_959_8 <= 0;
      __tmp_959_9 <= 0;
      __tmp_959_10 <= 0;
      __tmp_959_11 <= 0;
      __tmp_959_12 <= 0;
      __tmp_1293_1 <= 0;
      __tmp_1293_2 <= 0;
      __tmp_1293_3 <= 0;
      __tmp_1293_4 <= 0;
      __tmp_1293_5 <= 0;
      __tmp_1293_6 <= 0;
      __tmp_1293_7 <= 0;
      __tmp_1293_8 <= 0;
      __tmp_1293_9 <= 0;
      __tmp_1293_10 <= 0;
      __tmp_1293_11 <= 0;
      __tmp_1293_12 <= 0;
      __tmp_1295_1 <= 0;
      __tmp_1295_2 <= 0;
      __tmp_1295_3 <= 0;
      __tmp_1295_4 <= 0;
      __tmp_1295_5 <= 0;
      __tmp_1295_6 <= 0;
      __tmp_1295_7 <= 0;
      __tmp_1295_8 <= 0;
      __tmp_1295_9 <= 0;
      __tmp_1295_10 <= 0;
      __tmp_1295_11 <= 0;
      __tmp_1295_12 <= 0;
      __tmp_1297_1 <= 0;
      __tmp_1297_2 <= 0;
      __tmp_1297_3 <= 0;
      __tmp_1297_4 <= 0;
      __tmp_1297_5 <= 0;
      __tmp_1297_6 <= 0;
      __tmp_1297_7 <= 0;
      __tmp_1297_8 <= 0;
      __tmp_1297_9 <= 0;
      __tmp_1297_10 <= 0;
      __tmp_1297_11 <= 0;
      __tmp_1297_12 <= 0;
    end else begin
      _mul_rshift_clip_3_x_idle <= _mul_rshift_clip_3_x_idle;
      _mul_rshift_clip_3_x_source_ram_rvalid <= 0;
      _mul_rshift_clip_3_y_idle <= _mul_rshift_clip_3_y_idle;
      _mul_rshift_clip_3_y_source_ram_rvalid <= 0;
      _mul_rshift_clip_3_rshift_idle <= _mul_rshift_clip_3_rshift_idle;
      _mul_rshift_clip_3_rshift_source_ram_rvalid <= 0;
      _mul_rshift_clip_3_z_sink_wenable <= 0;
      _times_mul_odata_reg_41 <= _times_mul_odata_41;
      __delay_data_764 <= mul_rshift_clip_3_rshift_data;
      __delay_data_765 <= __delay_data_764;
      __delay_data_766 <= __delay_data_765;
      __delay_data_767 <= __delay_data_766;
      _sra_data_42 <= _times_data_41 >>> __delay_data_767;
      _greaterthan_data_43 <= _sra_data_42 > 8'sd127;
      _lessthan_data_47 <= _sra_data_42 < -8'sd127;
      _greatereq_data_51 <= _sra_data_42 >= 1'sd0;
      __delay_data_768 <= _sra_data_42;
      _cond_data_45 <= (_greaterthan_data_43)? 8'sd127 : __delay_data_768;
      _cond_data_49 <= (_lessthan_data_47)? -8'sd127 : __delay_data_768;
      __delay_data_769 <= _greatereq_data_51;
      _cond_data_53 <= (__delay_data_769)? _cond_data_45 : _cond_data_49;
      if(_substream_mul_rshift_clip_3_x_data_cond_763_39) begin
        __variable_wdata_38 <= _plus_data_762;
      end 
      if(_substream_mul_rshift_clip_3_y_data_cond_763_40) begin
        __variable_wdata_39 <= __delay_data_1368;
      end 
      if(_substream_mul_rshift_clip_3_rshift_data_cond_763_41) begin
        __variable_wdata_40 <= __delay_data_1396;
      end 
      __tmp_955_1 <= _tmp_955;
      __tmp_955_2 <= __tmp_955_1;
      __tmp_955_3 <= __tmp_955_2;
      __tmp_955_4 <= __tmp_955_3;
      __tmp_955_5 <= __tmp_955_4;
      __tmp_955_6 <= __tmp_955_5;
      __tmp_955_7 <= __tmp_955_6;
      __tmp_955_8 <= __tmp_955_7;
      __tmp_955_9 <= __tmp_955_8;
      __tmp_955_10 <= __tmp_955_9;
      __tmp_955_11 <= __tmp_955_10;
      __tmp_955_12 <= __tmp_955_11;
      __tmp_957_1 <= _tmp_957;
      __tmp_957_2 <= __tmp_957_1;
      __tmp_957_3 <= __tmp_957_2;
      __tmp_957_4 <= __tmp_957_3;
      __tmp_957_5 <= __tmp_957_4;
      __tmp_957_6 <= __tmp_957_5;
      __tmp_957_7 <= __tmp_957_6;
      __tmp_957_8 <= __tmp_957_7;
      __tmp_957_9 <= __tmp_957_8;
      __tmp_957_10 <= __tmp_957_9;
      __tmp_957_11 <= __tmp_957_10;
      __tmp_957_12 <= __tmp_957_11;
      __tmp_959_1 <= _tmp_959;
      __tmp_959_2 <= __tmp_959_1;
      __tmp_959_3 <= __tmp_959_2;
      __tmp_959_4 <= __tmp_959_3;
      __tmp_959_5 <= __tmp_959_4;
      __tmp_959_6 <= __tmp_959_5;
      __tmp_959_7 <= __tmp_959_6;
      __tmp_959_8 <= __tmp_959_7;
      __tmp_959_9 <= __tmp_959_8;
      __tmp_959_10 <= __tmp_959_9;
      __tmp_959_11 <= __tmp_959_10;
      __tmp_959_12 <= __tmp_959_11;
      if(_substream_mul_rshift_clip_3_x_data_cond_884_51) begin
        __variable_wdata_38 <= _plus_data_883;
      end 
      if(_substream_mul_rshift_clip_3_y_data_cond_884_52) begin
        __variable_wdata_39 <= __delay_data_1505;
      end 
      if(_substream_mul_rshift_clip_3_rshift_data_cond_884_53) begin
        __variable_wdata_40 <= __delay_data_1527;
      end 
      __tmp_1293_1 <= _tmp_1293;
      __tmp_1293_2 <= __tmp_1293_1;
      __tmp_1293_3 <= __tmp_1293_2;
      __tmp_1293_4 <= __tmp_1293_3;
      __tmp_1293_5 <= __tmp_1293_4;
      __tmp_1293_6 <= __tmp_1293_5;
      __tmp_1293_7 <= __tmp_1293_6;
      __tmp_1293_8 <= __tmp_1293_7;
      __tmp_1293_9 <= __tmp_1293_8;
      __tmp_1293_10 <= __tmp_1293_9;
      __tmp_1293_11 <= __tmp_1293_10;
      __tmp_1293_12 <= __tmp_1293_11;
      __tmp_1295_1 <= _tmp_1295;
      __tmp_1295_2 <= __tmp_1295_1;
      __tmp_1295_3 <= __tmp_1295_2;
      __tmp_1295_4 <= __tmp_1295_3;
      __tmp_1295_5 <= __tmp_1295_4;
      __tmp_1295_6 <= __tmp_1295_5;
      __tmp_1295_7 <= __tmp_1295_6;
      __tmp_1295_8 <= __tmp_1295_7;
      __tmp_1295_9 <= __tmp_1295_8;
      __tmp_1295_10 <= __tmp_1295_9;
      __tmp_1295_11 <= __tmp_1295_10;
      __tmp_1295_12 <= __tmp_1295_11;
      __tmp_1297_1 <= _tmp_1297;
      __tmp_1297_2 <= __tmp_1297_1;
      __tmp_1297_3 <= __tmp_1297_2;
      __tmp_1297_4 <= __tmp_1297_3;
      __tmp_1297_5 <= __tmp_1297_4;
      __tmp_1297_6 <= __tmp_1297_5;
      __tmp_1297_7 <= __tmp_1297_6;
      __tmp_1297_8 <= __tmp_1297_7;
      __tmp_1297_9 <= __tmp_1297_8;
      __tmp_1297_10 <= __tmp_1297_9;
      __tmp_1297_11 <= __tmp_1297_10;
      __tmp_1297_12 <= __tmp_1297_11;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_clip_3_fsm <= _mul_rshift_clip_3_fsm_init;
      _mul_rshift_clip_3_source_busy <= 0;
      _substream_mul_rshift_clip_3_x_data_cond_763_39 <= 0;
      _substream_mul_rshift_clip_3_y_data_cond_763_40 <= 0;
      _substream_mul_rshift_clip_3_rshift_data_cond_763_41 <= 0;
      _mul_rshift_clip_3_sink_busy <= 0;
      _mul_rshift_clip_3_sink_wait_count <= 0;
      _substream_mul_rshift_clip_3_x_data_cond_884_51 <= 0;
      _substream_mul_rshift_clip_3_y_data_cond_884_52 <= 0;
      _substream_mul_rshift_clip_3_rshift_data_cond_884_53 <= 0;
    end else begin
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_rshift_clip_3_source_busy <= 1;
      end 
      if(__tmp_795_34) begin
        _substream_mul_rshift_clip_3_x_data_cond_763_39 <= 1;
      end 
      if(__tmp_797_34) begin
        _substream_mul_rshift_clip_3_y_data_cond_763_40 <= 1;
      end 
      if(__tmp_799_34) begin
        _substream_mul_rshift_clip_3_rshift_data_cond_763_41 <= 1;
      end 
      if(_stream_conv2d_16_fsm == 3) begin
        _mul_rshift_clip_3_source_busy <= 0;
      end 
      if(__tmp_949_31) begin
        _substream_mul_rshift_clip_3_x_data_cond_763_39 <= 0;
      end 
      if(__tmp_951_31) begin
        _substream_mul_rshift_clip_3_y_data_cond_763_40 <= 0;
      end 
      if(__tmp_953_31) begin
        _substream_mul_rshift_clip_3_rshift_data_cond_763_41 <= 0;
      end 
      if((_mul_rshift_clip_3_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_955_12) begin
        _mul_rshift_clip_3_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_rshift_clip_3_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_957_12) begin
        _mul_rshift_clip_3_sink_wait_count <= _mul_rshift_clip_3_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_959_12) begin
        _mul_rshift_clip_3_sink_wait_count <= _mul_rshift_clip_3_sink_wait_count + 1;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) begin
        _mul_rshift_clip_3_source_busy <= 1;
      end 
      if(__tmp_1245_28) begin
        _substream_mul_rshift_clip_3_x_data_cond_884_51 <= 1;
      end 
      if(__tmp_1247_28) begin
        _substream_mul_rshift_clip_3_y_data_cond_884_52 <= 1;
      end 
      if(__tmp_1249_28) begin
        _substream_mul_rshift_clip_3_rshift_data_cond_884_53 <= 1;
      end 
      if(_stream_matmul_29_fsm == 3) begin
        _mul_rshift_clip_3_source_busy <= 0;
      end 
      if(__tmp_1287_25) begin
        _substream_mul_rshift_clip_3_x_data_cond_884_51 <= 0;
      end 
      if(__tmp_1289_25) begin
        _substream_mul_rshift_clip_3_y_data_cond_884_52 <= 0;
      end 
      if(__tmp_1291_25) begin
        _substream_mul_rshift_clip_3_rshift_data_cond_884_53 <= 0;
      end 
      if((_mul_rshift_clip_3_sink_wait_count == 1) && !((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) && __tmp_1293_12) begin
        _mul_rshift_clip_3_sink_busy <= 0;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) begin
        _mul_rshift_clip_3_sink_busy <= 1;
      end 
      if(!((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) && __tmp_1295_12) begin
        _mul_rshift_clip_3_sink_wait_count <= _mul_rshift_clip_3_sink_wait_count - 1;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag && !__tmp_1297_12) begin
        _mul_rshift_clip_3_sink_wait_count <= _mul_rshift_clip_3_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_4_x_idle <= 1;
      _mul_4_x_source_ram_rvalid <= 0;
      _mul_4_y_idle <= 1;
      _mul_4_y_source_ram_rvalid <= 0;
      _mul_4_rshift_idle <= 1;
      _mul_4_rshift_source_ram_rvalid <= 0;
      _mul_4_z_sink_wenable <= 0;
      _greaterthan_data_57 <= 0;
      _minus_data_59 <= 0;
      __delay_data_594 <= 0;
      __delay_data_597 <= 0;
      __delay_data_600 <= 0;
      _sll_data_61 <= 0;
      __delay_data_593 <= 0;
      __delay_data_595 <= 0;
      __delay_data_598 <= 0;
      __delay_data_601 <= 0;
      _cond_data_67 <= 0;
      __delay_data_596 <= 0;
      __delay_data_599 <= 0;
      __delay_data_602 <= 0;
      __muladd_madd_odata_reg_69 <= 0;
      __delay_data_603 <= 0;
      __delay_data_604 <= 0;
      __delay_data_605 <= 0;
      __delay_data_606 <= 0;
      _sra_data_70 <= 0;
      __variable_wdata_54 <= 0;
      __variable_wdata_55 <= 0;
      __variable_wdata_56 <= 0;
      __tmp_809_1 <= 0;
      __tmp_809_2 <= 0;
      __tmp_809_3 <= 0;
      __tmp_809_4 <= 0;
      __tmp_809_5 <= 0;
      __tmp_809_6 <= 0;
      __tmp_809_7 <= 0;
      __tmp_809_8 <= 0;
      __tmp_809_9 <= 0;
      __tmp_809_10 <= 0;
      __tmp_809_11 <= 0;
      __tmp_809_12 <= 0;
      __tmp_811_1 <= 0;
      __tmp_811_2 <= 0;
      __tmp_811_3 <= 0;
      __tmp_811_4 <= 0;
      __tmp_811_5 <= 0;
      __tmp_811_6 <= 0;
      __tmp_811_7 <= 0;
      __tmp_811_8 <= 0;
      __tmp_811_9 <= 0;
      __tmp_811_10 <= 0;
      __tmp_811_11 <= 0;
      __tmp_811_12 <= 0;
      __tmp_813_1 <= 0;
      __tmp_813_2 <= 0;
      __tmp_813_3 <= 0;
      __tmp_813_4 <= 0;
      __tmp_813_5 <= 0;
      __tmp_813_6 <= 0;
      __tmp_813_7 <= 0;
      __tmp_813_8 <= 0;
      __tmp_813_9 <= 0;
      __tmp_813_10 <= 0;
      __tmp_813_11 <= 0;
      __tmp_813_12 <= 0;
      __tmp_1259_1 <= 0;
      __tmp_1259_2 <= 0;
      __tmp_1259_3 <= 0;
      __tmp_1259_4 <= 0;
      __tmp_1259_5 <= 0;
      __tmp_1259_6 <= 0;
      __tmp_1259_7 <= 0;
      __tmp_1259_8 <= 0;
      __tmp_1259_9 <= 0;
      __tmp_1259_10 <= 0;
      __tmp_1259_11 <= 0;
      __tmp_1259_12 <= 0;
      __tmp_1261_1 <= 0;
      __tmp_1261_2 <= 0;
      __tmp_1261_3 <= 0;
      __tmp_1261_4 <= 0;
      __tmp_1261_5 <= 0;
      __tmp_1261_6 <= 0;
      __tmp_1261_7 <= 0;
      __tmp_1261_8 <= 0;
      __tmp_1261_9 <= 0;
      __tmp_1261_10 <= 0;
      __tmp_1261_11 <= 0;
      __tmp_1261_12 <= 0;
      __tmp_1263_1 <= 0;
      __tmp_1263_2 <= 0;
      __tmp_1263_3 <= 0;
      __tmp_1263_4 <= 0;
      __tmp_1263_5 <= 0;
      __tmp_1263_6 <= 0;
      __tmp_1263_7 <= 0;
      __tmp_1263_8 <= 0;
      __tmp_1263_9 <= 0;
      __tmp_1263_10 <= 0;
      __tmp_1263_11 <= 0;
      __tmp_1263_12 <= 0;
    end else begin
      _mul_4_x_idle <= _mul_4_x_idle;
      _mul_4_x_source_ram_rvalid <= 0;
      _mul_4_y_idle <= _mul_4_y_idle;
      _mul_4_y_source_ram_rvalid <= 0;
      _mul_4_rshift_idle <= _mul_4_rshift_idle;
      _mul_4_rshift_source_ram_rvalid <= 0;
      _mul_4_z_sink_wenable <= 0;
      _greaterthan_data_57 <= mul_4_rshift_data > 1'sd0;
      _minus_data_59 <= mul_4_rshift_data - 2'sd1;
      __delay_data_594 <= mul_4_x_data;
      __delay_data_597 <= mul_4_y_data;
      __delay_data_600 <= mul_4_rshift_data;
      _sll_data_61 <= 2'sd1 << _minus_data_59;
      __delay_data_593 <= _greaterthan_data_57;
      __delay_data_595 <= __delay_data_594;
      __delay_data_598 <= __delay_data_597;
      __delay_data_601 <= __delay_data_600;
      _cond_data_67 <= (__delay_data_593)? _sll_data_61 : 1'sd0;
      __delay_data_596 <= __delay_data_595;
      __delay_data_599 <= __delay_data_598;
      __delay_data_602 <= __delay_data_601;
      __muladd_madd_odata_reg_69 <= __muladd_madd_odata_69;
      __delay_data_603 <= __delay_data_602;
      __delay_data_604 <= __delay_data_603;
      __delay_data_605 <= __delay_data_604;
      __delay_data_606 <= __delay_data_605;
      _sra_data_70 <= __muladd_data_69 >>> __delay_data_606;
      if(_substream_mul_4_x_data_cond_592_0) begin
        __variable_wdata_54 <= _cond_data_575;
      end 
      if(_substream_mul_4_y_data_cond_592_1) begin
        __variable_wdata_55 <= __delay_data_955;
      end 
      if(_substream_mul_4_rshift_data_cond_592_2) begin
        __variable_wdata_56 <= __delay_data_961;
      end 
      __tmp_809_1 <= _tmp_809;
      __tmp_809_2 <= __tmp_809_1;
      __tmp_809_3 <= __tmp_809_2;
      __tmp_809_4 <= __tmp_809_3;
      __tmp_809_5 <= __tmp_809_4;
      __tmp_809_6 <= __tmp_809_5;
      __tmp_809_7 <= __tmp_809_6;
      __tmp_809_8 <= __tmp_809_7;
      __tmp_809_9 <= __tmp_809_8;
      __tmp_809_10 <= __tmp_809_9;
      __tmp_809_11 <= __tmp_809_10;
      __tmp_809_12 <= __tmp_809_11;
      __tmp_811_1 <= _tmp_811;
      __tmp_811_2 <= __tmp_811_1;
      __tmp_811_3 <= __tmp_811_2;
      __tmp_811_4 <= __tmp_811_3;
      __tmp_811_5 <= __tmp_811_4;
      __tmp_811_6 <= __tmp_811_5;
      __tmp_811_7 <= __tmp_811_6;
      __tmp_811_8 <= __tmp_811_7;
      __tmp_811_9 <= __tmp_811_8;
      __tmp_811_10 <= __tmp_811_9;
      __tmp_811_11 <= __tmp_811_10;
      __tmp_811_12 <= __tmp_811_11;
      __tmp_813_1 <= _tmp_813;
      __tmp_813_2 <= __tmp_813_1;
      __tmp_813_3 <= __tmp_813_2;
      __tmp_813_4 <= __tmp_813_3;
      __tmp_813_5 <= __tmp_813_4;
      __tmp_813_6 <= __tmp_813_5;
      __tmp_813_7 <= __tmp_813_6;
      __tmp_813_8 <= __tmp_813_7;
      __tmp_813_9 <= __tmp_813_8;
      __tmp_813_10 <= __tmp_813_9;
      __tmp_813_11 <= __tmp_813_10;
      __tmp_813_12 <= __tmp_813_11;
      if(_substream_mul_4_x_data_cond_874_44) begin
        __variable_wdata_54 <= _cond_data_873;
      end 
      if(_substream_mul_4_y_data_cond_874_45) begin
        __variable_wdata_55 <= __delay_data_1426;
      end 
      if(_substream_mul_4_rshift_data_cond_874_46) begin
        __variable_wdata_56 <= __delay_data_1428;
      end 
      __tmp_1259_1 <= _tmp_1259;
      __tmp_1259_2 <= __tmp_1259_1;
      __tmp_1259_3 <= __tmp_1259_2;
      __tmp_1259_4 <= __tmp_1259_3;
      __tmp_1259_5 <= __tmp_1259_4;
      __tmp_1259_6 <= __tmp_1259_5;
      __tmp_1259_7 <= __tmp_1259_6;
      __tmp_1259_8 <= __tmp_1259_7;
      __tmp_1259_9 <= __tmp_1259_8;
      __tmp_1259_10 <= __tmp_1259_9;
      __tmp_1259_11 <= __tmp_1259_10;
      __tmp_1259_12 <= __tmp_1259_11;
      __tmp_1261_1 <= _tmp_1261;
      __tmp_1261_2 <= __tmp_1261_1;
      __tmp_1261_3 <= __tmp_1261_2;
      __tmp_1261_4 <= __tmp_1261_3;
      __tmp_1261_5 <= __tmp_1261_4;
      __tmp_1261_6 <= __tmp_1261_5;
      __tmp_1261_7 <= __tmp_1261_6;
      __tmp_1261_8 <= __tmp_1261_7;
      __tmp_1261_9 <= __tmp_1261_8;
      __tmp_1261_10 <= __tmp_1261_9;
      __tmp_1261_11 <= __tmp_1261_10;
      __tmp_1261_12 <= __tmp_1261_11;
      __tmp_1263_1 <= _tmp_1263;
      __tmp_1263_2 <= __tmp_1263_1;
      __tmp_1263_3 <= __tmp_1263_2;
      __tmp_1263_4 <= __tmp_1263_3;
      __tmp_1263_5 <= __tmp_1263_4;
      __tmp_1263_6 <= __tmp_1263_5;
      __tmp_1263_7 <= __tmp_1263_6;
      __tmp_1263_8 <= __tmp_1263_7;
      __tmp_1263_9 <= __tmp_1263_8;
      __tmp_1263_10 <= __tmp_1263_9;
      __tmp_1263_11 <= __tmp_1263_10;
      __tmp_1263_12 <= __tmp_1263_11;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_4_fsm <= _mul_4_fsm_init;
      _mul_4_source_busy <= 0;
      _substream_mul_4_x_data_cond_592_0 <= 0;
      _substream_mul_4_y_data_cond_592_1 <= 0;
      _substream_mul_4_rshift_data_cond_592_2 <= 0;
      _mul_4_sink_busy <= 0;
      _mul_4_sink_wait_count <= 0;
      _substream_mul_4_x_data_cond_874_44 <= 0;
      _substream_mul_4_y_data_cond_874_45 <= 0;
      _substream_mul_4_rshift_data_cond_874_46 <= 0;
    end else begin
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_4_source_busy <= 1;
      end 
      if(__tmp_715_12) begin
        _substream_mul_4_x_data_cond_592_0 <= 1;
      end 
      if(__tmp_717_12) begin
        _substream_mul_4_y_data_cond_592_1 <= 1;
      end 
      if(__tmp_719_12) begin
        _substream_mul_4_rshift_data_cond_592_2 <= 1;
      end 
      if(_stream_conv2d_16_fsm == 3) begin
        _mul_4_source_busy <= 0;
      end 
      if(__tmp_803_9) begin
        _substream_mul_4_x_data_cond_592_0 <= 0;
      end 
      if(__tmp_805_9) begin
        _substream_mul_4_y_data_cond_592_1 <= 0;
      end 
      if(__tmp_807_9) begin
        _substream_mul_4_rshift_data_cond_592_2 <= 0;
      end 
      if((_mul_4_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_809_12) begin
        _mul_4_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_4_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_811_12) begin
        _mul_4_sink_wait_count <= _mul_4_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_813_12) begin
        _mul_4_sink_wait_count <= _mul_4_sink_wait_count + 1;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) begin
        _mul_4_source_busy <= 1;
      end 
      if(__tmp_1229_8) begin
        _substream_mul_4_x_data_cond_874_44 <= 1;
      end 
      if(__tmp_1231_8) begin
        _substream_mul_4_y_data_cond_874_45 <= 1;
      end 
      if(__tmp_1233_8) begin
        _substream_mul_4_rshift_data_cond_874_46 <= 1;
      end 
      if(_stream_matmul_29_fsm == 3) begin
        _mul_4_source_busy <= 0;
      end 
      if(__tmp_1253_5) begin
        _substream_mul_4_x_data_cond_874_44 <= 0;
      end 
      if(__tmp_1255_5) begin
        _substream_mul_4_y_data_cond_874_45 <= 0;
      end 
      if(__tmp_1257_5) begin
        _substream_mul_4_rshift_data_cond_874_46 <= 0;
      end 
      if((_mul_4_sink_wait_count == 1) && !((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) && __tmp_1259_12) begin
        _mul_4_sink_busy <= 0;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) begin
        _mul_4_sink_busy <= 1;
      end 
      if(!((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) && __tmp_1261_12) begin
        _mul_4_sink_wait_count <= _mul_4_sink_wait_count - 1;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag && !__tmp_1263_12) begin
        _mul_4_sink_wait_count <= _mul_4_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_5_x_idle <= 1;
      _mul_5_x_source_ram_rvalid <= 0;
      _mul_5_y_idle <= 1;
      _mul_5_y_source_ram_rvalid <= 0;
      _mul_5_rshift_idle <= 1;
      _mul_5_rshift_source_ram_rvalid <= 0;
      _mul_5_z_sink_wenable <= 0;
      _greaterthan_data_74 <= 0;
      _minus_data_76 <= 0;
      __delay_data_611 <= 0;
      __delay_data_614 <= 0;
      __delay_data_617 <= 0;
      _sll_data_78 <= 0;
      __delay_data_610 <= 0;
      __delay_data_612 <= 0;
      __delay_data_615 <= 0;
      __delay_data_618 <= 0;
      _cond_data_84 <= 0;
      __delay_data_613 <= 0;
      __delay_data_616 <= 0;
      __delay_data_619 <= 0;
      __muladd_madd_odata_reg_86 <= 0;
      __delay_data_620 <= 0;
      __delay_data_621 <= 0;
      __delay_data_622 <= 0;
      __delay_data_623 <= 0;
      _sra_data_87 <= 0;
      __variable_wdata_71 <= 0;
      __variable_wdata_72 <= 0;
      __variable_wdata_73 <= 0;
      __tmp_821_1 <= 0;
      __tmp_821_2 <= 0;
      __tmp_821_3 <= 0;
      __tmp_821_4 <= 0;
      __tmp_821_5 <= 0;
      __tmp_821_6 <= 0;
      __tmp_821_7 <= 0;
      __tmp_821_8 <= 0;
      __tmp_821_9 <= 0;
      __tmp_821_10 <= 0;
      __tmp_821_11 <= 0;
      __tmp_821_12 <= 0;
      __tmp_823_1 <= 0;
      __tmp_823_2 <= 0;
      __tmp_823_3 <= 0;
      __tmp_823_4 <= 0;
      __tmp_823_5 <= 0;
      __tmp_823_6 <= 0;
      __tmp_823_7 <= 0;
      __tmp_823_8 <= 0;
      __tmp_823_9 <= 0;
      __tmp_823_10 <= 0;
      __tmp_823_11 <= 0;
      __tmp_823_12 <= 0;
      __tmp_825_1 <= 0;
      __tmp_825_2 <= 0;
      __tmp_825_3 <= 0;
      __tmp_825_4 <= 0;
      __tmp_825_5 <= 0;
      __tmp_825_6 <= 0;
      __tmp_825_7 <= 0;
      __tmp_825_8 <= 0;
      __tmp_825_9 <= 0;
      __tmp_825_10 <= 0;
      __tmp_825_11 <= 0;
      __tmp_825_12 <= 0;
    end else begin
      _mul_5_x_idle <= _mul_5_x_idle;
      _mul_5_x_source_ram_rvalid <= 0;
      _mul_5_y_idle <= _mul_5_y_idle;
      _mul_5_y_source_ram_rvalid <= 0;
      _mul_5_rshift_idle <= _mul_5_rshift_idle;
      _mul_5_rshift_source_ram_rvalid <= 0;
      _mul_5_z_sink_wenable <= 0;
      _greaterthan_data_74 <= mul_5_rshift_data > 1'sd0;
      _minus_data_76 <= mul_5_rshift_data - 2'sd1;
      __delay_data_611 <= mul_5_x_data;
      __delay_data_614 <= mul_5_y_data;
      __delay_data_617 <= mul_5_rshift_data;
      _sll_data_78 <= 2'sd1 << _minus_data_76;
      __delay_data_610 <= _greaterthan_data_74;
      __delay_data_612 <= __delay_data_611;
      __delay_data_615 <= __delay_data_614;
      __delay_data_618 <= __delay_data_617;
      _cond_data_84 <= (__delay_data_610)? _sll_data_78 : 1'sd0;
      __delay_data_613 <= __delay_data_612;
      __delay_data_616 <= __delay_data_615;
      __delay_data_619 <= __delay_data_618;
      __muladd_madd_odata_reg_86 <= __muladd_madd_odata_86;
      __delay_data_620 <= __delay_data_619;
      __delay_data_621 <= __delay_data_620;
      __delay_data_622 <= __delay_data_621;
      __delay_data_623 <= __delay_data_622;
      _sra_data_87 <= __muladd_data_86 >>> __delay_data_623;
      if(_substream_mul_5_x_data_cond_609_3) begin
        __variable_wdata_71 <= _cond_data_577;
      end 
      if(_substream_mul_5_y_data_cond_609_4) begin
        __variable_wdata_72 <= __delay_data_1006;
      end 
      if(_substream_mul_5_rshift_data_cond_609_5) begin
        __variable_wdata_73 <= __delay_data_1012;
      end 
      __tmp_821_1 <= _tmp_821;
      __tmp_821_2 <= __tmp_821_1;
      __tmp_821_3 <= __tmp_821_2;
      __tmp_821_4 <= __tmp_821_3;
      __tmp_821_5 <= __tmp_821_4;
      __tmp_821_6 <= __tmp_821_5;
      __tmp_821_7 <= __tmp_821_6;
      __tmp_821_8 <= __tmp_821_7;
      __tmp_821_9 <= __tmp_821_8;
      __tmp_821_10 <= __tmp_821_9;
      __tmp_821_11 <= __tmp_821_10;
      __tmp_821_12 <= __tmp_821_11;
      __tmp_823_1 <= _tmp_823;
      __tmp_823_2 <= __tmp_823_1;
      __tmp_823_3 <= __tmp_823_2;
      __tmp_823_4 <= __tmp_823_3;
      __tmp_823_5 <= __tmp_823_4;
      __tmp_823_6 <= __tmp_823_5;
      __tmp_823_7 <= __tmp_823_6;
      __tmp_823_8 <= __tmp_823_7;
      __tmp_823_9 <= __tmp_823_8;
      __tmp_823_10 <= __tmp_823_9;
      __tmp_823_11 <= __tmp_823_10;
      __tmp_823_12 <= __tmp_823_11;
      __tmp_825_1 <= _tmp_825;
      __tmp_825_2 <= __tmp_825_1;
      __tmp_825_3 <= __tmp_825_2;
      __tmp_825_4 <= __tmp_825_3;
      __tmp_825_5 <= __tmp_825_4;
      __tmp_825_6 <= __tmp_825_5;
      __tmp_825_7 <= __tmp_825_6;
      __tmp_825_8 <= __tmp_825_7;
      __tmp_825_9 <= __tmp_825_8;
      __tmp_825_10 <= __tmp_825_9;
      __tmp_825_11 <= __tmp_825_10;
      __tmp_825_12 <= __tmp_825_11;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_5_fsm <= _mul_5_fsm_init;
      _mul_5_source_busy <= 0;
      _substream_mul_5_x_data_cond_609_3 <= 0;
      _substream_mul_5_y_data_cond_609_4 <= 0;
      _substream_mul_5_rshift_data_cond_609_5 <= 0;
      _mul_5_sink_busy <= 0;
      _mul_5_sink_wait_count <= 0;
    end else begin
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_5_source_busy <= 1;
      end 
      if(__tmp_721_12) begin
        _substream_mul_5_x_data_cond_609_3 <= 1;
      end 
      if(__tmp_723_12) begin
        _substream_mul_5_y_data_cond_609_4 <= 1;
      end 
      if(__tmp_725_12) begin
        _substream_mul_5_rshift_data_cond_609_5 <= 1;
      end 
      if(_stream_conv2d_16_fsm == 3) begin
        _mul_5_source_busy <= 0;
      end 
      if(__tmp_815_9) begin
        _substream_mul_5_x_data_cond_609_3 <= 0;
      end 
      if(__tmp_817_9) begin
        _substream_mul_5_y_data_cond_609_4 <= 0;
      end 
      if(__tmp_819_9) begin
        _substream_mul_5_rshift_data_cond_609_5 <= 0;
      end 
      if((_mul_5_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_821_12) begin
        _mul_5_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_5_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_823_12) begin
        _mul_5_sink_wait_count <= _mul_5_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_825_12) begin
        _mul_5_sink_wait_count <= _mul_5_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_6_x_idle <= 1;
      _mul_6_x_source_ram_rvalid <= 0;
      _mul_6_y_idle <= 1;
      _mul_6_y_source_ram_rvalid <= 0;
      _mul_6_rshift_idle <= 1;
      _mul_6_rshift_source_ram_rvalid <= 0;
      _mul_6_z_sink_wenable <= 0;
      _greaterthan_data_91 <= 0;
      _minus_data_93 <= 0;
      __delay_data_628 <= 0;
      __delay_data_631 <= 0;
      __delay_data_634 <= 0;
      _sll_data_95 <= 0;
      __delay_data_627 <= 0;
      __delay_data_629 <= 0;
      __delay_data_632 <= 0;
      __delay_data_635 <= 0;
      _cond_data_101 <= 0;
      __delay_data_630 <= 0;
      __delay_data_633 <= 0;
      __delay_data_636 <= 0;
      __muladd_madd_odata_reg_103 <= 0;
      __delay_data_637 <= 0;
      __delay_data_638 <= 0;
      __delay_data_639 <= 0;
      __delay_data_640 <= 0;
      _sra_data_104 <= 0;
      __variable_wdata_88 <= 0;
      __variable_wdata_89 <= 0;
      __variable_wdata_90 <= 0;
      __tmp_833_1 <= 0;
      __tmp_833_2 <= 0;
      __tmp_833_3 <= 0;
      __tmp_833_4 <= 0;
      __tmp_833_5 <= 0;
      __tmp_833_6 <= 0;
      __tmp_833_7 <= 0;
      __tmp_833_8 <= 0;
      __tmp_833_9 <= 0;
      __tmp_833_10 <= 0;
      __tmp_833_11 <= 0;
      __tmp_833_12 <= 0;
      __tmp_835_1 <= 0;
      __tmp_835_2 <= 0;
      __tmp_835_3 <= 0;
      __tmp_835_4 <= 0;
      __tmp_835_5 <= 0;
      __tmp_835_6 <= 0;
      __tmp_835_7 <= 0;
      __tmp_835_8 <= 0;
      __tmp_835_9 <= 0;
      __tmp_835_10 <= 0;
      __tmp_835_11 <= 0;
      __tmp_835_12 <= 0;
      __tmp_837_1 <= 0;
      __tmp_837_2 <= 0;
      __tmp_837_3 <= 0;
      __tmp_837_4 <= 0;
      __tmp_837_5 <= 0;
      __tmp_837_6 <= 0;
      __tmp_837_7 <= 0;
      __tmp_837_8 <= 0;
      __tmp_837_9 <= 0;
      __tmp_837_10 <= 0;
      __tmp_837_11 <= 0;
      __tmp_837_12 <= 0;
    end else begin
      _mul_6_x_idle <= _mul_6_x_idle;
      _mul_6_x_source_ram_rvalid <= 0;
      _mul_6_y_idle <= _mul_6_y_idle;
      _mul_6_y_source_ram_rvalid <= 0;
      _mul_6_rshift_idle <= _mul_6_rshift_idle;
      _mul_6_rshift_source_ram_rvalid <= 0;
      _mul_6_z_sink_wenable <= 0;
      _greaterthan_data_91 <= mul_6_rshift_data > 1'sd0;
      _minus_data_93 <= mul_6_rshift_data - 2'sd1;
      __delay_data_628 <= mul_6_x_data;
      __delay_data_631 <= mul_6_y_data;
      __delay_data_634 <= mul_6_rshift_data;
      _sll_data_95 <= 2'sd1 << _minus_data_93;
      __delay_data_627 <= _greaterthan_data_91;
      __delay_data_629 <= __delay_data_628;
      __delay_data_632 <= __delay_data_631;
      __delay_data_635 <= __delay_data_634;
      _cond_data_101 <= (__delay_data_627)? _sll_data_95 : 1'sd0;
      __delay_data_630 <= __delay_data_629;
      __delay_data_633 <= __delay_data_632;
      __delay_data_636 <= __delay_data_635;
      __muladd_madd_odata_reg_103 <= __muladd_madd_odata_103;
      __delay_data_637 <= __delay_data_636;
      __delay_data_638 <= __delay_data_637;
      __delay_data_639 <= __delay_data_638;
      __delay_data_640 <= __delay_data_639;
      _sra_data_104 <= __muladd_data_103 >>> __delay_data_640;
      if(_substream_mul_6_x_data_cond_626_6) begin
        __variable_wdata_88 <= _cond_data_579;
      end 
      if(_substream_mul_6_y_data_cond_626_7) begin
        __variable_wdata_89 <= __delay_data_1054;
      end 
      if(_substream_mul_6_rshift_data_cond_626_8) begin
        __variable_wdata_90 <= __delay_data_1060;
      end 
      __tmp_833_1 <= _tmp_833;
      __tmp_833_2 <= __tmp_833_1;
      __tmp_833_3 <= __tmp_833_2;
      __tmp_833_4 <= __tmp_833_3;
      __tmp_833_5 <= __tmp_833_4;
      __tmp_833_6 <= __tmp_833_5;
      __tmp_833_7 <= __tmp_833_6;
      __tmp_833_8 <= __tmp_833_7;
      __tmp_833_9 <= __tmp_833_8;
      __tmp_833_10 <= __tmp_833_9;
      __tmp_833_11 <= __tmp_833_10;
      __tmp_833_12 <= __tmp_833_11;
      __tmp_835_1 <= _tmp_835;
      __tmp_835_2 <= __tmp_835_1;
      __tmp_835_3 <= __tmp_835_2;
      __tmp_835_4 <= __tmp_835_3;
      __tmp_835_5 <= __tmp_835_4;
      __tmp_835_6 <= __tmp_835_5;
      __tmp_835_7 <= __tmp_835_6;
      __tmp_835_8 <= __tmp_835_7;
      __tmp_835_9 <= __tmp_835_8;
      __tmp_835_10 <= __tmp_835_9;
      __tmp_835_11 <= __tmp_835_10;
      __tmp_835_12 <= __tmp_835_11;
      __tmp_837_1 <= _tmp_837;
      __tmp_837_2 <= __tmp_837_1;
      __tmp_837_3 <= __tmp_837_2;
      __tmp_837_4 <= __tmp_837_3;
      __tmp_837_5 <= __tmp_837_4;
      __tmp_837_6 <= __tmp_837_5;
      __tmp_837_7 <= __tmp_837_6;
      __tmp_837_8 <= __tmp_837_7;
      __tmp_837_9 <= __tmp_837_8;
      __tmp_837_10 <= __tmp_837_9;
      __tmp_837_11 <= __tmp_837_10;
      __tmp_837_12 <= __tmp_837_11;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_6_fsm <= _mul_6_fsm_init;
      _mul_6_source_busy <= 0;
      _substream_mul_6_x_data_cond_626_6 <= 0;
      _substream_mul_6_y_data_cond_626_7 <= 0;
      _substream_mul_6_rshift_data_cond_626_8 <= 0;
      _mul_6_sink_busy <= 0;
      _mul_6_sink_wait_count <= 0;
    end else begin
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_6_source_busy <= 1;
      end 
      if(__tmp_727_12) begin
        _substream_mul_6_x_data_cond_626_6 <= 1;
      end 
      if(__tmp_729_12) begin
        _substream_mul_6_y_data_cond_626_7 <= 1;
      end 
      if(__tmp_731_12) begin
        _substream_mul_6_rshift_data_cond_626_8 <= 1;
      end 
      if(_stream_conv2d_16_fsm == 3) begin
        _mul_6_source_busy <= 0;
      end 
      if(__tmp_827_9) begin
        _substream_mul_6_x_data_cond_626_6 <= 0;
      end 
      if(__tmp_829_9) begin
        _substream_mul_6_y_data_cond_626_7 <= 0;
      end 
      if(__tmp_831_9) begin
        _substream_mul_6_rshift_data_cond_626_8 <= 0;
      end 
      if((_mul_6_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_833_12) begin
        _mul_6_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_6_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_835_12) begin
        _mul_6_sink_wait_count <= _mul_6_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_837_12) begin
        _mul_6_sink_wait_count <= _mul_6_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_7_x_idle <= 1;
      _mul_7_x_source_ram_rvalid <= 0;
      _mul_7_y_idle <= 1;
      _mul_7_y_source_ram_rvalid <= 0;
      _mul_7_rshift_idle <= 1;
      _mul_7_rshift_source_ram_rvalid <= 0;
      _mul_7_z_sink_wenable <= 0;
      _greaterthan_data_108 <= 0;
      _minus_data_110 <= 0;
      __delay_data_645 <= 0;
      __delay_data_648 <= 0;
      __delay_data_651 <= 0;
      _sll_data_112 <= 0;
      __delay_data_644 <= 0;
      __delay_data_646 <= 0;
      __delay_data_649 <= 0;
      __delay_data_652 <= 0;
      _cond_data_118 <= 0;
      __delay_data_647 <= 0;
      __delay_data_650 <= 0;
      __delay_data_653 <= 0;
      __muladd_madd_odata_reg_120 <= 0;
      __delay_data_654 <= 0;
      __delay_data_655 <= 0;
      __delay_data_656 <= 0;
      __delay_data_657 <= 0;
      _sra_data_121 <= 0;
      __variable_wdata_105 <= 0;
      __variable_wdata_106 <= 0;
      __variable_wdata_107 <= 0;
      __tmp_845_1 <= 0;
      __tmp_845_2 <= 0;
      __tmp_845_3 <= 0;
      __tmp_845_4 <= 0;
      __tmp_845_5 <= 0;
      __tmp_845_6 <= 0;
      __tmp_845_7 <= 0;
      __tmp_845_8 <= 0;
      __tmp_845_9 <= 0;
      __tmp_845_10 <= 0;
      __tmp_845_11 <= 0;
      __tmp_845_12 <= 0;
      __tmp_847_1 <= 0;
      __tmp_847_2 <= 0;
      __tmp_847_3 <= 0;
      __tmp_847_4 <= 0;
      __tmp_847_5 <= 0;
      __tmp_847_6 <= 0;
      __tmp_847_7 <= 0;
      __tmp_847_8 <= 0;
      __tmp_847_9 <= 0;
      __tmp_847_10 <= 0;
      __tmp_847_11 <= 0;
      __tmp_847_12 <= 0;
      __tmp_849_1 <= 0;
      __tmp_849_2 <= 0;
      __tmp_849_3 <= 0;
      __tmp_849_4 <= 0;
      __tmp_849_5 <= 0;
      __tmp_849_6 <= 0;
      __tmp_849_7 <= 0;
      __tmp_849_8 <= 0;
      __tmp_849_9 <= 0;
      __tmp_849_10 <= 0;
      __tmp_849_11 <= 0;
      __tmp_849_12 <= 0;
    end else begin
      _mul_7_x_idle <= _mul_7_x_idle;
      _mul_7_x_source_ram_rvalid <= 0;
      _mul_7_y_idle <= _mul_7_y_idle;
      _mul_7_y_source_ram_rvalid <= 0;
      _mul_7_rshift_idle <= _mul_7_rshift_idle;
      _mul_7_rshift_source_ram_rvalid <= 0;
      _mul_7_z_sink_wenable <= 0;
      _greaterthan_data_108 <= mul_7_rshift_data > 1'sd0;
      _minus_data_110 <= mul_7_rshift_data - 2'sd1;
      __delay_data_645 <= mul_7_x_data;
      __delay_data_648 <= mul_7_y_data;
      __delay_data_651 <= mul_7_rshift_data;
      _sll_data_112 <= 2'sd1 << _minus_data_110;
      __delay_data_644 <= _greaterthan_data_108;
      __delay_data_646 <= __delay_data_645;
      __delay_data_649 <= __delay_data_648;
      __delay_data_652 <= __delay_data_651;
      _cond_data_118 <= (__delay_data_644)? _sll_data_112 : 1'sd0;
      __delay_data_647 <= __delay_data_646;
      __delay_data_650 <= __delay_data_649;
      __delay_data_653 <= __delay_data_652;
      __muladd_madd_odata_reg_120 <= __muladd_madd_odata_120;
      __delay_data_654 <= __delay_data_653;
      __delay_data_655 <= __delay_data_654;
      __delay_data_656 <= __delay_data_655;
      __delay_data_657 <= __delay_data_656;
      _sra_data_121 <= __muladd_data_120 >>> __delay_data_657;
      if(_substream_mul_7_x_data_cond_643_9) begin
        __variable_wdata_105 <= _cond_data_581;
      end 
      if(_substream_mul_7_y_data_cond_643_10) begin
        __variable_wdata_106 <= __delay_data_1089;
      end 
      if(_substream_mul_7_rshift_data_cond_643_11) begin
        __variable_wdata_107 <= __delay_data_1095;
      end 
      __tmp_845_1 <= _tmp_845;
      __tmp_845_2 <= __tmp_845_1;
      __tmp_845_3 <= __tmp_845_2;
      __tmp_845_4 <= __tmp_845_3;
      __tmp_845_5 <= __tmp_845_4;
      __tmp_845_6 <= __tmp_845_5;
      __tmp_845_7 <= __tmp_845_6;
      __tmp_845_8 <= __tmp_845_7;
      __tmp_845_9 <= __tmp_845_8;
      __tmp_845_10 <= __tmp_845_9;
      __tmp_845_11 <= __tmp_845_10;
      __tmp_845_12 <= __tmp_845_11;
      __tmp_847_1 <= _tmp_847;
      __tmp_847_2 <= __tmp_847_1;
      __tmp_847_3 <= __tmp_847_2;
      __tmp_847_4 <= __tmp_847_3;
      __tmp_847_5 <= __tmp_847_4;
      __tmp_847_6 <= __tmp_847_5;
      __tmp_847_7 <= __tmp_847_6;
      __tmp_847_8 <= __tmp_847_7;
      __tmp_847_9 <= __tmp_847_8;
      __tmp_847_10 <= __tmp_847_9;
      __tmp_847_11 <= __tmp_847_10;
      __tmp_847_12 <= __tmp_847_11;
      __tmp_849_1 <= _tmp_849;
      __tmp_849_2 <= __tmp_849_1;
      __tmp_849_3 <= __tmp_849_2;
      __tmp_849_4 <= __tmp_849_3;
      __tmp_849_5 <= __tmp_849_4;
      __tmp_849_6 <= __tmp_849_5;
      __tmp_849_7 <= __tmp_849_6;
      __tmp_849_8 <= __tmp_849_7;
      __tmp_849_9 <= __tmp_849_8;
      __tmp_849_10 <= __tmp_849_9;
      __tmp_849_11 <= __tmp_849_10;
      __tmp_849_12 <= __tmp_849_11;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_7_fsm <= _mul_7_fsm_init;
      _mul_7_source_busy <= 0;
      _substream_mul_7_x_data_cond_643_9 <= 0;
      _substream_mul_7_y_data_cond_643_10 <= 0;
      _substream_mul_7_rshift_data_cond_643_11 <= 0;
      _mul_7_sink_busy <= 0;
      _mul_7_sink_wait_count <= 0;
    end else begin
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_7_source_busy <= 1;
      end 
      if(__tmp_733_12) begin
        _substream_mul_7_x_data_cond_643_9 <= 1;
      end 
      if(__tmp_735_12) begin
        _substream_mul_7_y_data_cond_643_10 <= 1;
      end 
      if(__tmp_737_12) begin
        _substream_mul_7_rshift_data_cond_643_11 <= 1;
      end 
      if(_stream_conv2d_16_fsm == 3) begin
        _mul_7_source_busy <= 0;
      end 
      if(__tmp_839_9) begin
        _substream_mul_7_x_data_cond_643_9 <= 0;
      end 
      if(__tmp_841_9) begin
        _substream_mul_7_y_data_cond_643_10 <= 0;
      end 
      if(__tmp_843_9) begin
        _substream_mul_7_rshift_data_cond_643_11 <= 0;
      end 
      if((_mul_7_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_845_12) begin
        _mul_7_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_7_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_847_12) begin
        _mul_7_sink_wait_count <= _mul_7_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_849_12) begin
        _mul_7_sink_wait_count <= _mul_7_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_8_x_idle <= 1;
      _mul_8_x_source_ram_rvalid <= 0;
      _mul_8_y_idle <= 1;
      _mul_8_y_source_ram_rvalid <= 0;
      _mul_8_rshift_idle <= 1;
      _mul_8_rshift_source_ram_rvalid <= 0;
      _mul_8_z_sink_wenable <= 0;
      _greaterthan_data_125 <= 0;
      _minus_data_127 <= 0;
      __delay_data_662 <= 0;
      __delay_data_665 <= 0;
      __delay_data_668 <= 0;
      _sll_data_129 <= 0;
      __delay_data_661 <= 0;
      __delay_data_663 <= 0;
      __delay_data_666 <= 0;
      __delay_data_669 <= 0;
      _cond_data_135 <= 0;
      __delay_data_664 <= 0;
      __delay_data_667 <= 0;
      __delay_data_670 <= 0;
      __muladd_madd_odata_reg_137 <= 0;
      __delay_data_671 <= 0;
      __delay_data_672 <= 0;
      __delay_data_673 <= 0;
      __delay_data_674 <= 0;
      _sra_data_138 <= 0;
      __variable_wdata_122 <= 0;
      __variable_wdata_123 <= 0;
      __variable_wdata_124 <= 0;
      __tmp_857_1 <= 0;
      __tmp_857_2 <= 0;
      __tmp_857_3 <= 0;
      __tmp_857_4 <= 0;
      __tmp_857_5 <= 0;
      __tmp_857_6 <= 0;
      __tmp_857_7 <= 0;
      __tmp_857_8 <= 0;
      __tmp_857_9 <= 0;
      __tmp_857_10 <= 0;
      __tmp_857_11 <= 0;
      __tmp_857_12 <= 0;
      __tmp_859_1 <= 0;
      __tmp_859_2 <= 0;
      __tmp_859_3 <= 0;
      __tmp_859_4 <= 0;
      __tmp_859_5 <= 0;
      __tmp_859_6 <= 0;
      __tmp_859_7 <= 0;
      __tmp_859_8 <= 0;
      __tmp_859_9 <= 0;
      __tmp_859_10 <= 0;
      __tmp_859_11 <= 0;
      __tmp_859_12 <= 0;
      __tmp_861_1 <= 0;
      __tmp_861_2 <= 0;
      __tmp_861_3 <= 0;
      __tmp_861_4 <= 0;
      __tmp_861_5 <= 0;
      __tmp_861_6 <= 0;
      __tmp_861_7 <= 0;
      __tmp_861_8 <= 0;
      __tmp_861_9 <= 0;
      __tmp_861_10 <= 0;
      __tmp_861_11 <= 0;
      __tmp_861_12 <= 0;
    end else begin
      _mul_8_x_idle <= _mul_8_x_idle;
      _mul_8_x_source_ram_rvalid <= 0;
      _mul_8_y_idle <= _mul_8_y_idle;
      _mul_8_y_source_ram_rvalid <= 0;
      _mul_8_rshift_idle <= _mul_8_rshift_idle;
      _mul_8_rshift_source_ram_rvalid <= 0;
      _mul_8_z_sink_wenable <= 0;
      _greaterthan_data_125 <= mul_8_rshift_data > 1'sd0;
      _minus_data_127 <= mul_8_rshift_data - 2'sd1;
      __delay_data_662 <= mul_8_x_data;
      __delay_data_665 <= mul_8_y_data;
      __delay_data_668 <= mul_8_rshift_data;
      _sll_data_129 <= 2'sd1 << _minus_data_127;
      __delay_data_661 <= _greaterthan_data_125;
      __delay_data_663 <= __delay_data_662;
      __delay_data_666 <= __delay_data_665;
      __delay_data_669 <= __delay_data_668;
      _cond_data_135 <= (__delay_data_661)? _sll_data_129 : 1'sd0;
      __delay_data_664 <= __delay_data_663;
      __delay_data_667 <= __delay_data_666;
      __delay_data_670 <= __delay_data_669;
      __muladd_madd_odata_reg_137 <= __muladd_madd_odata_137;
      __delay_data_671 <= __delay_data_670;
      __delay_data_672 <= __delay_data_671;
      __delay_data_673 <= __delay_data_672;
      __delay_data_674 <= __delay_data_673;
      _sra_data_138 <= __muladd_data_137 >>> __delay_data_674;
      if(_substream_mul_8_x_data_cond_660_12) begin
        __variable_wdata_122 <= _cond_data_583;
      end 
      if(_substream_mul_8_y_data_cond_660_13) begin
        __variable_wdata_123 <= __delay_data_1124;
      end 
      if(_substream_mul_8_rshift_data_cond_660_14) begin
        __variable_wdata_124 <= __delay_data_1130;
      end 
      __tmp_857_1 <= _tmp_857;
      __tmp_857_2 <= __tmp_857_1;
      __tmp_857_3 <= __tmp_857_2;
      __tmp_857_4 <= __tmp_857_3;
      __tmp_857_5 <= __tmp_857_4;
      __tmp_857_6 <= __tmp_857_5;
      __tmp_857_7 <= __tmp_857_6;
      __tmp_857_8 <= __tmp_857_7;
      __tmp_857_9 <= __tmp_857_8;
      __tmp_857_10 <= __tmp_857_9;
      __tmp_857_11 <= __tmp_857_10;
      __tmp_857_12 <= __tmp_857_11;
      __tmp_859_1 <= _tmp_859;
      __tmp_859_2 <= __tmp_859_1;
      __tmp_859_3 <= __tmp_859_2;
      __tmp_859_4 <= __tmp_859_3;
      __tmp_859_5 <= __tmp_859_4;
      __tmp_859_6 <= __tmp_859_5;
      __tmp_859_7 <= __tmp_859_6;
      __tmp_859_8 <= __tmp_859_7;
      __tmp_859_9 <= __tmp_859_8;
      __tmp_859_10 <= __tmp_859_9;
      __tmp_859_11 <= __tmp_859_10;
      __tmp_859_12 <= __tmp_859_11;
      __tmp_861_1 <= _tmp_861;
      __tmp_861_2 <= __tmp_861_1;
      __tmp_861_3 <= __tmp_861_2;
      __tmp_861_4 <= __tmp_861_3;
      __tmp_861_5 <= __tmp_861_4;
      __tmp_861_6 <= __tmp_861_5;
      __tmp_861_7 <= __tmp_861_6;
      __tmp_861_8 <= __tmp_861_7;
      __tmp_861_9 <= __tmp_861_8;
      __tmp_861_10 <= __tmp_861_9;
      __tmp_861_11 <= __tmp_861_10;
      __tmp_861_12 <= __tmp_861_11;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_8_fsm <= _mul_8_fsm_init;
      _mul_8_source_busy <= 0;
      _substream_mul_8_x_data_cond_660_12 <= 0;
      _substream_mul_8_y_data_cond_660_13 <= 0;
      _substream_mul_8_rshift_data_cond_660_14 <= 0;
      _mul_8_sink_busy <= 0;
      _mul_8_sink_wait_count <= 0;
    end else begin
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_8_source_busy <= 1;
      end 
      if(__tmp_739_12) begin
        _substream_mul_8_x_data_cond_660_12 <= 1;
      end 
      if(__tmp_741_12) begin
        _substream_mul_8_y_data_cond_660_13 <= 1;
      end 
      if(__tmp_743_12) begin
        _substream_mul_8_rshift_data_cond_660_14 <= 1;
      end 
      if(_stream_conv2d_16_fsm == 3) begin
        _mul_8_source_busy <= 0;
      end 
      if(__tmp_851_9) begin
        _substream_mul_8_x_data_cond_660_12 <= 0;
      end 
      if(__tmp_853_9) begin
        _substream_mul_8_y_data_cond_660_13 <= 0;
      end 
      if(__tmp_855_9) begin
        _substream_mul_8_rshift_data_cond_660_14 <= 0;
      end 
      if((_mul_8_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_857_12) begin
        _mul_8_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_8_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_859_12) begin
        _mul_8_sink_wait_count <= _mul_8_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_861_12) begin
        _mul_8_sink_wait_count <= _mul_8_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_9_x_idle <= 1;
      _mul_9_x_source_ram_rvalid <= 0;
      _mul_9_y_idle <= 1;
      _mul_9_y_source_ram_rvalid <= 0;
      _mul_9_rshift_idle <= 1;
      _mul_9_rshift_source_ram_rvalid <= 0;
      _mul_9_z_sink_wenable <= 0;
      _greaterthan_data_142 <= 0;
      _minus_data_144 <= 0;
      __delay_data_679 <= 0;
      __delay_data_682 <= 0;
      __delay_data_685 <= 0;
      _sll_data_146 <= 0;
      __delay_data_678 <= 0;
      __delay_data_680 <= 0;
      __delay_data_683 <= 0;
      __delay_data_686 <= 0;
      _cond_data_152 <= 0;
      __delay_data_681 <= 0;
      __delay_data_684 <= 0;
      __delay_data_687 <= 0;
      __muladd_madd_odata_reg_154 <= 0;
      __delay_data_688 <= 0;
      __delay_data_689 <= 0;
      __delay_data_690 <= 0;
      __delay_data_691 <= 0;
      _sra_data_155 <= 0;
      __variable_wdata_139 <= 0;
      __variable_wdata_140 <= 0;
      __variable_wdata_141 <= 0;
      __tmp_869_1 <= 0;
      __tmp_869_2 <= 0;
      __tmp_869_3 <= 0;
      __tmp_869_4 <= 0;
      __tmp_869_5 <= 0;
      __tmp_869_6 <= 0;
      __tmp_869_7 <= 0;
      __tmp_869_8 <= 0;
      __tmp_869_9 <= 0;
      __tmp_869_10 <= 0;
      __tmp_869_11 <= 0;
      __tmp_869_12 <= 0;
      __tmp_871_1 <= 0;
      __tmp_871_2 <= 0;
      __tmp_871_3 <= 0;
      __tmp_871_4 <= 0;
      __tmp_871_5 <= 0;
      __tmp_871_6 <= 0;
      __tmp_871_7 <= 0;
      __tmp_871_8 <= 0;
      __tmp_871_9 <= 0;
      __tmp_871_10 <= 0;
      __tmp_871_11 <= 0;
      __tmp_871_12 <= 0;
      __tmp_873_1 <= 0;
      __tmp_873_2 <= 0;
      __tmp_873_3 <= 0;
      __tmp_873_4 <= 0;
      __tmp_873_5 <= 0;
      __tmp_873_6 <= 0;
      __tmp_873_7 <= 0;
      __tmp_873_8 <= 0;
      __tmp_873_9 <= 0;
      __tmp_873_10 <= 0;
      __tmp_873_11 <= 0;
      __tmp_873_12 <= 0;
    end else begin
      _mul_9_x_idle <= _mul_9_x_idle;
      _mul_9_x_source_ram_rvalid <= 0;
      _mul_9_y_idle <= _mul_9_y_idle;
      _mul_9_y_source_ram_rvalid <= 0;
      _mul_9_rshift_idle <= _mul_9_rshift_idle;
      _mul_9_rshift_source_ram_rvalid <= 0;
      _mul_9_z_sink_wenable <= 0;
      _greaterthan_data_142 <= mul_9_rshift_data > 1'sd0;
      _minus_data_144 <= mul_9_rshift_data - 2'sd1;
      __delay_data_679 <= mul_9_x_data;
      __delay_data_682 <= mul_9_y_data;
      __delay_data_685 <= mul_9_rshift_data;
      _sll_data_146 <= 2'sd1 << _minus_data_144;
      __delay_data_678 <= _greaterthan_data_142;
      __delay_data_680 <= __delay_data_679;
      __delay_data_683 <= __delay_data_682;
      __delay_data_686 <= __delay_data_685;
      _cond_data_152 <= (__delay_data_678)? _sll_data_146 : 1'sd0;
      __delay_data_681 <= __delay_data_680;
      __delay_data_684 <= __delay_data_683;
      __delay_data_687 <= __delay_data_686;
      __muladd_madd_odata_reg_154 <= __muladd_madd_odata_154;
      __delay_data_688 <= __delay_data_687;
      __delay_data_689 <= __delay_data_688;
      __delay_data_690 <= __delay_data_689;
      __delay_data_691 <= __delay_data_690;
      _sra_data_155 <= __muladd_data_154 >>> __delay_data_691;
      if(_substream_mul_9_x_data_cond_677_15) begin
        __variable_wdata_139 <= _cond_data_585;
      end 
      if(_substream_mul_9_y_data_cond_677_16) begin
        __variable_wdata_140 <= __delay_data_1159;
      end 
      if(_substream_mul_9_rshift_data_cond_677_17) begin
        __variable_wdata_141 <= __delay_data_1165;
      end 
      __tmp_869_1 <= _tmp_869;
      __tmp_869_2 <= __tmp_869_1;
      __tmp_869_3 <= __tmp_869_2;
      __tmp_869_4 <= __tmp_869_3;
      __tmp_869_5 <= __tmp_869_4;
      __tmp_869_6 <= __tmp_869_5;
      __tmp_869_7 <= __tmp_869_6;
      __tmp_869_8 <= __tmp_869_7;
      __tmp_869_9 <= __tmp_869_8;
      __tmp_869_10 <= __tmp_869_9;
      __tmp_869_11 <= __tmp_869_10;
      __tmp_869_12 <= __tmp_869_11;
      __tmp_871_1 <= _tmp_871;
      __tmp_871_2 <= __tmp_871_1;
      __tmp_871_3 <= __tmp_871_2;
      __tmp_871_4 <= __tmp_871_3;
      __tmp_871_5 <= __tmp_871_4;
      __tmp_871_6 <= __tmp_871_5;
      __tmp_871_7 <= __tmp_871_6;
      __tmp_871_8 <= __tmp_871_7;
      __tmp_871_9 <= __tmp_871_8;
      __tmp_871_10 <= __tmp_871_9;
      __tmp_871_11 <= __tmp_871_10;
      __tmp_871_12 <= __tmp_871_11;
      __tmp_873_1 <= _tmp_873;
      __tmp_873_2 <= __tmp_873_1;
      __tmp_873_3 <= __tmp_873_2;
      __tmp_873_4 <= __tmp_873_3;
      __tmp_873_5 <= __tmp_873_4;
      __tmp_873_6 <= __tmp_873_5;
      __tmp_873_7 <= __tmp_873_6;
      __tmp_873_8 <= __tmp_873_7;
      __tmp_873_9 <= __tmp_873_8;
      __tmp_873_10 <= __tmp_873_9;
      __tmp_873_11 <= __tmp_873_10;
      __tmp_873_12 <= __tmp_873_11;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_9_fsm <= _mul_9_fsm_init;
      _mul_9_source_busy <= 0;
      _substream_mul_9_x_data_cond_677_15 <= 0;
      _substream_mul_9_y_data_cond_677_16 <= 0;
      _substream_mul_9_rshift_data_cond_677_17 <= 0;
      _mul_9_sink_busy <= 0;
      _mul_9_sink_wait_count <= 0;
    end else begin
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_9_source_busy <= 1;
      end 
      if(__tmp_745_12) begin
        _substream_mul_9_x_data_cond_677_15 <= 1;
      end 
      if(__tmp_747_12) begin
        _substream_mul_9_y_data_cond_677_16 <= 1;
      end 
      if(__tmp_749_12) begin
        _substream_mul_9_rshift_data_cond_677_17 <= 1;
      end 
      if(_stream_conv2d_16_fsm == 3) begin
        _mul_9_source_busy <= 0;
      end 
      if(__tmp_863_9) begin
        _substream_mul_9_x_data_cond_677_15 <= 0;
      end 
      if(__tmp_865_9) begin
        _substream_mul_9_y_data_cond_677_16 <= 0;
      end 
      if(__tmp_867_9) begin
        _substream_mul_9_rshift_data_cond_677_17 <= 0;
      end 
      if((_mul_9_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_869_12) begin
        _mul_9_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_9_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_871_12) begin
        _mul_9_sink_wait_count <= _mul_9_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_873_12) begin
        _mul_9_sink_wait_count <= _mul_9_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_10_x_idle <= 1;
      _mul_10_x_source_ram_rvalid <= 0;
      _mul_10_y_idle <= 1;
      _mul_10_y_source_ram_rvalid <= 0;
      _mul_10_rshift_idle <= 1;
      _mul_10_rshift_source_ram_rvalid <= 0;
      _mul_10_z_sink_wenable <= 0;
      _greaterthan_data_159 <= 0;
      _minus_data_161 <= 0;
      __delay_data_696 <= 0;
      __delay_data_699 <= 0;
      __delay_data_702 <= 0;
      _sll_data_163 <= 0;
      __delay_data_695 <= 0;
      __delay_data_697 <= 0;
      __delay_data_700 <= 0;
      __delay_data_703 <= 0;
      _cond_data_169 <= 0;
      __delay_data_698 <= 0;
      __delay_data_701 <= 0;
      __delay_data_704 <= 0;
      __muladd_madd_odata_reg_171 <= 0;
      __delay_data_705 <= 0;
      __delay_data_706 <= 0;
      __delay_data_707 <= 0;
      __delay_data_708 <= 0;
      _sra_data_172 <= 0;
      __variable_wdata_156 <= 0;
      __variable_wdata_157 <= 0;
      __variable_wdata_158 <= 0;
      __tmp_881_1 <= 0;
      __tmp_881_2 <= 0;
      __tmp_881_3 <= 0;
      __tmp_881_4 <= 0;
      __tmp_881_5 <= 0;
      __tmp_881_6 <= 0;
      __tmp_881_7 <= 0;
      __tmp_881_8 <= 0;
      __tmp_881_9 <= 0;
      __tmp_881_10 <= 0;
      __tmp_881_11 <= 0;
      __tmp_881_12 <= 0;
      __tmp_883_1 <= 0;
      __tmp_883_2 <= 0;
      __tmp_883_3 <= 0;
      __tmp_883_4 <= 0;
      __tmp_883_5 <= 0;
      __tmp_883_6 <= 0;
      __tmp_883_7 <= 0;
      __tmp_883_8 <= 0;
      __tmp_883_9 <= 0;
      __tmp_883_10 <= 0;
      __tmp_883_11 <= 0;
      __tmp_883_12 <= 0;
      __tmp_885_1 <= 0;
      __tmp_885_2 <= 0;
      __tmp_885_3 <= 0;
      __tmp_885_4 <= 0;
      __tmp_885_5 <= 0;
      __tmp_885_6 <= 0;
      __tmp_885_7 <= 0;
      __tmp_885_8 <= 0;
      __tmp_885_9 <= 0;
      __tmp_885_10 <= 0;
      __tmp_885_11 <= 0;
      __tmp_885_12 <= 0;
    end else begin
      _mul_10_x_idle <= _mul_10_x_idle;
      _mul_10_x_source_ram_rvalid <= 0;
      _mul_10_y_idle <= _mul_10_y_idle;
      _mul_10_y_source_ram_rvalid <= 0;
      _mul_10_rshift_idle <= _mul_10_rshift_idle;
      _mul_10_rshift_source_ram_rvalid <= 0;
      _mul_10_z_sink_wenable <= 0;
      _greaterthan_data_159 <= mul_10_rshift_data > 1'sd0;
      _minus_data_161 <= mul_10_rshift_data - 2'sd1;
      __delay_data_696 <= mul_10_x_data;
      __delay_data_699 <= mul_10_y_data;
      __delay_data_702 <= mul_10_rshift_data;
      _sll_data_163 <= 2'sd1 << _minus_data_161;
      __delay_data_695 <= _greaterthan_data_159;
      __delay_data_697 <= __delay_data_696;
      __delay_data_700 <= __delay_data_699;
      __delay_data_703 <= __delay_data_702;
      _cond_data_169 <= (__delay_data_695)? _sll_data_163 : 1'sd0;
      __delay_data_698 <= __delay_data_697;
      __delay_data_701 <= __delay_data_700;
      __delay_data_704 <= __delay_data_703;
      __muladd_madd_odata_reg_171 <= __muladd_madd_odata_171;
      __delay_data_705 <= __delay_data_704;
      __delay_data_706 <= __delay_data_705;
      __delay_data_707 <= __delay_data_706;
      __delay_data_708 <= __delay_data_707;
      _sra_data_172 <= __muladd_data_171 >>> __delay_data_708;
      if(_substream_mul_10_x_data_cond_694_18) begin
        __variable_wdata_156 <= _cond_data_587;
      end 
      if(_substream_mul_10_y_data_cond_694_19) begin
        __variable_wdata_157 <= __delay_data_1193;
      end 
      if(_substream_mul_10_rshift_data_cond_694_20) begin
        __variable_wdata_158 <= __delay_data_1199;
      end 
      __tmp_881_1 <= _tmp_881;
      __tmp_881_2 <= __tmp_881_1;
      __tmp_881_3 <= __tmp_881_2;
      __tmp_881_4 <= __tmp_881_3;
      __tmp_881_5 <= __tmp_881_4;
      __tmp_881_6 <= __tmp_881_5;
      __tmp_881_7 <= __tmp_881_6;
      __tmp_881_8 <= __tmp_881_7;
      __tmp_881_9 <= __tmp_881_8;
      __tmp_881_10 <= __tmp_881_9;
      __tmp_881_11 <= __tmp_881_10;
      __tmp_881_12 <= __tmp_881_11;
      __tmp_883_1 <= _tmp_883;
      __tmp_883_2 <= __tmp_883_1;
      __tmp_883_3 <= __tmp_883_2;
      __tmp_883_4 <= __tmp_883_3;
      __tmp_883_5 <= __tmp_883_4;
      __tmp_883_6 <= __tmp_883_5;
      __tmp_883_7 <= __tmp_883_6;
      __tmp_883_8 <= __tmp_883_7;
      __tmp_883_9 <= __tmp_883_8;
      __tmp_883_10 <= __tmp_883_9;
      __tmp_883_11 <= __tmp_883_10;
      __tmp_883_12 <= __tmp_883_11;
      __tmp_885_1 <= _tmp_885;
      __tmp_885_2 <= __tmp_885_1;
      __tmp_885_3 <= __tmp_885_2;
      __tmp_885_4 <= __tmp_885_3;
      __tmp_885_5 <= __tmp_885_4;
      __tmp_885_6 <= __tmp_885_5;
      __tmp_885_7 <= __tmp_885_6;
      __tmp_885_8 <= __tmp_885_7;
      __tmp_885_9 <= __tmp_885_8;
      __tmp_885_10 <= __tmp_885_9;
      __tmp_885_11 <= __tmp_885_10;
      __tmp_885_12 <= __tmp_885_11;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_10_fsm <= _mul_10_fsm_init;
      _mul_10_source_busy <= 0;
      _substream_mul_10_x_data_cond_694_18 <= 0;
      _substream_mul_10_y_data_cond_694_19 <= 0;
      _substream_mul_10_rshift_data_cond_694_20 <= 0;
      _mul_10_sink_busy <= 0;
      _mul_10_sink_wait_count <= 0;
    end else begin
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_10_source_busy <= 1;
      end 
      if(__tmp_751_12) begin
        _substream_mul_10_x_data_cond_694_18 <= 1;
      end 
      if(__tmp_753_12) begin
        _substream_mul_10_y_data_cond_694_19 <= 1;
      end 
      if(__tmp_755_12) begin
        _substream_mul_10_rshift_data_cond_694_20 <= 1;
      end 
      if(_stream_conv2d_16_fsm == 3) begin
        _mul_10_source_busy <= 0;
      end 
      if(__tmp_875_9) begin
        _substream_mul_10_x_data_cond_694_18 <= 0;
      end 
      if(__tmp_877_9) begin
        _substream_mul_10_y_data_cond_694_19 <= 0;
      end 
      if(__tmp_879_9) begin
        _substream_mul_10_rshift_data_cond_694_20 <= 0;
      end 
      if((_mul_10_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_881_12) begin
        _mul_10_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_10_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_883_12) begin
        _mul_10_sink_wait_count <= _mul_10_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_885_12) begin
        _mul_10_sink_wait_count <= _mul_10_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_11_x_idle <= 1;
      _mul_11_x_source_ram_rvalid <= 0;
      _mul_11_y_idle <= 1;
      _mul_11_y_source_ram_rvalid <= 0;
      _mul_11_rshift_idle <= 1;
      _mul_11_rshift_source_ram_rvalid <= 0;
      _mul_11_z_sink_wenable <= 0;
      _greaterthan_data_176 <= 0;
      _minus_data_178 <= 0;
      __delay_data_713 <= 0;
      __delay_data_716 <= 0;
      __delay_data_719 <= 0;
      _sll_data_180 <= 0;
      __delay_data_712 <= 0;
      __delay_data_714 <= 0;
      __delay_data_717 <= 0;
      __delay_data_720 <= 0;
      _cond_data_186 <= 0;
      __delay_data_715 <= 0;
      __delay_data_718 <= 0;
      __delay_data_721 <= 0;
      __muladd_madd_odata_reg_188 <= 0;
      __delay_data_722 <= 0;
      __delay_data_723 <= 0;
      __delay_data_724 <= 0;
      __delay_data_725 <= 0;
      _sra_data_189 <= 0;
      __variable_wdata_173 <= 0;
      __variable_wdata_174 <= 0;
      __variable_wdata_175 <= 0;
      __tmp_893_1 <= 0;
      __tmp_893_2 <= 0;
      __tmp_893_3 <= 0;
      __tmp_893_4 <= 0;
      __tmp_893_5 <= 0;
      __tmp_893_6 <= 0;
      __tmp_893_7 <= 0;
      __tmp_893_8 <= 0;
      __tmp_893_9 <= 0;
      __tmp_893_10 <= 0;
      __tmp_893_11 <= 0;
      __tmp_893_12 <= 0;
      __tmp_895_1 <= 0;
      __tmp_895_2 <= 0;
      __tmp_895_3 <= 0;
      __tmp_895_4 <= 0;
      __tmp_895_5 <= 0;
      __tmp_895_6 <= 0;
      __tmp_895_7 <= 0;
      __tmp_895_8 <= 0;
      __tmp_895_9 <= 0;
      __tmp_895_10 <= 0;
      __tmp_895_11 <= 0;
      __tmp_895_12 <= 0;
      __tmp_897_1 <= 0;
      __tmp_897_2 <= 0;
      __tmp_897_3 <= 0;
      __tmp_897_4 <= 0;
      __tmp_897_5 <= 0;
      __tmp_897_6 <= 0;
      __tmp_897_7 <= 0;
      __tmp_897_8 <= 0;
      __tmp_897_9 <= 0;
      __tmp_897_10 <= 0;
      __tmp_897_11 <= 0;
      __tmp_897_12 <= 0;
    end else begin
      _mul_11_x_idle <= _mul_11_x_idle;
      _mul_11_x_source_ram_rvalid <= 0;
      _mul_11_y_idle <= _mul_11_y_idle;
      _mul_11_y_source_ram_rvalid <= 0;
      _mul_11_rshift_idle <= _mul_11_rshift_idle;
      _mul_11_rshift_source_ram_rvalid <= 0;
      _mul_11_z_sink_wenable <= 0;
      _greaterthan_data_176 <= mul_11_rshift_data > 1'sd0;
      _minus_data_178 <= mul_11_rshift_data - 2'sd1;
      __delay_data_713 <= mul_11_x_data;
      __delay_data_716 <= mul_11_y_data;
      __delay_data_719 <= mul_11_rshift_data;
      _sll_data_180 <= 2'sd1 << _minus_data_178;
      __delay_data_712 <= _greaterthan_data_176;
      __delay_data_714 <= __delay_data_713;
      __delay_data_717 <= __delay_data_716;
      __delay_data_720 <= __delay_data_719;
      _cond_data_186 <= (__delay_data_712)? _sll_data_180 : 1'sd0;
      __delay_data_715 <= __delay_data_714;
      __delay_data_718 <= __delay_data_717;
      __delay_data_721 <= __delay_data_720;
      __muladd_madd_odata_reg_188 <= __muladd_madd_odata_188;
      __delay_data_722 <= __delay_data_721;
      __delay_data_723 <= __delay_data_722;
      __delay_data_724 <= __delay_data_723;
      __delay_data_725 <= __delay_data_724;
      _sra_data_189 <= __muladd_data_188 >>> __delay_data_725;
      if(_substream_mul_11_x_data_cond_711_21) begin
        __variable_wdata_173 <= _cond_data_589;
      end 
      if(_substream_mul_11_y_data_cond_711_22) begin
        __variable_wdata_174 <= __delay_data_1227;
      end 
      if(_substream_mul_11_rshift_data_cond_711_23) begin
        __variable_wdata_175 <= __delay_data_1233;
      end 
      __tmp_893_1 <= _tmp_893;
      __tmp_893_2 <= __tmp_893_1;
      __tmp_893_3 <= __tmp_893_2;
      __tmp_893_4 <= __tmp_893_3;
      __tmp_893_5 <= __tmp_893_4;
      __tmp_893_6 <= __tmp_893_5;
      __tmp_893_7 <= __tmp_893_6;
      __tmp_893_8 <= __tmp_893_7;
      __tmp_893_9 <= __tmp_893_8;
      __tmp_893_10 <= __tmp_893_9;
      __tmp_893_11 <= __tmp_893_10;
      __tmp_893_12 <= __tmp_893_11;
      __tmp_895_1 <= _tmp_895;
      __tmp_895_2 <= __tmp_895_1;
      __tmp_895_3 <= __tmp_895_2;
      __tmp_895_4 <= __tmp_895_3;
      __tmp_895_5 <= __tmp_895_4;
      __tmp_895_6 <= __tmp_895_5;
      __tmp_895_7 <= __tmp_895_6;
      __tmp_895_8 <= __tmp_895_7;
      __tmp_895_9 <= __tmp_895_8;
      __tmp_895_10 <= __tmp_895_9;
      __tmp_895_11 <= __tmp_895_10;
      __tmp_895_12 <= __tmp_895_11;
      __tmp_897_1 <= _tmp_897;
      __tmp_897_2 <= __tmp_897_1;
      __tmp_897_3 <= __tmp_897_2;
      __tmp_897_4 <= __tmp_897_3;
      __tmp_897_5 <= __tmp_897_4;
      __tmp_897_6 <= __tmp_897_5;
      __tmp_897_7 <= __tmp_897_6;
      __tmp_897_8 <= __tmp_897_7;
      __tmp_897_9 <= __tmp_897_8;
      __tmp_897_10 <= __tmp_897_9;
      __tmp_897_11 <= __tmp_897_10;
      __tmp_897_12 <= __tmp_897_11;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_11_fsm <= _mul_11_fsm_init;
      _mul_11_source_busy <= 0;
      _substream_mul_11_x_data_cond_711_21 <= 0;
      _substream_mul_11_y_data_cond_711_22 <= 0;
      _substream_mul_11_rshift_data_cond_711_23 <= 0;
      _mul_11_sink_busy <= 0;
      _mul_11_sink_wait_count <= 0;
    end else begin
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_11_source_busy <= 1;
      end 
      if(__tmp_757_12) begin
        _substream_mul_11_x_data_cond_711_21 <= 1;
      end 
      if(__tmp_759_12) begin
        _substream_mul_11_y_data_cond_711_22 <= 1;
      end 
      if(__tmp_761_12) begin
        _substream_mul_11_rshift_data_cond_711_23 <= 1;
      end 
      if(_stream_conv2d_16_fsm == 3) begin
        _mul_11_source_busy <= 0;
      end 
      if(__tmp_887_9) begin
        _substream_mul_11_x_data_cond_711_21 <= 0;
      end 
      if(__tmp_889_9) begin
        _substream_mul_11_y_data_cond_711_22 <= 0;
      end 
      if(__tmp_891_9) begin
        _substream_mul_11_rshift_data_cond_711_23 <= 0;
      end 
      if((_mul_11_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_893_12) begin
        _mul_11_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_11_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_895_12) begin
        _mul_11_sink_wait_count <= _mul_11_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_897_12) begin
        _mul_11_sink_wait_count <= _mul_11_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_12_x_idle <= 1;
      _mul_12_x_source_ram_rvalid <= 0;
      _mul_12_y_idle <= 1;
      _mul_12_y_source_ram_rvalid <= 0;
      _mul_12_rshift_idle <= 1;
      _mul_12_rshift_source_ram_rvalid <= 0;
      _mul_12_z_sink_wenable <= 0;
      _greaterthan_data_193 <= 0;
      _minus_data_195 <= 0;
      __delay_data_730 <= 0;
      __delay_data_733 <= 0;
      __delay_data_736 <= 0;
      _sll_data_197 <= 0;
      __delay_data_729 <= 0;
      __delay_data_731 <= 0;
      __delay_data_734 <= 0;
      __delay_data_737 <= 0;
      _cond_data_203 <= 0;
      __delay_data_732 <= 0;
      __delay_data_735 <= 0;
      __delay_data_738 <= 0;
      __muladd_madd_odata_reg_205 <= 0;
      __delay_data_739 <= 0;
      __delay_data_740 <= 0;
      __delay_data_741 <= 0;
      __delay_data_742 <= 0;
      _sra_data_206 <= 0;
      __variable_wdata_190 <= 0;
      __variable_wdata_191 <= 0;
      __variable_wdata_192 <= 0;
      __tmp_905_1 <= 0;
      __tmp_905_2 <= 0;
      __tmp_905_3 <= 0;
      __tmp_905_4 <= 0;
      __tmp_905_5 <= 0;
      __tmp_905_6 <= 0;
      __tmp_905_7 <= 0;
      __tmp_905_8 <= 0;
      __tmp_905_9 <= 0;
      __tmp_905_10 <= 0;
      __tmp_905_11 <= 0;
      __tmp_905_12 <= 0;
      __tmp_907_1 <= 0;
      __tmp_907_2 <= 0;
      __tmp_907_3 <= 0;
      __tmp_907_4 <= 0;
      __tmp_907_5 <= 0;
      __tmp_907_6 <= 0;
      __tmp_907_7 <= 0;
      __tmp_907_8 <= 0;
      __tmp_907_9 <= 0;
      __tmp_907_10 <= 0;
      __tmp_907_11 <= 0;
      __tmp_907_12 <= 0;
      __tmp_909_1 <= 0;
      __tmp_909_2 <= 0;
      __tmp_909_3 <= 0;
      __tmp_909_4 <= 0;
      __tmp_909_5 <= 0;
      __tmp_909_6 <= 0;
      __tmp_909_7 <= 0;
      __tmp_909_8 <= 0;
      __tmp_909_9 <= 0;
      __tmp_909_10 <= 0;
      __tmp_909_11 <= 0;
      __tmp_909_12 <= 0;
    end else begin
      _mul_12_x_idle <= _mul_12_x_idle;
      _mul_12_x_source_ram_rvalid <= 0;
      _mul_12_y_idle <= _mul_12_y_idle;
      _mul_12_y_source_ram_rvalid <= 0;
      _mul_12_rshift_idle <= _mul_12_rshift_idle;
      _mul_12_rshift_source_ram_rvalid <= 0;
      _mul_12_z_sink_wenable <= 0;
      _greaterthan_data_193 <= mul_12_rshift_data > 1'sd0;
      _minus_data_195 <= mul_12_rshift_data - 2'sd1;
      __delay_data_730 <= mul_12_x_data;
      __delay_data_733 <= mul_12_y_data;
      __delay_data_736 <= mul_12_rshift_data;
      _sll_data_197 <= 2'sd1 << _minus_data_195;
      __delay_data_729 <= _greaterthan_data_193;
      __delay_data_731 <= __delay_data_730;
      __delay_data_734 <= __delay_data_733;
      __delay_data_737 <= __delay_data_736;
      _cond_data_203 <= (__delay_data_729)? _sll_data_197 : 1'sd0;
      __delay_data_732 <= __delay_data_731;
      __delay_data_735 <= __delay_data_734;
      __delay_data_738 <= __delay_data_737;
      __muladd_madd_odata_reg_205 <= __muladd_madd_odata_205;
      __delay_data_739 <= __delay_data_738;
      __delay_data_740 <= __delay_data_739;
      __delay_data_741 <= __delay_data_740;
      __delay_data_742 <= __delay_data_741;
      _sra_data_206 <= __muladd_data_205 >>> __delay_data_742;
      if(_substream_mul_12_x_data_cond_728_24) begin
        __variable_wdata_190 <= _cond_data_591;
      end 
      if(_substream_mul_12_y_data_cond_728_25) begin
        __variable_wdata_191 <= __delay_data_1261;
      end 
      if(_substream_mul_12_rshift_data_cond_728_26) begin
        __variable_wdata_192 <= __delay_data_1267;
      end 
      __tmp_905_1 <= _tmp_905;
      __tmp_905_2 <= __tmp_905_1;
      __tmp_905_3 <= __tmp_905_2;
      __tmp_905_4 <= __tmp_905_3;
      __tmp_905_5 <= __tmp_905_4;
      __tmp_905_6 <= __tmp_905_5;
      __tmp_905_7 <= __tmp_905_6;
      __tmp_905_8 <= __tmp_905_7;
      __tmp_905_9 <= __tmp_905_8;
      __tmp_905_10 <= __tmp_905_9;
      __tmp_905_11 <= __tmp_905_10;
      __tmp_905_12 <= __tmp_905_11;
      __tmp_907_1 <= _tmp_907;
      __tmp_907_2 <= __tmp_907_1;
      __tmp_907_3 <= __tmp_907_2;
      __tmp_907_4 <= __tmp_907_3;
      __tmp_907_5 <= __tmp_907_4;
      __tmp_907_6 <= __tmp_907_5;
      __tmp_907_7 <= __tmp_907_6;
      __tmp_907_8 <= __tmp_907_7;
      __tmp_907_9 <= __tmp_907_8;
      __tmp_907_10 <= __tmp_907_9;
      __tmp_907_11 <= __tmp_907_10;
      __tmp_907_12 <= __tmp_907_11;
      __tmp_909_1 <= _tmp_909;
      __tmp_909_2 <= __tmp_909_1;
      __tmp_909_3 <= __tmp_909_2;
      __tmp_909_4 <= __tmp_909_3;
      __tmp_909_5 <= __tmp_909_4;
      __tmp_909_6 <= __tmp_909_5;
      __tmp_909_7 <= __tmp_909_6;
      __tmp_909_8 <= __tmp_909_7;
      __tmp_909_9 <= __tmp_909_8;
      __tmp_909_10 <= __tmp_909_9;
      __tmp_909_11 <= __tmp_909_10;
      __tmp_909_12 <= __tmp_909_11;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_12_fsm <= _mul_12_fsm_init;
      _mul_12_source_busy <= 0;
      _substream_mul_12_x_data_cond_728_24 <= 0;
      _substream_mul_12_y_data_cond_728_25 <= 0;
      _substream_mul_12_rshift_data_cond_728_26 <= 0;
      _mul_12_sink_busy <= 0;
      _mul_12_sink_wait_count <= 0;
    end else begin
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_12_source_busy <= 1;
      end 
      if(__tmp_763_12) begin
        _substream_mul_12_x_data_cond_728_24 <= 1;
      end 
      if(__tmp_765_12) begin
        _substream_mul_12_y_data_cond_728_25 <= 1;
      end 
      if(__tmp_767_12) begin
        _substream_mul_12_rshift_data_cond_728_26 <= 1;
      end 
      if(_stream_conv2d_16_fsm == 3) begin
        _mul_12_source_busy <= 0;
      end 
      if(__tmp_899_9) begin
        _substream_mul_12_x_data_cond_728_24 <= 0;
      end 
      if(__tmp_901_9) begin
        _substream_mul_12_y_data_cond_728_25 <= 0;
      end 
      if(__tmp_903_9) begin
        _substream_mul_12_rshift_data_cond_728_26 <= 0;
      end 
      if((_mul_12_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_905_12) begin
        _mul_12_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _mul_12_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_907_12) begin
        _mul_12_sink_wait_count <= _mul_12_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_909_12) begin
        _mul_12_sink_wait_count <= _mul_12_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_13_x_idle <= 1;
      __reduce_max_13_x_source_ram_rvalid <= 0;
      __reduce_max_13_data_sink_wenable <= 0;
      __reduce_max_13_valid_sink_wenable <= 0;
      _reducemax_data_211 <= -9'sd128;
      _reducemax_count_211 <= 0;
      _pulse_data_213 <= 1'sd0;
      _pulse_count_213 <= 0;
      __variable_wdata_207 <= 0;
      __variable_wdata_208 <= 0;
      __tmp_1056_1 <= 0;
      __tmp_1056_2 <= 0;
      __tmp_1056_3 <= 0;
      __tmp_1056_4 <= 0;
      __tmp_1056_5 <= 0;
      __tmp_1058_1 <= 0;
      __tmp_1058_2 <= 0;
      __tmp_1058_3 <= 0;
      __tmp_1058_4 <= 0;
      __tmp_1058_5 <= 0;
      __tmp_1060_1 <= 0;
      __tmp_1060_2 <= 0;
      __tmp_1060_3 <= 0;
      __tmp_1060_4 <= 0;
      __tmp_1060_5 <= 0;
    end else begin
      __reduce_max_13_x_idle <= __reduce_max_13_x_idle;
      __reduce_max_13_x_source_ram_rvalid <= 0;
      __reduce_max_13_data_sink_wenable <= 0;
      __reduce_max_13_valid_sink_wenable <= 0;
      _reducemax_data_211 <= (_reducemax_data_211 < _reduce_max_13_x_data)? _reduce_max_13_x_data : _reducemax_data_211;
      _reducemax_count_211 <= (_reducemax_count_211 >= _reduce_max_13_size_data - 1)? 0 : _reducemax_count_211 + 1;
      if(__reduce_max_13_reduce_reset) begin
        _reducemax_data_211 <= (-9'sd128 < _reduce_max_13_x_data)? _reduce_max_13_x_data : -9'sd128;
      end 
      if(__reduce_max_13_reduce_reset) begin
        _reducemax_count_211 <= 0;
      end 
      if(_reducemax_count_211 == 0) begin
        _reducemax_data_211 <= (-9'sd128 < _reduce_max_13_x_data)? _reduce_max_13_x_data : -9'sd128;
      end 
      _pulse_data_213 <= _pulse_count_213 >= _reduce_max_13_size_data - 1;
      _pulse_count_213 <= (_pulse_count_213 >= _reduce_max_13_size_data - 1)? 0 : _pulse_count_213 + 1;
      if(__reduce_max_13_reduce_reset) begin
        _pulse_data_213 <= _pulse_count_213 >= _reduce_max_13_size_data - 1;
      end 
      if(__reduce_max_13_reduce_reset) begin
        _pulse_count_213 <= 0;
      end 
      if(_pulse_count_213 == 0) begin
        _pulse_data_213 <= _pulse_count_213 >= _reduce_max_13_size_data - 1;
      end 
      if(_substream__reduce_max_13_x_data_cond_792_42) begin
        __variable_wdata_207 <= _cond_data_791;
      end 
      if(_substream__reduce_max_13_size_data_cond_792_43) begin
        __variable_wdata_208 <= __delay_data_1416;
      end 
      __tmp_1056_1 <= _tmp_1056;
      __tmp_1056_2 <= __tmp_1056_1;
      __tmp_1056_3 <= __tmp_1056_2;
      __tmp_1056_4 <= __tmp_1056_3;
      __tmp_1056_5 <= __tmp_1056_4;
      __tmp_1058_1 <= _tmp_1058;
      __tmp_1058_2 <= __tmp_1058_1;
      __tmp_1058_3 <= __tmp_1058_2;
      __tmp_1058_4 <= __tmp_1058_3;
      __tmp_1058_5 <= __tmp_1058_4;
      __tmp_1060_1 <= _tmp_1060;
      __tmp_1060_2 <= __tmp_1060_1;
      __tmp_1060_3 <= __tmp_1060_2;
      __tmp_1060_4 <= __tmp_1060_3;
      __tmp_1060_5 <= __tmp_1060_4;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_13_fsm <= __reduce_max_13_fsm_init;
      __reduce_max_13_source_busy <= 0;
      __reduce_max_13_reduce_reset <= 1;
      _substream__reduce_max_13_x_data_cond_792_42 <= 0;
      _substream__reduce_max_13_size_data_cond_792_43 <= 0;
      __reduce_max_13_sink_busy <= 0;
      __reduce_max_13_sink_wait_count <= 0;
    end else begin
      if((_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag) begin
        __reduce_max_13_source_busy <= 1;
      end 
      if(__tmp_1042_9) begin
        __reduce_max_13_reduce_reset <= 0;
      end 
      if(__tmp_1044_7) begin
        _substream__reduce_max_13_x_data_cond_792_42 <= 1;
      end 
      if(__tmp_1046_7) begin
        _substream__reduce_max_13_size_data_cond_792_43 <= 1;
      end 
      if(_stream_max_pool_serial_18_fsm == 3) begin
        __reduce_max_13_source_busy <= 0;
      end 
      if(__tmp_1050_5) begin
        __reduce_max_13_reduce_reset <= 1;
      end 
      if(__tmp_1052_4) begin
        _substream__reduce_max_13_x_data_cond_792_42 <= 0;
      end 
      if(__tmp_1054_4) begin
        _substream__reduce_max_13_size_data_cond_792_43 <= 0;
      end 
      if((__reduce_max_13_sink_wait_count == 1) && !((_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag) && __tmp_1056_5) begin
        __reduce_max_13_sink_busy <= 0;
      end 
      if((_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag) begin
        __reduce_max_13_sink_busy <= 1;
      end 
      if(!((_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag) && __tmp_1058_5) begin
        __reduce_max_13_sink_wait_count <= __reduce_max_13_sink_wait_count - 1;
      end 
      if((_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag && !__tmp_1060_5) begin
        __reduce_max_13_sink_wait_count <= __reduce_max_13_sink_wait_count + 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_6_idle <= 1;
      _stream_conv2d_16_source_6_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_8_idle <= 1;
      _stream_conv2d_16_source_8_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_10_idle <= 1;
      _stream_conv2d_16_source_10_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_12_idle <= 1;
      _stream_conv2d_16_source_12_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_14_idle <= 1;
      _stream_conv2d_16_source_14_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_19_idle <= 1;
      _stream_conv2d_16_source_19_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_20_idle <= 1;
      _stream_conv2d_16_source_20_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_21_idle <= 1;
      _stream_conv2d_16_source_21_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_22_idle <= 1;
      _stream_conv2d_16_source_22_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_23_idle <= 1;
      _stream_conv2d_16_source_23_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_24_idle <= 1;
      _stream_conv2d_16_source_24_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_25_idle <= 1;
      _stream_conv2d_16_source_25_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_26_idle <= 1;
      _stream_conv2d_16_source_26_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_27_idle <= 1;
      _stream_conv2d_16_source_27_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_28_idle <= 1;
      _stream_conv2d_16_source_28_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_29_idle <= 1;
      _stream_conv2d_16_source_29_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_30_idle <= 1;
      _stream_conv2d_16_source_30_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_31_idle <= 1;
      _stream_conv2d_16_source_31_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_32_idle <= 1;
      _stream_conv2d_16_source_32_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_33_idle <= 1;
      _stream_conv2d_16_source_33_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_34_idle <= 1;
      _stream_conv2d_16_source_34_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_35_idle <= 1;
      _stream_conv2d_16_source_35_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_36_idle <= 1;
      _stream_conv2d_16_source_36_source_ram_rvalid <= 0;
      _stream_conv2d_16_sink_37_sink_wenable <= 0;
      _stream_conv2d_16_sink_38_sink_wenable <= 0;
      _cond_data_235 <= 0;
      _cond_data_242 <= 0;
      _cond_data_249 <= 0;
      _cond_data_256 <= 0;
      _cond_data_263 <= 0;
      _eq_data_277 <= 0;
      _eq_data_281 <= 0;
      _eq_data_284 <= 0;
      _eq_data_287 <= 0;
      _eq_data_291 <= 0;
      _eq_data_294 <= 0;
      _eq_data_297 <= 0;
      _eq_data_301 <= 0;
      _eq_data_304 <= 0;
      _eq_data_307 <= 0;
      _eq_data_311 <= 0;
      _eq_data_314 <= 0;
      _eq_data_317 <= 0;
      _eq_data_321 <= 0;
      _eq_data_324 <= 0;
      _eq_data_327 <= 0;
      _eq_data_331 <= 0;
      _eq_data_334 <= 0;
      _eq_data_337 <= 0;
      _eq_data_341 <= 0;
      _eq_data_344 <= 0;
      _eq_data_347 <= 0;
      _eq_data_351 <= 0;
      _eq_data_354 <= 0;
      _eq_data_357 <= 0;
      _eq_data_361 <= 0;
      _eq_data_364 <= 0;
      _eq_data_367 <= 0;
      _eq_data_371 <= 0;
      _eq_data_374 <= 0;
      _eq_data_377 <= 0;
      _eq_data_381 <= 0;
      _eq_data_384 <= 0;
      _eq_data_387 <= 0;
      _eq_data_391 <= 0;
      _eq_data_394 <= 0;
      _eq_data_397 <= 0;
      _eq_data_401 <= 0;
      _eq_data_404 <= 0;
      _eq_data_407 <= 0;
      _eq_data_411 <= 0;
      _eq_data_414 <= 0;
      _eq_data_417 <= 0;
      _eq_data_421 <= 0;
      _eq_data_424 <= 0;
      _eq_data_427 <= 0;
      _eq_data_431 <= 0;
      _eq_data_434 <= 0;
      _eq_data_437 <= 0;
      _eq_data_441 <= 0;
      _eq_data_444 <= 0;
      _eq_data_447 <= 0;
      _eq_data_451 <= 0;
      _eq_data_454 <= 0;
      __delay_data_898 <= 0;
      __delay_data_900 <= 0;
      __delay_data_904 <= 0;
      __delay_data_907 <= 0;
      __delay_data_909 <= 0;
      __delay_data_913 <= 0;
      __delay_data_916 <= 0;
      __delay_data_918 <= 0;
      __delay_data_922 <= 0;
      __delay_data_940 <= 0;
      __delay_data_947 <= 0;
      __delay_data_948 <= 0;
      __delay_data_992 <= 0;
      __delay_data_999 <= 0;
      __delay_data_1040 <= 0;
      __delay_data_1047 <= 0;
      __delay_data_1075 <= 0;
      __delay_data_1082 <= 0;
      __delay_data_1110 <= 0;
      __delay_data_1117 <= 0;
      __delay_data_1145 <= 0;
      __delay_data_1152 <= 0;
      __delay_data_1179 <= 0;
      __delay_data_1186 <= 0;
      __delay_data_1213 <= 0;
      __delay_data_1220 <= 0;
      __delay_data_1247 <= 0;
      __delay_data_1254 <= 0;
      __delay_data_1268 <= 0;
      __delay_data_1289 <= 0;
      __delay_data_1339 <= 0;
      _cond_data_279 <= 0;
      _cond_data_289 <= 0;
      _cond_data_299 <= 0;
      _cond_data_309 <= 0;
      _cond_data_319 <= 0;
      _cond_data_329 <= 0;
      _cond_data_339 <= 0;
      _cond_data_349 <= 0;
      _cond_data_359 <= 0;
      _plus_data_607 <= 0;
      _plus_data_624 <= 0;
      _plus_data_641 <= 0;
      _plus_data_658 <= 0;
      _plus_data_675 <= 0;
      _plus_data_692 <= 0;
      _plus_data_709 <= 0;
      _plus_data_726 <= 0;
      _plus_data_743 <= 0;
      _plus_data_759 <= 0;
      _plus_data_770 <= 0;
      __delay_data_899 <= 0;
      __delay_data_901 <= 0;
      __delay_data_902 <= 0;
      __delay_data_905 <= 0;
      __delay_data_908 <= 0;
      __delay_data_910 <= 0;
      __delay_data_911 <= 0;
      __delay_data_914 <= 0;
      __delay_data_917 <= 0;
      __delay_data_919 <= 0;
      __delay_data_920 <= 0;
      __delay_data_923 <= 0;
      __delay_data_925 <= 0;
      __delay_data_928 <= 0;
      __delay_data_933 <= 0;
      __delay_data_941 <= 0;
      __delay_data_949 <= 0;
      __delay_data_962 <= 0;
      __delay_data_963 <= 0;
      __delay_data_964 <= 0;
      __delay_data_967 <= 0;
      __delay_data_968 <= 0;
      __delay_data_969 <= 0;
      __delay_data_972 <= 0;
      __delay_data_973 <= 0;
      __delay_data_974 <= 0;
      __delay_data_977 <= 0;
      __delay_data_980 <= 0;
      __delay_data_985 <= 0;
      __delay_data_993 <= 0;
      __delay_data_1000 <= 0;
      __delay_data_1013 <= 0;
      __delay_data_1014 <= 0;
      __delay_data_1017 <= 0;
      __delay_data_1018 <= 0;
      __delay_data_1021 <= 0;
      __delay_data_1022 <= 0;
      __delay_data_1025 <= 0;
      __delay_data_1028 <= 0;
      __delay_data_1033 <= 0;
      __delay_data_1041 <= 0;
      __delay_data_1048 <= 0;
      __delay_data_1061 <= 0;
      __delay_data_1064 <= 0;
      __delay_data_1069 <= 0;
      __delay_data_1076 <= 0;
      __delay_data_1083 <= 0;
      __delay_data_1096 <= 0;
      __delay_data_1099 <= 0;
      __delay_data_1104 <= 0;
      __delay_data_1111 <= 0;
      __delay_data_1118 <= 0;
      __delay_data_1131 <= 0;
      __delay_data_1134 <= 0;
      __delay_data_1139 <= 0;
      __delay_data_1146 <= 0;
      __delay_data_1153 <= 0;
      __delay_data_1166 <= 0;
      __delay_data_1169 <= 0;
      __delay_data_1173 <= 0;
      __delay_data_1180 <= 0;
      __delay_data_1187 <= 0;
      __delay_data_1200 <= 0;
      __delay_data_1203 <= 0;
      __delay_data_1207 <= 0;
      __delay_data_1214 <= 0;
      __delay_data_1221 <= 0;
      __delay_data_1234 <= 0;
      __delay_data_1237 <= 0;
      __delay_data_1241 <= 0;
      __delay_data_1248 <= 0;
      __delay_data_1255 <= 0;
      __delay_data_1290 <= 0;
      __delay_data_1311 <= 0;
      __delay_data_1340 <= 0;
      _cond_data_283 <= 0;
      _cond_data_293 <= 0;
      _cond_data_303 <= 0;
      _cond_data_313 <= 0;
      _cond_data_323 <= 0;
      _cond_data_333 <= 0;
      _cond_data_343 <= 0;
      _cond_data_353 <= 0;
      _cond_data_363 <= 0;
      __delay_data_903 <= 0;
      __delay_data_906 <= 0;
      __delay_data_912 <= 0;
      __delay_data_915 <= 0;
      __delay_data_921 <= 0;
      __delay_data_924 <= 0;
      __delay_data_926 <= 0;
      __delay_data_929 <= 0;
      __delay_data_934 <= 0;
      __delay_data_942 <= 0;
      __delay_data_950 <= 0;
      __delay_data_956 <= 0;
      __delay_data_965 <= 0;
      __delay_data_966 <= 0;
      __delay_data_970 <= 0;
      __delay_data_971 <= 0;
      __delay_data_975 <= 0;
      __delay_data_976 <= 0;
      __delay_data_978 <= 0;
      __delay_data_981 <= 0;
      __delay_data_986 <= 0;
      __delay_data_994 <= 0;
      __delay_data_1001 <= 0;
      __delay_data_1007 <= 0;
      __delay_data_1015 <= 0;
      __delay_data_1016 <= 0;
      __delay_data_1019 <= 0;
      __delay_data_1020 <= 0;
      __delay_data_1023 <= 0;
      __delay_data_1024 <= 0;
      __delay_data_1026 <= 0;
      __delay_data_1029 <= 0;
      __delay_data_1034 <= 0;
      __delay_data_1042 <= 0;
      __delay_data_1049 <= 0;
      __delay_data_1055 <= 0;
      __delay_data_1062 <= 0;
      __delay_data_1065 <= 0;
      __delay_data_1070 <= 0;
      __delay_data_1077 <= 0;
      __delay_data_1084 <= 0;
      __delay_data_1090 <= 0;
      __delay_data_1097 <= 0;
      __delay_data_1100 <= 0;
      __delay_data_1105 <= 0;
      __delay_data_1112 <= 0;
      __delay_data_1119 <= 0;
      __delay_data_1125 <= 0;
      __delay_data_1132 <= 0;
      __delay_data_1135 <= 0;
      __delay_data_1140 <= 0;
      __delay_data_1147 <= 0;
      __delay_data_1154 <= 0;
      __delay_data_1160 <= 0;
      __delay_data_1167 <= 0;
      __delay_data_1170 <= 0;
      __delay_data_1174 <= 0;
      __delay_data_1181 <= 0;
      __delay_data_1188 <= 0;
      __delay_data_1194 <= 0;
      __delay_data_1201 <= 0;
      __delay_data_1204 <= 0;
      __delay_data_1208 <= 0;
      __delay_data_1215 <= 0;
      __delay_data_1222 <= 0;
      __delay_data_1228 <= 0;
      __delay_data_1235 <= 0;
      __delay_data_1238 <= 0;
      __delay_data_1242 <= 0;
      __delay_data_1249 <= 0;
      __delay_data_1256 <= 0;
      __delay_data_1262 <= 0;
      __delay_data_1269 <= 0;
      __delay_data_1291 <= 0;
      __delay_data_1312 <= 0;
      __delay_data_1341 <= 0;
      __delay_data_1369 <= 0;
      _cond_data_286 <= 0;
      _cond_data_296 <= 0;
      _cond_data_306 <= 0;
      _cond_data_316 <= 0;
      _cond_data_326 <= 0;
      _cond_data_336 <= 0;
      _cond_data_346 <= 0;
      _cond_data_356 <= 0;
      _cond_data_366 <= 0;
      __delay_data_927 <= 0;
      __delay_data_930 <= 0;
      __delay_data_935 <= 0;
      __delay_data_943 <= 0;
      __delay_data_951 <= 0;
      __delay_data_957 <= 0;
      __delay_data_979 <= 0;
      __delay_data_982 <= 0;
      __delay_data_987 <= 0;
      __delay_data_995 <= 0;
      __delay_data_1002 <= 0;
      __delay_data_1008 <= 0;
      __delay_data_1027 <= 0;
      __delay_data_1030 <= 0;
      __delay_data_1035 <= 0;
      __delay_data_1043 <= 0;
      __delay_data_1050 <= 0;
      __delay_data_1056 <= 0;
      __delay_data_1063 <= 0;
      __delay_data_1066 <= 0;
      __delay_data_1071 <= 0;
      __delay_data_1078 <= 0;
      __delay_data_1085 <= 0;
      __delay_data_1091 <= 0;
      __delay_data_1098 <= 0;
      __delay_data_1101 <= 0;
      __delay_data_1106 <= 0;
      __delay_data_1113 <= 0;
      __delay_data_1120 <= 0;
      __delay_data_1126 <= 0;
      __delay_data_1133 <= 0;
      __delay_data_1136 <= 0;
      __delay_data_1141 <= 0;
      __delay_data_1148 <= 0;
      __delay_data_1155 <= 0;
      __delay_data_1161 <= 0;
      __delay_data_1168 <= 0;
      __delay_data_1171 <= 0;
      __delay_data_1175 <= 0;
      __delay_data_1182 <= 0;
      __delay_data_1189 <= 0;
      __delay_data_1195 <= 0;
      __delay_data_1202 <= 0;
      __delay_data_1205 <= 0;
      __delay_data_1209 <= 0;
      __delay_data_1216 <= 0;
      __delay_data_1223 <= 0;
      __delay_data_1229 <= 0;
      __delay_data_1236 <= 0;
      __delay_data_1239 <= 0;
      __delay_data_1243 <= 0;
      __delay_data_1250 <= 0;
      __delay_data_1257 <= 0;
      __delay_data_1263 <= 0;
      __delay_data_1270 <= 0;
      __delay_data_1292 <= 0;
      __delay_data_1313 <= 0;
      __delay_data_1342 <= 0;
      __delay_data_1370 <= 0;
      _cond_data_369 <= 0;
      _cond_data_379 <= 0;
      _cond_data_389 <= 0;
      _cond_data_399 <= 0;
      _cond_data_409 <= 0;
      _cond_data_419 <= 0;
      _cond_data_429 <= 0;
      _cond_data_439 <= 0;
      _cond_data_449 <= 0;
      __delay_data_931 <= 0;
      __delay_data_932 <= 0;
      __delay_data_936 <= 0;
      __delay_data_938 <= 0;
      __delay_data_944 <= 0;
      __delay_data_952 <= 0;
      __delay_data_958 <= 0;
      __delay_data_983 <= 0;
      __delay_data_984 <= 0;
      __delay_data_988 <= 0;
      __delay_data_990 <= 0;
      __delay_data_996 <= 0;
      __delay_data_1003 <= 0;
      __delay_data_1009 <= 0;
      __delay_data_1031 <= 0;
      __delay_data_1032 <= 0;
      __delay_data_1036 <= 0;
      __delay_data_1038 <= 0;
      __delay_data_1044 <= 0;
      __delay_data_1051 <= 0;
      __delay_data_1057 <= 0;
      __delay_data_1067 <= 0;
      __delay_data_1068 <= 0;
      __delay_data_1072 <= 0;
      __delay_data_1079 <= 0;
      __delay_data_1086 <= 0;
      __delay_data_1092 <= 0;
      __delay_data_1102 <= 0;
      __delay_data_1103 <= 0;
      __delay_data_1107 <= 0;
      __delay_data_1114 <= 0;
      __delay_data_1121 <= 0;
      __delay_data_1127 <= 0;
      __delay_data_1137 <= 0;
      __delay_data_1138 <= 0;
      __delay_data_1142 <= 0;
      __delay_data_1149 <= 0;
      __delay_data_1156 <= 0;
      __delay_data_1162 <= 0;
      __delay_data_1172 <= 0;
      __delay_data_1176 <= 0;
      __delay_data_1183 <= 0;
      __delay_data_1190 <= 0;
      __delay_data_1196 <= 0;
      __delay_data_1206 <= 0;
      __delay_data_1210 <= 0;
      __delay_data_1217 <= 0;
      __delay_data_1224 <= 0;
      __delay_data_1230 <= 0;
      __delay_data_1240 <= 0;
      __delay_data_1244 <= 0;
      __delay_data_1251 <= 0;
      __delay_data_1258 <= 0;
      __delay_data_1264 <= 0;
      __delay_data_1271 <= 0;
      __delay_data_1293 <= 0;
      __delay_data_1314 <= 0;
      __delay_data_1343 <= 0;
      __delay_data_1371 <= 0;
      _cond_data_373 <= 0;
      _cond_data_383 <= 0;
      _cond_data_393 <= 0;
      _cond_data_403 <= 0;
      _cond_data_413 <= 0;
      _cond_data_423 <= 0;
      _cond_data_433 <= 0;
      _cond_data_443 <= 0;
      _cond_data_453 <= 0;
      __delay_data_937 <= 0;
      __delay_data_939 <= 0;
      __delay_data_945 <= 0;
      __delay_data_953 <= 0;
      __delay_data_959 <= 0;
      __delay_data_989 <= 0;
      __delay_data_991 <= 0;
      __delay_data_997 <= 0;
      __delay_data_1004 <= 0;
      __delay_data_1010 <= 0;
      __delay_data_1037 <= 0;
      __delay_data_1039 <= 0;
      __delay_data_1045 <= 0;
      __delay_data_1052 <= 0;
      __delay_data_1058 <= 0;
      __delay_data_1073 <= 0;
      __delay_data_1074 <= 0;
      __delay_data_1080 <= 0;
      __delay_data_1087 <= 0;
      __delay_data_1093 <= 0;
      __delay_data_1108 <= 0;
      __delay_data_1109 <= 0;
      __delay_data_1115 <= 0;
      __delay_data_1122 <= 0;
      __delay_data_1128 <= 0;
      __delay_data_1143 <= 0;
      __delay_data_1144 <= 0;
      __delay_data_1150 <= 0;
      __delay_data_1157 <= 0;
      __delay_data_1163 <= 0;
      __delay_data_1177 <= 0;
      __delay_data_1178 <= 0;
      __delay_data_1184 <= 0;
      __delay_data_1191 <= 0;
      __delay_data_1197 <= 0;
      __delay_data_1211 <= 0;
      __delay_data_1212 <= 0;
      __delay_data_1218 <= 0;
      __delay_data_1225 <= 0;
      __delay_data_1231 <= 0;
      __delay_data_1245 <= 0;
      __delay_data_1246 <= 0;
      __delay_data_1252 <= 0;
      __delay_data_1259 <= 0;
      __delay_data_1265 <= 0;
      __delay_data_1272 <= 0;
      __delay_data_1294 <= 0;
      __delay_data_1315 <= 0;
      __delay_data_1344 <= 0;
      __delay_data_1372 <= 0;
      _cond_data_376 <= 0;
      _cond_data_386 <= 0;
      _cond_data_396 <= 0;
      _cond_data_406 <= 0;
      _cond_data_416 <= 0;
      _cond_data_426 <= 0;
      _cond_data_436 <= 0;
      _cond_data_446 <= 0;
      _cond_data_456 <= 0;
      __delay_data_946 <= 0;
      __delay_data_954 <= 0;
      __delay_data_960 <= 0;
      __delay_data_998 <= 0;
      __delay_data_1005 <= 0;
      __delay_data_1011 <= 0;
      __delay_data_1046 <= 0;
      __delay_data_1053 <= 0;
      __delay_data_1059 <= 0;
      __delay_data_1081 <= 0;
      __delay_data_1088 <= 0;
      __delay_data_1094 <= 0;
      __delay_data_1116 <= 0;
      __delay_data_1123 <= 0;
      __delay_data_1129 <= 0;
      __delay_data_1151 <= 0;
      __delay_data_1158 <= 0;
      __delay_data_1164 <= 0;
      __delay_data_1185 <= 0;
      __delay_data_1192 <= 0;
      __delay_data_1198 <= 0;
      __delay_data_1219 <= 0;
      __delay_data_1226 <= 0;
      __delay_data_1232 <= 0;
      __delay_data_1253 <= 0;
      __delay_data_1260 <= 0;
      __delay_data_1266 <= 0;
      __delay_data_1273 <= 0;
      __delay_data_1295 <= 0;
      __delay_data_1316 <= 0;
      __delay_data_1345 <= 0;
      __delay_data_1373 <= 0;
      _cond_data_575 <= 0;
      _cond_data_577 <= 0;
      _cond_data_579 <= 0;
      _cond_data_581 <= 0;
      _cond_data_583 <= 0;
      _cond_data_585 <= 0;
      _cond_data_587 <= 0;
      _cond_data_589 <= 0;
      _cond_data_591 <= 0;
      __delay_data_955 <= 0;
      __delay_data_961 <= 0;
      __delay_data_1006 <= 0;
      __delay_data_1012 <= 0;
      __delay_data_1054 <= 0;
      __delay_data_1060 <= 0;
      __delay_data_1089 <= 0;
      __delay_data_1095 <= 0;
      __delay_data_1124 <= 0;
      __delay_data_1130 <= 0;
      __delay_data_1159 <= 0;
      __delay_data_1165 <= 0;
      __delay_data_1193 <= 0;
      __delay_data_1199 <= 0;
      __delay_data_1227 <= 0;
      __delay_data_1233 <= 0;
      __delay_data_1261 <= 0;
      __delay_data_1267 <= 0;
      __delay_data_1274 <= 0;
      __delay_data_1296 <= 0;
      __delay_data_1317 <= 0;
      __delay_data_1346 <= 0;
      __delay_data_1374 <= 0;
      __delay_data_1275 <= 0;
      __delay_data_1297 <= 0;
      __delay_data_1318 <= 0;
      __delay_data_1347 <= 0;
      __delay_data_1375 <= 0;
      __delay_data_1276 <= 0;
      __delay_data_1298 <= 0;
      __delay_data_1319 <= 0;
      __delay_data_1348 <= 0;
      __delay_data_1376 <= 0;
      __delay_data_1277 <= 0;
      __delay_data_1299 <= 0;
      __delay_data_1320 <= 0;
      __delay_data_1349 <= 0;
      __delay_data_1377 <= 0;
      __delay_data_1278 <= 0;
      __delay_data_1300 <= 0;
      __delay_data_1321 <= 0;
      __delay_data_1350 <= 0;
      __delay_data_1378 <= 0;
      __delay_data_1279 <= 0;
      __delay_data_1301 <= 0;
      __delay_data_1322 <= 0;
      __delay_data_1351 <= 0;
      __delay_data_1379 <= 0;
      __delay_data_1280 <= 0;
      __delay_data_1302 <= 0;
      __delay_data_1323 <= 0;
      __delay_data_1352 <= 0;
      __delay_data_1380 <= 0;
      __delay_data_1281 <= 0;
      __delay_data_1303 <= 0;
      __delay_data_1324 <= 0;
      __delay_data_1353 <= 0;
      __delay_data_1381 <= 0;
      __delay_data_1282 <= 0;
      __delay_data_1304 <= 0;
      __delay_data_1325 <= 0;
      __delay_data_1354 <= 0;
      __delay_data_1382 <= 0;
      __delay_data_1283 <= 0;
      __delay_data_1305 <= 0;
      __delay_data_1326 <= 0;
      __delay_data_1355 <= 0;
      __delay_data_1383 <= 0;
      __substreamoutput_data_608 <= 0;
      __substreamoutput_data_625 <= 0;
      __substreamoutput_data_642 <= 0;
      __substreamoutput_data_659 <= 0;
      __substreamoutput_data_676 <= 0;
      __substreamoutput_data_693 <= 0;
      __substreamoutput_data_710 <= 0;
      __substreamoutput_data_727 <= 0;
      __substreamoutput_data_744 <= 0;
      __delay_data_1284 <= 0;
      __delay_data_1306 <= 0;
      __delay_data_1327 <= 0;
      __delay_data_1356 <= 0;
      __delay_data_1384 <= 0;
      __delay_data_1285 <= 0;
      __delay_data_1307 <= 0;
      __delay_data_1328 <= 0;
      __delay_data_1357 <= 0;
      __delay_data_1385 <= 0;
      __delay_data_1286 <= 0;
      __delay_data_1308 <= 0;
      __delay_data_1329 <= 0;
      __delay_data_1358 <= 0;
      __delay_data_1386 <= 0;
      __delay_data_1287 <= 0;
      __delay_data_1309 <= 0;
      __delay_data_1330 <= 0;
      __delay_data_1359 <= 0;
      __delay_data_1387 <= 0;
      __substreamoutput_data_746 <= 0;
      __delay_data_1288 <= 0;
      __delay_data_1310 <= 0;
      __delay_data_1331 <= 0;
      __delay_data_1360 <= 0;
      __delay_data_1388 <= 0;
      __delay_data_1332 <= 0;
      __delay_data_1361 <= 0;
      __delay_data_1389 <= 0;
      __delay_data_1333 <= 0;
      __delay_data_1362 <= 0;
      __delay_data_1390 <= 0;
      __delay_data_1334 <= 0;
      __delay_data_1363 <= 0;
      __delay_data_1391 <= 0;
      __delay_data_1335 <= 0;
      __delay_data_1364 <= 0;
      __delay_data_1392 <= 0;
      __delay_data_1336 <= 0;
      __delay_data_1365 <= 0;
      __delay_data_1393 <= 0;
      __delay_data_1337 <= 0;
      __delay_data_1366 <= 0;
      __delay_data_1394 <= 0;
      __substreamoutput_data_760 <= 0;
      __substreamoutput_data_761 <= 0;
      __delay_data_1338 <= 0;
      __delay_data_1367 <= 0;
      __delay_data_1395 <= 0;
      _plus_data_762 <= 0;
      __delay_data_1368 <= 0;
      __delay_data_1396 <= 0;
      __delay_data_1398 <= 0;
      __delay_data_1399 <= 0;
      __delay_data_1400 <= 0;
      __delay_data_1401 <= 0;
      __delay_data_1402 <= 0;
      __delay_data_1403 <= 0;
      __delay_data_1404 <= 0;
      __delay_data_1405 <= 0;
      __delay_data_1406 <= 0;
      __delay_data_1407 <= 0;
      __substreamoutput_data_771 <= 0;
      __delay_data_1408 <= 0;
      _greaterthan_data_773 <= 0;
      __delay_data_1397 <= 0;
      __delay_data_1409 <= 0;
      _cond_data_775 <= 0;
      __delay_data_1410 <= 0;
      _set_flag_457 <= 0;
      _stream_conv2d_16_constant_0_next_constant_data <= 0;
      __variable_wdata_214 <= 0;
      _set_flag_458 <= 0;
      _stream_conv2d_16_constant_1_next_constant_data <= 0;
      __variable_wdata_215 <= 0;
      _set_flag_459 <= 0;
      _stream_conv2d_16_constant_2_next_constant_data <= 0;
      __variable_wdata_216 <= 0;
      _set_flag_460 <= 0;
      _stream_conv2d_16_constant_3_next_constant_data <= 0;
      __variable_wdata_217 <= 0;
      _set_flag_461 <= 0;
      _stream_conv2d_16_constant_4_next_constant_data <= 0;
      __variable_wdata_218 <= 0;
      _set_flag_462 <= 0;
      _stream_conv2d_16_constant_5_next_constant_data <= 0;
      __variable_wdata_229 <= 0;
      _set_flag_463 <= 0;
      _stream_conv2d_16_source_6_source_mode <= 3'b0;
      _stream_conv2d_16_source_6_source_offset <= 0;
      _source_stream_conv2d_16_source_6_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_6_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_6_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_6_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_6_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_6_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_6_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_6_pat_stride_3 <= 0;
      _stream_conv2d_16_source_6_source_ram_sel <= 0;
      __tmp_472_1 <= 0;
      __variable_wdata_230 <= 0;
      _stream_conv2d_16_source_6_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_6_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_6_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_6_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_6_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_6_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_6_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_6_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_6_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_6_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_6_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_6_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_6_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_6_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_6_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_6_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_6_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_6_source_ram_raddr <= 0;
      _stream_conv2d_16_source_6_source_ram_renable <= 0;
      _set_flag_473 <= 0;
      _stream_conv2d_16_constant_7_next_constant_data <= 0;
      __variable_wdata_236 <= 0;
      _set_flag_474 <= 0;
      _stream_conv2d_16_source_8_source_mode <= 3'b0;
      _stream_conv2d_16_source_8_source_offset <= 0;
      _source_stream_conv2d_16_source_8_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_8_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_8_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_8_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_8_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_8_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_8_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_8_pat_stride_3 <= 0;
      _stream_conv2d_16_source_8_source_ram_sel <= 0;
      __tmp_483_1 <= 0;
      __variable_wdata_237 <= 0;
      _stream_conv2d_16_source_8_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_8_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_8_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_8_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_8_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_8_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_8_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_8_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_8_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_8_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_8_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_8_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_8_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_8_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_8_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_8_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_8_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_8_source_ram_raddr <= 0;
      _stream_conv2d_16_source_8_source_ram_renable <= 0;
      _set_flag_484 <= 0;
      _stream_conv2d_16_constant_9_next_constant_data <= 0;
      __variable_wdata_243 <= 0;
      _set_flag_485 <= 0;
      _stream_conv2d_16_source_10_source_mode <= 3'b0;
      _stream_conv2d_16_source_10_source_empty_data <= 0;
      __variable_wdata_244 <= 0;
      _set_flag_486 <= 0;
      _stream_conv2d_16_constant_11_next_constant_data <= 0;
      __variable_wdata_250 <= 0;
      _set_flag_487 <= 0;
      _stream_conv2d_16_source_12_source_mode <= 3'b0;
      _stream_conv2d_16_source_12_source_empty_data <= 0;
      __variable_wdata_251 <= 0;
      _set_flag_488 <= 0;
      _stream_conv2d_16_constant_13_next_constant_data <= 0;
      __variable_wdata_257 <= 0;
      _set_flag_489 <= 0;
      _stream_conv2d_16_source_14_source_mode <= 3'b0;
      _stream_conv2d_16_source_14_source_empty_data <= 0;
      __variable_wdata_258 <= 0;
      _set_flag_490 <= 0;
      _stream_conv2d_16_constant_15_next_constant_data <= 0;
      __variable_wdata_264 <= 0;
      _set_flag_491 <= 0;
      _stream_conv2d_16_constant_16_next_constant_data <= 0;
      __variable_wdata_265 <= 0;
      _set_flag_492 <= 0;
      _stream_conv2d_16_constant_17_next_constant_data <= 0;
      __variable_wdata_266 <= 0;
      _set_flag_493 <= 0;
      _stream_conv2d_16_constant_18_next_constant_data <= 0;
      __variable_wdata_267 <= 0;
      _set_flag_494 <= 0;
      _stream_conv2d_16_source_19_source_mode <= 3'b0;
      _stream_conv2d_16_source_19_source_offset <= 0;
      _source_stream_conv2d_16_source_19_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_19_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_19_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_19_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_19_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_19_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_19_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_19_pat_stride_3 <= 0;
      _stream_conv2d_16_source_19_source_ram_sel <= 0;
      __tmp_503_1 <= 0;
      __variable_wdata_268 <= 0;
      _stream_conv2d_16_source_19_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_19_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_19_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_19_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_19_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_19_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_19_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_19_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_19_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_19_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_19_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_19_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_19_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_19_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_19_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_19_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_19_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_19_source_ram_raddr <= 0;
      _stream_conv2d_16_source_19_source_ram_renable <= 0;
      _set_flag_504 <= 0;
      _stream_conv2d_16_source_20_source_mode <= 3'b0;
      _stream_conv2d_16_source_20_source_offset <= 0;
      _source_stream_conv2d_16_source_20_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_20_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_20_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_20_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_20_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_20_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_20_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_20_pat_stride_3 <= 0;
      _stream_conv2d_16_source_20_source_ram_sel <= 0;
      __tmp_513_1 <= 0;
      __variable_wdata_269 <= 0;
      _stream_conv2d_16_source_20_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_20_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_20_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_20_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_20_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_20_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_20_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_20_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_20_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_20_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_20_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_20_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_20_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_20_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_20_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_20_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_20_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_20_source_ram_raddr <= 0;
      _stream_conv2d_16_source_20_source_ram_renable <= 0;
      _set_flag_514 <= 0;
      _stream_conv2d_16_source_21_source_mode <= 3'b0;
      _stream_conv2d_16_source_21_source_offset <= 0;
      _source_stream_conv2d_16_source_21_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_21_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_21_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_21_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_21_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_21_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_21_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_21_pat_stride_3 <= 0;
      _stream_conv2d_16_source_21_source_ram_sel <= 0;
      __tmp_523_1 <= 0;
      __variable_wdata_270 <= 0;
      _stream_conv2d_16_source_21_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_21_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_21_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_21_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_21_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_21_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_21_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_21_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_21_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_21_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_21_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_21_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_21_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_21_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_21_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_21_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_21_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_21_source_ram_raddr <= 0;
      _stream_conv2d_16_source_21_source_ram_renable <= 0;
      _set_flag_524 <= 0;
      _stream_conv2d_16_source_22_source_mode <= 3'b0;
      _stream_conv2d_16_source_22_source_offset <= 0;
      _source_stream_conv2d_16_source_22_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_22_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_22_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_22_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_22_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_22_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_22_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_22_pat_stride_3 <= 0;
      _stream_conv2d_16_source_22_source_ram_sel <= 0;
      __tmp_533_1 <= 0;
      __variable_wdata_271 <= 0;
      _stream_conv2d_16_source_22_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_22_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_22_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_22_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_22_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_22_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_22_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_22_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_22_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_22_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_22_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_22_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_22_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_22_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_22_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_22_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_22_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_22_source_ram_raddr <= 0;
      _stream_conv2d_16_source_22_source_ram_renable <= 0;
      _set_flag_534 <= 0;
      _stream_conv2d_16_source_23_source_mode <= 3'b0;
      _stream_conv2d_16_source_23_source_offset <= 0;
      _source_stream_conv2d_16_source_23_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_23_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_23_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_23_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_23_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_23_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_23_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_23_pat_stride_3 <= 0;
      _stream_conv2d_16_source_23_source_ram_sel <= 0;
      __tmp_543_1 <= 0;
      __variable_wdata_272 <= 0;
      _stream_conv2d_16_source_23_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_23_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_23_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_23_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_23_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_23_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_23_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_23_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_23_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_23_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_23_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_23_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_23_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_23_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_23_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_23_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_23_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_23_source_ram_raddr <= 0;
      _stream_conv2d_16_source_23_source_ram_renable <= 0;
      _set_flag_544 <= 0;
      _stream_conv2d_16_source_24_source_mode <= 3'b0;
      _stream_conv2d_16_source_24_source_offset <= 0;
      _source_stream_conv2d_16_source_24_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_24_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_24_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_24_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_24_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_24_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_24_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_24_pat_stride_3 <= 0;
      _stream_conv2d_16_source_24_source_ram_sel <= 0;
      __tmp_553_1 <= 0;
      __variable_wdata_273 <= 0;
      _stream_conv2d_16_source_24_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_24_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_24_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_24_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_24_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_24_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_24_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_24_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_24_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_24_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_24_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_24_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_24_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_24_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_24_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_24_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_24_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_24_source_ram_raddr <= 0;
      _stream_conv2d_16_source_24_source_ram_renable <= 0;
      _set_flag_554 <= 0;
      _stream_conv2d_16_source_25_source_mode <= 3'b0;
      _stream_conv2d_16_source_25_source_offset <= 0;
      _source_stream_conv2d_16_source_25_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_25_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_25_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_25_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_25_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_25_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_25_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_25_pat_stride_3 <= 0;
      _stream_conv2d_16_source_25_source_ram_sel <= 0;
      __tmp_563_1 <= 0;
      __variable_wdata_274 <= 0;
      _stream_conv2d_16_source_25_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_25_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_25_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_25_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_25_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_25_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_25_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_25_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_25_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_25_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_25_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_25_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_25_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_25_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_25_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_25_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_25_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_25_source_ram_raddr <= 0;
      _stream_conv2d_16_source_25_source_ram_renable <= 0;
      _set_flag_564 <= 0;
      _stream_conv2d_16_source_26_source_mode <= 3'b0;
      _stream_conv2d_16_source_26_source_offset <= 0;
      _source_stream_conv2d_16_source_26_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_26_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_26_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_26_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_26_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_26_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_26_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_26_pat_stride_3 <= 0;
      _stream_conv2d_16_source_26_source_ram_sel <= 0;
      __tmp_573_1 <= 0;
      __variable_wdata_275 <= 0;
      _stream_conv2d_16_source_26_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_26_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_26_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_26_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_26_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_26_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_26_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_26_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_26_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_26_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_26_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_26_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_26_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_26_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_26_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_26_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_26_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_26_source_ram_raddr <= 0;
      _stream_conv2d_16_source_26_source_ram_renable <= 0;
      _set_flag_574 <= 0;
      _stream_conv2d_16_source_27_source_mode <= 3'b0;
      _stream_conv2d_16_source_27_source_offset <= 0;
      _source_stream_conv2d_16_source_27_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_27_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_27_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_27_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_27_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_27_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_27_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_27_pat_stride_3 <= 0;
      _stream_conv2d_16_source_27_source_ram_sel <= 0;
      __tmp_583_1 <= 0;
      __variable_wdata_276 <= 0;
      _stream_conv2d_16_source_27_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_27_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_27_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_27_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_27_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_27_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_27_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_27_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_27_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_27_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_27_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_27_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_27_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_27_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_27_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_27_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_27_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_27_source_ram_raddr <= 0;
      _stream_conv2d_16_source_27_source_ram_renable <= 0;
      _set_flag_584 <= 0;
      _stream_conv2d_16_source_28_source_mode <= 3'b0;
      _stream_conv2d_16_source_28_source_offset <= 0;
      _source_stream_conv2d_16_source_28_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_28_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_28_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_28_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_28_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_28_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_28_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_28_pat_stride_3 <= 0;
      _stream_conv2d_16_source_28_source_ram_sel <= 0;
      __tmp_597_1 <= 0;
      __variable_wdata_502 <= 0;
      _stream_conv2d_16_source_28_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_28_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_28_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_28_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_28_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_28_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_28_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_28_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_28_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_28_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_28_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_28_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_28_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_28_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_28_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_28_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_28_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_28_source_ram_raddr <= 0;
      _stream_conv2d_16_source_28_source_ram_renable <= 0;
      _set_flag_598 <= 0;
      _stream_conv2d_16_source_29_source_mode <= 3'b0;
      _stream_conv2d_16_source_29_source_offset <= 0;
      _source_stream_conv2d_16_source_29_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_29_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_29_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_29_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_29_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_29_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_29_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_29_pat_stride_3 <= 0;
      _stream_conv2d_16_source_29_source_ram_sel <= 0;
      __tmp_611_1 <= 0;
      __variable_wdata_503 <= 0;
      _stream_conv2d_16_source_29_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_29_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_29_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_29_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_29_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_29_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_29_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_29_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_29_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_29_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_29_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_29_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_29_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_29_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_29_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_29_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_29_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_29_source_ram_raddr <= 0;
      _stream_conv2d_16_source_29_source_ram_renable <= 0;
      _set_flag_612 <= 0;
      _stream_conv2d_16_source_30_source_mode <= 3'b0;
      _stream_conv2d_16_source_30_source_offset <= 0;
      _source_stream_conv2d_16_source_30_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_30_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_30_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_30_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_30_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_30_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_30_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_30_pat_stride_3 <= 0;
      _stream_conv2d_16_source_30_source_ram_sel <= 0;
      __tmp_625_1 <= 0;
      __variable_wdata_504 <= 0;
      _stream_conv2d_16_source_30_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_30_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_30_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_30_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_30_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_30_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_30_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_30_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_30_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_30_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_30_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_30_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_30_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_30_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_30_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_30_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_30_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_30_source_ram_raddr <= 0;
      _stream_conv2d_16_source_30_source_ram_renable <= 0;
      _set_flag_626 <= 0;
      _stream_conv2d_16_source_31_source_mode <= 3'b0;
      _stream_conv2d_16_source_31_source_offset <= 0;
      _source_stream_conv2d_16_source_31_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_31_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_31_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_31_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_31_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_31_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_31_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_31_pat_stride_3 <= 0;
      _stream_conv2d_16_source_31_source_ram_sel <= 0;
      __tmp_639_1 <= 0;
      __variable_wdata_505 <= 0;
      _stream_conv2d_16_source_31_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_31_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_31_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_31_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_31_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_31_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_31_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_31_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_31_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_31_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_31_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_31_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_31_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_31_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_31_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_31_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_31_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_31_source_ram_raddr <= 0;
      _stream_conv2d_16_source_31_source_ram_renable <= 0;
      _set_flag_640 <= 0;
      _stream_conv2d_16_source_32_source_mode <= 3'b0;
      _stream_conv2d_16_source_32_source_offset <= 0;
      _source_stream_conv2d_16_source_32_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_32_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_32_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_32_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_32_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_32_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_32_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_32_pat_stride_3 <= 0;
      _stream_conv2d_16_source_32_source_ram_sel <= 0;
      __tmp_653_1 <= 0;
      __variable_wdata_506 <= 0;
      _stream_conv2d_16_source_32_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_32_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_32_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_32_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_32_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_32_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_32_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_32_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_32_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_32_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_32_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_32_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_32_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_32_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_32_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_32_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_32_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_32_source_ram_raddr <= 0;
      _stream_conv2d_16_source_32_source_ram_renable <= 0;
      _set_flag_654 <= 0;
      _stream_conv2d_16_source_33_source_mode <= 3'b0;
      _stream_conv2d_16_source_33_source_offset <= 0;
      _source_stream_conv2d_16_source_33_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_33_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_33_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_33_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_33_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_33_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_33_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_33_pat_stride_3 <= 0;
      _stream_conv2d_16_source_33_source_ram_sel <= 0;
      __tmp_667_1 <= 0;
      __variable_wdata_507 <= 0;
      _stream_conv2d_16_source_33_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_33_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_33_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_33_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_33_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_33_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_33_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_33_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_33_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_33_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_33_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_33_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_33_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_33_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_33_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_33_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_33_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_33_source_ram_raddr <= 0;
      _stream_conv2d_16_source_33_source_ram_renable <= 0;
      _set_flag_668 <= 0;
      _stream_conv2d_16_source_34_source_mode <= 3'b0;
      _stream_conv2d_16_source_34_source_offset <= 0;
      _source_stream_conv2d_16_source_34_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_34_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_34_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_34_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_34_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_34_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_34_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_34_pat_stride_3 <= 0;
      _stream_conv2d_16_source_34_source_ram_sel <= 0;
      __tmp_681_1 <= 0;
      __variable_wdata_508 <= 0;
      _stream_conv2d_16_source_34_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_34_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_34_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_34_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_34_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_34_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_34_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_34_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_34_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_34_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_34_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_34_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_34_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_34_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_34_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_34_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_34_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_34_source_ram_raddr <= 0;
      _stream_conv2d_16_source_34_source_ram_renable <= 0;
      _set_flag_682 <= 0;
      _stream_conv2d_16_source_35_source_mode <= 3'b0;
      _stream_conv2d_16_source_35_source_offset <= 0;
      _source_stream_conv2d_16_source_35_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_35_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_35_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_35_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_35_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_35_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_35_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_35_pat_stride_3 <= 0;
      _stream_conv2d_16_source_35_source_ram_sel <= 0;
      __tmp_695_1 <= 0;
      __variable_wdata_509 <= 0;
      _stream_conv2d_16_source_35_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_35_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_35_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_35_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_35_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_35_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_35_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_35_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_35_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_35_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_35_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_35_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_35_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_35_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_35_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_35_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_35_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_35_source_ram_raddr <= 0;
      _stream_conv2d_16_source_35_source_ram_renable <= 0;
      _set_flag_696 <= 0;
      _stream_conv2d_16_source_36_source_mode <= 3'b0;
      _stream_conv2d_16_source_36_source_offset <= 0;
      _source_stream_conv2d_16_source_36_pat_size_0 <= 0;
      _source_stream_conv2d_16_source_36_pat_stride_0 <= 0;
      _source_stream_conv2d_16_source_36_pat_size_1 <= 0;
      _source_stream_conv2d_16_source_36_pat_stride_1 <= 0;
      _source_stream_conv2d_16_source_36_pat_size_2 <= 0;
      _source_stream_conv2d_16_source_36_pat_stride_2 <= 0;
      _source_stream_conv2d_16_source_36_pat_size_3 <= 0;
      _source_stream_conv2d_16_source_36_pat_stride_3 <= 0;
      _stream_conv2d_16_source_36_source_ram_sel <= 0;
      __tmp_709_1 <= 0;
      __variable_wdata_510 <= 0;
      _stream_conv2d_16_source_36_source_offset_buf <= 0;
      _source_stream_conv2d_16_source_36_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_16_source_36_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_16_source_36_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_16_source_36_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_16_source_36_pat_count_0 <= 0;
      _source_stream_conv2d_16_source_36_pat_count_1 <= 0;
      _source_stream_conv2d_16_source_36_pat_count_2 <= 0;
      _source_stream_conv2d_16_source_36_pat_count_3 <= 0;
      _source_stream_conv2d_16_source_36_pat_size_buf_0 <= 0;
      _source_stream_conv2d_16_source_36_pat_size_buf_1 <= 0;
      _source_stream_conv2d_16_source_36_pat_size_buf_2 <= 0;
      _source_stream_conv2d_16_source_36_pat_size_buf_3 <= 0;
      _source_stream_conv2d_16_source_36_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_16_source_36_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_16_source_36_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_16_source_36_pat_stride_buf_3 <= 0;
      _stream_conv2d_16_source_36_source_ram_raddr <= 0;
      _stream_conv2d_16_source_36_source_ram_renable <= 0;
      _set_flag_710 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_1 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_2 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_3 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_4 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_5 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_6 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_7 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_8 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_9 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_10 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_11 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_12 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_13 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_14 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_15 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_16 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_17 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_18 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_19 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_20 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_21 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_22 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_23 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_24 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_25 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_26 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_27 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_28 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_29 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_30 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_31 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_32 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_33 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_34 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_35 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_36 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_37 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_38 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_39 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_40 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_41 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_42 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_43 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_44 <= 0;
      __stream_conv2d_16_sink_37_sink_offset_0_45 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_1 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_2 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_3 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_4 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_5 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_6 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_7 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_8 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_9 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_10 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_11 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_12 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_13 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_14 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_15 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_16 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_17 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_18 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_19 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_20 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_21 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_22 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_23 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_24 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_25 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_26 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_27 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_28 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_29 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_30 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_31 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_32 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_33 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_34 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_35 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_36 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_37 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_38 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_39 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_40 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_41 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_42 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_43 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_44 <= 0;
      __stream_conv2d_16_sink_37_sink_size_1_45 <= 0;
      __stream_seq_14_cond_2_1 <= 0;
      __stream_seq_14_cond_2_2 <= 0;
      __stream_seq_14_cond_2_3 <= 0;
      __stream_seq_14_cond_2_4 <= 0;
      __stream_seq_14_cond_2_5 <= 0;
      __stream_seq_14_cond_2_6 <= 0;
      __stream_seq_14_cond_2_7 <= 0;
      __stream_seq_14_cond_2_8 <= 0;
      __stream_seq_14_cond_2_9 <= 0;
      __stream_seq_14_cond_2_10 <= 0;
      __stream_seq_14_cond_2_11 <= 0;
      __stream_seq_14_cond_2_12 <= 0;
      __stream_seq_14_cond_2_13 <= 0;
      __stream_seq_14_cond_2_14 <= 0;
      __stream_seq_14_cond_2_15 <= 0;
      __stream_seq_14_cond_2_16 <= 0;
      __stream_seq_14_cond_2_17 <= 0;
      __stream_seq_14_cond_2_18 <= 0;
      __stream_seq_14_cond_2_19 <= 0;
      __stream_seq_14_cond_2_20 <= 0;
      __stream_seq_14_cond_2_21 <= 0;
      __stream_seq_14_cond_2_22 <= 0;
      __stream_seq_14_cond_2_23 <= 0;
      __stream_seq_14_cond_2_24 <= 0;
      __stream_seq_14_cond_2_25 <= 0;
      __stream_seq_14_cond_2_26 <= 0;
      __stream_seq_14_cond_2_27 <= 0;
      __stream_seq_14_cond_2_28 <= 0;
      __stream_seq_14_cond_2_29 <= 0;
      __stream_seq_14_cond_2_30 <= 0;
      __stream_seq_14_cond_2_31 <= 0;
      __stream_seq_14_cond_2_32 <= 0;
      __stream_seq_14_cond_2_33 <= 0;
      __stream_seq_14_cond_2_34 <= 0;
      __stream_seq_14_cond_2_35 <= 0;
      __stream_seq_14_cond_2_36 <= 0;
      __stream_seq_14_cond_2_37 <= 0;
      __stream_seq_14_cond_2_38 <= 0;
      __stream_seq_14_cond_2_39 <= 0;
      __stream_seq_14_cond_2_40 <= 0;
      __stream_seq_14_cond_2_41 <= 0;
      __stream_seq_14_cond_2_42 <= 0;
      __stream_seq_14_cond_2_43 <= 0;
      __stream_seq_14_cond_2_44 <= 0;
      __stream_seq_14_cond_2_45 <= 0;
      _stream_conv2d_16_sink_37_sink_mode <= 3'b0;
      _stream_conv2d_16_sink_37_sink_offset <= 0;
      _stream_conv2d_16_sink_37_sink_size <= 0;
      _stream_conv2d_16_sink_37_sink_stride <= 0;
      __set_flag_710_1 <= 0;
      __set_flag_710_2 <= 0;
      __set_flag_710_3 <= 0;
      __set_flag_710_4 <= 0;
      __set_flag_710_5 <= 0;
      __set_flag_710_6 <= 0;
      __set_flag_710_7 <= 0;
      __set_flag_710_8 <= 0;
      __set_flag_710_9 <= 0;
      __set_flag_710_10 <= 0;
      __set_flag_710_11 <= 0;
      __set_flag_710_12 <= 0;
      __set_flag_710_13 <= 0;
      __set_flag_710_14 <= 0;
      __set_flag_710_15 <= 0;
      __set_flag_710_16 <= 0;
      __set_flag_710_17 <= 0;
      __set_flag_710_18 <= 0;
      __set_flag_710_19 <= 0;
      __set_flag_710_20 <= 0;
      __set_flag_710_21 <= 0;
      __set_flag_710_22 <= 0;
      __set_flag_710_23 <= 0;
      __set_flag_710_24 <= 0;
      __set_flag_710_25 <= 0;
      __set_flag_710_26 <= 0;
      __set_flag_710_27 <= 0;
      __set_flag_710_28 <= 0;
      __set_flag_710_29 <= 0;
      __set_flag_710_30 <= 0;
      __set_flag_710_31 <= 0;
      __set_flag_710_32 <= 0;
      __set_flag_710_33 <= 0;
      __set_flag_710_34 <= 0;
      __set_flag_710_35 <= 0;
      __set_flag_710_36 <= 0;
      __set_flag_710_37 <= 0;
      __set_flag_710_38 <= 0;
      __set_flag_710_39 <= 0;
      __set_flag_710_40 <= 0;
      __set_flag_710_41 <= 0;
      __set_flag_710_42 <= 0;
      __set_flag_710_43 <= 0;
      __set_flag_710_44 <= 0;
      __set_flag_710_45 <= 0;
      _stream_conv2d_16_sink_37_sink_ram_sel <= 0;
      __stream_conv2d_16_start_1 <= 0;
      __stream_conv2d_16_start_2 <= 0;
      __stream_conv2d_16_start_3 <= 0;
      __stream_conv2d_16_start_4 <= 0;
      __stream_conv2d_16_start_5 <= 0;
      __stream_conv2d_16_start_6 <= 0;
      __stream_conv2d_16_start_7 <= 0;
      __stream_conv2d_16_start_8 <= 0;
      __stream_conv2d_16_start_9 <= 0;
      __stream_conv2d_16_start_10 <= 0;
      __stream_conv2d_16_start_11 <= 0;
      __stream_conv2d_16_start_12 <= 0;
      __stream_conv2d_16_start_13 <= 0;
      __stream_conv2d_16_start_14 <= 0;
      __stream_conv2d_16_start_15 <= 0;
      __stream_conv2d_16_start_16 <= 0;
      __stream_conv2d_16_start_17 <= 0;
      __stream_conv2d_16_start_18 <= 0;
      __stream_conv2d_16_start_19 <= 0;
      __stream_conv2d_16_start_20 <= 0;
      __stream_conv2d_16_start_21 <= 0;
      __stream_conv2d_16_start_22 <= 0;
      __stream_conv2d_16_start_23 <= 0;
      __stream_conv2d_16_start_24 <= 0;
      __stream_conv2d_16_start_25 <= 0;
      __stream_conv2d_16_start_26 <= 0;
      __stream_conv2d_16_start_27 <= 0;
      __stream_conv2d_16_start_28 <= 0;
      __stream_conv2d_16_start_29 <= 0;
      __stream_conv2d_16_start_30 <= 0;
      __stream_conv2d_16_start_31 <= 0;
      __stream_conv2d_16_start_32 <= 0;
      __stream_conv2d_16_start_33 <= 0;
      __stream_conv2d_16_start_34 <= 0;
      __stream_conv2d_16_start_35 <= 0;
      __stream_conv2d_16_start_36 <= 0;
      __stream_conv2d_16_start_37 <= 0;
      __stream_conv2d_16_start_38 <= 0;
      __stream_conv2d_16_start_39 <= 0;
      __stream_conv2d_16_start_40 <= 0;
      __stream_conv2d_16_start_41 <= 0;
      __stream_conv2d_16_start_42 <= 0;
      __stream_conv2d_16_start_43 <= 0;
      __stream_conv2d_16_start_44 <= 0;
      __stream_conv2d_16_start_45 <= 0;
      __stream_conv2d_16_start_46 <= 0;
      _stream_conv2d_16_sink_37_sink_waddr <= 0;
      _stream_conv2d_16_sink_37_sink_count <= 0;
      _stream_conv2d_16_sink_37_sink_offset_buf <= 0;
      _stream_conv2d_16_sink_37_sink_stride_buf <= 0;
      _stream_conv2d_16_sink_37_sink_wdata <= 0;
      __tmp_713_1 <= 0;
      __tmp_713_2 <= 0;
      __tmp_713_3 <= 0;
      __tmp_713_4 <= 0;
      __tmp_713_5 <= 0;
      __tmp_715_1 <= 0;
      __tmp_715_2 <= 0;
      __tmp_715_3 <= 0;
      __tmp_715_4 <= 0;
      __tmp_715_5 <= 0;
      __tmp_715_6 <= 0;
      __tmp_715_7 <= 0;
      __tmp_715_8 <= 0;
      __tmp_715_9 <= 0;
      __tmp_715_10 <= 0;
      __tmp_715_11 <= 0;
      __tmp_715_12 <= 0;
      __tmp_717_1 <= 0;
      __tmp_717_2 <= 0;
      __tmp_717_3 <= 0;
      __tmp_717_4 <= 0;
      __tmp_717_5 <= 0;
      __tmp_717_6 <= 0;
      __tmp_717_7 <= 0;
      __tmp_717_8 <= 0;
      __tmp_717_9 <= 0;
      __tmp_717_10 <= 0;
      __tmp_717_11 <= 0;
      __tmp_717_12 <= 0;
      __tmp_719_1 <= 0;
      __tmp_719_2 <= 0;
      __tmp_719_3 <= 0;
      __tmp_719_4 <= 0;
      __tmp_719_5 <= 0;
      __tmp_719_6 <= 0;
      __tmp_719_7 <= 0;
      __tmp_719_8 <= 0;
      __tmp_719_9 <= 0;
      __tmp_719_10 <= 0;
      __tmp_719_11 <= 0;
      __tmp_719_12 <= 0;
      __tmp_721_1 <= 0;
      __tmp_721_2 <= 0;
      __tmp_721_3 <= 0;
      __tmp_721_4 <= 0;
      __tmp_721_5 <= 0;
      __tmp_721_6 <= 0;
      __tmp_721_7 <= 0;
      __tmp_721_8 <= 0;
      __tmp_721_9 <= 0;
      __tmp_721_10 <= 0;
      __tmp_721_11 <= 0;
      __tmp_721_12 <= 0;
      __tmp_723_1 <= 0;
      __tmp_723_2 <= 0;
      __tmp_723_3 <= 0;
      __tmp_723_4 <= 0;
      __tmp_723_5 <= 0;
      __tmp_723_6 <= 0;
      __tmp_723_7 <= 0;
      __tmp_723_8 <= 0;
      __tmp_723_9 <= 0;
      __tmp_723_10 <= 0;
      __tmp_723_11 <= 0;
      __tmp_723_12 <= 0;
      __tmp_725_1 <= 0;
      __tmp_725_2 <= 0;
      __tmp_725_3 <= 0;
      __tmp_725_4 <= 0;
      __tmp_725_5 <= 0;
      __tmp_725_6 <= 0;
      __tmp_725_7 <= 0;
      __tmp_725_8 <= 0;
      __tmp_725_9 <= 0;
      __tmp_725_10 <= 0;
      __tmp_725_11 <= 0;
      __tmp_725_12 <= 0;
      __tmp_727_1 <= 0;
      __tmp_727_2 <= 0;
      __tmp_727_3 <= 0;
      __tmp_727_4 <= 0;
      __tmp_727_5 <= 0;
      __tmp_727_6 <= 0;
      __tmp_727_7 <= 0;
      __tmp_727_8 <= 0;
      __tmp_727_9 <= 0;
      __tmp_727_10 <= 0;
      __tmp_727_11 <= 0;
      __tmp_727_12 <= 0;
      __tmp_729_1 <= 0;
      __tmp_729_2 <= 0;
      __tmp_729_3 <= 0;
      __tmp_729_4 <= 0;
      __tmp_729_5 <= 0;
      __tmp_729_6 <= 0;
      __tmp_729_7 <= 0;
      __tmp_729_8 <= 0;
      __tmp_729_9 <= 0;
      __tmp_729_10 <= 0;
      __tmp_729_11 <= 0;
      __tmp_729_12 <= 0;
      __tmp_731_1 <= 0;
      __tmp_731_2 <= 0;
      __tmp_731_3 <= 0;
      __tmp_731_4 <= 0;
      __tmp_731_5 <= 0;
      __tmp_731_6 <= 0;
      __tmp_731_7 <= 0;
      __tmp_731_8 <= 0;
      __tmp_731_9 <= 0;
      __tmp_731_10 <= 0;
      __tmp_731_11 <= 0;
      __tmp_731_12 <= 0;
      __tmp_733_1 <= 0;
      __tmp_733_2 <= 0;
      __tmp_733_3 <= 0;
      __tmp_733_4 <= 0;
      __tmp_733_5 <= 0;
      __tmp_733_6 <= 0;
      __tmp_733_7 <= 0;
      __tmp_733_8 <= 0;
      __tmp_733_9 <= 0;
      __tmp_733_10 <= 0;
      __tmp_733_11 <= 0;
      __tmp_733_12 <= 0;
      __tmp_735_1 <= 0;
      __tmp_735_2 <= 0;
      __tmp_735_3 <= 0;
      __tmp_735_4 <= 0;
      __tmp_735_5 <= 0;
      __tmp_735_6 <= 0;
      __tmp_735_7 <= 0;
      __tmp_735_8 <= 0;
      __tmp_735_9 <= 0;
      __tmp_735_10 <= 0;
      __tmp_735_11 <= 0;
      __tmp_735_12 <= 0;
      __tmp_737_1 <= 0;
      __tmp_737_2 <= 0;
      __tmp_737_3 <= 0;
      __tmp_737_4 <= 0;
      __tmp_737_5 <= 0;
      __tmp_737_6 <= 0;
      __tmp_737_7 <= 0;
      __tmp_737_8 <= 0;
      __tmp_737_9 <= 0;
      __tmp_737_10 <= 0;
      __tmp_737_11 <= 0;
      __tmp_737_12 <= 0;
      __tmp_739_1 <= 0;
      __tmp_739_2 <= 0;
      __tmp_739_3 <= 0;
      __tmp_739_4 <= 0;
      __tmp_739_5 <= 0;
      __tmp_739_6 <= 0;
      __tmp_739_7 <= 0;
      __tmp_739_8 <= 0;
      __tmp_739_9 <= 0;
      __tmp_739_10 <= 0;
      __tmp_739_11 <= 0;
      __tmp_739_12 <= 0;
      __tmp_741_1 <= 0;
      __tmp_741_2 <= 0;
      __tmp_741_3 <= 0;
      __tmp_741_4 <= 0;
      __tmp_741_5 <= 0;
      __tmp_741_6 <= 0;
      __tmp_741_7 <= 0;
      __tmp_741_8 <= 0;
      __tmp_741_9 <= 0;
      __tmp_741_10 <= 0;
      __tmp_741_11 <= 0;
      __tmp_741_12 <= 0;
      __tmp_743_1 <= 0;
      __tmp_743_2 <= 0;
      __tmp_743_3 <= 0;
      __tmp_743_4 <= 0;
      __tmp_743_5 <= 0;
      __tmp_743_6 <= 0;
      __tmp_743_7 <= 0;
      __tmp_743_8 <= 0;
      __tmp_743_9 <= 0;
      __tmp_743_10 <= 0;
      __tmp_743_11 <= 0;
      __tmp_743_12 <= 0;
      __tmp_745_1 <= 0;
      __tmp_745_2 <= 0;
      __tmp_745_3 <= 0;
      __tmp_745_4 <= 0;
      __tmp_745_5 <= 0;
      __tmp_745_6 <= 0;
      __tmp_745_7 <= 0;
      __tmp_745_8 <= 0;
      __tmp_745_9 <= 0;
      __tmp_745_10 <= 0;
      __tmp_745_11 <= 0;
      __tmp_745_12 <= 0;
      __tmp_747_1 <= 0;
      __tmp_747_2 <= 0;
      __tmp_747_3 <= 0;
      __tmp_747_4 <= 0;
      __tmp_747_5 <= 0;
      __tmp_747_6 <= 0;
      __tmp_747_7 <= 0;
      __tmp_747_8 <= 0;
      __tmp_747_9 <= 0;
      __tmp_747_10 <= 0;
      __tmp_747_11 <= 0;
      __tmp_747_12 <= 0;
      __tmp_749_1 <= 0;
      __tmp_749_2 <= 0;
      __tmp_749_3 <= 0;
      __tmp_749_4 <= 0;
      __tmp_749_5 <= 0;
      __tmp_749_6 <= 0;
      __tmp_749_7 <= 0;
      __tmp_749_8 <= 0;
      __tmp_749_9 <= 0;
      __tmp_749_10 <= 0;
      __tmp_749_11 <= 0;
      __tmp_749_12 <= 0;
      __tmp_751_1 <= 0;
      __tmp_751_2 <= 0;
      __tmp_751_3 <= 0;
      __tmp_751_4 <= 0;
      __tmp_751_5 <= 0;
      __tmp_751_6 <= 0;
      __tmp_751_7 <= 0;
      __tmp_751_8 <= 0;
      __tmp_751_9 <= 0;
      __tmp_751_10 <= 0;
      __tmp_751_11 <= 0;
      __tmp_751_12 <= 0;
      __tmp_753_1 <= 0;
      __tmp_753_2 <= 0;
      __tmp_753_3 <= 0;
      __tmp_753_4 <= 0;
      __tmp_753_5 <= 0;
      __tmp_753_6 <= 0;
      __tmp_753_7 <= 0;
      __tmp_753_8 <= 0;
      __tmp_753_9 <= 0;
      __tmp_753_10 <= 0;
      __tmp_753_11 <= 0;
      __tmp_753_12 <= 0;
      __tmp_755_1 <= 0;
      __tmp_755_2 <= 0;
      __tmp_755_3 <= 0;
      __tmp_755_4 <= 0;
      __tmp_755_5 <= 0;
      __tmp_755_6 <= 0;
      __tmp_755_7 <= 0;
      __tmp_755_8 <= 0;
      __tmp_755_9 <= 0;
      __tmp_755_10 <= 0;
      __tmp_755_11 <= 0;
      __tmp_755_12 <= 0;
      __tmp_757_1 <= 0;
      __tmp_757_2 <= 0;
      __tmp_757_3 <= 0;
      __tmp_757_4 <= 0;
      __tmp_757_5 <= 0;
      __tmp_757_6 <= 0;
      __tmp_757_7 <= 0;
      __tmp_757_8 <= 0;
      __tmp_757_9 <= 0;
      __tmp_757_10 <= 0;
      __tmp_757_11 <= 0;
      __tmp_757_12 <= 0;
      __tmp_759_1 <= 0;
      __tmp_759_2 <= 0;
      __tmp_759_3 <= 0;
      __tmp_759_4 <= 0;
      __tmp_759_5 <= 0;
      __tmp_759_6 <= 0;
      __tmp_759_7 <= 0;
      __tmp_759_8 <= 0;
      __tmp_759_9 <= 0;
      __tmp_759_10 <= 0;
      __tmp_759_11 <= 0;
      __tmp_759_12 <= 0;
      __tmp_761_1 <= 0;
      __tmp_761_2 <= 0;
      __tmp_761_3 <= 0;
      __tmp_761_4 <= 0;
      __tmp_761_5 <= 0;
      __tmp_761_6 <= 0;
      __tmp_761_7 <= 0;
      __tmp_761_8 <= 0;
      __tmp_761_9 <= 0;
      __tmp_761_10 <= 0;
      __tmp_761_11 <= 0;
      __tmp_761_12 <= 0;
      __tmp_763_1 <= 0;
      __tmp_763_2 <= 0;
      __tmp_763_3 <= 0;
      __tmp_763_4 <= 0;
      __tmp_763_5 <= 0;
      __tmp_763_6 <= 0;
      __tmp_763_7 <= 0;
      __tmp_763_8 <= 0;
      __tmp_763_9 <= 0;
      __tmp_763_10 <= 0;
      __tmp_763_11 <= 0;
      __tmp_763_12 <= 0;
      __tmp_765_1 <= 0;
      __tmp_765_2 <= 0;
      __tmp_765_3 <= 0;
      __tmp_765_4 <= 0;
      __tmp_765_5 <= 0;
      __tmp_765_6 <= 0;
      __tmp_765_7 <= 0;
      __tmp_765_8 <= 0;
      __tmp_765_9 <= 0;
      __tmp_765_10 <= 0;
      __tmp_765_11 <= 0;
      __tmp_765_12 <= 0;
      __tmp_767_1 <= 0;
      __tmp_767_2 <= 0;
      __tmp_767_3 <= 0;
      __tmp_767_4 <= 0;
      __tmp_767_5 <= 0;
      __tmp_767_6 <= 0;
      __tmp_767_7 <= 0;
      __tmp_767_8 <= 0;
      __tmp_767_9 <= 0;
      __tmp_767_10 <= 0;
      __tmp_767_11 <= 0;
      __tmp_767_12 <= 0;
      __tmp_769_1 <= 0;
      __tmp_769_2 <= 0;
      __tmp_769_3 <= 0;
      __tmp_769_4 <= 0;
      __tmp_769_5 <= 0;
      __tmp_769_6 <= 0;
      __tmp_769_7 <= 0;
      __tmp_769_8 <= 0;
      __tmp_769_9 <= 0;
      __tmp_769_10 <= 0;
      __tmp_769_11 <= 0;
      __tmp_769_12 <= 0;
      __tmp_769_13 <= 0;
      __tmp_769_14 <= 0;
      __tmp_769_15 <= 0;
      __tmp_769_16 <= 0;
      __tmp_769_17 <= 0;
      __tmp_769_18 <= 0;
      __tmp_769_19 <= 0;
      __tmp_769_20 <= 0;
      __tmp_769_21 <= 0;
      __tmp_769_22 <= 0;
      __tmp_771_1 <= 0;
      __tmp_771_2 <= 0;
      __tmp_771_3 <= 0;
      __tmp_771_4 <= 0;
      __tmp_771_5 <= 0;
      __tmp_771_6 <= 0;
      __tmp_771_7 <= 0;
      __tmp_771_8 <= 0;
      __tmp_771_9 <= 0;
      __tmp_771_10 <= 0;
      __tmp_771_11 <= 0;
      __tmp_771_12 <= 0;
      __tmp_771_13 <= 0;
      __tmp_771_14 <= 0;
      __tmp_771_15 <= 0;
      __tmp_771_16 <= 0;
      __tmp_771_17 <= 0;
      __tmp_771_18 <= 0;
      __tmp_771_19 <= 0;
      __tmp_771_20 <= 0;
      __tmp_771_21 <= 0;
      __tmp_771_22 <= 0;
      __tmp_773_1 <= 0;
      __tmp_773_2 <= 0;
      __tmp_773_3 <= 0;
      __tmp_773_4 <= 0;
      __tmp_773_5 <= 0;
      __tmp_773_6 <= 0;
      __tmp_773_7 <= 0;
      __tmp_773_8 <= 0;
      __tmp_773_9 <= 0;
      __tmp_773_10 <= 0;
      __tmp_773_11 <= 0;
      __tmp_773_12 <= 0;
      __tmp_773_13 <= 0;
      __tmp_773_14 <= 0;
      __tmp_773_15 <= 0;
      __tmp_773_16 <= 0;
      __tmp_773_17 <= 0;
      __tmp_773_18 <= 0;
      __tmp_773_19 <= 0;
      __tmp_773_20 <= 0;
      __tmp_773_21 <= 0;
      __tmp_773_22 <= 0;
      __tmp_775_1 <= 0;
      __tmp_775_2 <= 0;
      __tmp_775_3 <= 0;
      __tmp_775_4 <= 0;
      __tmp_775_5 <= 0;
      __tmp_775_6 <= 0;
      __tmp_775_7 <= 0;
      __tmp_775_8 <= 0;
      __tmp_775_9 <= 0;
      __tmp_775_10 <= 0;
      __tmp_775_11 <= 0;
      __tmp_775_12 <= 0;
      __tmp_775_13 <= 0;
      __tmp_775_14 <= 0;
      __tmp_775_15 <= 0;
      __tmp_775_16 <= 0;
      __tmp_775_17 <= 0;
      __tmp_775_18 <= 0;
      __tmp_775_19 <= 0;
      __tmp_775_20 <= 0;
      __tmp_775_21 <= 0;
      __tmp_775_22 <= 0;
      __tmp_777_1 <= 0;
      __tmp_777_2 <= 0;
      __tmp_777_3 <= 0;
      __tmp_777_4 <= 0;
      __tmp_777_5 <= 0;
      __tmp_777_6 <= 0;
      __tmp_777_7 <= 0;
      __tmp_777_8 <= 0;
      __tmp_777_9 <= 0;
      __tmp_777_10 <= 0;
      __tmp_777_11 <= 0;
      __tmp_777_12 <= 0;
      __tmp_777_13 <= 0;
      __tmp_777_14 <= 0;
      __tmp_777_15 <= 0;
      __tmp_777_16 <= 0;
      __tmp_777_17 <= 0;
      __tmp_777_18 <= 0;
      __tmp_777_19 <= 0;
      __tmp_777_20 <= 0;
      __tmp_777_21 <= 0;
      __tmp_777_22 <= 0;
      __tmp_779_1 <= 0;
      __tmp_779_2 <= 0;
      __tmp_779_3 <= 0;
      __tmp_779_4 <= 0;
      __tmp_779_5 <= 0;
      __tmp_779_6 <= 0;
      __tmp_779_7 <= 0;
      __tmp_779_8 <= 0;
      __tmp_779_9 <= 0;
      __tmp_779_10 <= 0;
      __tmp_779_11 <= 0;
      __tmp_779_12 <= 0;
      __tmp_779_13 <= 0;
      __tmp_779_14 <= 0;
      __tmp_779_15 <= 0;
      __tmp_779_16 <= 0;
      __tmp_779_17 <= 0;
      __tmp_779_18 <= 0;
      __tmp_779_19 <= 0;
      __tmp_779_20 <= 0;
      __tmp_779_21 <= 0;
      __tmp_779_22 <= 0;
      __tmp_781_1 <= 0;
      __tmp_781_2 <= 0;
      __tmp_781_3 <= 0;
      __tmp_781_4 <= 0;
      __tmp_781_5 <= 0;
      __tmp_781_6 <= 0;
      __tmp_781_7 <= 0;
      __tmp_781_8 <= 0;
      __tmp_781_9 <= 0;
      __tmp_781_10 <= 0;
      __tmp_781_11 <= 0;
      __tmp_781_12 <= 0;
      __tmp_781_13 <= 0;
      __tmp_781_14 <= 0;
      __tmp_781_15 <= 0;
      __tmp_781_16 <= 0;
      __tmp_781_17 <= 0;
      __tmp_781_18 <= 0;
      __tmp_781_19 <= 0;
      __tmp_781_20 <= 0;
      __tmp_781_21 <= 0;
      __tmp_781_22 <= 0;
      __tmp_783_1 <= 0;
      __tmp_783_2 <= 0;
      __tmp_783_3 <= 0;
      __tmp_783_4 <= 0;
      __tmp_783_5 <= 0;
      __tmp_783_6 <= 0;
      __tmp_783_7 <= 0;
      __tmp_783_8 <= 0;
      __tmp_783_9 <= 0;
      __tmp_783_10 <= 0;
      __tmp_783_11 <= 0;
      __tmp_783_12 <= 0;
      __tmp_783_13 <= 0;
      __tmp_783_14 <= 0;
      __tmp_783_15 <= 0;
      __tmp_783_16 <= 0;
      __tmp_783_17 <= 0;
      __tmp_783_18 <= 0;
      __tmp_783_19 <= 0;
      __tmp_783_20 <= 0;
      __tmp_783_21 <= 0;
      __tmp_783_22 <= 0;
      __tmp_785_1 <= 0;
      __tmp_785_2 <= 0;
      __tmp_785_3 <= 0;
      __tmp_785_4 <= 0;
      __tmp_785_5 <= 0;
      __tmp_785_6 <= 0;
      __tmp_785_7 <= 0;
      __tmp_785_8 <= 0;
      __tmp_785_9 <= 0;
      __tmp_785_10 <= 0;
      __tmp_785_11 <= 0;
      __tmp_785_12 <= 0;
      __tmp_785_13 <= 0;
      __tmp_785_14 <= 0;
      __tmp_785_15 <= 0;
      __tmp_785_16 <= 0;
      __tmp_785_17 <= 0;
      __tmp_785_18 <= 0;
      __tmp_785_19 <= 0;
      __tmp_785_20 <= 0;
      __tmp_785_21 <= 0;
      __tmp_785_22 <= 0;
      __tmp_787_1 <= 0;
      __tmp_787_2 <= 0;
      __tmp_787_3 <= 0;
      __tmp_787_4 <= 0;
      __tmp_787_5 <= 0;
      __tmp_787_6 <= 0;
      __tmp_787_7 <= 0;
      __tmp_787_8 <= 0;
      __tmp_787_9 <= 0;
      __tmp_787_10 <= 0;
      __tmp_787_11 <= 0;
      __tmp_787_12 <= 0;
      __tmp_787_13 <= 0;
      __tmp_787_14 <= 0;
      __tmp_787_15 <= 0;
      __tmp_787_16 <= 0;
      __tmp_787_17 <= 0;
      __tmp_787_18 <= 0;
      __tmp_787_19 <= 0;
      __tmp_787_20 <= 0;
      __tmp_787_21 <= 0;
      __tmp_787_22 <= 0;
      __tmp_787_23 <= 0;
      __tmp_787_24 <= 0;
      __tmp_787_25 <= 0;
      __tmp_787_26 <= 0;
      __tmp_787_27 <= 0;
      __tmp_787_28 <= 0;
      __tmp_789_1 <= 0;
      __tmp_789_2 <= 0;
      __tmp_789_3 <= 0;
      __tmp_789_4 <= 0;
      __tmp_789_5 <= 0;
      __tmp_789_6 <= 0;
      __tmp_789_7 <= 0;
      __tmp_789_8 <= 0;
      __tmp_789_9 <= 0;
      __tmp_789_10 <= 0;
      __tmp_789_11 <= 0;
      __tmp_789_12 <= 0;
      __tmp_789_13 <= 0;
      __tmp_789_14 <= 0;
      __tmp_789_15 <= 0;
      __tmp_789_16 <= 0;
      __tmp_789_17 <= 0;
      __tmp_789_18 <= 0;
      __tmp_789_19 <= 0;
      __tmp_789_20 <= 0;
      __tmp_789_21 <= 0;
      __tmp_789_22 <= 0;
      __tmp_789_23 <= 0;
      __tmp_789_24 <= 0;
      __tmp_789_25 <= 0;
      __tmp_789_26 <= 0;
      __tmp_791_1 <= 0;
      __tmp_791_2 <= 0;
      __tmp_791_3 <= 0;
      __tmp_791_4 <= 0;
      __tmp_791_5 <= 0;
      __tmp_791_6 <= 0;
      __tmp_791_7 <= 0;
      __tmp_791_8 <= 0;
      __tmp_791_9 <= 0;
      __tmp_791_10 <= 0;
      __tmp_791_11 <= 0;
      __tmp_791_12 <= 0;
      __tmp_791_13 <= 0;
      __tmp_791_14 <= 0;
      __tmp_791_15 <= 0;
      __tmp_791_16 <= 0;
      __tmp_791_17 <= 0;
      __tmp_791_18 <= 0;
      __tmp_791_19 <= 0;
      __tmp_791_20 <= 0;
      __tmp_791_21 <= 0;
      __tmp_791_22 <= 0;
      __tmp_791_23 <= 0;
      __tmp_791_24 <= 0;
      __tmp_791_25 <= 0;
      __tmp_791_26 <= 0;
      __tmp_793_1 <= 0;
      __tmp_793_2 <= 0;
      __tmp_793_3 <= 0;
      __tmp_793_4 <= 0;
      __tmp_793_5 <= 0;
      __tmp_793_6 <= 0;
      __tmp_793_7 <= 0;
      __tmp_793_8 <= 0;
      __tmp_793_9 <= 0;
      __tmp_793_10 <= 0;
      __tmp_793_11 <= 0;
      __tmp_793_12 <= 0;
      __tmp_793_13 <= 0;
      __tmp_793_14 <= 0;
      __tmp_793_15 <= 0;
      __tmp_793_16 <= 0;
      __tmp_793_17 <= 0;
      __tmp_793_18 <= 0;
      __tmp_793_19 <= 0;
      __tmp_793_20 <= 0;
      __tmp_793_21 <= 0;
      __tmp_793_22 <= 0;
      __tmp_793_23 <= 0;
      __tmp_793_24 <= 0;
      __tmp_793_25 <= 0;
      __tmp_793_26 <= 0;
      __tmp_795_1 <= 0;
      __tmp_795_2 <= 0;
      __tmp_795_3 <= 0;
      __tmp_795_4 <= 0;
      __tmp_795_5 <= 0;
      __tmp_795_6 <= 0;
      __tmp_795_7 <= 0;
      __tmp_795_8 <= 0;
      __tmp_795_9 <= 0;
      __tmp_795_10 <= 0;
      __tmp_795_11 <= 0;
      __tmp_795_12 <= 0;
      __tmp_795_13 <= 0;
      __tmp_795_14 <= 0;
      __tmp_795_15 <= 0;
      __tmp_795_16 <= 0;
      __tmp_795_17 <= 0;
      __tmp_795_18 <= 0;
      __tmp_795_19 <= 0;
      __tmp_795_20 <= 0;
      __tmp_795_21 <= 0;
      __tmp_795_22 <= 0;
      __tmp_795_23 <= 0;
      __tmp_795_24 <= 0;
      __tmp_795_25 <= 0;
      __tmp_795_26 <= 0;
      __tmp_795_27 <= 0;
      __tmp_795_28 <= 0;
      __tmp_795_29 <= 0;
      __tmp_795_30 <= 0;
      __tmp_795_31 <= 0;
      __tmp_795_32 <= 0;
      __tmp_795_33 <= 0;
      __tmp_795_34 <= 0;
      __tmp_797_1 <= 0;
      __tmp_797_2 <= 0;
      __tmp_797_3 <= 0;
      __tmp_797_4 <= 0;
      __tmp_797_5 <= 0;
      __tmp_797_6 <= 0;
      __tmp_797_7 <= 0;
      __tmp_797_8 <= 0;
      __tmp_797_9 <= 0;
      __tmp_797_10 <= 0;
      __tmp_797_11 <= 0;
      __tmp_797_12 <= 0;
      __tmp_797_13 <= 0;
      __tmp_797_14 <= 0;
      __tmp_797_15 <= 0;
      __tmp_797_16 <= 0;
      __tmp_797_17 <= 0;
      __tmp_797_18 <= 0;
      __tmp_797_19 <= 0;
      __tmp_797_20 <= 0;
      __tmp_797_21 <= 0;
      __tmp_797_22 <= 0;
      __tmp_797_23 <= 0;
      __tmp_797_24 <= 0;
      __tmp_797_25 <= 0;
      __tmp_797_26 <= 0;
      __tmp_797_27 <= 0;
      __tmp_797_28 <= 0;
      __tmp_797_29 <= 0;
      __tmp_797_30 <= 0;
      __tmp_797_31 <= 0;
      __tmp_797_32 <= 0;
      __tmp_797_33 <= 0;
      __tmp_797_34 <= 0;
      __tmp_799_1 <= 0;
      __tmp_799_2 <= 0;
      __tmp_799_3 <= 0;
      __tmp_799_4 <= 0;
      __tmp_799_5 <= 0;
      __tmp_799_6 <= 0;
      __tmp_799_7 <= 0;
      __tmp_799_8 <= 0;
      __tmp_799_9 <= 0;
      __tmp_799_10 <= 0;
      __tmp_799_11 <= 0;
      __tmp_799_12 <= 0;
      __tmp_799_13 <= 0;
      __tmp_799_14 <= 0;
      __tmp_799_15 <= 0;
      __tmp_799_16 <= 0;
      __tmp_799_17 <= 0;
      __tmp_799_18 <= 0;
      __tmp_799_19 <= 0;
      __tmp_799_20 <= 0;
      __tmp_799_21 <= 0;
      __tmp_799_22 <= 0;
      __tmp_799_23 <= 0;
      __tmp_799_24 <= 0;
      __tmp_799_25 <= 0;
      __tmp_799_26 <= 0;
      __tmp_799_27 <= 0;
      __tmp_799_28 <= 0;
      __tmp_799_29 <= 0;
      __tmp_799_30 <= 0;
      __tmp_799_31 <= 0;
      __tmp_799_32 <= 0;
      __tmp_799_33 <= 0;
      __tmp_799_34 <= 0;
      __tmp_801_1 <= 0;
      __tmp_803_1 <= 0;
      __tmp_803_2 <= 0;
      __tmp_803_3 <= 0;
      __tmp_803_4 <= 0;
      __tmp_803_5 <= 0;
      __tmp_803_6 <= 0;
      __tmp_803_7 <= 0;
      __tmp_803_8 <= 0;
      __tmp_803_9 <= 0;
      __tmp_805_1 <= 0;
      __tmp_805_2 <= 0;
      __tmp_805_3 <= 0;
      __tmp_805_4 <= 0;
      __tmp_805_5 <= 0;
      __tmp_805_6 <= 0;
      __tmp_805_7 <= 0;
      __tmp_805_8 <= 0;
      __tmp_805_9 <= 0;
      __tmp_807_1 <= 0;
      __tmp_807_2 <= 0;
      __tmp_807_3 <= 0;
      __tmp_807_4 <= 0;
      __tmp_807_5 <= 0;
      __tmp_807_6 <= 0;
      __tmp_807_7 <= 0;
      __tmp_807_8 <= 0;
      __tmp_807_9 <= 0;
      __tmp_815_1 <= 0;
      __tmp_815_2 <= 0;
      __tmp_815_3 <= 0;
      __tmp_815_4 <= 0;
      __tmp_815_5 <= 0;
      __tmp_815_6 <= 0;
      __tmp_815_7 <= 0;
      __tmp_815_8 <= 0;
      __tmp_815_9 <= 0;
      __tmp_817_1 <= 0;
      __tmp_817_2 <= 0;
      __tmp_817_3 <= 0;
      __tmp_817_4 <= 0;
      __tmp_817_5 <= 0;
      __tmp_817_6 <= 0;
      __tmp_817_7 <= 0;
      __tmp_817_8 <= 0;
      __tmp_817_9 <= 0;
      __tmp_819_1 <= 0;
      __tmp_819_2 <= 0;
      __tmp_819_3 <= 0;
      __tmp_819_4 <= 0;
      __tmp_819_5 <= 0;
      __tmp_819_6 <= 0;
      __tmp_819_7 <= 0;
      __tmp_819_8 <= 0;
      __tmp_819_9 <= 0;
      __tmp_827_1 <= 0;
      __tmp_827_2 <= 0;
      __tmp_827_3 <= 0;
      __tmp_827_4 <= 0;
      __tmp_827_5 <= 0;
      __tmp_827_6 <= 0;
      __tmp_827_7 <= 0;
      __tmp_827_8 <= 0;
      __tmp_827_9 <= 0;
      __tmp_829_1 <= 0;
      __tmp_829_2 <= 0;
      __tmp_829_3 <= 0;
      __tmp_829_4 <= 0;
      __tmp_829_5 <= 0;
      __tmp_829_6 <= 0;
      __tmp_829_7 <= 0;
      __tmp_829_8 <= 0;
      __tmp_829_9 <= 0;
      __tmp_831_1 <= 0;
      __tmp_831_2 <= 0;
      __tmp_831_3 <= 0;
      __tmp_831_4 <= 0;
      __tmp_831_5 <= 0;
      __tmp_831_6 <= 0;
      __tmp_831_7 <= 0;
      __tmp_831_8 <= 0;
      __tmp_831_9 <= 0;
      __tmp_839_1 <= 0;
      __tmp_839_2 <= 0;
      __tmp_839_3 <= 0;
      __tmp_839_4 <= 0;
      __tmp_839_5 <= 0;
      __tmp_839_6 <= 0;
      __tmp_839_7 <= 0;
      __tmp_839_8 <= 0;
      __tmp_839_9 <= 0;
      __tmp_841_1 <= 0;
      __tmp_841_2 <= 0;
      __tmp_841_3 <= 0;
      __tmp_841_4 <= 0;
      __tmp_841_5 <= 0;
      __tmp_841_6 <= 0;
      __tmp_841_7 <= 0;
      __tmp_841_8 <= 0;
      __tmp_841_9 <= 0;
      __tmp_843_1 <= 0;
      __tmp_843_2 <= 0;
      __tmp_843_3 <= 0;
      __tmp_843_4 <= 0;
      __tmp_843_5 <= 0;
      __tmp_843_6 <= 0;
      __tmp_843_7 <= 0;
      __tmp_843_8 <= 0;
      __tmp_843_9 <= 0;
      __tmp_851_1 <= 0;
      __tmp_851_2 <= 0;
      __tmp_851_3 <= 0;
      __tmp_851_4 <= 0;
      __tmp_851_5 <= 0;
      __tmp_851_6 <= 0;
      __tmp_851_7 <= 0;
      __tmp_851_8 <= 0;
      __tmp_851_9 <= 0;
      __tmp_853_1 <= 0;
      __tmp_853_2 <= 0;
      __tmp_853_3 <= 0;
      __tmp_853_4 <= 0;
      __tmp_853_5 <= 0;
      __tmp_853_6 <= 0;
      __tmp_853_7 <= 0;
      __tmp_853_8 <= 0;
      __tmp_853_9 <= 0;
      __tmp_855_1 <= 0;
      __tmp_855_2 <= 0;
      __tmp_855_3 <= 0;
      __tmp_855_4 <= 0;
      __tmp_855_5 <= 0;
      __tmp_855_6 <= 0;
      __tmp_855_7 <= 0;
      __tmp_855_8 <= 0;
      __tmp_855_9 <= 0;
      __tmp_863_1 <= 0;
      __tmp_863_2 <= 0;
      __tmp_863_3 <= 0;
      __tmp_863_4 <= 0;
      __tmp_863_5 <= 0;
      __tmp_863_6 <= 0;
      __tmp_863_7 <= 0;
      __tmp_863_8 <= 0;
      __tmp_863_9 <= 0;
      __tmp_865_1 <= 0;
      __tmp_865_2 <= 0;
      __tmp_865_3 <= 0;
      __tmp_865_4 <= 0;
      __tmp_865_5 <= 0;
      __tmp_865_6 <= 0;
      __tmp_865_7 <= 0;
      __tmp_865_8 <= 0;
      __tmp_865_9 <= 0;
      __tmp_867_1 <= 0;
      __tmp_867_2 <= 0;
      __tmp_867_3 <= 0;
      __tmp_867_4 <= 0;
      __tmp_867_5 <= 0;
      __tmp_867_6 <= 0;
      __tmp_867_7 <= 0;
      __tmp_867_8 <= 0;
      __tmp_867_9 <= 0;
      __tmp_875_1 <= 0;
      __tmp_875_2 <= 0;
      __tmp_875_3 <= 0;
      __tmp_875_4 <= 0;
      __tmp_875_5 <= 0;
      __tmp_875_6 <= 0;
      __tmp_875_7 <= 0;
      __tmp_875_8 <= 0;
      __tmp_875_9 <= 0;
      __tmp_877_1 <= 0;
      __tmp_877_2 <= 0;
      __tmp_877_3 <= 0;
      __tmp_877_4 <= 0;
      __tmp_877_5 <= 0;
      __tmp_877_6 <= 0;
      __tmp_877_7 <= 0;
      __tmp_877_8 <= 0;
      __tmp_877_9 <= 0;
      __tmp_879_1 <= 0;
      __tmp_879_2 <= 0;
      __tmp_879_3 <= 0;
      __tmp_879_4 <= 0;
      __tmp_879_5 <= 0;
      __tmp_879_6 <= 0;
      __tmp_879_7 <= 0;
      __tmp_879_8 <= 0;
      __tmp_879_9 <= 0;
      __tmp_887_1 <= 0;
      __tmp_887_2 <= 0;
      __tmp_887_3 <= 0;
      __tmp_887_4 <= 0;
      __tmp_887_5 <= 0;
      __tmp_887_6 <= 0;
      __tmp_887_7 <= 0;
      __tmp_887_8 <= 0;
      __tmp_887_9 <= 0;
      __tmp_889_1 <= 0;
      __tmp_889_2 <= 0;
      __tmp_889_3 <= 0;
      __tmp_889_4 <= 0;
      __tmp_889_5 <= 0;
      __tmp_889_6 <= 0;
      __tmp_889_7 <= 0;
      __tmp_889_8 <= 0;
      __tmp_889_9 <= 0;
      __tmp_891_1 <= 0;
      __tmp_891_2 <= 0;
      __tmp_891_3 <= 0;
      __tmp_891_4 <= 0;
      __tmp_891_5 <= 0;
      __tmp_891_6 <= 0;
      __tmp_891_7 <= 0;
      __tmp_891_8 <= 0;
      __tmp_891_9 <= 0;
      __tmp_899_1 <= 0;
      __tmp_899_2 <= 0;
      __tmp_899_3 <= 0;
      __tmp_899_4 <= 0;
      __tmp_899_5 <= 0;
      __tmp_899_6 <= 0;
      __tmp_899_7 <= 0;
      __tmp_899_8 <= 0;
      __tmp_899_9 <= 0;
      __tmp_901_1 <= 0;
      __tmp_901_2 <= 0;
      __tmp_901_3 <= 0;
      __tmp_901_4 <= 0;
      __tmp_901_5 <= 0;
      __tmp_901_6 <= 0;
      __tmp_901_7 <= 0;
      __tmp_901_8 <= 0;
      __tmp_901_9 <= 0;
      __tmp_903_1 <= 0;
      __tmp_903_2 <= 0;
      __tmp_903_3 <= 0;
      __tmp_903_4 <= 0;
      __tmp_903_5 <= 0;
      __tmp_903_6 <= 0;
      __tmp_903_7 <= 0;
      __tmp_903_8 <= 0;
      __tmp_903_9 <= 0;
      __tmp_911_1 <= 0;
      __tmp_911_2 <= 0;
      __tmp_911_3 <= 0;
      __tmp_911_4 <= 0;
      __tmp_911_5 <= 0;
      __tmp_911_6 <= 0;
      __tmp_911_7 <= 0;
      __tmp_911_8 <= 0;
      __tmp_911_9 <= 0;
      __tmp_911_10 <= 0;
      __tmp_911_11 <= 0;
      __tmp_911_12 <= 0;
      __tmp_911_13 <= 0;
      __tmp_911_14 <= 0;
      __tmp_911_15 <= 0;
      __tmp_911_16 <= 0;
      __tmp_911_17 <= 0;
      __tmp_911_18 <= 0;
      __tmp_911_19 <= 0;
      __tmp_913_1 <= 0;
      __tmp_913_2 <= 0;
      __tmp_913_3 <= 0;
      __tmp_913_4 <= 0;
      __tmp_913_5 <= 0;
      __tmp_913_6 <= 0;
      __tmp_913_7 <= 0;
      __tmp_913_8 <= 0;
      __tmp_913_9 <= 0;
      __tmp_913_10 <= 0;
      __tmp_913_11 <= 0;
      __tmp_913_12 <= 0;
      __tmp_913_13 <= 0;
      __tmp_913_14 <= 0;
      __tmp_913_15 <= 0;
      __tmp_913_16 <= 0;
      __tmp_913_17 <= 0;
      __tmp_913_18 <= 0;
      __tmp_913_19 <= 0;
      __tmp_915_1 <= 0;
      __tmp_915_2 <= 0;
      __tmp_915_3 <= 0;
      __tmp_915_4 <= 0;
      __tmp_915_5 <= 0;
      __tmp_915_6 <= 0;
      __tmp_915_7 <= 0;
      __tmp_915_8 <= 0;
      __tmp_915_9 <= 0;
      __tmp_915_10 <= 0;
      __tmp_915_11 <= 0;
      __tmp_915_12 <= 0;
      __tmp_915_13 <= 0;
      __tmp_915_14 <= 0;
      __tmp_915_15 <= 0;
      __tmp_915_16 <= 0;
      __tmp_915_17 <= 0;
      __tmp_915_18 <= 0;
      __tmp_915_19 <= 0;
      __tmp_917_1 <= 0;
      __tmp_917_2 <= 0;
      __tmp_917_3 <= 0;
      __tmp_917_4 <= 0;
      __tmp_917_5 <= 0;
      __tmp_917_6 <= 0;
      __tmp_917_7 <= 0;
      __tmp_917_8 <= 0;
      __tmp_917_9 <= 0;
      __tmp_917_10 <= 0;
      __tmp_917_11 <= 0;
      __tmp_917_12 <= 0;
      __tmp_917_13 <= 0;
      __tmp_917_14 <= 0;
      __tmp_917_15 <= 0;
      __tmp_917_16 <= 0;
      __tmp_917_17 <= 0;
      __tmp_917_18 <= 0;
      __tmp_917_19 <= 0;
      __tmp_919_1 <= 0;
      __tmp_919_2 <= 0;
      __tmp_919_3 <= 0;
      __tmp_919_4 <= 0;
      __tmp_919_5 <= 0;
      __tmp_919_6 <= 0;
      __tmp_919_7 <= 0;
      __tmp_919_8 <= 0;
      __tmp_919_9 <= 0;
      __tmp_919_10 <= 0;
      __tmp_919_11 <= 0;
      __tmp_919_12 <= 0;
      __tmp_919_13 <= 0;
      __tmp_919_14 <= 0;
      __tmp_919_15 <= 0;
      __tmp_919_16 <= 0;
      __tmp_919_17 <= 0;
      __tmp_919_18 <= 0;
      __tmp_919_19 <= 0;
      __tmp_921_1 <= 0;
      __tmp_921_2 <= 0;
      __tmp_921_3 <= 0;
      __tmp_921_4 <= 0;
      __tmp_921_5 <= 0;
      __tmp_921_6 <= 0;
      __tmp_921_7 <= 0;
      __tmp_921_8 <= 0;
      __tmp_921_9 <= 0;
      __tmp_921_10 <= 0;
      __tmp_921_11 <= 0;
      __tmp_921_12 <= 0;
      __tmp_921_13 <= 0;
      __tmp_921_14 <= 0;
      __tmp_921_15 <= 0;
      __tmp_921_16 <= 0;
      __tmp_921_17 <= 0;
      __tmp_921_18 <= 0;
      __tmp_921_19 <= 0;
      __tmp_923_1 <= 0;
      __tmp_923_2 <= 0;
      __tmp_923_3 <= 0;
      __tmp_923_4 <= 0;
      __tmp_923_5 <= 0;
      __tmp_923_6 <= 0;
      __tmp_923_7 <= 0;
      __tmp_923_8 <= 0;
      __tmp_923_9 <= 0;
      __tmp_923_10 <= 0;
      __tmp_923_11 <= 0;
      __tmp_923_12 <= 0;
      __tmp_923_13 <= 0;
      __tmp_923_14 <= 0;
      __tmp_923_15 <= 0;
      __tmp_923_16 <= 0;
      __tmp_923_17 <= 0;
      __tmp_923_18 <= 0;
      __tmp_923_19 <= 0;
      __tmp_925_1 <= 0;
      __tmp_925_2 <= 0;
      __tmp_925_3 <= 0;
      __tmp_925_4 <= 0;
      __tmp_925_5 <= 0;
      __tmp_925_6 <= 0;
      __tmp_925_7 <= 0;
      __tmp_925_8 <= 0;
      __tmp_925_9 <= 0;
      __tmp_925_10 <= 0;
      __tmp_925_11 <= 0;
      __tmp_925_12 <= 0;
      __tmp_925_13 <= 0;
      __tmp_925_14 <= 0;
      __tmp_925_15 <= 0;
      __tmp_925_16 <= 0;
      __tmp_925_17 <= 0;
      __tmp_925_18 <= 0;
      __tmp_925_19 <= 0;
      __tmp_927_1 <= 0;
      __tmp_927_2 <= 0;
      __tmp_927_3 <= 0;
      __tmp_927_4 <= 0;
      __tmp_927_5 <= 0;
      __tmp_927_6 <= 0;
      __tmp_927_7 <= 0;
      __tmp_927_8 <= 0;
      __tmp_927_9 <= 0;
      __tmp_927_10 <= 0;
      __tmp_927_11 <= 0;
      __tmp_927_12 <= 0;
      __tmp_927_13 <= 0;
      __tmp_927_14 <= 0;
      __tmp_927_15 <= 0;
      __tmp_927_16 <= 0;
      __tmp_927_17 <= 0;
      __tmp_927_18 <= 0;
      __tmp_927_19 <= 0;
      __tmp_935_1 <= 0;
      __tmp_935_2 <= 0;
      __tmp_935_3 <= 0;
      __tmp_935_4 <= 0;
      __tmp_935_5 <= 0;
      __tmp_935_6 <= 0;
      __tmp_935_7 <= 0;
      __tmp_935_8 <= 0;
      __tmp_935_9 <= 0;
      __tmp_935_10 <= 0;
      __tmp_935_11 <= 0;
      __tmp_935_12 <= 0;
      __tmp_935_13 <= 0;
      __tmp_935_14 <= 0;
      __tmp_935_15 <= 0;
      __tmp_935_16 <= 0;
      __tmp_935_17 <= 0;
      __tmp_935_18 <= 0;
      __tmp_935_19 <= 0;
      __tmp_935_20 <= 0;
      __tmp_935_21 <= 0;
      __tmp_935_22 <= 0;
      __tmp_935_23 <= 0;
      __tmp_935_24 <= 0;
      __tmp_937_1 <= 0;
      __tmp_937_2 <= 0;
      __tmp_937_3 <= 0;
      __tmp_937_4 <= 0;
      __tmp_937_5 <= 0;
      __tmp_937_6 <= 0;
      __tmp_937_7 <= 0;
      __tmp_937_8 <= 0;
      __tmp_937_9 <= 0;
      __tmp_937_10 <= 0;
      __tmp_937_11 <= 0;
      __tmp_937_12 <= 0;
      __tmp_937_13 <= 0;
      __tmp_937_14 <= 0;
      __tmp_937_15 <= 0;
      __tmp_937_16 <= 0;
      __tmp_937_17 <= 0;
      __tmp_937_18 <= 0;
      __tmp_937_19 <= 0;
      __tmp_937_20 <= 0;
      __tmp_937_21 <= 0;
      __tmp_937_22 <= 0;
      __tmp_937_23 <= 0;
      __tmp_939_1 <= 0;
      __tmp_939_2 <= 0;
      __tmp_939_3 <= 0;
      __tmp_939_4 <= 0;
      __tmp_939_5 <= 0;
      __tmp_939_6 <= 0;
      __tmp_939_7 <= 0;
      __tmp_939_8 <= 0;
      __tmp_939_9 <= 0;
      __tmp_939_10 <= 0;
      __tmp_939_11 <= 0;
      __tmp_939_12 <= 0;
      __tmp_939_13 <= 0;
      __tmp_939_14 <= 0;
      __tmp_939_15 <= 0;
      __tmp_939_16 <= 0;
      __tmp_939_17 <= 0;
      __tmp_939_18 <= 0;
      __tmp_939_19 <= 0;
      __tmp_939_20 <= 0;
      __tmp_939_21 <= 0;
      __tmp_939_22 <= 0;
      __tmp_939_23 <= 0;
      __tmp_941_1 <= 0;
      __tmp_941_2 <= 0;
      __tmp_941_3 <= 0;
      __tmp_941_4 <= 0;
      __tmp_941_5 <= 0;
      __tmp_941_6 <= 0;
      __tmp_941_7 <= 0;
      __tmp_941_8 <= 0;
      __tmp_941_9 <= 0;
      __tmp_941_10 <= 0;
      __tmp_941_11 <= 0;
      __tmp_941_12 <= 0;
      __tmp_941_13 <= 0;
      __tmp_941_14 <= 0;
      __tmp_941_15 <= 0;
      __tmp_941_16 <= 0;
      __tmp_941_17 <= 0;
      __tmp_941_18 <= 0;
      __tmp_941_19 <= 0;
      __tmp_941_20 <= 0;
      __tmp_941_21 <= 0;
      __tmp_941_22 <= 0;
      __tmp_941_23 <= 0;
      __tmp_949_1 <= 0;
      __tmp_949_2 <= 0;
      __tmp_949_3 <= 0;
      __tmp_949_4 <= 0;
      __tmp_949_5 <= 0;
      __tmp_949_6 <= 0;
      __tmp_949_7 <= 0;
      __tmp_949_8 <= 0;
      __tmp_949_9 <= 0;
      __tmp_949_10 <= 0;
      __tmp_949_11 <= 0;
      __tmp_949_12 <= 0;
      __tmp_949_13 <= 0;
      __tmp_949_14 <= 0;
      __tmp_949_15 <= 0;
      __tmp_949_16 <= 0;
      __tmp_949_17 <= 0;
      __tmp_949_18 <= 0;
      __tmp_949_19 <= 0;
      __tmp_949_20 <= 0;
      __tmp_949_21 <= 0;
      __tmp_949_22 <= 0;
      __tmp_949_23 <= 0;
      __tmp_949_24 <= 0;
      __tmp_949_25 <= 0;
      __tmp_949_26 <= 0;
      __tmp_949_27 <= 0;
      __tmp_949_28 <= 0;
      __tmp_949_29 <= 0;
      __tmp_949_30 <= 0;
      __tmp_949_31 <= 0;
      __tmp_951_1 <= 0;
      __tmp_951_2 <= 0;
      __tmp_951_3 <= 0;
      __tmp_951_4 <= 0;
      __tmp_951_5 <= 0;
      __tmp_951_6 <= 0;
      __tmp_951_7 <= 0;
      __tmp_951_8 <= 0;
      __tmp_951_9 <= 0;
      __tmp_951_10 <= 0;
      __tmp_951_11 <= 0;
      __tmp_951_12 <= 0;
      __tmp_951_13 <= 0;
      __tmp_951_14 <= 0;
      __tmp_951_15 <= 0;
      __tmp_951_16 <= 0;
      __tmp_951_17 <= 0;
      __tmp_951_18 <= 0;
      __tmp_951_19 <= 0;
      __tmp_951_20 <= 0;
      __tmp_951_21 <= 0;
      __tmp_951_22 <= 0;
      __tmp_951_23 <= 0;
      __tmp_951_24 <= 0;
      __tmp_951_25 <= 0;
      __tmp_951_26 <= 0;
      __tmp_951_27 <= 0;
      __tmp_951_28 <= 0;
      __tmp_951_29 <= 0;
      __tmp_951_30 <= 0;
      __tmp_951_31 <= 0;
      __tmp_953_1 <= 0;
      __tmp_953_2 <= 0;
      __tmp_953_3 <= 0;
      __tmp_953_4 <= 0;
      __tmp_953_5 <= 0;
      __tmp_953_6 <= 0;
      __tmp_953_7 <= 0;
      __tmp_953_8 <= 0;
      __tmp_953_9 <= 0;
      __tmp_953_10 <= 0;
      __tmp_953_11 <= 0;
      __tmp_953_12 <= 0;
      __tmp_953_13 <= 0;
      __tmp_953_14 <= 0;
      __tmp_953_15 <= 0;
      __tmp_953_16 <= 0;
      __tmp_953_17 <= 0;
      __tmp_953_18 <= 0;
      __tmp_953_19 <= 0;
      __tmp_953_20 <= 0;
      __tmp_953_21 <= 0;
      __tmp_953_22 <= 0;
      __tmp_953_23 <= 0;
      __tmp_953_24 <= 0;
      __tmp_953_25 <= 0;
      __tmp_953_26 <= 0;
      __tmp_953_27 <= 0;
      __tmp_953_28 <= 0;
      __tmp_953_29 <= 0;
      __tmp_953_30 <= 0;
      __tmp_953_31 <= 0;
      __tmp_961_1 <= 0;
      __tmp_961_2 <= 0;
      __tmp_961_3 <= 0;
      __tmp_961_4 <= 0;
      __tmp_961_5 <= 0;
      __tmp_961_6 <= 0;
      __tmp_961_7 <= 0;
      __tmp_961_8 <= 0;
      __tmp_961_9 <= 0;
      __tmp_961_10 <= 0;
      __tmp_961_11 <= 0;
      __tmp_961_12 <= 0;
      __tmp_961_13 <= 0;
      __tmp_961_14 <= 0;
      __tmp_961_15 <= 0;
      __tmp_961_16 <= 0;
      __tmp_961_17 <= 0;
      __tmp_961_18 <= 0;
      __tmp_961_19 <= 0;
      __tmp_961_20 <= 0;
      __tmp_961_21 <= 0;
      __tmp_961_22 <= 0;
      __tmp_961_23 <= 0;
      __tmp_961_24 <= 0;
      __tmp_961_25 <= 0;
      __tmp_961_26 <= 0;
      __tmp_961_27 <= 0;
      __tmp_961_28 <= 0;
      __tmp_961_29 <= 0;
      __tmp_961_30 <= 0;
      __tmp_961_31 <= 0;
      __tmp_961_32 <= 0;
      __tmp_961_33 <= 0;
      __tmp_961_34 <= 0;
      __tmp_961_35 <= 0;
      __tmp_961_36 <= 0;
      __tmp_961_37 <= 0;
      __tmp_961_38 <= 0;
      __tmp_961_39 <= 0;
      __tmp_961_40 <= 0;
      __tmp_961_41 <= 0;
      __tmp_961_42 <= 0;
      __tmp_961_43 <= 0;
      __tmp_961_44 <= 0;
      __tmp_961_45 <= 0;
      __tmp_961_46 <= 0;
      __tmp_963_1 <= 0;
      __tmp_963_2 <= 0;
      __tmp_963_3 <= 0;
      __tmp_963_4 <= 0;
      __tmp_963_5 <= 0;
      __tmp_963_6 <= 0;
      __tmp_963_7 <= 0;
      __tmp_963_8 <= 0;
      __tmp_963_9 <= 0;
      __tmp_963_10 <= 0;
      __tmp_963_11 <= 0;
      __tmp_963_12 <= 0;
      __tmp_963_13 <= 0;
      __tmp_963_14 <= 0;
      __tmp_963_15 <= 0;
      __tmp_963_16 <= 0;
      __tmp_963_17 <= 0;
      __tmp_963_18 <= 0;
      __tmp_963_19 <= 0;
      __tmp_963_20 <= 0;
      __tmp_963_21 <= 0;
      __tmp_963_22 <= 0;
      __tmp_963_23 <= 0;
      __tmp_963_24 <= 0;
      __tmp_963_25 <= 0;
      __tmp_963_26 <= 0;
      __tmp_963_27 <= 0;
      __tmp_963_28 <= 0;
      __tmp_963_29 <= 0;
      __tmp_963_30 <= 0;
      __tmp_963_31 <= 0;
      __tmp_963_32 <= 0;
      __tmp_963_33 <= 0;
      __tmp_963_34 <= 0;
      __tmp_963_35 <= 0;
      __tmp_963_36 <= 0;
      __tmp_963_37 <= 0;
      __tmp_963_38 <= 0;
      __tmp_963_39 <= 0;
      __tmp_963_40 <= 0;
      __tmp_963_41 <= 0;
      __tmp_963_42 <= 0;
      __tmp_963_43 <= 0;
      __tmp_963_44 <= 0;
      __tmp_963_45 <= 0;
      __tmp_963_46 <= 0;
      __tmp_965_1 <= 0;
      __tmp_965_2 <= 0;
      __tmp_965_3 <= 0;
      __tmp_965_4 <= 0;
      __tmp_965_5 <= 0;
      __tmp_965_6 <= 0;
      __tmp_965_7 <= 0;
      __tmp_965_8 <= 0;
      __tmp_965_9 <= 0;
      __tmp_965_10 <= 0;
      __tmp_965_11 <= 0;
      __tmp_965_12 <= 0;
      __tmp_965_13 <= 0;
      __tmp_965_14 <= 0;
      __tmp_965_15 <= 0;
      __tmp_965_16 <= 0;
      __tmp_965_17 <= 0;
      __tmp_965_18 <= 0;
      __tmp_965_19 <= 0;
      __tmp_965_20 <= 0;
      __tmp_965_21 <= 0;
      __tmp_965_22 <= 0;
      __tmp_965_23 <= 0;
      __tmp_965_24 <= 0;
      __tmp_965_25 <= 0;
      __tmp_965_26 <= 0;
      __tmp_965_27 <= 0;
      __tmp_965_28 <= 0;
      __tmp_965_29 <= 0;
      __tmp_965_30 <= 0;
      __tmp_965_31 <= 0;
      __tmp_965_32 <= 0;
      __tmp_965_33 <= 0;
      __tmp_965_34 <= 0;
      __tmp_965_35 <= 0;
      __tmp_965_36 <= 0;
      __tmp_965_37 <= 0;
      __tmp_965_38 <= 0;
      __tmp_965_39 <= 0;
      __tmp_965_40 <= 0;
      __tmp_965_41 <= 0;
      __tmp_965_42 <= 0;
      __tmp_965_43 <= 0;
      __tmp_965_44 <= 0;
      __tmp_965_45 <= 0;
      __tmp_965_46 <= 0;
      __tmp_967_1 <= 0;
      __tmp_967_2 <= 0;
      __tmp_967_3 <= 0;
      __tmp_967_4 <= 0;
      __tmp_967_5 <= 0;
      __tmp_967_6 <= 0;
      __tmp_967_7 <= 0;
      __tmp_967_8 <= 0;
      __tmp_967_9 <= 0;
      __tmp_967_10 <= 0;
      __tmp_967_11 <= 0;
      __tmp_967_12 <= 0;
      __tmp_967_13 <= 0;
      __tmp_967_14 <= 0;
      __tmp_967_15 <= 0;
      __tmp_967_16 <= 0;
      __tmp_967_17 <= 0;
      __tmp_967_18 <= 0;
      __tmp_967_19 <= 0;
      __tmp_967_20 <= 0;
      __tmp_967_21 <= 0;
      __tmp_967_22 <= 0;
      __tmp_967_23 <= 0;
      __tmp_967_24 <= 0;
      __tmp_967_25 <= 0;
      __tmp_967_26 <= 0;
      __tmp_967_27 <= 0;
      __tmp_967_28 <= 0;
      __tmp_967_29 <= 0;
      __tmp_967_30 <= 0;
      __tmp_967_31 <= 0;
      __tmp_967_32 <= 0;
      __tmp_967_33 <= 0;
      __tmp_967_34 <= 0;
      __tmp_967_35 <= 0;
      __tmp_967_36 <= 0;
      __tmp_967_37 <= 0;
      __tmp_967_38 <= 0;
      __tmp_967_39 <= 0;
      __tmp_967_40 <= 0;
      __tmp_967_41 <= 0;
      __tmp_967_42 <= 0;
      __tmp_967_43 <= 0;
      __tmp_967_44 <= 0;
      __tmp_967_45 <= 0;
      __tmp_967_46 <= 0;
      __tmp_969_1 <= 0;
      __tmp_969_2 <= 0;
      __tmp_969_3 <= 0;
      __tmp_969_4 <= 0;
      __tmp_969_5 <= 0;
      __tmp_969_6 <= 0;
      __tmp_969_7 <= 0;
      __tmp_969_8 <= 0;
      __tmp_969_9 <= 0;
      __tmp_969_10 <= 0;
      __tmp_969_11 <= 0;
      __tmp_969_12 <= 0;
      __tmp_969_13 <= 0;
      __tmp_969_14 <= 0;
      __tmp_969_15 <= 0;
      __tmp_969_16 <= 0;
      __tmp_969_17 <= 0;
      __tmp_969_18 <= 0;
      __tmp_969_19 <= 0;
      __tmp_969_20 <= 0;
      __tmp_969_21 <= 0;
      __tmp_969_22 <= 0;
      __tmp_969_23 <= 0;
      __tmp_969_24 <= 0;
      __tmp_969_25 <= 0;
      __tmp_969_26 <= 0;
      __tmp_969_27 <= 0;
      __tmp_969_28 <= 0;
      __tmp_969_29 <= 0;
      __tmp_969_30 <= 0;
      __tmp_969_31 <= 0;
      __tmp_969_32 <= 0;
      __tmp_969_33 <= 0;
      __tmp_969_34 <= 0;
      __tmp_969_35 <= 0;
      __tmp_969_36 <= 0;
      __tmp_969_37 <= 0;
      __tmp_969_38 <= 0;
      __tmp_969_39 <= 0;
      __tmp_969_40 <= 0;
      __tmp_969_41 <= 0;
      __tmp_969_42 <= 0;
    end else begin
      if(__stream_seq_14_cond_2_45) begin
        _stream_conv2d_16_sink_37_sink_mode <= 3'b1;
        _stream_conv2d_16_sink_37_sink_offset <= __stream_conv2d_16_sink_37_sink_offset_0_45;
        _stream_conv2d_16_sink_37_sink_size <= __stream_conv2d_16_sink_37_sink_size_1_45;
        _stream_conv2d_16_sink_37_sink_stride <= 1;
      end 
      __stream_conv2d_16_sink_37_sink_offset_0_45 <= __stream_conv2d_16_sink_37_sink_offset_0_44;
      __stream_conv2d_16_sink_37_sink_size_1_45 <= __stream_conv2d_16_sink_37_sink_size_1_44;
      __stream_seq_14_cond_2_45 <= __stream_seq_14_cond_2_44;
      __stream_conv2d_16_sink_37_sink_offset_0_44 <= __stream_conv2d_16_sink_37_sink_offset_0_43;
      __stream_conv2d_16_sink_37_sink_size_1_44 <= __stream_conv2d_16_sink_37_sink_size_1_43;
      __stream_seq_14_cond_2_44 <= __stream_seq_14_cond_2_43;
      __stream_conv2d_16_sink_37_sink_offset_0_43 <= __stream_conv2d_16_sink_37_sink_offset_0_42;
      __stream_conv2d_16_sink_37_sink_size_1_43 <= __stream_conv2d_16_sink_37_sink_size_1_42;
      __stream_seq_14_cond_2_43 <= __stream_seq_14_cond_2_42;
      __stream_conv2d_16_sink_37_sink_offset_0_42 <= __stream_conv2d_16_sink_37_sink_offset_0_41;
      __stream_conv2d_16_sink_37_sink_size_1_42 <= __stream_conv2d_16_sink_37_sink_size_1_41;
      __stream_seq_14_cond_2_42 <= __stream_seq_14_cond_2_41;
      __stream_conv2d_16_sink_37_sink_offset_0_41 <= __stream_conv2d_16_sink_37_sink_offset_0_40;
      __stream_conv2d_16_sink_37_sink_size_1_41 <= __stream_conv2d_16_sink_37_sink_size_1_40;
      __stream_seq_14_cond_2_41 <= __stream_seq_14_cond_2_40;
      __stream_conv2d_16_sink_37_sink_offset_0_40 <= __stream_conv2d_16_sink_37_sink_offset_0_39;
      __stream_conv2d_16_sink_37_sink_size_1_40 <= __stream_conv2d_16_sink_37_sink_size_1_39;
      __stream_seq_14_cond_2_40 <= __stream_seq_14_cond_2_39;
      __stream_conv2d_16_sink_37_sink_offset_0_39 <= __stream_conv2d_16_sink_37_sink_offset_0_38;
      __stream_conv2d_16_sink_37_sink_size_1_39 <= __stream_conv2d_16_sink_37_sink_size_1_38;
      __stream_seq_14_cond_2_39 <= __stream_seq_14_cond_2_38;
      __stream_conv2d_16_sink_37_sink_offset_0_38 <= __stream_conv2d_16_sink_37_sink_offset_0_37;
      __stream_conv2d_16_sink_37_sink_size_1_38 <= __stream_conv2d_16_sink_37_sink_size_1_37;
      __stream_seq_14_cond_2_38 <= __stream_seq_14_cond_2_37;
      __stream_conv2d_16_sink_37_sink_offset_0_37 <= __stream_conv2d_16_sink_37_sink_offset_0_36;
      __stream_conv2d_16_sink_37_sink_size_1_37 <= __stream_conv2d_16_sink_37_sink_size_1_36;
      __stream_seq_14_cond_2_37 <= __stream_seq_14_cond_2_36;
      __stream_conv2d_16_sink_37_sink_offset_0_36 <= __stream_conv2d_16_sink_37_sink_offset_0_35;
      __stream_conv2d_16_sink_37_sink_size_1_36 <= __stream_conv2d_16_sink_37_sink_size_1_35;
      __stream_seq_14_cond_2_36 <= __stream_seq_14_cond_2_35;
      __stream_conv2d_16_sink_37_sink_offset_0_35 <= __stream_conv2d_16_sink_37_sink_offset_0_34;
      __stream_conv2d_16_sink_37_sink_size_1_35 <= __stream_conv2d_16_sink_37_sink_size_1_34;
      __stream_seq_14_cond_2_35 <= __stream_seq_14_cond_2_34;
      __stream_conv2d_16_sink_37_sink_offset_0_34 <= __stream_conv2d_16_sink_37_sink_offset_0_33;
      __stream_conv2d_16_sink_37_sink_size_1_34 <= __stream_conv2d_16_sink_37_sink_size_1_33;
      __stream_seq_14_cond_2_34 <= __stream_seq_14_cond_2_33;
      __stream_conv2d_16_sink_37_sink_offset_0_33 <= __stream_conv2d_16_sink_37_sink_offset_0_32;
      __stream_conv2d_16_sink_37_sink_size_1_33 <= __stream_conv2d_16_sink_37_sink_size_1_32;
      __stream_seq_14_cond_2_33 <= __stream_seq_14_cond_2_32;
      __stream_conv2d_16_sink_37_sink_offset_0_32 <= __stream_conv2d_16_sink_37_sink_offset_0_31;
      __stream_conv2d_16_sink_37_sink_size_1_32 <= __stream_conv2d_16_sink_37_sink_size_1_31;
      __stream_seq_14_cond_2_32 <= __stream_seq_14_cond_2_31;
      __stream_conv2d_16_sink_37_sink_offset_0_31 <= __stream_conv2d_16_sink_37_sink_offset_0_30;
      __stream_conv2d_16_sink_37_sink_size_1_31 <= __stream_conv2d_16_sink_37_sink_size_1_30;
      __stream_seq_14_cond_2_31 <= __stream_seq_14_cond_2_30;
      __stream_conv2d_16_sink_37_sink_offset_0_30 <= __stream_conv2d_16_sink_37_sink_offset_0_29;
      __stream_conv2d_16_sink_37_sink_size_1_30 <= __stream_conv2d_16_sink_37_sink_size_1_29;
      __stream_seq_14_cond_2_30 <= __stream_seq_14_cond_2_29;
      __stream_conv2d_16_sink_37_sink_offset_0_29 <= __stream_conv2d_16_sink_37_sink_offset_0_28;
      __stream_conv2d_16_sink_37_sink_size_1_29 <= __stream_conv2d_16_sink_37_sink_size_1_28;
      __stream_seq_14_cond_2_29 <= __stream_seq_14_cond_2_28;
      __stream_conv2d_16_sink_37_sink_offset_0_28 <= __stream_conv2d_16_sink_37_sink_offset_0_27;
      __stream_conv2d_16_sink_37_sink_size_1_28 <= __stream_conv2d_16_sink_37_sink_size_1_27;
      __stream_seq_14_cond_2_28 <= __stream_seq_14_cond_2_27;
      __stream_conv2d_16_sink_37_sink_offset_0_27 <= __stream_conv2d_16_sink_37_sink_offset_0_26;
      __stream_conv2d_16_sink_37_sink_size_1_27 <= __stream_conv2d_16_sink_37_sink_size_1_26;
      __stream_seq_14_cond_2_27 <= __stream_seq_14_cond_2_26;
      __stream_conv2d_16_sink_37_sink_offset_0_26 <= __stream_conv2d_16_sink_37_sink_offset_0_25;
      __stream_conv2d_16_sink_37_sink_size_1_26 <= __stream_conv2d_16_sink_37_sink_size_1_25;
      __stream_seq_14_cond_2_26 <= __stream_seq_14_cond_2_25;
      __stream_conv2d_16_sink_37_sink_offset_0_25 <= __stream_conv2d_16_sink_37_sink_offset_0_24;
      __stream_conv2d_16_sink_37_sink_size_1_25 <= __stream_conv2d_16_sink_37_sink_size_1_24;
      __stream_seq_14_cond_2_25 <= __stream_seq_14_cond_2_24;
      __stream_conv2d_16_sink_37_sink_offset_0_24 <= __stream_conv2d_16_sink_37_sink_offset_0_23;
      __stream_conv2d_16_sink_37_sink_size_1_24 <= __stream_conv2d_16_sink_37_sink_size_1_23;
      __stream_seq_14_cond_2_24 <= __stream_seq_14_cond_2_23;
      __stream_conv2d_16_sink_37_sink_offset_0_23 <= __stream_conv2d_16_sink_37_sink_offset_0_22;
      __stream_conv2d_16_sink_37_sink_size_1_23 <= __stream_conv2d_16_sink_37_sink_size_1_22;
      __stream_seq_14_cond_2_23 <= __stream_seq_14_cond_2_22;
      __stream_conv2d_16_sink_37_sink_offset_0_22 <= __stream_conv2d_16_sink_37_sink_offset_0_21;
      __stream_conv2d_16_sink_37_sink_size_1_22 <= __stream_conv2d_16_sink_37_sink_size_1_21;
      __stream_seq_14_cond_2_22 <= __stream_seq_14_cond_2_21;
      __stream_conv2d_16_sink_37_sink_offset_0_21 <= __stream_conv2d_16_sink_37_sink_offset_0_20;
      __stream_conv2d_16_sink_37_sink_size_1_21 <= __stream_conv2d_16_sink_37_sink_size_1_20;
      __stream_seq_14_cond_2_21 <= __stream_seq_14_cond_2_20;
      __stream_conv2d_16_sink_37_sink_offset_0_20 <= __stream_conv2d_16_sink_37_sink_offset_0_19;
      __stream_conv2d_16_sink_37_sink_size_1_20 <= __stream_conv2d_16_sink_37_sink_size_1_19;
      __stream_seq_14_cond_2_20 <= __stream_seq_14_cond_2_19;
      __stream_conv2d_16_sink_37_sink_offset_0_19 <= __stream_conv2d_16_sink_37_sink_offset_0_18;
      __stream_conv2d_16_sink_37_sink_size_1_19 <= __stream_conv2d_16_sink_37_sink_size_1_18;
      __stream_seq_14_cond_2_19 <= __stream_seq_14_cond_2_18;
      __stream_conv2d_16_sink_37_sink_offset_0_18 <= __stream_conv2d_16_sink_37_sink_offset_0_17;
      __stream_conv2d_16_sink_37_sink_size_1_18 <= __stream_conv2d_16_sink_37_sink_size_1_17;
      __stream_seq_14_cond_2_18 <= __stream_seq_14_cond_2_17;
      __stream_conv2d_16_sink_37_sink_offset_0_17 <= __stream_conv2d_16_sink_37_sink_offset_0_16;
      __stream_conv2d_16_sink_37_sink_size_1_17 <= __stream_conv2d_16_sink_37_sink_size_1_16;
      __stream_seq_14_cond_2_17 <= __stream_seq_14_cond_2_16;
      __stream_conv2d_16_sink_37_sink_offset_0_16 <= __stream_conv2d_16_sink_37_sink_offset_0_15;
      __stream_conv2d_16_sink_37_sink_size_1_16 <= __stream_conv2d_16_sink_37_sink_size_1_15;
      __stream_seq_14_cond_2_16 <= __stream_seq_14_cond_2_15;
      __stream_conv2d_16_sink_37_sink_offset_0_15 <= __stream_conv2d_16_sink_37_sink_offset_0_14;
      __stream_conv2d_16_sink_37_sink_size_1_15 <= __stream_conv2d_16_sink_37_sink_size_1_14;
      __stream_seq_14_cond_2_15 <= __stream_seq_14_cond_2_14;
      __stream_conv2d_16_sink_37_sink_offset_0_14 <= __stream_conv2d_16_sink_37_sink_offset_0_13;
      __stream_conv2d_16_sink_37_sink_size_1_14 <= __stream_conv2d_16_sink_37_sink_size_1_13;
      __stream_seq_14_cond_2_14 <= __stream_seq_14_cond_2_13;
      __stream_conv2d_16_sink_37_sink_offset_0_13 <= __stream_conv2d_16_sink_37_sink_offset_0_12;
      __stream_conv2d_16_sink_37_sink_size_1_13 <= __stream_conv2d_16_sink_37_sink_size_1_12;
      __stream_seq_14_cond_2_13 <= __stream_seq_14_cond_2_12;
      __stream_conv2d_16_sink_37_sink_offset_0_12 <= __stream_conv2d_16_sink_37_sink_offset_0_11;
      __stream_conv2d_16_sink_37_sink_size_1_12 <= __stream_conv2d_16_sink_37_sink_size_1_11;
      __stream_seq_14_cond_2_12 <= __stream_seq_14_cond_2_11;
      __stream_conv2d_16_sink_37_sink_offset_0_11 <= __stream_conv2d_16_sink_37_sink_offset_0_10;
      __stream_conv2d_16_sink_37_sink_size_1_11 <= __stream_conv2d_16_sink_37_sink_size_1_10;
      __stream_seq_14_cond_2_11 <= __stream_seq_14_cond_2_10;
      __stream_conv2d_16_sink_37_sink_offset_0_10 <= __stream_conv2d_16_sink_37_sink_offset_0_9;
      __stream_conv2d_16_sink_37_sink_size_1_10 <= __stream_conv2d_16_sink_37_sink_size_1_9;
      __stream_seq_14_cond_2_10 <= __stream_seq_14_cond_2_9;
      __stream_conv2d_16_sink_37_sink_offset_0_9 <= __stream_conv2d_16_sink_37_sink_offset_0_8;
      __stream_conv2d_16_sink_37_sink_size_1_9 <= __stream_conv2d_16_sink_37_sink_size_1_8;
      __stream_seq_14_cond_2_9 <= __stream_seq_14_cond_2_8;
      __stream_conv2d_16_sink_37_sink_offset_0_8 <= __stream_conv2d_16_sink_37_sink_offset_0_7;
      __stream_conv2d_16_sink_37_sink_size_1_8 <= __stream_conv2d_16_sink_37_sink_size_1_7;
      __stream_seq_14_cond_2_8 <= __stream_seq_14_cond_2_7;
      __stream_conv2d_16_sink_37_sink_offset_0_7 <= __stream_conv2d_16_sink_37_sink_offset_0_6;
      __stream_conv2d_16_sink_37_sink_size_1_7 <= __stream_conv2d_16_sink_37_sink_size_1_6;
      __stream_seq_14_cond_2_7 <= __stream_seq_14_cond_2_6;
      __stream_conv2d_16_sink_37_sink_offset_0_6 <= __stream_conv2d_16_sink_37_sink_offset_0_5;
      __stream_conv2d_16_sink_37_sink_size_1_6 <= __stream_conv2d_16_sink_37_sink_size_1_5;
      __stream_seq_14_cond_2_6 <= __stream_seq_14_cond_2_5;
      __stream_conv2d_16_sink_37_sink_offset_0_5 <= __stream_conv2d_16_sink_37_sink_offset_0_4;
      __stream_conv2d_16_sink_37_sink_size_1_5 <= __stream_conv2d_16_sink_37_sink_size_1_4;
      __stream_seq_14_cond_2_5 <= __stream_seq_14_cond_2_4;
      __stream_conv2d_16_sink_37_sink_offset_0_4 <= __stream_conv2d_16_sink_37_sink_offset_0_3;
      __stream_conv2d_16_sink_37_sink_size_1_4 <= __stream_conv2d_16_sink_37_sink_size_1_3;
      __stream_seq_14_cond_2_4 <= __stream_seq_14_cond_2_3;
      __stream_conv2d_16_sink_37_sink_offset_0_3 <= __stream_conv2d_16_sink_37_sink_offset_0_2;
      __stream_conv2d_16_sink_37_sink_size_1_3 <= __stream_conv2d_16_sink_37_sink_size_1_2;
      __stream_seq_14_cond_2_3 <= __stream_seq_14_cond_2_2;
      __stream_conv2d_16_sink_37_sink_offset_0_2 <= __stream_conv2d_16_sink_37_sink_offset_0_1;
      __stream_conv2d_16_sink_37_sink_size_1_2 <= __stream_conv2d_16_sink_37_sink_size_1_1;
      __stream_seq_14_cond_2_2 <= __stream_seq_14_cond_2_1;
      _stream_conv2d_16_source_6_idle <= _stream_conv2d_16_source_6_idle;
      _stream_conv2d_16_source_6_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_8_idle <= _stream_conv2d_16_source_8_idle;
      _stream_conv2d_16_source_8_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_10_idle <= _stream_conv2d_16_source_10_idle;
      _stream_conv2d_16_source_10_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_12_idle <= _stream_conv2d_16_source_12_idle;
      _stream_conv2d_16_source_12_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_14_idle <= _stream_conv2d_16_source_14_idle;
      _stream_conv2d_16_source_14_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_19_idle <= _stream_conv2d_16_source_19_idle;
      _stream_conv2d_16_source_19_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_20_idle <= _stream_conv2d_16_source_20_idle;
      _stream_conv2d_16_source_20_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_21_idle <= _stream_conv2d_16_source_21_idle;
      _stream_conv2d_16_source_21_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_22_idle <= _stream_conv2d_16_source_22_idle;
      _stream_conv2d_16_source_22_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_23_idle <= _stream_conv2d_16_source_23_idle;
      _stream_conv2d_16_source_23_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_24_idle <= _stream_conv2d_16_source_24_idle;
      _stream_conv2d_16_source_24_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_25_idle <= _stream_conv2d_16_source_25_idle;
      _stream_conv2d_16_source_25_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_26_idle <= _stream_conv2d_16_source_26_idle;
      _stream_conv2d_16_source_26_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_27_idle <= _stream_conv2d_16_source_27_idle;
      _stream_conv2d_16_source_27_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_28_idle <= _stream_conv2d_16_source_28_idle;
      _stream_conv2d_16_source_28_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_29_idle <= _stream_conv2d_16_source_29_idle;
      _stream_conv2d_16_source_29_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_30_idle <= _stream_conv2d_16_source_30_idle;
      _stream_conv2d_16_source_30_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_31_idle <= _stream_conv2d_16_source_31_idle;
      _stream_conv2d_16_source_31_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_32_idle <= _stream_conv2d_16_source_32_idle;
      _stream_conv2d_16_source_32_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_33_idle <= _stream_conv2d_16_source_33_idle;
      _stream_conv2d_16_source_33_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_34_idle <= _stream_conv2d_16_source_34_idle;
      _stream_conv2d_16_source_34_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_35_idle <= _stream_conv2d_16_source_35_idle;
      _stream_conv2d_16_source_35_source_ram_rvalid <= 0;
      _stream_conv2d_16_source_36_idle <= _stream_conv2d_16_source_36_idle;
      _stream_conv2d_16_source_36_source_ram_rvalid <= 0;
      _stream_conv2d_16_sink_37_sink_wenable <= 0;
      _stream_conv2d_16_sink_38_sink_wenable <= 0;
      _cond_data_235 <= (stream_conv2d_16_constant_5_data)? _reinterpretcast_data_234 : _reinterpretcast_data_234;
      _cond_data_242 <= (stream_conv2d_16_constant_7_data)? _reinterpretcast_data_241 : _reinterpretcast_data_241;
      _cond_data_249 <= (stream_conv2d_16_constant_9_data)? _reinterpretcast_data_248 : _reinterpretcast_data_248;
      _cond_data_256 <= (stream_conv2d_16_constant_11_data)? _reinterpretcast_data_255 : _reinterpretcast_data_255;
      _cond_data_263 <= (stream_conv2d_16_constant_13_data)? _reinterpretcast_data_262 : _reinterpretcast_data_262;
      _eq_data_277 <= stream_conv2d_16_constant_1_data == 3'sd2;
      _eq_data_281 <= stream_conv2d_16_constant_1_data == 2'sd1;
      _eq_data_284 <= stream_conv2d_16_constant_1_data == 1'sd0;
      _eq_data_287 <= stream_conv2d_16_constant_1_data == 3'sd2;
      _eq_data_291 <= stream_conv2d_16_constant_1_data == 2'sd1;
      _eq_data_294 <= stream_conv2d_16_constant_1_data == 1'sd0;
      _eq_data_297 <= stream_conv2d_16_constant_1_data == 3'sd2;
      _eq_data_301 <= stream_conv2d_16_constant_1_data == 2'sd1;
      _eq_data_304 <= stream_conv2d_16_constant_1_data == 1'sd0;
      _eq_data_307 <= stream_conv2d_16_constant_1_data == 3'sd2;
      _eq_data_311 <= stream_conv2d_16_constant_1_data == 2'sd1;
      _eq_data_314 <= stream_conv2d_16_constant_1_data == 1'sd0;
      _eq_data_317 <= stream_conv2d_16_constant_1_data == 3'sd2;
      _eq_data_321 <= stream_conv2d_16_constant_1_data == 2'sd1;
      _eq_data_324 <= stream_conv2d_16_constant_1_data == 1'sd0;
      _eq_data_327 <= stream_conv2d_16_constant_1_data == 3'sd2;
      _eq_data_331 <= stream_conv2d_16_constant_1_data == 2'sd1;
      _eq_data_334 <= stream_conv2d_16_constant_1_data == 1'sd0;
      _eq_data_337 <= stream_conv2d_16_constant_1_data == 3'sd2;
      _eq_data_341 <= stream_conv2d_16_constant_1_data == 2'sd1;
      _eq_data_344 <= stream_conv2d_16_constant_1_data == 1'sd0;
      _eq_data_347 <= stream_conv2d_16_constant_1_data == 3'sd2;
      _eq_data_351 <= stream_conv2d_16_constant_1_data == 2'sd1;
      _eq_data_354 <= stream_conv2d_16_constant_1_data == 1'sd0;
      _eq_data_357 <= stream_conv2d_16_constant_1_data == 3'sd2;
      _eq_data_361 <= stream_conv2d_16_constant_1_data == 2'sd1;
      _eq_data_364 <= stream_conv2d_16_constant_1_data == 1'sd0;
      _eq_data_367 <= stream_conv2d_16_constant_2_data == 3'sd2;
      _eq_data_371 <= stream_conv2d_16_constant_2_data == 2'sd1;
      _eq_data_374 <= stream_conv2d_16_constant_2_data == 1'sd0;
      _eq_data_377 <= stream_conv2d_16_constant_2_data == 3'sd2;
      _eq_data_381 <= stream_conv2d_16_constant_2_data == 2'sd1;
      _eq_data_384 <= stream_conv2d_16_constant_2_data == 1'sd0;
      _eq_data_387 <= stream_conv2d_16_constant_2_data == 3'sd2;
      _eq_data_391 <= stream_conv2d_16_constant_2_data == 2'sd1;
      _eq_data_394 <= stream_conv2d_16_constant_2_data == 1'sd0;
      _eq_data_397 <= stream_conv2d_16_constant_2_data == 3'sd2;
      _eq_data_401 <= stream_conv2d_16_constant_2_data == 2'sd1;
      _eq_data_404 <= stream_conv2d_16_constant_2_data == 1'sd0;
      _eq_data_407 <= stream_conv2d_16_constant_2_data == 3'sd2;
      _eq_data_411 <= stream_conv2d_16_constant_2_data == 2'sd1;
      _eq_data_414 <= stream_conv2d_16_constant_2_data == 1'sd0;
      _eq_data_417 <= stream_conv2d_16_constant_2_data == 3'sd2;
      _eq_data_421 <= stream_conv2d_16_constant_2_data == 2'sd1;
      _eq_data_424 <= stream_conv2d_16_constant_2_data == 1'sd0;
      _eq_data_427 <= stream_conv2d_16_constant_2_data == 3'sd2;
      _eq_data_431 <= stream_conv2d_16_constant_2_data == 2'sd1;
      _eq_data_434 <= stream_conv2d_16_constant_2_data == 1'sd0;
      _eq_data_437 <= stream_conv2d_16_constant_2_data == 3'sd2;
      _eq_data_441 <= stream_conv2d_16_constant_2_data == 2'sd1;
      _eq_data_444 <= stream_conv2d_16_constant_2_data == 1'sd0;
      _eq_data_447 <= stream_conv2d_16_constant_2_data == 3'sd2;
      _eq_data_451 <= stream_conv2d_16_constant_2_data == 2'sd1;
      _eq_data_454 <= stream_conv2d_16_constant_2_data == 1'sd0;
      __delay_data_898 <= stream_conv2d_16_source_21_data;
      __delay_data_900 <= stream_conv2d_16_source_20_data;
      __delay_data_904 <= stream_conv2d_16_source_19_data;
      __delay_data_907 <= stream_conv2d_16_source_24_data;
      __delay_data_909 <= stream_conv2d_16_source_23_data;
      __delay_data_913 <= stream_conv2d_16_source_22_data;
      __delay_data_916 <= stream_conv2d_16_source_27_data;
      __delay_data_918 <= stream_conv2d_16_source_26_data;
      __delay_data_922 <= stream_conv2d_16_source_25_data;
      __delay_data_940 <= _pointer_data_556;
      __delay_data_947 <= stream_conv2d_16_constant_15_data;
      __delay_data_948 <= _reinterpretcast_data_547;
      __delay_data_992 <= _pointer_data_558;
      __delay_data_999 <= _reinterpretcast_data_548;
      __delay_data_1040 <= _pointer_data_560;
      __delay_data_1047 <= _reinterpretcast_data_549;
      __delay_data_1075 <= _pointer_data_562;
      __delay_data_1082 <= _reinterpretcast_data_550;
      __delay_data_1110 <= _pointer_data_564;
      __delay_data_1117 <= _reinterpretcast_data_551;
      __delay_data_1145 <= _pointer_data_566;
      __delay_data_1152 <= _reinterpretcast_data_552;
      __delay_data_1179 <= _pointer_data_568;
      __delay_data_1186 <= _reinterpretcast_data_553;
      __delay_data_1213 <= _pointer_data_570;
      __delay_data_1220 <= _reinterpretcast_data_554;
      __delay_data_1247 <= _pointer_data_572;
      __delay_data_1254 <= _reinterpretcast_data_555;
      __delay_data_1268 <= stream_conv2d_16_constant_16_data;
      __delay_data_1289 <= stream_conv2d_16_constant_0_data;
      __delay_data_1339 <= stream_conv2d_16_constant_17_data;
      _cond_data_279 <= (_eq_data_277)? __delay_data_898 : 1'sd0;
      _cond_data_289 <= (_eq_data_287)? __delay_data_904 : 1'sd0;
      _cond_data_299 <= (_eq_data_297)? __delay_data_900 : 1'sd0;
      _cond_data_309 <= (_eq_data_307)? __delay_data_907 : 1'sd0;
      _cond_data_319 <= (_eq_data_317)? __delay_data_913 : 1'sd0;
      _cond_data_329 <= (_eq_data_327)? __delay_data_909 : 1'sd0;
      _cond_data_339 <= (_eq_data_337)? __delay_data_916 : 1'sd0;
      _cond_data_349 <= (_eq_data_347)? __delay_data_922 : 1'sd0;
      _cond_data_359 <= (_eq_data_357)? __delay_data_918 : 1'sd0;
      _plus_data_607 <= _cond_data_249 + __delay_data_947;
      _plus_data_624 <= _cond_data_249 + __delay_data_947;
      _plus_data_641 <= _cond_data_249 + __delay_data_947;
      _plus_data_658 <= _cond_data_249 + __delay_data_947;
      _plus_data_675 <= _cond_data_249 + __delay_data_947;
      _plus_data_692 <= _cond_data_249 + __delay_data_947;
      _plus_data_709 <= _cond_data_249 + __delay_data_947;
      _plus_data_726 <= _cond_data_249 + __delay_data_947;
      _plus_data_743 <= _cond_data_249 + __delay_data_947;
      _plus_data_759 <= _cond_data_256 + __delay_data_1268;
      _plus_data_770 <= _cond_data_263 + __delay_data_1339;
      __delay_data_899 <= _eq_data_281;
      __delay_data_901 <= __delay_data_900;
      __delay_data_902 <= _eq_data_284;
      __delay_data_905 <= __delay_data_904;
      __delay_data_908 <= _eq_data_311;
      __delay_data_910 <= __delay_data_909;
      __delay_data_911 <= _eq_data_314;
      __delay_data_914 <= __delay_data_913;
      __delay_data_917 <= _eq_data_341;
      __delay_data_919 <= __delay_data_918;
      __delay_data_920 <= _eq_data_344;
      __delay_data_923 <= __delay_data_922;
      __delay_data_925 <= _eq_data_367;
      __delay_data_928 <= _eq_data_371;
      __delay_data_933 <= _eq_data_374;
      __delay_data_941 <= __delay_data_940;
      __delay_data_949 <= __delay_data_948;
      __delay_data_962 <= _eq_data_291;
      __delay_data_963 <= __delay_data_898;
      __delay_data_964 <= _eq_data_294;
      __delay_data_967 <= _eq_data_321;
      __delay_data_968 <= __delay_data_907;
      __delay_data_969 <= _eq_data_324;
      __delay_data_972 <= _eq_data_351;
      __delay_data_973 <= __delay_data_916;
      __delay_data_974 <= _eq_data_354;
      __delay_data_977 <= _eq_data_397;
      __delay_data_980 <= _eq_data_401;
      __delay_data_985 <= _eq_data_404;
      __delay_data_993 <= __delay_data_992;
      __delay_data_1000 <= __delay_data_999;
      __delay_data_1013 <= _eq_data_301;
      __delay_data_1014 <= _eq_data_304;
      __delay_data_1017 <= _eq_data_331;
      __delay_data_1018 <= _eq_data_334;
      __delay_data_1021 <= _eq_data_361;
      __delay_data_1022 <= _eq_data_364;
      __delay_data_1025 <= _eq_data_427;
      __delay_data_1028 <= _eq_data_431;
      __delay_data_1033 <= _eq_data_434;
      __delay_data_1041 <= __delay_data_1040;
      __delay_data_1048 <= __delay_data_1047;
      __delay_data_1061 <= _eq_data_377;
      __delay_data_1064 <= _eq_data_381;
      __delay_data_1069 <= _eq_data_384;
      __delay_data_1076 <= __delay_data_1075;
      __delay_data_1083 <= __delay_data_1082;
      __delay_data_1096 <= _eq_data_407;
      __delay_data_1099 <= _eq_data_411;
      __delay_data_1104 <= _eq_data_414;
      __delay_data_1111 <= __delay_data_1110;
      __delay_data_1118 <= __delay_data_1117;
      __delay_data_1131 <= _eq_data_437;
      __delay_data_1134 <= _eq_data_441;
      __delay_data_1139 <= _eq_data_444;
      __delay_data_1146 <= __delay_data_1145;
      __delay_data_1153 <= __delay_data_1152;
      __delay_data_1166 <= _eq_data_387;
      __delay_data_1169 <= _eq_data_391;
      __delay_data_1173 <= _eq_data_394;
      __delay_data_1180 <= __delay_data_1179;
      __delay_data_1187 <= __delay_data_1186;
      __delay_data_1200 <= _eq_data_417;
      __delay_data_1203 <= _eq_data_421;
      __delay_data_1207 <= _eq_data_424;
      __delay_data_1214 <= __delay_data_1213;
      __delay_data_1221 <= __delay_data_1220;
      __delay_data_1234 <= _eq_data_447;
      __delay_data_1237 <= _eq_data_451;
      __delay_data_1241 <= _eq_data_454;
      __delay_data_1248 <= __delay_data_1247;
      __delay_data_1255 <= __delay_data_1254;
      __delay_data_1290 <= __delay_data_1289;
      __delay_data_1311 <= _cond_data_235;
      __delay_data_1340 <= _cond_data_242;
      _cond_data_283 <= (__delay_data_899)? __delay_data_901 : _cond_data_279;
      _cond_data_293 <= (__delay_data_962)? __delay_data_963 : _cond_data_289;
      _cond_data_303 <= (__delay_data_1013)? __delay_data_905 : _cond_data_299;
      _cond_data_313 <= (__delay_data_908)? __delay_data_910 : _cond_data_309;
      _cond_data_323 <= (__delay_data_967)? __delay_data_968 : _cond_data_319;
      _cond_data_333 <= (__delay_data_1017)? __delay_data_914 : _cond_data_329;
      _cond_data_343 <= (__delay_data_917)? __delay_data_919 : _cond_data_339;
      _cond_data_353 <= (__delay_data_972)? __delay_data_973 : _cond_data_349;
      _cond_data_363 <= (__delay_data_1021)? __delay_data_923 : _cond_data_359;
      __delay_data_903 <= __delay_data_902;
      __delay_data_906 <= __delay_data_905;
      __delay_data_912 <= __delay_data_911;
      __delay_data_915 <= __delay_data_914;
      __delay_data_921 <= __delay_data_920;
      __delay_data_924 <= __delay_data_923;
      __delay_data_926 <= __delay_data_925;
      __delay_data_929 <= __delay_data_928;
      __delay_data_934 <= __delay_data_933;
      __delay_data_942 <= __delay_data_941;
      __delay_data_950 <= __delay_data_949;
      __delay_data_956 <= _plus_data_607;
      __delay_data_965 <= __delay_data_964;
      __delay_data_966 <= __delay_data_901;
      __delay_data_970 <= __delay_data_969;
      __delay_data_971 <= __delay_data_910;
      __delay_data_975 <= __delay_data_974;
      __delay_data_976 <= __delay_data_919;
      __delay_data_978 <= __delay_data_977;
      __delay_data_981 <= __delay_data_980;
      __delay_data_986 <= __delay_data_985;
      __delay_data_994 <= __delay_data_993;
      __delay_data_1001 <= __delay_data_1000;
      __delay_data_1007 <= _plus_data_624;
      __delay_data_1015 <= __delay_data_1014;
      __delay_data_1016 <= __delay_data_963;
      __delay_data_1019 <= __delay_data_1018;
      __delay_data_1020 <= __delay_data_968;
      __delay_data_1023 <= __delay_data_1022;
      __delay_data_1024 <= __delay_data_973;
      __delay_data_1026 <= __delay_data_1025;
      __delay_data_1029 <= __delay_data_1028;
      __delay_data_1034 <= __delay_data_1033;
      __delay_data_1042 <= __delay_data_1041;
      __delay_data_1049 <= __delay_data_1048;
      __delay_data_1055 <= _plus_data_641;
      __delay_data_1062 <= __delay_data_1061;
      __delay_data_1065 <= __delay_data_1064;
      __delay_data_1070 <= __delay_data_1069;
      __delay_data_1077 <= __delay_data_1076;
      __delay_data_1084 <= __delay_data_1083;
      __delay_data_1090 <= _plus_data_658;
      __delay_data_1097 <= __delay_data_1096;
      __delay_data_1100 <= __delay_data_1099;
      __delay_data_1105 <= __delay_data_1104;
      __delay_data_1112 <= __delay_data_1111;
      __delay_data_1119 <= __delay_data_1118;
      __delay_data_1125 <= _plus_data_675;
      __delay_data_1132 <= __delay_data_1131;
      __delay_data_1135 <= __delay_data_1134;
      __delay_data_1140 <= __delay_data_1139;
      __delay_data_1147 <= __delay_data_1146;
      __delay_data_1154 <= __delay_data_1153;
      __delay_data_1160 <= _plus_data_692;
      __delay_data_1167 <= __delay_data_1166;
      __delay_data_1170 <= __delay_data_1169;
      __delay_data_1174 <= __delay_data_1173;
      __delay_data_1181 <= __delay_data_1180;
      __delay_data_1188 <= __delay_data_1187;
      __delay_data_1194 <= _plus_data_709;
      __delay_data_1201 <= __delay_data_1200;
      __delay_data_1204 <= __delay_data_1203;
      __delay_data_1208 <= __delay_data_1207;
      __delay_data_1215 <= __delay_data_1214;
      __delay_data_1222 <= __delay_data_1221;
      __delay_data_1228 <= _plus_data_726;
      __delay_data_1235 <= __delay_data_1234;
      __delay_data_1238 <= __delay_data_1237;
      __delay_data_1242 <= __delay_data_1241;
      __delay_data_1249 <= __delay_data_1248;
      __delay_data_1256 <= __delay_data_1255;
      __delay_data_1262 <= _plus_data_743;
      __delay_data_1269 <= _plus_data_759;
      __delay_data_1291 <= __delay_data_1290;
      __delay_data_1312 <= __delay_data_1311;
      __delay_data_1341 <= __delay_data_1340;
      __delay_data_1369 <= _plus_data_770;
      _cond_data_286 <= (__delay_data_903)? __delay_data_906 : _cond_data_283;
      _cond_data_296 <= (__delay_data_965)? __delay_data_966 : _cond_data_293;
      _cond_data_306 <= (__delay_data_1015)? __delay_data_1016 : _cond_data_303;
      _cond_data_316 <= (__delay_data_912)? __delay_data_915 : _cond_data_313;
      _cond_data_326 <= (__delay_data_970)? __delay_data_971 : _cond_data_323;
      _cond_data_336 <= (__delay_data_1019)? __delay_data_1020 : _cond_data_333;
      _cond_data_346 <= (__delay_data_921)? __delay_data_924 : _cond_data_343;
      _cond_data_356 <= (__delay_data_975)? __delay_data_976 : _cond_data_353;
      _cond_data_366 <= (__delay_data_1023)? __delay_data_1024 : _cond_data_363;
      __delay_data_927 <= __delay_data_926;
      __delay_data_930 <= __delay_data_929;
      __delay_data_935 <= __delay_data_934;
      __delay_data_943 <= __delay_data_942;
      __delay_data_951 <= __delay_data_950;
      __delay_data_957 <= __delay_data_956;
      __delay_data_979 <= __delay_data_978;
      __delay_data_982 <= __delay_data_981;
      __delay_data_987 <= __delay_data_986;
      __delay_data_995 <= __delay_data_994;
      __delay_data_1002 <= __delay_data_1001;
      __delay_data_1008 <= __delay_data_1007;
      __delay_data_1027 <= __delay_data_1026;
      __delay_data_1030 <= __delay_data_1029;
      __delay_data_1035 <= __delay_data_1034;
      __delay_data_1043 <= __delay_data_1042;
      __delay_data_1050 <= __delay_data_1049;
      __delay_data_1056 <= __delay_data_1055;
      __delay_data_1063 <= __delay_data_1062;
      __delay_data_1066 <= __delay_data_1065;
      __delay_data_1071 <= __delay_data_1070;
      __delay_data_1078 <= __delay_data_1077;
      __delay_data_1085 <= __delay_data_1084;
      __delay_data_1091 <= __delay_data_1090;
      __delay_data_1098 <= __delay_data_1097;
      __delay_data_1101 <= __delay_data_1100;
      __delay_data_1106 <= __delay_data_1105;
      __delay_data_1113 <= __delay_data_1112;
      __delay_data_1120 <= __delay_data_1119;
      __delay_data_1126 <= __delay_data_1125;
      __delay_data_1133 <= __delay_data_1132;
      __delay_data_1136 <= __delay_data_1135;
      __delay_data_1141 <= __delay_data_1140;
      __delay_data_1148 <= __delay_data_1147;
      __delay_data_1155 <= __delay_data_1154;
      __delay_data_1161 <= __delay_data_1160;
      __delay_data_1168 <= __delay_data_1167;
      __delay_data_1171 <= __delay_data_1170;
      __delay_data_1175 <= __delay_data_1174;
      __delay_data_1182 <= __delay_data_1181;
      __delay_data_1189 <= __delay_data_1188;
      __delay_data_1195 <= __delay_data_1194;
      __delay_data_1202 <= __delay_data_1201;
      __delay_data_1205 <= __delay_data_1204;
      __delay_data_1209 <= __delay_data_1208;
      __delay_data_1216 <= __delay_data_1215;
      __delay_data_1223 <= __delay_data_1222;
      __delay_data_1229 <= __delay_data_1228;
      __delay_data_1236 <= __delay_data_1235;
      __delay_data_1239 <= __delay_data_1238;
      __delay_data_1243 <= __delay_data_1242;
      __delay_data_1250 <= __delay_data_1249;
      __delay_data_1257 <= __delay_data_1256;
      __delay_data_1263 <= __delay_data_1262;
      __delay_data_1270 <= __delay_data_1269;
      __delay_data_1292 <= __delay_data_1291;
      __delay_data_1313 <= __delay_data_1312;
      __delay_data_1342 <= __delay_data_1341;
      __delay_data_1370 <= __delay_data_1369;
      _cond_data_369 <= (__delay_data_927)? _cond_data_346 : 1'sd0;
      _cond_data_379 <= (__delay_data_1063)? _cond_data_286 : 1'sd0;
      _cond_data_389 <= (__delay_data_1168)? _cond_data_316 : 1'sd0;
      _cond_data_399 <= (__delay_data_979)? _cond_data_356 : 1'sd0;
      _cond_data_409 <= (__delay_data_1098)? _cond_data_296 : 1'sd0;
      _cond_data_419 <= (__delay_data_1202)? _cond_data_326 : 1'sd0;
      _cond_data_429 <= (__delay_data_1027)? _cond_data_366 : 1'sd0;
      _cond_data_439 <= (__delay_data_1133)? _cond_data_306 : 1'sd0;
      _cond_data_449 <= (__delay_data_1236)? _cond_data_336 : 1'sd0;
      __delay_data_931 <= __delay_data_930;
      __delay_data_932 <= _cond_data_316;
      __delay_data_936 <= __delay_data_935;
      __delay_data_938 <= _cond_data_286;
      __delay_data_944 <= __delay_data_943;
      __delay_data_952 <= __delay_data_951;
      __delay_data_958 <= __delay_data_957;
      __delay_data_983 <= __delay_data_982;
      __delay_data_984 <= _cond_data_326;
      __delay_data_988 <= __delay_data_987;
      __delay_data_990 <= _cond_data_296;
      __delay_data_996 <= __delay_data_995;
      __delay_data_1003 <= __delay_data_1002;
      __delay_data_1009 <= __delay_data_1008;
      __delay_data_1031 <= __delay_data_1030;
      __delay_data_1032 <= _cond_data_336;
      __delay_data_1036 <= __delay_data_1035;
      __delay_data_1038 <= _cond_data_306;
      __delay_data_1044 <= __delay_data_1043;
      __delay_data_1051 <= __delay_data_1050;
      __delay_data_1057 <= __delay_data_1056;
      __delay_data_1067 <= __delay_data_1066;
      __delay_data_1068 <= _cond_data_346;
      __delay_data_1072 <= __delay_data_1071;
      __delay_data_1079 <= __delay_data_1078;
      __delay_data_1086 <= __delay_data_1085;
      __delay_data_1092 <= __delay_data_1091;
      __delay_data_1102 <= __delay_data_1101;
      __delay_data_1103 <= _cond_data_356;
      __delay_data_1107 <= __delay_data_1106;
      __delay_data_1114 <= __delay_data_1113;
      __delay_data_1121 <= __delay_data_1120;
      __delay_data_1127 <= __delay_data_1126;
      __delay_data_1137 <= __delay_data_1136;
      __delay_data_1138 <= _cond_data_366;
      __delay_data_1142 <= __delay_data_1141;
      __delay_data_1149 <= __delay_data_1148;
      __delay_data_1156 <= __delay_data_1155;
      __delay_data_1162 <= __delay_data_1161;
      __delay_data_1172 <= __delay_data_1171;
      __delay_data_1176 <= __delay_data_1175;
      __delay_data_1183 <= __delay_data_1182;
      __delay_data_1190 <= __delay_data_1189;
      __delay_data_1196 <= __delay_data_1195;
      __delay_data_1206 <= __delay_data_1205;
      __delay_data_1210 <= __delay_data_1209;
      __delay_data_1217 <= __delay_data_1216;
      __delay_data_1224 <= __delay_data_1223;
      __delay_data_1230 <= __delay_data_1229;
      __delay_data_1240 <= __delay_data_1239;
      __delay_data_1244 <= __delay_data_1243;
      __delay_data_1251 <= __delay_data_1250;
      __delay_data_1258 <= __delay_data_1257;
      __delay_data_1264 <= __delay_data_1263;
      __delay_data_1271 <= __delay_data_1270;
      __delay_data_1293 <= __delay_data_1292;
      __delay_data_1314 <= __delay_data_1313;
      __delay_data_1343 <= __delay_data_1342;
      __delay_data_1371 <= __delay_data_1370;
      _cond_data_373 <= (__delay_data_931)? __delay_data_932 : _cond_data_369;
      _cond_data_383 <= (__delay_data_1067)? __delay_data_1068 : _cond_data_379;
      _cond_data_393 <= (__delay_data_1172)? __delay_data_938 : _cond_data_389;
      _cond_data_403 <= (__delay_data_983)? __delay_data_984 : _cond_data_399;
      _cond_data_413 <= (__delay_data_1102)? __delay_data_1103 : _cond_data_409;
      _cond_data_423 <= (__delay_data_1206)? __delay_data_990 : _cond_data_419;
      _cond_data_433 <= (__delay_data_1031)? __delay_data_1032 : _cond_data_429;
      _cond_data_443 <= (__delay_data_1137)? __delay_data_1138 : _cond_data_439;
      _cond_data_453 <= (__delay_data_1240)? __delay_data_1038 : _cond_data_449;
      __delay_data_937 <= __delay_data_936;
      __delay_data_939 <= __delay_data_938;
      __delay_data_945 <= __delay_data_944;
      __delay_data_953 <= __delay_data_952;
      __delay_data_959 <= __delay_data_958;
      __delay_data_989 <= __delay_data_988;
      __delay_data_991 <= __delay_data_990;
      __delay_data_997 <= __delay_data_996;
      __delay_data_1004 <= __delay_data_1003;
      __delay_data_1010 <= __delay_data_1009;
      __delay_data_1037 <= __delay_data_1036;
      __delay_data_1039 <= __delay_data_1038;
      __delay_data_1045 <= __delay_data_1044;
      __delay_data_1052 <= __delay_data_1051;
      __delay_data_1058 <= __delay_data_1057;
      __delay_data_1073 <= __delay_data_1072;
      __delay_data_1074 <= __delay_data_932;
      __delay_data_1080 <= __delay_data_1079;
      __delay_data_1087 <= __delay_data_1086;
      __delay_data_1093 <= __delay_data_1092;
      __delay_data_1108 <= __delay_data_1107;
      __delay_data_1109 <= __delay_data_984;
      __delay_data_1115 <= __delay_data_1114;
      __delay_data_1122 <= __delay_data_1121;
      __delay_data_1128 <= __delay_data_1127;
      __delay_data_1143 <= __delay_data_1142;
      __delay_data_1144 <= __delay_data_1032;
      __delay_data_1150 <= __delay_data_1149;
      __delay_data_1157 <= __delay_data_1156;
      __delay_data_1163 <= __delay_data_1162;
      __delay_data_1177 <= __delay_data_1176;
      __delay_data_1178 <= __delay_data_1068;
      __delay_data_1184 <= __delay_data_1183;
      __delay_data_1191 <= __delay_data_1190;
      __delay_data_1197 <= __delay_data_1196;
      __delay_data_1211 <= __delay_data_1210;
      __delay_data_1212 <= __delay_data_1103;
      __delay_data_1218 <= __delay_data_1217;
      __delay_data_1225 <= __delay_data_1224;
      __delay_data_1231 <= __delay_data_1230;
      __delay_data_1245 <= __delay_data_1244;
      __delay_data_1246 <= __delay_data_1138;
      __delay_data_1252 <= __delay_data_1251;
      __delay_data_1259 <= __delay_data_1258;
      __delay_data_1265 <= __delay_data_1264;
      __delay_data_1272 <= __delay_data_1271;
      __delay_data_1294 <= __delay_data_1293;
      __delay_data_1315 <= __delay_data_1314;
      __delay_data_1344 <= __delay_data_1343;
      __delay_data_1372 <= __delay_data_1371;
      _cond_data_376 <= (__delay_data_937)? __delay_data_939 : _cond_data_373;
      _cond_data_386 <= (__delay_data_1073)? __delay_data_1074 : _cond_data_383;
      _cond_data_396 <= (__delay_data_1177)? __delay_data_1178 : _cond_data_393;
      _cond_data_406 <= (__delay_data_989)? __delay_data_991 : _cond_data_403;
      _cond_data_416 <= (__delay_data_1108)? __delay_data_1109 : _cond_data_413;
      _cond_data_426 <= (__delay_data_1211)? __delay_data_1212 : _cond_data_423;
      _cond_data_436 <= (__delay_data_1037)? __delay_data_1039 : _cond_data_433;
      _cond_data_446 <= (__delay_data_1143)? __delay_data_1144 : _cond_data_443;
      _cond_data_456 <= (__delay_data_1245)? __delay_data_1246 : _cond_data_453;
      __delay_data_946 <= __delay_data_945;
      __delay_data_954 <= __delay_data_953;
      __delay_data_960 <= __delay_data_959;
      __delay_data_998 <= __delay_data_997;
      __delay_data_1005 <= __delay_data_1004;
      __delay_data_1011 <= __delay_data_1010;
      __delay_data_1046 <= __delay_data_1045;
      __delay_data_1053 <= __delay_data_1052;
      __delay_data_1059 <= __delay_data_1058;
      __delay_data_1081 <= __delay_data_1080;
      __delay_data_1088 <= __delay_data_1087;
      __delay_data_1094 <= __delay_data_1093;
      __delay_data_1116 <= __delay_data_1115;
      __delay_data_1123 <= __delay_data_1122;
      __delay_data_1129 <= __delay_data_1128;
      __delay_data_1151 <= __delay_data_1150;
      __delay_data_1158 <= __delay_data_1157;
      __delay_data_1164 <= __delay_data_1163;
      __delay_data_1185 <= __delay_data_1184;
      __delay_data_1192 <= __delay_data_1191;
      __delay_data_1198 <= __delay_data_1197;
      __delay_data_1219 <= __delay_data_1218;
      __delay_data_1226 <= __delay_data_1225;
      __delay_data_1232 <= __delay_data_1231;
      __delay_data_1253 <= __delay_data_1252;
      __delay_data_1260 <= __delay_data_1259;
      __delay_data_1266 <= __delay_data_1265;
      __delay_data_1273 <= __delay_data_1272;
      __delay_data_1295 <= __delay_data_1294;
      __delay_data_1316 <= __delay_data_1315;
      __delay_data_1345 <= __delay_data_1344;
      __delay_data_1373 <= __delay_data_1372;
      _cond_data_575 <= (__delay_data_946)? 1'sd0 : _reinterpretcast_data_493;
      _cond_data_577 <= (__delay_data_998)? 1'sd0 : _reinterpretcast_data_494;
      _cond_data_579 <= (__delay_data_1046)? 1'sd0 : _reinterpretcast_data_495;
      _cond_data_581 <= (__delay_data_1081)? 1'sd0 : _reinterpretcast_data_496;
      _cond_data_583 <= (__delay_data_1116)? 1'sd0 : _reinterpretcast_data_497;
      _cond_data_585 <= (__delay_data_1151)? 1'sd0 : _reinterpretcast_data_498;
      _cond_data_587 <= (__delay_data_1185)? 1'sd0 : _reinterpretcast_data_499;
      _cond_data_589 <= (__delay_data_1219)? 1'sd0 : _reinterpretcast_data_500;
      _cond_data_591 <= (__delay_data_1253)? 1'sd0 : _reinterpretcast_data_501;
      __delay_data_955 <= __delay_data_954;
      __delay_data_961 <= __delay_data_960;
      __delay_data_1006 <= __delay_data_1005;
      __delay_data_1012 <= __delay_data_1011;
      __delay_data_1054 <= __delay_data_1053;
      __delay_data_1060 <= __delay_data_1059;
      __delay_data_1089 <= __delay_data_1088;
      __delay_data_1095 <= __delay_data_1094;
      __delay_data_1124 <= __delay_data_1123;
      __delay_data_1130 <= __delay_data_1129;
      __delay_data_1159 <= __delay_data_1158;
      __delay_data_1165 <= __delay_data_1164;
      __delay_data_1193 <= __delay_data_1192;
      __delay_data_1199 <= __delay_data_1198;
      __delay_data_1227 <= __delay_data_1226;
      __delay_data_1233 <= __delay_data_1232;
      __delay_data_1261 <= __delay_data_1260;
      __delay_data_1267 <= __delay_data_1266;
      __delay_data_1274 <= __delay_data_1273;
      __delay_data_1296 <= __delay_data_1295;
      __delay_data_1317 <= __delay_data_1316;
      __delay_data_1346 <= __delay_data_1345;
      __delay_data_1374 <= __delay_data_1373;
      __delay_data_1275 <= __delay_data_1274;
      __delay_data_1297 <= __delay_data_1296;
      __delay_data_1318 <= __delay_data_1317;
      __delay_data_1347 <= __delay_data_1346;
      __delay_data_1375 <= __delay_data_1374;
      __delay_data_1276 <= __delay_data_1275;
      __delay_data_1298 <= __delay_data_1297;
      __delay_data_1319 <= __delay_data_1318;
      __delay_data_1348 <= __delay_data_1347;
      __delay_data_1376 <= __delay_data_1375;
      __delay_data_1277 <= __delay_data_1276;
      __delay_data_1299 <= __delay_data_1298;
      __delay_data_1320 <= __delay_data_1319;
      __delay_data_1349 <= __delay_data_1348;
      __delay_data_1377 <= __delay_data_1376;
      __delay_data_1278 <= __delay_data_1277;
      __delay_data_1300 <= __delay_data_1299;
      __delay_data_1321 <= __delay_data_1320;
      __delay_data_1350 <= __delay_data_1349;
      __delay_data_1378 <= __delay_data_1377;
      __delay_data_1279 <= __delay_data_1278;
      __delay_data_1301 <= __delay_data_1300;
      __delay_data_1322 <= __delay_data_1321;
      __delay_data_1351 <= __delay_data_1350;
      __delay_data_1379 <= __delay_data_1378;
      __delay_data_1280 <= __delay_data_1279;
      __delay_data_1302 <= __delay_data_1301;
      __delay_data_1323 <= __delay_data_1322;
      __delay_data_1352 <= __delay_data_1351;
      __delay_data_1380 <= __delay_data_1379;
      __delay_data_1281 <= __delay_data_1280;
      __delay_data_1303 <= __delay_data_1302;
      __delay_data_1324 <= __delay_data_1323;
      __delay_data_1353 <= __delay_data_1352;
      __delay_data_1381 <= __delay_data_1380;
      __delay_data_1282 <= __delay_data_1281;
      __delay_data_1304 <= __delay_data_1303;
      __delay_data_1325 <= __delay_data_1324;
      __delay_data_1354 <= __delay_data_1353;
      __delay_data_1382 <= __delay_data_1381;
      __delay_data_1283 <= __delay_data_1282;
      __delay_data_1305 <= __delay_data_1304;
      __delay_data_1326 <= __delay_data_1325;
      __delay_data_1355 <= __delay_data_1354;
      __delay_data_1383 <= __delay_data_1382;
      __substreamoutput_data_608 <= mul_4_z_data;
      __substreamoutput_data_625 <= mul_5_z_data;
      __substreamoutput_data_642 <= mul_6_z_data;
      __substreamoutput_data_659 <= mul_7_z_data;
      __substreamoutput_data_676 <= mul_8_z_data;
      __substreamoutput_data_693 <= mul_9_z_data;
      __substreamoutput_data_710 <= mul_10_z_data;
      __substreamoutput_data_727 <= mul_11_z_data;
      __substreamoutput_data_744 <= mul_12_z_data;
      __delay_data_1284 <= __delay_data_1283;
      __delay_data_1306 <= __delay_data_1305;
      __delay_data_1327 <= __delay_data_1326;
      __delay_data_1356 <= __delay_data_1355;
      __delay_data_1384 <= __delay_data_1383;
      __delay_data_1285 <= __delay_data_1284;
      __delay_data_1307 <= __delay_data_1306;
      __delay_data_1328 <= __delay_data_1327;
      __delay_data_1357 <= __delay_data_1356;
      __delay_data_1385 <= __delay_data_1384;
      __delay_data_1286 <= __delay_data_1285;
      __delay_data_1308 <= __delay_data_1307;
      __delay_data_1329 <= __delay_data_1328;
      __delay_data_1358 <= __delay_data_1357;
      __delay_data_1386 <= __delay_data_1385;
      __delay_data_1287 <= __delay_data_1286;
      __delay_data_1309 <= __delay_data_1308;
      __delay_data_1330 <= __delay_data_1329;
      __delay_data_1359 <= __delay_data_1358;
      __delay_data_1387 <= __delay_data_1386;
      __substreamoutput_data_746 <= add_tree_2_sum_data;
      __delay_data_1288 <= __delay_data_1287;
      __delay_data_1310 <= __delay_data_1309;
      __delay_data_1331 <= __delay_data_1330;
      __delay_data_1360 <= __delay_data_1359;
      __delay_data_1388 <= __delay_data_1387;
      __delay_data_1332 <= __delay_data_1331;
      __delay_data_1361 <= __delay_data_1360;
      __delay_data_1389 <= __delay_data_1388;
      __delay_data_1333 <= __delay_data_1332;
      __delay_data_1362 <= __delay_data_1361;
      __delay_data_1390 <= __delay_data_1389;
      __delay_data_1334 <= __delay_data_1333;
      __delay_data_1363 <= __delay_data_1362;
      __delay_data_1391 <= __delay_data_1390;
      __delay_data_1335 <= __delay_data_1334;
      __delay_data_1364 <= __delay_data_1363;
      __delay_data_1392 <= __delay_data_1391;
      __delay_data_1336 <= __delay_data_1335;
      __delay_data_1365 <= __delay_data_1364;
      __delay_data_1393 <= __delay_data_1392;
      __delay_data_1337 <= __delay_data_1336;
      __delay_data_1366 <= __delay_data_1365;
      __delay_data_1394 <= __delay_data_1393;
      __substreamoutput_data_760 <= acc_0_sum_data;
      __substreamoutput_data_761 <= acc_0_valid_data;
      __delay_data_1338 <= __delay_data_1337;
      __delay_data_1367 <= __delay_data_1366;
      __delay_data_1395 <= __delay_data_1394;
      _plus_data_762 <= __substreamoutput_data_760 + __delay_data_1338;
      __delay_data_1368 <= __delay_data_1367;
      __delay_data_1396 <= __delay_data_1395;
      __delay_data_1398 <= __substreamoutput_data_761;
      __delay_data_1399 <= __delay_data_1398;
      __delay_data_1400 <= __delay_data_1399;
      __delay_data_1401 <= __delay_data_1400;
      __delay_data_1402 <= __delay_data_1401;
      __delay_data_1403 <= __delay_data_1402;
      __delay_data_1404 <= __delay_data_1403;
      __delay_data_1405 <= __delay_data_1404;
      __delay_data_1406 <= __delay_data_1405;
      __delay_data_1407 <= __delay_data_1406;
      __substreamoutput_data_771 <= mul_rshift_clip_3_z_data;
      __delay_data_1408 <= __delay_data_1407;
      _greaterthan_data_773 <= __substreamoutput_data_771 > 1'sd0;
      __delay_data_1397 <= __substreamoutput_data_771;
      __delay_data_1409 <= __delay_data_1408;
      _cond_data_775 <= (_greaterthan_data_773)? __delay_data_1397 : 1'sd0;
      __delay_data_1410 <= __delay_data_1409;
      _set_flag_457 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_457 <= 1;
      end 
      if(_set_flag_457) begin
        _stream_conv2d_16_constant_0_next_constant_data <= cparam_conv2d_16_stream_reduce_size;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_214 <= _stream_conv2d_16_constant_0_next_constant_data;
      end 
      _set_flag_458 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_458 <= 1;
      end 
      if(_set_flag_458) begin
        _stream_conv2d_16_constant_1_next_constant_data <= conv2d_16_col_select;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_215 <= _stream_conv2d_16_constant_1_next_constant_data;
      end 
      _set_flag_459 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_459 <= 1;
      end 
      if(_set_flag_459) begin
        _stream_conv2d_16_constant_2_next_constant_data <= conv2d_16_row_select_buf;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_216 <= _stream_conv2d_16_constant_2_next_constant_data;
      end 
      _set_flag_460 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_460 <= 1;
      end 
      if(_set_flag_460) begin
        _stream_conv2d_16_constant_3_next_constant_data <= conv2d_16_stream_pad_masks;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_217 <= _stream_conv2d_16_constant_3_next_constant_data;
      end 
      _set_flag_461 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_461 <= 1;
      end 
      if(_set_flag_461) begin
        _stream_conv2d_16_constant_4_next_constant_data <= cparam_conv2d_16_stream_omit_mask;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_218 <= _stream_conv2d_16_constant_4_next_constant_data;
      end 
      _set_flag_462 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_462 <= 1;
      end 
      if(_set_flag_462) begin
        _stream_conv2d_16_constant_5_next_constant_data <= cparam_conv2d_16_bias_scala;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_229 <= _stream_conv2d_16_constant_5_next_constant_data;
      end 
      _set_flag_463 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_463 <= 1;
      end 
      if(_set_flag_463) begin
        _stream_conv2d_16_source_6_source_mode <= 3'b10;
        _stream_conv2d_16_source_6_source_offset <= (cparam_conv2d_16_bias_num == 1)? 0 : conv2d_16_och_count_buf;
      end 
      if(_set_flag_463) begin
        _source_stream_conv2d_16_source_6_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_6_pat_stride_0 <= 0;
      end 
      if(_set_flag_463) begin
        _source_stream_conv2d_16_source_6_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_6_pat_stride_1 <= (cparam_conv2d_16_bias_num == 1)? 0 : 1;
      end 
      if(_set_flag_463) begin
        _source_stream_conv2d_16_source_6_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_6_pat_stride_2 <= 0;
      end 
      if(_set_flag_463) begin
        _source_stream_conv2d_16_source_6_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_6_pat_stride_3 <= 0;
      end 
      if(_set_flag_463) begin
        _stream_conv2d_16_source_6_source_ram_sel <= 1;
      end 
      __tmp_472_1 <= _tmp_472;
      if(__tmp_472_1) begin
        _stream_conv2d_16_source_6_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_6_source_ram_rvalid) begin
        __variable_wdata_230 <= _stream_conv2d_16_source_6_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _stream_conv2d_16_source_6_idle <= 0;
        _stream_conv2d_16_source_6_source_offset_buf <= _stream_conv2d_16_source_6_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_count_0 <= _source_stream_conv2d_16_source_6_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_count_1 <= _source_stream_conv2d_16_source_6_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_count_2 <= _source_stream_conv2d_16_source_6_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_count_3 <= _source_stream_conv2d_16_source_6_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_size_buf_0 <= _source_stream_conv2d_16_source_6_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_size_buf_1 <= _source_stream_conv2d_16_source_6_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_size_buf_2 <= _source_stream_conv2d_16_source_6_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_size_buf_3 <= _source_stream_conv2d_16_source_6_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_stride_buf_0 <= _source_stream_conv2d_16_source_6_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_stride_buf_1 <= _source_stream_conv2d_16_source_6_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_stride_buf_2 <= _source_stream_conv2d_16_source_6_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_6_pat_stride_buf_3 <= _source_stream_conv2d_16_source_6_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_6_source_pat_fsm_0 == 1) begin
        _stream_conv2d_16_source_6_source_ram_raddr <= _stream_conv2d_16_source_6_source_pat_all_offset;
        _stream_conv2d_16_source_6_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_6_source_pat_fsm_0 == 1) begin
        _source_stream_conv2d_16_source_6_pat_cur_offset_0 <= _source_stream_conv2d_16_source_6_pat_cur_offset_0 + _source_stream_conv2d_16_source_6_pat_stride_buf_0;
        _source_stream_conv2d_16_source_6_pat_count_0 <= _source_stream_conv2d_16_source_6_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_6_source_pat_fsm_0 == 1) && (_source_stream_conv2d_16_source_6_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_6_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_6_pat_count_0 <= _source_stream_conv2d_16_source_6_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_6_source_pat_fsm_0 == 1) && (_source_stream_conv2d_16_source_6_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_6_pat_cur_offset_1 <= _source_stream_conv2d_16_source_6_pat_cur_offset_1 + _source_stream_conv2d_16_source_6_pat_stride_buf_1;
        _source_stream_conv2d_16_source_6_pat_count_1 <= _source_stream_conv2d_16_source_6_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_6_source_pat_fsm_0 == 1) && (_source_stream_conv2d_16_source_6_pat_count_0 == 0) && (_source_stream_conv2d_16_source_6_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_6_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_6_pat_count_1 <= _source_stream_conv2d_16_source_6_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_6_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_16_source_6_pat_count_0 == 0) && (_source_stream_conv2d_16_source_6_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_6_pat_cur_offset_2 <= _source_stream_conv2d_16_source_6_pat_cur_offset_2 + _source_stream_conv2d_16_source_6_pat_stride_buf_2;
        _source_stream_conv2d_16_source_6_pat_count_2 <= _source_stream_conv2d_16_source_6_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_6_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_16_source_6_pat_count_0 == 0) && (_source_stream_conv2d_16_source_6_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_6_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_6_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_6_pat_count_2 <= _source_stream_conv2d_16_source_6_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_6_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_16_source_6_pat_count_0 == 0) && (_source_stream_conv2d_16_source_6_pat_count_1 == 0) && (_source_stream_conv2d_16_source_6_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_6_pat_cur_offset_3 <= _source_stream_conv2d_16_source_6_pat_cur_offset_3 + _source_stream_conv2d_16_source_6_pat_stride_buf_3;
        _source_stream_conv2d_16_source_6_pat_count_3 <= _source_stream_conv2d_16_source_6_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_6_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_16_source_6_pat_count_0 == 0) && (_source_stream_conv2d_16_source_6_pat_count_1 == 0) && (_source_stream_conv2d_16_source_6_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_6_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_6_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_6_pat_count_3 <= _source_stream_conv2d_16_source_6_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_6_source_pat_fsm_0 == 2) begin
        _stream_conv2d_16_source_6_source_ram_renable <= 0;
        _stream_conv2d_16_source_6_idle <= 1;
      end 
      _set_flag_473 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_473 <= 1;
      end 
      if(_set_flag_473) begin
        _stream_conv2d_16_constant_7_next_constant_data <= cparam_conv2d_16_scale_scala;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_236 <= _stream_conv2d_16_constant_7_next_constant_data;
      end 
      _set_flag_474 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_474 <= 1;
      end 
      if(_set_flag_474) begin
        _stream_conv2d_16_source_8_source_mode <= 3'b10;
        _stream_conv2d_16_source_8_source_offset <= (cparam_conv2d_16_scale_num == 1)? 0 : conv2d_16_och_count_buf;
      end 
      if(_set_flag_474) begin
        _source_stream_conv2d_16_source_8_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_8_pat_stride_0 <= 0;
      end 
      if(_set_flag_474) begin
        _source_stream_conv2d_16_source_8_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_8_pat_stride_1 <= (cparam_conv2d_16_scale_num == 1)? 0 : 1;
      end 
      if(_set_flag_474) begin
        _source_stream_conv2d_16_source_8_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_8_pat_stride_2 <= 0;
      end 
      if(_set_flag_474) begin
        _source_stream_conv2d_16_source_8_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_8_pat_stride_3 <= 0;
      end 
      if(_set_flag_474) begin
        _stream_conv2d_16_source_8_source_ram_sel <= 2;
      end 
      __tmp_483_1 <= _tmp_483;
      if(__tmp_483_1) begin
        _stream_conv2d_16_source_8_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_8_source_ram_rvalid) begin
        __variable_wdata_237 <= _stream_conv2d_16_source_8_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _stream_conv2d_16_source_8_idle <= 0;
        _stream_conv2d_16_source_8_source_offset_buf <= _stream_conv2d_16_source_8_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_count_0 <= _source_stream_conv2d_16_source_8_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_count_1 <= _source_stream_conv2d_16_source_8_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_count_2 <= _source_stream_conv2d_16_source_8_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_count_3 <= _source_stream_conv2d_16_source_8_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_size_buf_0 <= _source_stream_conv2d_16_source_8_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_size_buf_1 <= _source_stream_conv2d_16_source_8_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_size_buf_2 <= _source_stream_conv2d_16_source_8_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_size_buf_3 <= _source_stream_conv2d_16_source_8_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_stride_buf_0 <= _source_stream_conv2d_16_source_8_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_stride_buf_1 <= _source_stream_conv2d_16_source_8_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_stride_buf_2 <= _source_stream_conv2d_16_source_8_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_8_pat_stride_buf_3 <= _source_stream_conv2d_16_source_8_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_8_source_pat_fsm_1 == 1) begin
        _stream_conv2d_16_source_8_source_ram_raddr <= _stream_conv2d_16_source_8_source_pat_all_offset;
        _stream_conv2d_16_source_8_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_8_source_pat_fsm_1 == 1) begin
        _source_stream_conv2d_16_source_8_pat_cur_offset_0 <= _source_stream_conv2d_16_source_8_pat_cur_offset_0 + _source_stream_conv2d_16_source_8_pat_stride_buf_0;
        _source_stream_conv2d_16_source_8_pat_count_0 <= _source_stream_conv2d_16_source_8_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_8_source_pat_fsm_1 == 1) && (_source_stream_conv2d_16_source_8_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_8_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_8_pat_count_0 <= _source_stream_conv2d_16_source_8_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_8_source_pat_fsm_1 == 1) && (_source_stream_conv2d_16_source_8_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_8_pat_cur_offset_1 <= _source_stream_conv2d_16_source_8_pat_cur_offset_1 + _source_stream_conv2d_16_source_8_pat_stride_buf_1;
        _source_stream_conv2d_16_source_8_pat_count_1 <= _source_stream_conv2d_16_source_8_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_8_source_pat_fsm_1 == 1) && (_source_stream_conv2d_16_source_8_pat_count_0 == 0) && (_source_stream_conv2d_16_source_8_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_8_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_8_pat_count_1 <= _source_stream_conv2d_16_source_8_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_8_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_16_source_8_pat_count_0 == 0) && (_source_stream_conv2d_16_source_8_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_8_pat_cur_offset_2 <= _source_stream_conv2d_16_source_8_pat_cur_offset_2 + _source_stream_conv2d_16_source_8_pat_stride_buf_2;
        _source_stream_conv2d_16_source_8_pat_count_2 <= _source_stream_conv2d_16_source_8_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_8_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_16_source_8_pat_count_0 == 0) && (_source_stream_conv2d_16_source_8_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_8_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_8_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_8_pat_count_2 <= _source_stream_conv2d_16_source_8_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_8_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_16_source_8_pat_count_0 == 0) && (_source_stream_conv2d_16_source_8_pat_count_1 == 0) && (_source_stream_conv2d_16_source_8_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_8_pat_cur_offset_3 <= _source_stream_conv2d_16_source_8_pat_cur_offset_3 + _source_stream_conv2d_16_source_8_pat_stride_buf_3;
        _source_stream_conv2d_16_source_8_pat_count_3 <= _source_stream_conv2d_16_source_8_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_8_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_16_source_8_pat_count_0 == 0) && (_source_stream_conv2d_16_source_8_pat_count_1 == 0) && (_source_stream_conv2d_16_source_8_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_8_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_8_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_8_pat_count_3 <= _source_stream_conv2d_16_source_8_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_8_source_pat_fsm_1 == 2) begin
        _stream_conv2d_16_source_8_source_ram_renable <= 0;
        _stream_conv2d_16_source_8_idle <= 1;
      end 
      _set_flag_484 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_484 <= 1;
      end 
      if(_set_flag_484) begin
        _stream_conv2d_16_constant_9_next_constant_data <= 1;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_243 <= _stream_conv2d_16_constant_9_next_constant_data;
      end 
      _set_flag_485 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_485 <= 1;
      end 
      if(_set_flag_485) begin
        _stream_conv2d_16_source_10_source_mode <= 3'b0;
        _stream_conv2d_16_source_10_source_empty_data <= 0;
      end 
      if(_stream_conv2d_16_start && !(|(_stream_conv2d_16_source_10_source_mode & 3'b0))) begin
        _stream_conv2d_16_source_10_idle <= 1;
      end 
      if(_stream_conv2d_16_start && !(|(_stream_conv2d_16_source_10_source_mode & 3'b0))) begin
        __variable_wdata_244 <= _stream_conv2d_16_source_10_source_empty_data;
      end 
      _set_flag_486 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_486 <= 1;
      end 
      if(_set_flag_486) begin
        _stream_conv2d_16_constant_11_next_constant_data <= 1;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_250 <= _stream_conv2d_16_constant_11_next_constant_data;
      end 
      _set_flag_487 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_487 <= 1;
      end 
      if(_set_flag_487) begin
        _stream_conv2d_16_source_12_source_mode <= 3'b0;
        _stream_conv2d_16_source_12_source_empty_data <= 0;
      end 
      if(_stream_conv2d_16_start && !(|(_stream_conv2d_16_source_12_source_mode & 3'b0))) begin
        _stream_conv2d_16_source_12_idle <= 1;
      end 
      if(_stream_conv2d_16_start && !(|(_stream_conv2d_16_source_12_source_mode & 3'b0))) begin
        __variable_wdata_251 <= _stream_conv2d_16_source_12_source_empty_data;
      end 
      _set_flag_488 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_488 <= 1;
      end 
      if(_set_flag_488) begin
        _stream_conv2d_16_constant_13_next_constant_data <= 1;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_257 <= _stream_conv2d_16_constant_13_next_constant_data;
      end 
      _set_flag_489 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_489 <= 1;
      end 
      if(_set_flag_489) begin
        _stream_conv2d_16_source_14_source_mode <= 3'b0;
        _stream_conv2d_16_source_14_source_empty_data <= 0;
      end 
      if(_stream_conv2d_16_start && !(|(_stream_conv2d_16_source_14_source_mode & 3'b0))) begin
        _stream_conv2d_16_source_14_idle <= 1;
      end 
      if(_stream_conv2d_16_start && !(|(_stream_conv2d_16_source_14_source_mode & 3'b0))) begin
        __variable_wdata_258 <= _stream_conv2d_16_source_14_source_empty_data;
      end 
      _set_flag_490 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_490 <= 1;
      end 
      if(_set_flag_490) begin
        _stream_conv2d_16_constant_15_next_constant_data <= cparam_conv2d_16_cshamt_mul_value;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_264 <= _stream_conv2d_16_constant_15_next_constant_data;
      end 
      _set_flag_491 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_491 <= 1;
      end 
      if(_set_flag_491) begin
        _stream_conv2d_16_constant_16_next_constant_data <= cparam_conv2d_16_cshamt_sum_value;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_265 <= _stream_conv2d_16_constant_16_next_constant_data;
      end 
      _set_flag_492 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_492 <= 1;
      end 
      if(_set_flag_492) begin
        _stream_conv2d_16_constant_17_next_constant_data <= cparam_conv2d_16_cshamt_out_value;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_266 <= _stream_conv2d_16_constant_17_next_constant_data;
      end 
      _set_flag_493 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_493 <= 1;
      end 
      if(_set_flag_493) begin
        _stream_conv2d_16_constant_18_next_constant_data <= cparam_conv2d_16_act_func_index;
      end 
      if(_stream_conv2d_16_start) begin
        __variable_wdata_267 <= _stream_conv2d_16_constant_18_next_constant_data;
      end 
      _set_flag_494 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_494 <= 1;
      end 
      if(_set_flag_494) begin
        _stream_conv2d_16_source_19_source_mode <= 3'b10;
        _stream_conv2d_16_source_19_source_offset <= conv2d_16_stream_act_local_0 + conv2d_16_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_494) begin
        _source_stream_conv2d_16_source_19_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_19_pat_stride_0 <= 1;
      end 
      if(_set_flag_494) begin
        _source_stream_conv2d_16_source_19_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_19_pat_stride_1 <= 0;
      end 
      if(_set_flag_494) begin
        _source_stream_conv2d_16_source_19_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_19_pat_stride_2 <= 0;
      end 
      if(_set_flag_494) begin
        _source_stream_conv2d_16_source_19_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_19_pat_stride_3 <= 0;
      end 
      if(_set_flag_494) begin
        _stream_conv2d_16_source_19_source_ram_sel <= 3;
      end 
      __tmp_503_1 <= _tmp_503;
      if(__tmp_503_1) begin
        _stream_conv2d_16_source_19_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_19_source_ram_rvalid) begin
        __variable_wdata_268 <= _stream_conv2d_16_source_19_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _stream_conv2d_16_source_19_idle <= 0;
        _stream_conv2d_16_source_19_source_offset_buf <= _stream_conv2d_16_source_19_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_count_0 <= _source_stream_conv2d_16_source_19_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_count_1 <= _source_stream_conv2d_16_source_19_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_count_2 <= _source_stream_conv2d_16_source_19_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_count_3 <= _source_stream_conv2d_16_source_19_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_size_buf_0 <= _source_stream_conv2d_16_source_19_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_size_buf_1 <= _source_stream_conv2d_16_source_19_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_size_buf_2 <= _source_stream_conv2d_16_source_19_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_size_buf_3 <= _source_stream_conv2d_16_source_19_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_stride_buf_0 <= _source_stream_conv2d_16_source_19_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_stride_buf_1 <= _source_stream_conv2d_16_source_19_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_stride_buf_2 <= _source_stream_conv2d_16_source_19_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_19_pat_stride_buf_3 <= _source_stream_conv2d_16_source_19_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_19_source_pat_fsm_2 == 1) begin
        _stream_conv2d_16_source_19_source_ram_raddr <= _stream_conv2d_16_source_19_source_pat_all_offset;
        _stream_conv2d_16_source_19_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_19_source_pat_fsm_2 == 1) begin
        _source_stream_conv2d_16_source_19_pat_cur_offset_0 <= _source_stream_conv2d_16_source_19_pat_cur_offset_0 + _source_stream_conv2d_16_source_19_pat_stride_buf_0;
        _source_stream_conv2d_16_source_19_pat_count_0 <= _source_stream_conv2d_16_source_19_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_19_source_pat_fsm_2 == 1) && (_source_stream_conv2d_16_source_19_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_19_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_19_pat_count_0 <= _source_stream_conv2d_16_source_19_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_19_source_pat_fsm_2 == 1) && (_source_stream_conv2d_16_source_19_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_19_pat_cur_offset_1 <= _source_stream_conv2d_16_source_19_pat_cur_offset_1 + _source_stream_conv2d_16_source_19_pat_stride_buf_1;
        _source_stream_conv2d_16_source_19_pat_count_1 <= _source_stream_conv2d_16_source_19_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_19_source_pat_fsm_2 == 1) && (_source_stream_conv2d_16_source_19_pat_count_0 == 0) && (_source_stream_conv2d_16_source_19_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_19_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_19_pat_count_1 <= _source_stream_conv2d_16_source_19_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_19_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_16_source_19_pat_count_0 == 0) && (_source_stream_conv2d_16_source_19_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_19_pat_cur_offset_2 <= _source_stream_conv2d_16_source_19_pat_cur_offset_2 + _source_stream_conv2d_16_source_19_pat_stride_buf_2;
        _source_stream_conv2d_16_source_19_pat_count_2 <= _source_stream_conv2d_16_source_19_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_19_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_16_source_19_pat_count_0 == 0) && (_source_stream_conv2d_16_source_19_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_19_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_19_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_19_pat_count_2 <= _source_stream_conv2d_16_source_19_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_19_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_16_source_19_pat_count_0 == 0) && (_source_stream_conv2d_16_source_19_pat_count_1 == 0) && (_source_stream_conv2d_16_source_19_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_19_pat_cur_offset_3 <= _source_stream_conv2d_16_source_19_pat_cur_offset_3 + _source_stream_conv2d_16_source_19_pat_stride_buf_3;
        _source_stream_conv2d_16_source_19_pat_count_3 <= _source_stream_conv2d_16_source_19_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_19_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_16_source_19_pat_count_0 == 0) && (_source_stream_conv2d_16_source_19_pat_count_1 == 0) && (_source_stream_conv2d_16_source_19_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_19_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_19_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_19_pat_count_3 <= _source_stream_conv2d_16_source_19_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_19_source_pat_fsm_2 == 2) begin
        _stream_conv2d_16_source_19_source_ram_renable <= 0;
        _stream_conv2d_16_source_19_idle <= 1;
      end 
      _set_flag_504 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_504 <= 1;
      end 
      if(_set_flag_504) begin
        _stream_conv2d_16_source_20_source_mode <= 3'b10;
        _stream_conv2d_16_source_20_source_offset <= conv2d_16_stream_act_local_1 + conv2d_16_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_504) begin
        _source_stream_conv2d_16_source_20_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_504) begin
        _source_stream_conv2d_16_source_20_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_20_pat_stride_1 <= 0;
      end 
      if(_set_flag_504) begin
        _source_stream_conv2d_16_source_20_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_504) begin
        _source_stream_conv2d_16_source_20_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_504) begin
        _stream_conv2d_16_source_20_source_ram_sel <= 4;
      end 
      __tmp_513_1 <= _tmp_513;
      if(__tmp_513_1) begin
        _stream_conv2d_16_source_20_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_20_source_ram_rvalid) begin
        __variable_wdata_269 <= _stream_conv2d_16_source_20_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _stream_conv2d_16_source_20_idle <= 0;
        _stream_conv2d_16_source_20_source_offset_buf <= _stream_conv2d_16_source_20_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_count_0 <= _source_stream_conv2d_16_source_20_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_count_1 <= _source_stream_conv2d_16_source_20_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_count_2 <= _source_stream_conv2d_16_source_20_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_count_3 <= _source_stream_conv2d_16_source_20_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_size_buf_0 <= _source_stream_conv2d_16_source_20_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_size_buf_1 <= _source_stream_conv2d_16_source_20_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_size_buf_2 <= _source_stream_conv2d_16_source_20_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_size_buf_3 <= _source_stream_conv2d_16_source_20_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_stride_buf_0 <= _source_stream_conv2d_16_source_20_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_stride_buf_1 <= _source_stream_conv2d_16_source_20_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_stride_buf_2 <= _source_stream_conv2d_16_source_20_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_20_pat_stride_buf_3 <= _source_stream_conv2d_16_source_20_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_20_source_pat_fsm_3 == 1) begin
        _stream_conv2d_16_source_20_source_ram_raddr <= _stream_conv2d_16_source_20_source_pat_all_offset;
        _stream_conv2d_16_source_20_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_20_source_pat_fsm_3 == 1) begin
        _source_stream_conv2d_16_source_20_pat_cur_offset_0 <= _source_stream_conv2d_16_source_20_pat_cur_offset_0 + _source_stream_conv2d_16_source_20_pat_stride_buf_0;
        _source_stream_conv2d_16_source_20_pat_count_0 <= _source_stream_conv2d_16_source_20_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_20_source_pat_fsm_3 == 1) && (_source_stream_conv2d_16_source_20_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_20_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_20_pat_count_0 <= _source_stream_conv2d_16_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_20_source_pat_fsm_3 == 1) && (_source_stream_conv2d_16_source_20_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_20_pat_cur_offset_1 <= _source_stream_conv2d_16_source_20_pat_cur_offset_1 + _source_stream_conv2d_16_source_20_pat_stride_buf_1;
        _source_stream_conv2d_16_source_20_pat_count_1 <= _source_stream_conv2d_16_source_20_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_20_source_pat_fsm_3 == 1) && (_source_stream_conv2d_16_source_20_pat_count_0 == 0) && (_source_stream_conv2d_16_source_20_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_20_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_20_pat_count_1 <= _source_stream_conv2d_16_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_20_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_16_source_20_pat_count_0 == 0) && (_source_stream_conv2d_16_source_20_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_20_pat_cur_offset_2 <= _source_stream_conv2d_16_source_20_pat_cur_offset_2 + _source_stream_conv2d_16_source_20_pat_stride_buf_2;
        _source_stream_conv2d_16_source_20_pat_count_2 <= _source_stream_conv2d_16_source_20_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_20_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_16_source_20_pat_count_0 == 0) && (_source_stream_conv2d_16_source_20_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_20_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_20_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_20_pat_count_2 <= _source_stream_conv2d_16_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_20_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_16_source_20_pat_count_0 == 0) && (_source_stream_conv2d_16_source_20_pat_count_1 == 0) && (_source_stream_conv2d_16_source_20_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_20_pat_cur_offset_3 <= _source_stream_conv2d_16_source_20_pat_cur_offset_3 + _source_stream_conv2d_16_source_20_pat_stride_buf_3;
        _source_stream_conv2d_16_source_20_pat_count_3 <= _source_stream_conv2d_16_source_20_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_20_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_16_source_20_pat_count_0 == 0) && (_source_stream_conv2d_16_source_20_pat_count_1 == 0) && (_source_stream_conv2d_16_source_20_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_20_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_20_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_20_pat_count_3 <= _source_stream_conv2d_16_source_20_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_20_source_pat_fsm_3 == 2) begin
        _stream_conv2d_16_source_20_source_ram_renable <= 0;
        _stream_conv2d_16_source_20_idle <= 1;
      end 
      _set_flag_514 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_514 <= 1;
      end 
      if(_set_flag_514) begin
        _stream_conv2d_16_source_21_source_mode <= 3'b10;
        _stream_conv2d_16_source_21_source_offset <= conv2d_16_stream_act_local_2 + conv2d_16_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_514) begin
        _source_stream_conv2d_16_source_21_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_21_pat_stride_0 <= 1;
      end 
      if(_set_flag_514) begin
        _source_stream_conv2d_16_source_21_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_21_pat_stride_1 <= 0;
      end 
      if(_set_flag_514) begin
        _source_stream_conv2d_16_source_21_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_21_pat_stride_2 <= 0;
      end 
      if(_set_flag_514) begin
        _source_stream_conv2d_16_source_21_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_21_pat_stride_3 <= 0;
      end 
      if(_set_flag_514) begin
        _stream_conv2d_16_source_21_source_ram_sel <= 5;
      end 
      __tmp_523_1 <= _tmp_523;
      if(__tmp_523_1) begin
        _stream_conv2d_16_source_21_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_21_source_ram_rvalid) begin
        __variable_wdata_270 <= _stream_conv2d_16_source_21_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _stream_conv2d_16_source_21_idle <= 0;
        _stream_conv2d_16_source_21_source_offset_buf <= _stream_conv2d_16_source_21_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_count_0 <= _source_stream_conv2d_16_source_21_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_count_1 <= _source_stream_conv2d_16_source_21_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_count_2 <= _source_stream_conv2d_16_source_21_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_count_3 <= _source_stream_conv2d_16_source_21_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_size_buf_0 <= _source_stream_conv2d_16_source_21_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_size_buf_1 <= _source_stream_conv2d_16_source_21_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_size_buf_2 <= _source_stream_conv2d_16_source_21_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_size_buf_3 <= _source_stream_conv2d_16_source_21_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_stride_buf_0 <= _source_stream_conv2d_16_source_21_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_stride_buf_1 <= _source_stream_conv2d_16_source_21_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_stride_buf_2 <= _source_stream_conv2d_16_source_21_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_21_pat_stride_buf_3 <= _source_stream_conv2d_16_source_21_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_21_source_pat_fsm_4 == 1) begin
        _stream_conv2d_16_source_21_source_ram_raddr <= _stream_conv2d_16_source_21_source_pat_all_offset;
        _stream_conv2d_16_source_21_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_21_source_pat_fsm_4 == 1) begin
        _source_stream_conv2d_16_source_21_pat_cur_offset_0 <= _source_stream_conv2d_16_source_21_pat_cur_offset_0 + _source_stream_conv2d_16_source_21_pat_stride_buf_0;
        _source_stream_conv2d_16_source_21_pat_count_0 <= _source_stream_conv2d_16_source_21_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_21_source_pat_fsm_4 == 1) && (_source_stream_conv2d_16_source_21_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_21_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_21_pat_count_0 <= _source_stream_conv2d_16_source_21_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_21_source_pat_fsm_4 == 1) && (_source_stream_conv2d_16_source_21_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_21_pat_cur_offset_1 <= _source_stream_conv2d_16_source_21_pat_cur_offset_1 + _source_stream_conv2d_16_source_21_pat_stride_buf_1;
        _source_stream_conv2d_16_source_21_pat_count_1 <= _source_stream_conv2d_16_source_21_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_21_source_pat_fsm_4 == 1) && (_source_stream_conv2d_16_source_21_pat_count_0 == 0) && (_source_stream_conv2d_16_source_21_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_21_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_21_pat_count_1 <= _source_stream_conv2d_16_source_21_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_21_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_16_source_21_pat_count_0 == 0) && (_source_stream_conv2d_16_source_21_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_21_pat_cur_offset_2 <= _source_stream_conv2d_16_source_21_pat_cur_offset_2 + _source_stream_conv2d_16_source_21_pat_stride_buf_2;
        _source_stream_conv2d_16_source_21_pat_count_2 <= _source_stream_conv2d_16_source_21_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_21_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_16_source_21_pat_count_0 == 0) && (_source_stream_conv2d_16_source_21_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_21_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_21_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_21_pat_count_2 <= _source_stream_conv2d_16_source_21_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_21_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_16_source_21_pat_count_0 == 0) && (_source_stream_conv2d_16_source_21_pat_count_1 == 0) && (_source_stream_conv2d_16_source_21_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_21_pat_cur_offset_3 <= _source_stream_conv2d_16_source_21_pat_cur_offset_3 + _source_stream_conv2d_16_source_21_pat_stride_buf_3;
        _source_stream_conv2d_16_source_21_pat_count_3 <= _source_stream_conv2d_16_source_21_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_21_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_16_source_21_pat_count_0 == 0) && (_source_stream_conv2d_16_source_21_pat_count_1 == 0) && (_source_stream_conv2d_16_source_21_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_21_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_21_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_21_pat_count_3 <= _source_stream_conv2d_16_source_21_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_21_source_pat_fsm_4 == 2) begin
        _stream_conv2d_16_source_21_source_ram_renable <= 0;
        _stream_conv2d_16_source_21_idle <= 1;
      end 
      _set_flag_524 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_524 <= 1;
      end 
      if(_set_flag_524) begin
        _stream_conv2d_16_source_22_source_mode <= 3'b10;
        _stream_conv2d_16_source_22_source_offset <= conv2d_16_stream_act_local_3 + conv2d_16_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_524) begin
        _source_stream_conv2d_16_source_22_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_22_pat_stride_0 <= 1;
      end 
      if(_set_flag_524) begin
        _source_stream_conv2d_16_source_22_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_22_pat_stride_1 <= 0;
      end 
      if(_set_flag_524) begin
        _source_stream_conv2d_16_source_22_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_22_pat_stride_2 <= 0;
      end 
      if(_set_flag_524) begin
        _source_stream_conv2d_16_source_22_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_22_pat_stride_3 <= 0;
      end 
      if(_set_flag_524) begin
        _stream_conv2d_16_source_22_source_ram_sel <= 6;
      end 
      __tmp_533_1 <= _tmp_533;
      if(__tmp_533_1) begin
        _stream_conv2d_16_source_22_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_22_source_ram_rvalid) begin
        __variable_wdata_271 <= _stream_conv2d_16_source_22_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _stream_conv2d_16_source_22_idle <= 0;
        _stream_conv2d_16_source_22_source_offset_buf <= _stream_conv2d_16_source_22_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_count_0 <= _source_stream_conv2d_16_source_22_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_count_1 <= _source_stream_conv2d_16_source_22_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_count_2 <= _source_stream_conv2d_16_source_22_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_count_3 <= _source_stream_conv2d_16_source_22_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_size_buf_0 <= _source_stream_conv2d_16_source_22_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_size_buf_1 <= _source_stream_conv2d_16_source_22_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_size_buf_2 <= _source_stream_conv2d_16_source_22_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_size_buf_3 <= _source_stream_conv2d_16_source_22_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_stride_buf_0 <= _source_stream_conv2d_16_source_22_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_stride_buf_1 <= _source_stream_conv2d_16_source_22_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_stride_buf_2 <= _source_stream_conv2d_16_source_22_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_22_pat_stride_buf_3 <= _source_stream_conv2d_16_source_22_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_22_source_pat_fsm_5 == 1) begin
        _stream_conv2d_16_source_22_source_ram_raddr <= _stream_conv2d_16_source_22_source_pat_all_offset;
        _stream_conv2d_16_source_22_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_22_source_pat_fsm_5 == 1) begin
        _source_stream_conv2d_16_source_22_pat_cur_offset_0 <= _source_stream_conv2d_16_source_22_pat_cur_offset_0 + _source_stream_conv2d_16_source_22_pat_stride_buf_0;
        _source_stream_conv2d_16_source_22_pat_count_0 <= _source_stream_conv2d_16_source_22_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_22_source_pat_fsm_5 == 1) && (_source_stream_conv2d_16_source_22_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_22_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_22_pat_count_0 <= _source_stream_conv2d_16_source_22_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_22_source_pat_fsm_5 == 1) && (_source_stream_conv2d_16_source_22_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_22_pat_cur_offset_1 <= _source_stream_conv2d_16_source_22_pat_cur_offset_1 + _source_stream_conv2d_16_source_22_pat_stride_buf_1;
        _source_stream_conv2d_16_source_22_pat_count_1 <= _source_stream_conv2d_16_source_22_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_22_source_pat_fsm_5 == 1) && (_source_stream_conv2d_16_source_22_pat_count_0 == 0) && (_source_stream_conv2d_16_source_22_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_22_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_22_pat_count_1 <= _source_stream_conv2d_16_source_22_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_22_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_16_source_22_pat_count_0 == 0) && (_source_stream_conv2d_16_source_22_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_22_pat_cur_offset_2 <= _source_stream_conv2d_16_source_22_pat_cur_offset_2 + _source_stream_conv2d_16_source_22_pat_stride_buf_2;
        _source_stream_conv2d_16_source_22_pat_count_2 <= _source_stream_conv2d_16_source_22_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_22_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_16_source_22_pat_count_0 == 0) && (_source_stream_conv2d_16_source_22_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_22_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_22_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_22_pat_count_2 <= _source_stream_conv2d_16_source_22_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_22_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_16_source_22_pat_count_0 == 0) && (_source_stream_conv2d_16_source_22_pat_count_1 == 0) && (_source_stream_conv2d_16_source_22_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_22_pat_cur_offset_3 <= _source_stream_conv2d_16_source_22_pat_cur_offset_3 + _source_stream_conv2d_16_source_22_pat_stride_buf_3;
        _source_stream_conv2d_16_source_22_pat_count_3 <= _source_stream_conv2d_16_source_22_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_22_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_16_source_22_pat_count_0 == 0) && (_source_stream_conv2d_16_source_22_pat_count_1 == 0) && (_source_stream_conv2d_16_source_22_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_22_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_22_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_22_pat_count_3 <= _source_stream_conv2d_16_source_22_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_22_source_pat_fsm_5 == 2) begin
        _stream_conv2d_16_source_22_source_ram_renable <= 0;
        _stream_conv2d_16_source_22_idle <= 1;
      end 
      _set_flag_534 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_534 <= 1;
      end 
      if(_set_flag_534) begin
        _stream_conv2d_16_source_23_source_mode <= 3'b10;
        _stream_conv2d_16_source_23_source_offset <= conv2d_16_stream_act_local_4 + conv2d_16_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_534) begin
        _source_stream_conv2d_16_source_23_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_23_pat_stride_0 <= 1;
      end 
      if(_set_flag_534) begin
        _source_stream_conv2d_16_source_23_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_23_pat_stride_1 <= 0;
      end 
      if(_set_flag_534) begin
        _source_stream_conv2d_16_source_23_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_23_pat_stride_2 <= 0;
      end 
      if(_set_flag_534) begin
        _source_stream_conv2d_16_source_23_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_23_pat_stride_3 <= 0;
      end 
      if(_set_flag_534) begin
        _stream_conv2d_16_source_23_source_ram_sel <= 7;
      end 
      __tmp_543_1 <= _tmp_543;
      if(__tmp_543_1) begin
        _stream_conv2d_16_source_23_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_23_source_ram_rvalid) begin
        __variable_wdata_272 <= _stream_conv2d_16_source_23_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _stream_conv2d_16_source_23_idle <= 0;
        _stream_conv2d_16_source_23_source_offset_buf <= _stream_conv2d_16_source_23_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_count_0 <= _source_stream_conv2d_16_source_23_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_count_1 <= _source_stream_conv2d_16_source_23_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_count_2 <= _source_stream_conv2d_16_source_23_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_count_3 <= _source_stream_conv2d_16_source_23_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_size_buf_0 <= _source_stream_conv2d_16_source_23_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_size_buf_1 <= _source_stream_conv2d_16_source_23_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_size_buf_2 <= _source_stream_conv2d_16_source_23_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_size_buf_3 <= _source_stream_conv2d_16_source_23_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_stride_buf_0 <= _source_stream_conv2d_16_source_23_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_stride_buf_1 <= _source_stream_conv2d_16_source_23_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_stride_buf_2 <= _source_stream_conv2d_16_source_23_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_23_pat_stride_buf_3 <= _source_stream_conv2d_16_source_23_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_23_source_pat_fsm_6 == 1) begin
        _stream_conv2d_16_source_23_source_ram_raddr <= _stream_conv2d_16_source_23_source_pat_all_offset;
        _stream_conv2d_16_source_23_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_23_source_pat_fsm_6 == 1) begin
        _source_stream_conv2d_16_source_23_pat_cur_offset_0 <= _source_stream_conv2d_16_source_23_pat_cur_offset_0 + _source_stream_conv2d_16_source_23_pat_stride_buf_0;
        _source_stream_conv2d_16_source_23_pat_count_0 <= _source_stream_conv2d_16_source_23_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_23_source_pat_fsm_6 == 1) && (_source_stream_conv2d_16_source_23_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_23_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_23_pat_count_0 <= _source_stream_conv2d_16_source_23_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_23_source_pat_fsm_6 == 1) && (_source_stream_conv2d_16_source_23_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_23_pat_cur_offset_1 <= _source_stream_conv2d_16_source_23_pat_cur_offset_1 + _source_stream_conv2d_16_source_23_pat_stride_buf_1;
        _source_stream_conv2d_16_source_23_pat_count_1 <= _source_stream_conv2d_16_source_23_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_23_source_pat_fsm_6 == 1) && (_source_stream_conv2d_16_source_23_pat_count_0 == 0) && (_source_stream_conv2d_16_source_23_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_23_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_23_pat_count_1 <= _source_stream_conv2d_16_source_23_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_23_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_16_source_23_pat_count_0 == 0) && (_source_stream_conv2d_16_source_23_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_23_pat_cur_offset_2 <= _source_stream_conv2d_16_source_23_pat_cur_offset_2 + _source_stream_conv2d_16_source_23_pat_stride_buf_2;
        _source_stream_conv2d_16_source_23_pat_count_2 <= _source_stream_conv2d_16_source_23_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_23_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_16_source_23_pat_count_0 == 0) && (_source_stream_conv2d_16_source_23_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_23_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_23_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_23_pat_count_2 <= _source_stream_conv2d_16_source_23_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_23_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_16_source_23_pat_count_0 == 0) && (_source_stream_conv2d_16_source_23_pat_count_1 == 0) && (_source_stream_conv2d_16_source_23_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_23_pat_cur_offset_3 <= _source_stream_conv2d_16_source_23_pat_cur_offset_3 + _source_stream_conv2d_16_source_23_pat_stride_buf_3;
        _source_stream_conv2d_16_source_23_pat_count_3 <= _source_stream_conv2d_16_source_23_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_23_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_16_source_23_pat_count_0 == 0) && (_source_stream_conv2d_16_source_23_pat_count_1 == 0) && (_source_stream_conv2d_16_source_23_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_23_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_23_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_23_pat_count_3 <= _source_stream_conv2d_16_source_23_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_23_source_pat_fsm_6 == 2) begin
        _stream_conv2d_16_source_23_source_ram_renable <= 0;
        _stream_conv2d_16_source_23_idle <= 1;
      end 
      _set_flag_544 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_544 <= 1;
      end 
      if(_set_flag_544) begin
        _stream_conv2d_16_source_24_source_mode <= 3'b10;
        _stream_conv2d_16_source_24_source_offset <= conv2d_16_stream_act_local_5 + conv2d_16_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_544) begin
        _source_stream_conv2d_16_source_24_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_24_pat_stride_0 <= 1;
      end 
      if(_set_flag_544) begin
        _source_stream_conv2d_16_source_24_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_24_pat_stride_1 <= 0;
      end 
      if(_set_flag_544) begin
        _source_stream_conv2d_16_source_24_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_24_pat_stride_2 <= 0;
      end 
      if(_set_flag_544) begin
        _source_stream_conv2d_16_source_24_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_24_pat_stride_3 <= 0;
      end 
      if(_set_flag_544) begin
        _stream_conv2d_16_source_24_source_ram_sel <= 8;
      end 
      __tmp_553_1 <= _tmp_553;
      if(__tmp_553_1) begin
        _stream_conv2d_16_source_24_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_24_source_ram_rvalid) begin
        __variable_wdata_273 <= _stream_conv2d_16_source_24_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _stream_conv2d_16_source_24_idle <= 0;
        _stream_conv2d_16_source_24_source_offset_buf <= _stream_conv2d_16_source_24_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_count_0 <= _source_stream_conv2d_16_source_24_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_count_1 <= _source_stream_conv2d_16_source_24_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_count_2 <= _source_stream_conv2d_16_source_24_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_count_3 <= _source_stream_conv2d_16_source_24_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_size_buf_0 <= _source_stream_conv2d_16_source_24_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_size_buf_1 <= _source_stream_conv2d_16_source_24_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_size_buf_2 <= _source_stream_conv2d_16_source_24_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_size_buf_3 <= _source_stream_conv2d_16_source_24_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_stride_buf_0 <= _source_stream_conv2d_16_source_24_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_stride_buf_1 <= _source_stream_conv2d_16_source_24_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_stride_buf_2 <= _source_stream_conv2d_16_source_24_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_24_pat_stride_buf_3 <= _source_stream_conv2d_16_source_24_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_24_source_pat_fsm_7 == 1) begin
        _stream_conv2d_16_source_24_source_ram_raddr <= _stream_conv2d_16_source_24_source_pat_all_offset;
        _stream_conv2d_16_source_24_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_24_source_pat_fsm_7 == 1) begin
        _source_stream_conv2d_16_source_24_pat_cur_offset_0 <= _source_stream_conv2d_16_source_24_pat_cur_offset_0 + _source_stream_conv2d_16_source_24_pat_stride_buf_0;
        _source_stream_conv2d_16_source_24_pat_count_0 <= _source_stream_conv2d_16_source_24_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_24_source_pat_fsm_7 == 1) && (_source_stream_conv2d_16_source_24_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_24_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_24_pat_count_0 <= _source_stream_conv2d_16_source_24_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_24_source_pat_fsm_7 == 1) && (_source_stream_conv2d_16_source_24_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_24_pat_cur_offset_1 <= _source_stream_conv2d_16_source_24_pat_cur_offset_1 + _source_stream_conv2d_16_source_24_pat_stride_buf_1;
        _source_stream_conv2d_16_source_24_pat_count_1 <= _source_stream_conv2d_16_source_24_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_24_source_pat_fsm_7 == 1) && (_source_stream_conv2d_16_source_24_pat_count_0 == 0) && (_source_stream_conv2d_16_source_24_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_24_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_24_pat_count_1 <= _source_stream_conv2d_16_source_24_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_24_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_16_source_24_pat_count_0 == 0) && (_source_stream_conv2d_16_source_24_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_24_pat_cur_offset_2 <= _source_stream_conv2d_16_source_24_pat_cur_offset_2 + _source_stream_conv2d_16_source_24_pat_stride_buf_2;
        _source_stream_conv2d_16_source_24_pat_count_2 <= _source_stream_conv2d_16_source_24_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_24_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_16_source_24_pat_count_0 == 0) && (_source_stream_conv2d_16_source_24_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_24_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_24_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_24_pat_count_2 <= _source_stream_conv2d_16_source_24_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_24_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_16_source_24_pat_count_0 == 0) && (_source_stream_conv2d_16_source_24_pat_count_1 == 0) && (_source_stream_conv2d_16_source_24_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_24_pat_cur_offset_3 <= _source_stream_conv2d_16_source_24_pat_cur_offset_3 + _source_stream_conv2d_16_source_24_pat_stride_buf_3;
        _source_stream_conv2d_16_source_24_pat_count_3 <= _source_stream_conv2d_16_source_24_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_24_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_16_source_24_pat_count_0 == 0) && (_source_stream_conv2d_16_source_24_pat_count_1 == 0) && (_source_stream_conv2d_16_source_24_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_24_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_24_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_24_pat_count_3 <= _source_stream_conv2d_16_source_24_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_24_source_pat_fsm_7 == 2) begin
        _stream_conv2d_16_source_24_source_ram_renable <= 0;
        _stream_conv2d_16_source_24_idle <= 1;
      end 
      _set_flag_554 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_554 <= 1;
      end 
      if(_set_flag_554) begin
        _stream_conv2d_16_source_25_source_mode <= 3'b10;
        _stream_conv2d_16_source_25_source_offset <= conv2d_16_stream_act_local_6 + conv2d_16_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_554) begin
        _source_stream_conv2d_16_source_25_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_25_pat_stride_0 <= 1;
      end 
      if(_set_flag_554) begin
        _source_stream_conv2d_16_source_25_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_25_pat_stride_1 <= 0;
      end 
      if(_set_flag_554) begin
        _source_stream_conv2d_16_source_25_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_25_pat_stride_2 <= 0;
      end 
      if(_set_flag_554) begin
        _source_stream_conv2d_16_source_25_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_25_pat_stride_3 <= 0;
      end 
      if(_set_flag_554) begin
        _stream_conv2d_16_source_25_source_ram_sel <= 9;
      end 
      __tmp_563_1 <= _tmp_563;
      if(__tmp_563_1) begin
        _stream_conv2d_16_source_25_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_25_source_ram_rvalid) begin
        __variable_wdata_274 <= _stream_conv2d_16_source_25_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _stream_conv2d_16_source_25_idle <= 0;
        _stream_conv2d_16_source_25_source_offset_buf <= _stream_conv2d_16_source_25_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_count_0 <= _source_stream_conv2d_16_source_25_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_count_1 <= _source_stream_conv2d_16_source_25_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_count_2 <= _source_stream_conv2d_16_source_25_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_count_3 <= _source_stream_conv2d_16_source_25_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_size_buf_0 <= _source_stream_conv2d_16_source_25_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_size_buf_1 <= _source_stream_conv2d_16_source_25_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_size_buf_2 <= _source_stream_conv2d_16_source_25_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_size_buf_3 <= _source_stream_conv2d_16_source_25_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_stride_buf_0 <= _source_stream_conv2d_16_source_25_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_stride_buf_1 <= _source_stream_conv2d_16_source_25_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_stride_buf_2 <= _source_stream_conv2d_16_source_25_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_25_pat_stride_buf_3 <= _source_stream_conv2d_16_source_25_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_25_source_pat_fsm_8 == 1) begin
        _stream_conv2d_16_source_25_source_ram_raddr <= _stream_conv2d_16_source_25_source_pat_all_offset;
        _stream_conv2d_16_source_25_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_25_source_pat_fsm_8 == 1) begin
        _source_stream_conv2d_16_source_25_pat_cur_offset_0 <= _source_stream_conv2d_16_source_25_pat_cur_offset_0 + _source_stream_conv2d_16_source_25_pat_stride_buf_0;
        _source_stream_conv2d_16_source_25_pat_count_0 <= _source_stream_conv2d_16_source_25_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_25_source_pat_fsm_8 == 1) && (_source_stream_conv2d_16_source_25_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_25_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_25_pat_count_0 <= _source_stream_conv2d_16_source_25_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_25_source_pat_fsm_8 == 1) && (_source_stream_conv2d_16_source_25_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_25_pat_cur_offset_1 <= _source_stream_conv2d_16_source_25_pat_cur_offset_1 + _source_stream_conv2d_16_source_25_pat_stride_buf_1;
        _source_stream_conv2d_16_source_25_pat_count_1 <= _source_stream_conv2d_16_source_25_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_25_source_pat_fsm_8 == 1) && (_source_stream_conv2d_16_source_25_pat_count_0 == 0) && (_source_stream_conv2d_16_source_25_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_25_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_25_pat_count_1 <= _source_stream_conv2d_16_source_25_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_25_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_16_source_25_pat_count_0 == 0) && (_source_stream_conv2d_16_source_25_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_25_pat_cur_offset_2 <= _source_stream_conv2d_16_source_25_pat_cur_offset_2 + _source_stream_conv2d_16_source_25_pat_stride_buf_2;
        _source_stream_conv2d_16_source_25_pat_count_2 <= _source_stream_conv2d_16_source_25_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_25_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_16_source_25_pat_count_0 == 0) && (_source_stream_conv2d_16_source_25_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_25_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_25_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_25_pat_count_2 <= _source_stream_conv2d_16_source_25_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_25_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_16_source_25_pat_count_0 == 0) && (_source_stream_conv2d_16_source_25_pat_count_1 == 0) && (_source_stream_conv2d_16_source_25_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_25_pat_cur_offset_3 <= _source_stream_conv2d_16_source_25_pat_cur_offset_3 + _source_stream_conv2d_16_source_25_pat_stride_buf_3;
        _source_stream_conv2d_16_source_25_pat_count_3 <= _source_stream_conv2d_16_source_25_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_25_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_16_source_25_pat_count_0 == 0) && (_source_stream_conv2d_16_source_25_pat_count_1 == 0) && (_source_stream_conv2d_16_source_25_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_25_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_25_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_25_pat_count_3 <= _source_stream_conv2d_16_source_25_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_25_source_pat_fsm_8 == 2) begin
        _stream_conv2d_16_source_25_source_ram_renable <= 0;
        _stream_conv2d_16_source_25_idle <= 1;
      end 
      _set_flag_564 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_564 <= 1;
      end 
      if(_set_flag_564) begin
        _stream_conv2d_16_source_26_source_mode <= 3'b10;
        _stream_conv2d_16_source_26_source_offset <= conv2d_16_stream_act_local_7 + conv2d_16_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_564) begin
        _source_stream_conv2d_16_source_26_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_26_pat_stride_0 <= 1;
      end 
      if(_set_flag_564) begin
        _source_stream_conv2d_16_source_26_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_26_pat_stride_1 <= 0;
      end 
      if(_set_flag_564) begin
        _source_stream_conv2d_16_source_26_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_26_pat_stride_2 <= 0;
      end 
      if(_set_flag_564) begin
        _source_stream_conv2d_16_source_26_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_26_pat_stride_3 <= 0;
      end 
      if(_set_flag_564) begin
        _stream_conv2d_16_source_26_source_ram_sel <= 10;
      end 
      __tmp_573_1 <= _tmp_573;
      if(__tmp_573_1) begin
        _stream_conv2d_16_source_26_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_26_source_ram_rvalid) begin
        __variable_wdata_275 <= _stream_conv2d_16_source_26_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _stream_conv2d_16_source_26_idle <= 0;
        _stream_conv2d_16_source_26_source_offset_buf <= _stream_conv2d_16_source_26_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_count_0 <= _source_stream_conv2d_16_source_26_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_count_1 <= _source_stream_conv2d_16_source_26_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_count_2 <= _source_stream_conv2d_16_source_26_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_count_3 <= _source_stream_conv2d_16_source_26_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_size_buf_0 <= _source_stream_conv2d_16_source_26_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_size_buf_1 <= _source_stream_conv2d_16_source_26_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_size_buf_2 <= _source_stream_conv2d_16_source_26_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_size_buf_3 <= _source_stream_conv2d_16_source_26_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_stride_buf_0 <= _source_stream_conv2d_16_source_26_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_stride_buf_1 <= _source_stream_conv2d_16_source_26_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_stride_buf_2 <= _source_stream_conv2d_16_source_26_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_26_pat_stride_buf_3 <= _source_stream_conv2d_16_source_26_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_26_source_pat_fsm_9 == 1) begin
        _stream_conv2d_16_source_26_source_ram_raddr <= _stream_conv2d_16_source_26_source_pat_all_offset;
        _stream_conv2d_16_source_26_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_26_source_pat_fsm_9 == 1) begin
        _source_stream_conv2d_16_source_26_pat_cur_offset_0 <= _source_stream_conv2d_16_source_26_pat_cur_offset_0 + _source_stream_conv2d_16_source_26_pat_stride_buf_0;
        _source_stream_conv2d_16_source_26_pat_count_0 <= _source_stream_conv2d_16_source_26_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_26_source_pat_fsm_9 == 1) && (_source_stream_conv2d_16_source_26_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_26_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_26_pat_count_0 <= _source_stream_conv2d_16_source_26_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_26_source_pat_fsm_9 == 1) && (_source_stream_conv2d_16_source_26_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_26_pat_cur_offset_1 <= _source_stream_conv2d_16_source_26_pat_cur_offset_1 + _source_stream_conv2d_16_source_26_pat_stride_buf_1;
        _source_stream_conv2d_16_source_26_pat_count_1 <= _source_stream_conv2d_16_source_26_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_26_source_pat_fsm_9 == 1) && (_source_stream_conv2d_16_source_26_pat_count_0 == 0) && (_source_stream_conv2d_16_source_26_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_26_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_26_pat_count_1 <= _source_stream_conv2d_16_source_26_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_26_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_16_source_26_pat_count_0 == 0) && (_source_stream_conv2d_16_source_26_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_26_pat_cur_offset_2 <= _source_stream_conv2d_16_source_26_pat_cur_offset_2 + _source_stream_conv2d_16_source_26_pat_stride_buf_2;
        _source_stream_conv2d_16_source_26_pat_count_2 <= _source_stream_conv2d_16_source_26_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_26_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_16_source_26_pat_count_0 == 0) && (_source_stream_conv2d_16_source_26_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_26_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_26_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_26_pat_count_2 <= _source_stream_conv2d_16_source_26_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_26_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_16_source_26_pat_count_0 == 0) && (_source_stream_conv2d_16_source_26_pat_count_1 == 0) && (_source_stream_conv2d_16_source_26_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_26_pat_cur_offset_3 <= _source_stream_conv2d_16_source_26_pat_cur_offset_3 + _source_stream_conv2d_16_source_26_pat_stride_buf_3;
        _source_stream_conv2d_16_source_26_pat_count_3 <= _source_stream_conv2d_16_source_26_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_26_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_16_source_26_pat_count_0 == 0) && (_source_stream_conv2d_16_source_26_pat_count_1 == 0) && (_source_stream_conv2d_16_source_26_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_26_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_26_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_26_pat_count_3 <= _source_stream_conv2d_16_source_26_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_26_source_pat_fsm_9 == 2) begin
        _stream_conv2d_16_source_26_source_ram_renable <= 0;
        _stream_conv2d_16_source_26_idle <= 1;
      end 
      _set_flag_574 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_574 <= 1;
      end 
      if(_set_flag_574) begin
        _stream_conv2d_16_source_27_source_mode <= 3'b10;
        _stream_conv2d_16_source_27_source_offset <= conv2d_16_stream_act_local_8 + conv2d_16_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_574) begin
        _source_stream_conv2d_16_source_27_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_27_pat_stride_0 <= 1;
      end 
      if(_set_flag_574) begin
        _source_stream_conv2d_16_source_27_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_27_pat_stride_1 <= 0;
      end 
      if(_set_flag_574) begin
        _source_stream_conv2d_16_source_27_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_27_pat_stride_2 <= 0;
      end 
      if(_set_flag_574) begin
        _source_stream_conv2d_16_source_27_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_27_pat_stride_3 <= 0;
      end 
      if(_set_flag_574) begin
        _stream_conv2d_16_source_27_source_ram_sel <= 11;
      end 
      __tmp_583_1 <= _tmp_583;
      if(__tmp_583_1) begin
        _stream_conv2d_16_source_27_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_27_source_ram_rvalid) begin
        __variable_wdata_276 <= _stream_conv2d_16_source_27_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _stream_conv2d_16_source_27_idle <= 0;
        _stream_conv2d_16_source_27_source_offset_buf <= _stream_conv2d_16_source_27_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_count_0 <= _source_stream_conv2d_16_source_27_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_count_1 <= _source_stream_conv2d_16_source_27_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_count_2 <= _source_stream_conv2d_16_source_27_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_count_3 <= _source_stream_conv2d_16_source_27_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_size_buf_0 <= _source_stream_conv2d_16_source_27_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_size_buf_1 <= _source_stream_conv2d_16_source_27_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_size_buf_2 <= _source_stream_conv2d_16_source_27_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_size_buf_3 <= _source_stream_conv2d_16_source_27_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_stride_buf_0 <= _source_stream_conv2d_16_source_27_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_stride_buf_1 <= _source_stream_conv2d_16_source_27_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_stride_buf_2 <= _source_stream_conv2d_16_source_27_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_27_pat_stride_buf_3 <= _source_stream_conv2d_16_source_27_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_27_source_pat_fsm_10 == 1) begin
        _stream_conv2d_16_source_27_source_ram_raddr <= _stream_conv2d_16_source_27_source_pat_all_offset;
        _stream_conv2d_16_source_27_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_27_source_pat_fsm_10 == 1) begin
        _source_stream_conv2d_16_source_27_pat_cur_offset_0 <= _source_stream_conv2d_16_source_27_pat_cur_offset_0 + _source_stream_conv2d_16_source_27_pat_stride_buf_0;
        _source_stream_conv2d_16_source_27_pat_count_0 <= _source_stream_conv2d_16_source_27_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_27_source_pat_fsm_10 == 1) && (_source_stream_conv2d_16_source_27_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_27_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_27_pat_count_0 <= _source_stream_conv2d_16_source_27_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_27_source_pat_fsm_10 == 1) && (_source_stream_conv2d_16_source_27_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_27_pat_cur_offset_1 <= _source_stream_conv2d_16_source_27_pat_cur_offset_1 + _source_stream_conv2d_16_source_27_pat_stride_buf_1;
        _source_stream_conv2d_16_source_27_pat_count_1 <= _source_stream_conv2d_16_source_27_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_27_source_pat_fsm_10 == 1) && (_source_stream_conv2d_16_source_27_pat_count_0 == 0) && (_source_stream_conv2d_16_source_27_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_27_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_27_pat_count_1 <= _source_stream_conv2d_16_source_27_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_27_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_16_source_27_pat_count_0 == 0) && (_source_stream_conv2d_16_source_27_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_27_pat_cur_offset_2 <= _source_stream_conv2d_16_source_27_pat_cur_offset_2 + _source_stream_conv2d_16_source_27_pat_stride_buf_2;
        _source_stream_conv2d_16_source_27_pat_count_2 <= _source_stream_conv2d_16_source_27_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_27_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_16_source_27_pat_count_0 == 0) && (_source_stream_conv2d_16_source_27_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_27_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_27_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_27_pat_count_2 <= _source_stream_conv2d_16_source_27_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_27_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_16_source_27_pat_count_0 == 0) && (_source_stream_conv2d_16_source_27_pat_count_1 == 0) && (_source_stream_conv2d_16_source_27_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_27_pat_cur_offset_3 <= _source_stream_conv2d_16_source_27_pat_cur_offset_3 + _source_stream_conv2d_16_source_27_pat_stride_buf_3;
        _source_stream_conv2d_16_source_27_pat_count_3 <= _source_stream_conv2d_16_source_27_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_27_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_16_source_27_pat_count_0 == 0) && (_source_stream_conv2d_16_source_27_pat_count_1 == 0) && (_source_stream_conv2d_16_source_27_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_27_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_27_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_27_pat_count_3 <= _source_stream_conv2d_16_source_27_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_27_source_pat_fsm_10 == 2) begin
        _stream_conv2d_16_source_27_source_ram_renable <= 0;
        _stream_conv2d_16_source_27_idle <= 1;
      end 
      _set_flag_584 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_584 <= 1;
      end 
      if(_set_flag_584) begin
        _stream_conv2d_16_source_28_source_mode <= 3'b10;
        _stream_conv2d_16_source_28_source_offset <= conv2d_16_filter_page_comp_offset_buf;
      end 
      if(_set_flag_584) begin
        _source_stream_conv2d_16_source_28_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_28_pat_stride_0 <= 1;
      end 
      if(_set_flag_584) begin
        _source_stream_conv2d_16_source_28_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_28_pat_stride_1 <= cparam_conv2d_16_stream_aligned_reduce_size;
      end 
      if(_set_flag_584) begin
        _source_stream_conv2d_16_source_28_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_28_pat_stride_2 <= 0;
      end 
      if(_set_flag_584) begin
        _source_stream_conv2d_16_source_28_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_28_pat_stride_3 <= 0;
      end 
      if(_set_flag_584) begin
        _stream_conv2d_16_source_28_source_ram_sel <= 12;
      end 
      __tmp_597_1 <= _tmp_597;
      if(__tmp_597_1) begin
        _stream_conv2d_16_source_28_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_28_source_ram_rvalid) begin
        __variable_wdata_502 <= _stream_conv2d_16_source_28_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _stream_conv2d_16_source_28_idle <= 0;
        _stream_conv2d_16_source_28_source_offset_buf <= _stream_conv2d_16_source_28_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_count_0 <= _source_stream_conv2d_16_source_28_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_count_1 <= _source_stream_conv2d_16_source_28_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_count_2 <= _source_stream_conv2d_16_source_28_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_count_3 <= _source_stream_conv2d_16_source_28_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_size_buf_0 <= _source_stream_conv2d_16_source_28_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_size_buf_1 <= _source_stream_conv2d_16_source_28_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_size_buf_2 <= _source_stream_conv2d_16_source_28_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_size_buf_3 <= _source_stream_conv2d_16_source_28_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_stride_buf_0 <= _source_stream_conv2d_16_source_28_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_stride_buf_1 <= _source_stream_conv2d_16_source_28_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_stride_buf_2 <= _source_stream_conv2d_16_source_28_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_28_pat_stride_buf_3 <= _source_stream_conv2d_16_source_28_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_28_source_pat_fsm_11 == 1) begin
        _stream_conv2d_16_source_28_source_ram_raddr <= _stream_conv2d_16_source_28_source_pat_all_offset;
        _stream_conv2d_16_source_28_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_28_source_pat_fsm_11 == 1) begin
        _source_stream_conv2d_16_source_28_pat_cur_offset_0 <= _source_stream_conv2d_16_source_28_pat_cur_offset_0 + _source_stream_conv2d_16_source_28_pat_stride_buf_0;
        _source_stream_conv2d_16_source_28_pat_count_0 <= _source_stream_conv2d_16_source_28_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_28_source_pat_fsm_11 == 1) && (_source_stream_conv2d_16_source_28_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_28_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_28_pat_count_0 <= _source_stream_conv2d_16_source_28_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_28_source_pat_fsm_11 == 1) && (_source_stream_conv2d_16_source_28_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_28_pat_cur_offset_1 <= _source_stream_conv2d_16_source_28_pat_cur_offset_1 + _source_stream_conv2d_16_source_28_pat_stride_buf_1;
        _source_stream_conv2d_16_source_28_pat_count_1 <= _source_stream_conv2d_16_source_28_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_28_source_pat_fsm_11 == 1) && (_source_stream_conv2d_16_source_28_pat_count_0 == 0) && (_source_stream_conv2d_16_source_28_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_28_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_28_pat_count_1 <= _source_stream_conv2d_16_source_28_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_28_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_16_source_28_pat_count_0 == 0) && (_source_stream_conv2d_16_source_28_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_28_pat_cur_offset_2 <= _source_stream_conv2d_16_source_28_pat_cur_offset_2 + _source_stream_conv2d_16_source_28_pat_stride_buf_2;
        _source_stream_conv2d_16_source_28_pat_count_2 <= _source_stream_conv2d_16_source_28_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_28_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_16_source_28_pat_count_0 == 0) && (_source_stream_conv2d_16_source_28_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_28_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_28_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_28_pat_count_2 <= _source_stream_conv2d_16_source_28_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_28_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_16_source_28_pat_count_0 == 0) && (_source_stream_conv2d_16_source_28_pat_count_1 == 0) && (_source_stream_conv2d_16_source_28_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_28_pat_cur_offset_3 <= _source_stream_conv2d_16_source_28_pat_cur_offset_3 + _source_stream_conv2d_16_source_28_pat_stride_buf_3;
        _source_stream_conv2d_16_source_28_pat_count_3 <= _source_stream_conv2d_16_source_28_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_28_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_16_source_28_pat_count_0 == 0) && (_source_stream_conv2d_16_source_28_pat_count_1 == 0) && (_source_stream_conv2d_16_source_28_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_28_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_28_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_28_pat_count_3 <= _source_stream_conv2d_16_source_28_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_28_source_pat_fsm_11 == 2) begin
        _stream_conv2d_16_source_28_source_ram_renable <= 0;
        _stream_conv2d_16_source_28_idle <= 1;
      end 
      _set_flag_598 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_598 <= 1;
      end 
      if(_set_flag_598) begin
        _stream_conv2d_16_source_29_source_mode <= 3'b10;
        _stream_conv2d_16_source_29_source_offset <= conv2d_16_filter_page_comp_offset_buf;
      end 
      if(_set_flag_598) begin
        _source_stream_conv2d_16_source_29_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_29_pat_stride_0 <= 1;
      end 
      if(_set_flag_598) begin
        _source_stream_conv2d_16_source_29_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_29_pat_stride_1 <= cparam_conv2d_16_stream_aligned_reduce_size;
      end 
      if(_set_flag_598) begin
        _source_stream_conv2d_16_source_29_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_29_pat_stride_2 <= 0;
      end 
      if(_set_flag_598) begin
        _source_stream_conv2d_16_source_29_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_29_pat_stride_3 <= 0;
      end 
      if(_set_flag_598) begin
        _stream_conv2d_16_source_29_source_ram_sel <= 13;
      end 
      __tmp_611_1 <= _tmp_611;
      if(__tmp_611_1) begin
        _stream_conv2d_16_source_29_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_29_source_ram_rvalid) begin
        __variable_wdata_503 <= _stream_conv2d_16_source_29_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _stream_conv2d_16_source_29_idle <= 0;
        _stream_conv2d_16_source_29_source_offset_buf <= _stream_conv2d_16_source_29_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_count_0 <= _source_stream_conv2d_16_source_29_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_count_1 <= _source_stream_conv2d_16_source_29_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_count_2 <= _source_stream_conv2d_16_source_29_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_count_3 <= _source_stream_conv2d_16_source_29_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_size_buf_0 <= _source_stream_conv2d_16_source_29_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_size_buf_1 <= _source_stream_conv2d_16_source_29_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_size_buf_2 <= _source_stream_conv2d_16_source_29_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_size_buf_3 <= _source_stream_conv2d_16_source_29_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_stride_buf_0 <= _source_stream_conv2d_16_source_29_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_stride_buf_1 <= _source_stream_conv2d_16_source_29_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_stride_buf_2 <= _source_stream_conv2d_16_source_29_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_29_pat_stride_buf_3 <= _source_stream_conv2d_16_source_29_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_29_source_pat_fsm_12 == 1) begin
        _stream_conv2d_16_source_29_source_ram_raddr <= _stream_conv2d_16_source_29_source_pat_all_offset;
        _stream_conv2d_16_source_29_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_29_source_pat_fsm_12 == 1) begin
        _source_stream_conv2d_16_source_29_pat_cur_offset_0 <= _source_stream_conv2d_16_source_29_pat_cur_offset_0 + _source_stream_conv2d_16_source_29_pat_stride_buf_0;
        _source_stream_conv2d_16_source_29_pat_count_0 <= _source_stream_conv2d_16_source_29_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_29_source_pat_fsm_12 == 1) && (_source_stream_conv2d_16_source_29_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_29_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_29_pat_count_0 <= _source_stream_conv2d_16_source_29_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_29_source_pat_fsm_12 == 1) && (_source_stream_conv2d_16_source_29_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_29_pat_cur_offset_1 <= _source_stream_conv2d_16_source_29_pat_cur_offset_1 + _source_stream_conv2d_16_source_29_pat_stride_buf_1;
        _source_stream_conv2d_16_source_29_pat_count_1 <= _source_stream_conv2d_16_source_29_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_29_source_pat_fsm_12 == 1) && (_source_stream_conv2d_16_source_29_pat_count_0 == 0) && (_source_stream_conv2d_16_source_29_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_29_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_29_pat_count_1 <= _source_stream_conv2d_16_source_29_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_29_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_16_source_29_pat_count_0 == 0) && (_source_stream_conv2d_16_source_29_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_29_pat_cur_offset_2 <= _source_stream_conv2d_16_source_29_pat_cur_offset_2 + _source_stream_conv2d_16_source_29_pat_stride_buf_2;
        _source_stream_conv2d_16_source_29_pat_count_2 <= _source_stream_conv2d_16_source_29_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_29_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_16_source_29_pat_count_0 == 0) && (_source_stream_conv2d_16_source_29_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_29_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_29_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_29_pat_count_2 <= _source_stream_conv2d_16_source_29_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_29_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_16_source_29_pat_count_0 == 0) && (_source_stream_conv2d_16_source_29_pat_count_1 == 0) && (_source_stream_conv2d_16_source_29_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_29_pat_cur_offset_3 <= _source_stream_conv2d_16_source_29_pat_cur_offset_3 + _source_stream_conv2d_16_source_29_pat_stride_buf_3;
        _source_stream_conv2d_16_source_29_pat_count_3 <= _source_stream_conv2d_16_source_29_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_29_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_16_source_29_pat_count_0 == 0) && (_source_stream_conv2d_16_source_29_pat_count_1 == 0) && (_source_stream_conv2d_16_source_29_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_29_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_29_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_29_pat_count_3 <= _source_stream_conv2d_16_source_29_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_29_source_pat_fsm_12 == 2) begin
        _stream_conv2d_16_source_29_source_ram_renable <= 0;
        _stream_conv2d_16_source_29_idle <= 1;
      end 
      _set_flag_612 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_612 <= 1;
      end 
      if(_set_flag_612) begin
        _stream_conv2d_16_source_30_source_mode <= 3'b10;
        _stream_conv2d_16_source_30_source_offset <= conv2d_16_filter_page_comp_offset_buf;
      end 
      if(_set_flag_612) begin
        _source_stream_conv2d_16_source_30_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_30_pat_stride_0 <= 1;
      end 
      if(_set_flag_612) begin
        _source_stream_conv2d_16_source_30_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_30_pat_stride_1 <= cparam_conv2d_16_stream_aligned_reduce_size;
      end 
      if(_set_flag_612) begin
        _source_stream_conv2d_16_source_30_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_30_pat_stride_2 <= 0;
      end 
      if(_set_flag_612) begin
        _source_stream_conv2d_16_source_30_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_30_pat_stride_3 <= 0;
      end 
      if(_set_flag_612) begin
        _stream_conv2d_16_source_30_source_ram_sel <= 14;
      end 
      __tmp_625_1 <= _tmp_625;
      if(__tmp_625_1) begin
        _stream_conv2d_16_source_30_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_30_source_ram_rvalid) begin
        __variable_wdata_504 <= _stream_conv2d_16_source_30_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _stream_conv2d_16_source_30_idle <= 0;
        _stream_conv2d_16_source_30_source_offset_buf <= _stream_conv2d_16_source_30_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_count_0 <= _source_stream_conv2d_16_source_30_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_count_1 <= _source_stream_conv2d_16_source_30_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_count_2 <= _source_stream_conv2d_16_source_30_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_count_3 <= _source_stream_conv2d_16_source_30_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_size_buf_0 <= _source_stream_conv2d_16_source_30_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_size_buf_1 <= _source_stream_conv2d_16_source_30_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_size_buf_2 <= _source_stream_conv2d_16_source_30_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_size_buf_3 <= _source_stream_conv2d_16_source_30_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_stride_buf_0 <= _source_stream_conv2d_16_source_30_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_stride_buf_1 <= _source_stream_conv2d_16_source_30_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_stride_buf_2 <= _source_stream_conv2d_16_source_30_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_30_pat_stride_buf_3 <= _source_stream_conv2d_16_source_30_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_30_source_pat_fsm_13 == 1) begin
        _stream_conv2d_16_source_30_source_ram_raddr <= _stream_conv2d_16_source_30_source_pat_all_offset;
        _stream_conv2d_16_source_30_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_30_source_pat_fsm_13 == 1) begin
        _source_stream_conv2d_16_source_30_pat_cur_offset_0 <= _source_stream_conv2d_16_source_30_pat_cur_offset_0 + _source_stream_conv2d_16_source_30_pat_stride_buf_0;
        _source_stream_conv2d_16_source_30_pat_count_0 <= _source_stream_conv2d_16_source_30_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_30_source_pat_fsm_13 == 1) && (_source_stream_conv2d_16_source_30_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_30_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_30_pat_count_0 <= _source_stream_conv2d_16_source_30_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_30_source_pat_fsm_13 == 1) && (_source_stream_conv2d_16_source_30_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_30_pat_cur_offset_1 <= _source_stream_conv2d_16_source_30_pat_cur_offset_1 + _source_stream_conv2d_16_source_30_pat_stride_buf_1;
        _source_stream_conv2d_16_source_30_pat_count_1 <= _source_stream_conv2d_16_source_30_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_30_source_pat_fsm_13 == 1) && (_source_stream_conv2d_16_source_30_pat_count_0 == 0) && (_source_stream_conv2d_16_source_30_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_30_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_30_pat_count_1 <= _source_stream_conv2d_16_source_30_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_30_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_16_source_30_pat_count_0 == 0) && (_source_stream_conv2d_16_source_30_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_30_pat_cur_offset_2 <= _source_stream_conv2d_16_source_30_pat_cur_offset_2 + _source_stream_conv2d_16_source_30_pat_stride_buf_2;
        _source_stream_conv2d_16_source_30_pat_count_2 <= _source_stream_conv2d_16_source_30_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_30_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_16_source_30_pat_count_0 == 0) && (_source_stream_conv2d_16_source_30_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_30_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_30_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_30_pat_count_2 <= _source_stream_conv2d_16_source_30_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_30_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_16_source_30_pat_count_0 == 0) && (_source_stream_conv2d_16_source_30_pat_count_1 == 0) && (_source_stream_conv2d_16_source_30_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_30_pat_cur_offset_3 <= _source_stream_conv2d_16_source_30_pat_cur_offset_3 + _source_stream_conv2d_16_source_30_pat_stride_buf_3;
        _source_stream_conv2d_16_source_30_pat_count_3 <= _source_stream_conv2d_16_source_30_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_30_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_16_source_30_pat_count_0 == 0) && (_source_stream_conv2d_16_source_30_pat_count_1 == 0) && (_source_stream_conv2d_16_source_30_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_30_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_30_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_30_pat_count_3 <= _source_stream_conv2d_16_source_30_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_30_source_pat_fsm_13 == 2) begin
        _stream_conv2d_16_source_30_source_ram_renable <= 0;
        _stream_conv2d_16_source_30_idle <= 1;
      end 
      _set_flag_626 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_626 <= 1;
      end 
      if(_set_flag_626) begin
        _stream_conv2d_16_source_31_source_mode <= 3'b10;
        _stream_conv2d_16_source_31_source_offset <= conv2d_16_filter_page_comp_offset_buf;
      end 
      if(_set_flag_626) begin
        _source_stream_conv2d_16_source_31_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_31_pat_stride_0 <= 1;
      end 
      if(_set_flag_626) begin
        _source_stream_conv2d_16_source_31_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_31_pat_stride_1 <= cparam_conv2d_16_stream_aligned_reduce_size;
      end 
      if(_set_flag_626) begin
        _source_stream_conv2d_16_source_31_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_31_pat_stride_2 <= 0;
      end 
      if(_set_flag_626) begin
        _source_stream_conv2d_16_source_31_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_31_pat_stride_3 <= 0;
      end 
      if(_set_flag_626) begin
        _stream_conv2d_16_source_31_source_ram_sel <= 15;
      end 
      __tmp_639_1 <= _tmp_639;
      if(__tmp_639_1) begin
        _stream_conv2d_16_source_31_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_31_source_ram_rvalid) begin
        __variable_wdata_505 <= _stream_conv2d_16_source_31_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _stream_conv2d_16_source_31_idle <= 0;
        _stream_conv2d_16_source_31_source_offset_buf <= _stream_conv2d_16_source_31_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_count_0 <= _source_stream_conv2d_16_source_31_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_count_1 <= _source_stream_conv2d_16_source_31_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_count_2 <= _source_stream_conv2d_16_source_31_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_count_3 <= _source_stream_conv2d_16_source_31_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_size_buf_0 <= _source_stream_conv2d_16_source_31_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_size_buf_1 <= _source_stream_conv2d_16_source_31_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_size_buf_2 <= _source_stream_conv2d_16_source_31_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_size_buf_3 <= _source_stream_conv2d_16_source_31_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_stride_buf_0 <= _source_stream_conv2d_16_source_31_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_stride_buf_1 <= _source_stream_conv2d_16_source_31_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_stride_buf_2 <= _source_stream_conv2d_16_source_31_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_31_pat_stride_buf_3 <= _source_stream_conv2d_16_source_31_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_31_source_pat_fsm_14 == 1) begin
        _stream_conv2d_16_source_31_source_ram_raddr <= _stream_conv2d_16_source_31_source_pat_all_offset;
        _stream_conv2d_16_source_31_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_31_source_pat_fsm_14 == 1) begin
        _source_stream_conv2d_16_source_31_pat_cur_offset_0 <= _source_stream_conv2d_16_source_31_pat_cur_offset_0 + _source_stream_conv2d_16_source_31_pat_stride_buf_0;
        _source_stream_conv2d_16_source_31_pat_count_0 <= _source_stream_conv2d_16_source_31_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_31_source_pat_fsm_14 == 1) && (_source_stream_conv2d_16_source_31_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_31_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_31_pat_count_0 <= _source_stream_conv2d_16_source_31_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_31_source_pat_fsm_14 == 1) && (_source_stream_conv2d_16_source_31_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_31_pat_cur_offset_1 <= _source_stream_conv2d_16_source_31_pat_cur_offset_1 + _source_stream_conv2d_16_source_31_pat_stride_buf_1;
        _source_stream_conv2d_16_source_31_pat_count_1 <= _source_stream_conv2d_16_source_31_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_31_source_pat_fsm_14 == 1) && (_source_stream_conv2d_16_source_31_pat_count_0 == 0) && (_source_stream_conv2d_16_source_31_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_31_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_31_pat_count_1 <= _source_stream_conv2d_16_source_31_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_31_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_16_source_31_pat_count_0 == 0) && (_source_stream_conv2d_16_source_31_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_31_pat_cur_offset_2 <= _source_stream_conv2d_16_source_31_pat_cur_offset_2 + _source_stream_conv2d_16_source_31_pat_stride_buf_2;
        _source_stream_conv2d_16_source_31_pat_count_2 <= _source_stream_conv2d_16_source_31_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_31_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_16_source_31_pat_count_0 == 0) && (_source_stream_conv2d_16_source_31_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_31_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_31_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_31_pat_count_2 <= _source_stream_conv2d_16_source_31_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_31_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_16_source_31_pat_count_0 == 0) && (_source_stream_conv2d_16_source_31_pat_count_1 == 0) && (_source_stream_conv2d_16_source_31_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_31_pat_cur_offset_3 <= _source_stream_conv2d_16_source_31_pat_cur_offset_3 + _source_stream_conv2d_16_source_31_pat_stride_buf_3;
        _source_stream_conv2d_16_source_31_pat_count_3 <= _source_stream_conv2d_16_source_31_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_31_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_16_source_31_pat_count_0 == 0) && (_source_stream_conv2d_16_source_31_pat_count_1 == 0) && (_source_stream_conv2d_16_source_31_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_31_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_31_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_31_pat_count_3 <= _source_stream_conv2d_16_source_31_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_31_source_pat_fsm_14 == 2) begin
        _stream_conv2d_16_source_31_source_ram_renable <= 0;
        _stream_conv2d_16_source_31_idle <= 1;
      end 
      _set_flag_640 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_640 <= 1;
      end 
      if(_set_flag_640) begin
        _stream_conv2d_16_source_32_source_mode <= 3'b10;
        _stream_conv2d_16_source_32_source_offset <= conv2d_16_filter_page_comp_offset_buf;
      end 
      if(_set_flag_640) begin
        _source_stream_conv2d_16_source_32_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_32_pat_stride_0 <= 1;
      end 
      if(_set_flag_640) begin
        _source_stream_conv2d_16_source_32_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_32_pat_stride_1 <= cparam_conv2d_16_stream_aligned_reduce_size;
      end 
      if(_set_flag_640) begin
        _source_stream_conv2d_16_source_32_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_32_pat_stride_2 <= 0;
      end 
      if(_set_flag_640) begin
        _source_stream_conv2d_16_source_32_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_32_pat_stride_3 <= 0;
      end 
      if(_set_flag_640) begin
        _stream_conv2d_16_source_32_source_ram_sel <= 16;
      end 
      __tmp_653_1 <= _tmp_653;
      if(__tmp_653_1) begin
        _stream_conv2d_16_source_32_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_32_source_ram_rvalid) begin
        __variable_wdata_506 <= _stream_conv2d_16_source_32_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _stream_conv2d_16_source_32_idle <= 0;
        _stream_conv2d_16_source_32_source_offset_buf <= _stream_conv2d_16_source_32_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_count_0 <= _source_stream_conv2d_16_source_32_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_count_1 <= _source_stream_conv2d_16_source_32_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_count_2 <= _source_stream_conv2d_16_source_32_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_count_3 <= _source_stream_conv2d_16_source_32_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_size_buf_0 <= _source_stream_conv2d_16_source_32_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_size_buf_1 <= _source_stream_conv2d_16_source_32_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_size_buf_2 <= _source_stream_conv2d_16_source_32_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_size_buf_3 <= _source_stream_conv2d_16_source_32_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_stride_buf_0 <= _source_stream_conv2d_16_source_32_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_stride_buf_1 <= _source_stream_conv2d_16_source_32_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_stride_buf_2 <= _source_stream_conv2d_16_source_32_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_32_pat_stride_buf_3 <= _source_stream_conv2d_16_source_32_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_32_source_pat_fsm_15 == 1) begin
        _stream_conv2d_16_source_32_source_ram_raddr <= _stream_conv2d_16_source_32_source_pat_all_offset;
        _stream_conv2d_16_source_32_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_32_source_pat_fsm_15 == 1) begin
        _source_stream_conv2d_16_source_32_pat_cur_offset_0 <= _source_stream_conv2d_16_source_32_pat_cur_offset_0 + _source_stream_conv2d_16_source_32_pat_stride_buf_0;
        _source_stream_conv2d_16_source_32_pat_count_0 <= _source_stream_conv2d_16_source_32_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_32_source_pat_fsm_15 == 1) && (_source_stream_conv2d_16_source_32_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_32_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_32_pat_count_0 <= _source_stream_conv2d_16_source_32_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_32_source_pat_fsm_15 == 1) && (_source_stream_conv2d_16_source_32_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_32_pat_cur_offset_1 <= _source_stream_conv2d_16_source_32_pat_cur_offset_1 + _source_stream_conv2d_16_source_32_pat_stride_buf_1;
        _source_stream_conv2d_16_source_32_pat_count_1 <= _source_stream_conv2d_16_source_32_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_32_source_pat_fsm_15 == 1) && (_source_stream_conv2d_16_source_32_pat_count_0 == 0) && (_source_stream_conv2d_16_source_32_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_32_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_32_pat_count_1 <= _source_stream_conv2d_16_source_32_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_32_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_16_source_32_pat_count_0 == 0) && (_source_stream_conv2d_16_source_32_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_32_pat_cur_offset_2 <= _source_stream_conv2d_16_source_32_pat_cur_offset_2 + _source_stream_conv2d_16_source_32_pat_stride_buf_2;
        _source_stream_conv2d_16_source_32_pat_count_2 <= _source_stream_conv2d_16_source_32_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_32_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_16_source_32_pat_count_0 == 0) && (_source_stream_conv2d_16_source_32_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_32_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_32_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_32_pat_count_2 <= _source_stream_conv2d_16_source_32_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_32_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_16_source_32_pat_count_0 == 0) && (_source_stream_conv2d_16_source_32_pat_count_1 == 0) && (_source_stream_conv2d_16_source_32_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_32_pat_cur_offset_3 <= _source_stream_conv2d_16_source_32_pat_cur_offset_3 + _source_stream_conv2d_16_source_32_pat_stride_buf_3;
        _source_stream_conv2d_16_source_32_pat_count_3 <= _source_stream_conv2d_16_source_32_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_32_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_16_source_32_pat_count_0 == 0) && (_source_stream_conv2d_16_source_32_pat_count_1 == 0) && (_source_stream_conv2d_16_source_32_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_32_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_32_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_32_pat_count_3 <= _source_stream_conv2d_16_source_32_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_32_source_pat_fsm_15 == 2) begin
        _stream_conv2d_16_source_32_source_ram_renable <= 0;
        _stream_conv2d_16_source_32_idle <= 1;
      end 
      _set_flag_654 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_654 <= 1;
      end 
      if(_set_flag_654) begin
        _stream_conv2d_16_source_33_source_mode <= 3'b10;
        _stream_conv2d_16_source_33_source_offset <= conv2d_16_filter_page_comp_offset_buf;
      end 
      if(_set_flag_654) begin
        _source_stream_conv2d_16_source_33_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_33_pat_stride_0 <= 1;
      end 
      if(_set_flag_654) begin
        _source_stream_conv2d_16_source_33_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_33_pat_stride_1 <= cparam_conv2d_16_stream_aligned_reduce_size;
      end 
      if(_set_flag_654) begin
        _source_stream_conv2d_16_source_33_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_33_pat_stride_2 <= 0;
      end 
      if(_set_flag_654) begin
        _source_stream_conv2d_16_source_33_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_33_pat_stride_3 <= 0;
      end 
      if(_set_flag_654) begin
        _stream_conv2d_16_source_33_source_ram_sel <= 17;
      end 
      __tmp_667_1 <= _tmp_667;
      if(__tmp_667_1) begin
        _stream_conv2d_16_source_33_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_33_source_ram_rvalid) begin
        __variable_wdata_507 <= _stream_conv2d_16_source_33_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _stream_conv2d_16_source_33_idle <= 0;
        _stream_conv2d_16_source_33_source_offset_buf <= _stream_conv2d_16_source_33_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_count_0 <= _source_stream_conv2d_16_source_33_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_count_1 <= _source_stream_conv2d_16_source_33_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_count_2 <= _source_stream_conv2d_16_source_33_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_count_3 <= _source_stream_conv2d_16_source_33_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_size_buf_0 <= _source_stream_conv2d_16_source_33_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_size_buf_1 <= _source_stream_conv2d_16_source_33_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_size_buf_2 <= _source_stream_conv2d_16_source_33_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_size_buf_3 <= _source_stream_conv2d_16_source_33_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_stride_buf_0 <= _source_stream_conv2d_16_source_33_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_stride_buf_1 <= _source_stream_conv2d_16_source_33_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_stride_buf_2 <= _source_stream_conv2d_16_source_33_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_33_pat_stride_buf_3 <= _source_stream_conv2d_16_source_33_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_33_source_pat_fsm_16 == 1) begin
        _stream_conv2d_16_source_33_source_ram_raddr <= _stream_conv2d_16_source_33_source_pat_all_offset;
        _stream_conv2d_16_source_33_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_33_source_pat_fsm_16 == 1) begin
        _source_stream_conv2d_16_source_33_pat_cur_offset_0 <= _source_stream_conv2d_16_source_33_pat_cur_offset_0 + _source_stream_conv2d_16_source_33_pat_stride_buf_0;
        _source_stream_conv2d_16_source_33_pat_count_0 <= _source_stream_conv2d_16_source_33_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_33_source_pat_fsm_16 == 1) && (_source_stream_conv2d_16_source_33_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_33_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_33_pat_count_0 <= _source_stream_conv2d_16_source_33_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_33_source_pat_fsm_16 == 1) && (_source_stream_conv2d_16_source_33_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_33_pat_cur_offset_1 <= _source_stream_conv2d_16_source_33_pat_cur_offset_1 + _source_stream_conv2d_16_source_33_pat_stride_buf_1;
        _source_stream_conv2d_16_source_33_pat_count_1 <= _source_stream_conv2d_16_source_33_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_33_source_pat_fsm_16 == 1) && (_source_stream_conv2d_16_source_33_pat_count_0 == 0) && (_source_stream_conv2d_16_source_33_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_33_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_33_pat_count_1 <= _source_stream_conv2d_16_source_33_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_33_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_16_source_33_pat_count_0 == 0) && (_source_stream_conv2d_16_source_33_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_33_pat_cur_offset_2 <= _source_stream_conv2d_16_source_33_pat_cur_offset_2 + _source_stream_conv2d_16_source_33_pat_stride_buf_2;
        _source_stream_conv2d_16_source_33_pat_count_2 <= _source_stream_conv2d_16_source_33_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_33_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_16_source_33_pat_count_0 == 0) && (_source_stream_conv2d_16_source_33_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_33_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_33_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_33_pat_count_2 <= _source_stream_conv2d_16_source_33_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_33_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_16_source_33_pat_count_0 == 0) && (_source_stream_conv2d_16_source_33_pat_count_1 == 0) && (_source_stream_conv2d_16_source_33_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_33_pat_cur_offset_3 <= _source_stream_conv2d_16_source_33_pat_cur_offset_3 + _source_stream_conv2d_16_source_33_pat_stride_buf_3;
        _source_stream_conv2d_16_source_33_pat_count_3 <= _source_stream_conv2d_16_source_33_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_33_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_16_source_33_pat_count_0 == 0) && (_source_stream_conv2d_16_source_33_pat_count_1 == 0) && (_source_stream_conv2d_16_source_33_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_33_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_33_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_33_pat_count_3 <= _source_stream_conv2d_16_source_33_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_33_source_pat_fsm_16 == 2) begin
        _stream_conv2d_16_source_33_source_ram_renable <= 0;
        _stream_conv2d_16_source_33_idle <= 1;
      end 
      _set_flag_668 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_668 <= 1;
      end 
      if(_set_flag_668) begin
        _stream_conv2d_16_source_34_source_mode <= 3'b10;
        _stream_conv2d_16_source_34_source_offset <= conv2d_16_filter_page_comp_offset_buf;
      end 
      if(_set_flag_668) begin
        _source_stream_conv2d_16_source_34_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_34_pat_stride_0 <= 1;
      end 
      if(_set_flag_668) begin
        _source_stream_conv2d_16_source_34_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_34_pat_stride_1 <= cparam_conv2d_16_stream_aligned_reduce_size;
      end 
      if(_set_flag_668) begin
        _source_stream_conv2d_16_source_34_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_34_pat_stride_2 <= 0;
      end 
      if(_set_flag_668) begin
        _source_stream_conv2d_16_source_34_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_34_pat_stride_3 <= 0;
      end 
      if(_set_flag_668) begin
        _stream_conv2d_16_source_34_source_ram_sel <= 18;
      end 
      __tmp_681_1 <= _tmp_681;
      if(__tmp_681_1) begin
        _stream_conv2d_16_source_34_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_34_source_ram_rvalid) begin
        __variable_wdata_508 <= _stream_conv2d_16_source_34_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _stream_conv2d_16_source_34_idle <= 0;
        _stream_conv2d_16_source_34_source_offset_buf <= _stream_conv2d_16_source_34_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_count_0 <= _source_stream_conv2d_16_source_34_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_count_1 <= _source_stream_conv2d_16_source_34_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_count_2 <= _source_stream_conv2d_16_source_34_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_count_3 <= _source_stream_conv2d_16_source_34_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_size_buf_0 <= _source_stream_conv2d_16_source_34_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_size_buf_1 <= _source_stream_conv2d_16_source_34_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_size_buf_2 <= _source_stream_conv2d_16_source_34_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_size_buf_3 <= _source_stream_conv2d_16_source_34_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_stride_buf_0 <= _source_stream_conv2d_16_source_34_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_stride_buf_1 <= _source_stream_conv2d_16_source_34_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_stride_buf_2 <= _source_stream_conv2d_16_source_34_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_34_pat_stride_buf_3 <= _source_stream_conv2d_16_source_34_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_34_source_pat_fsm_17 == 1) begin
        _stream_conv2d_16_source_34_source_ram_raddr <= _stream_conv2d_16_source_34_source_pat_all_offset;
        _stream_conv2d_16_source_34_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_34_source_pat_fsm_17 == 1) begin
        _source_stream_conv2d_16_source_34_pat_cur_offset_0 <= _source_stream_conv2d_16_source_34_pat_cur_offset_0 + _source_stream_conv2d_16_source_34_pat_stride_buf_0;
        _source_stream_conv2d_16_source_34_pat_count_0 <= _source_stream_conv2d_16_source_34_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_34_source_pat_fsm_17 == 1) && (_source_stream_conv2d_16_source_34_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_34_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_34_pat_count_0 <= _source_stream_conv2d_16_source_34_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_34_source_pat_fsm_17 == 1) && (_source_stream_conv2d_16_source_34_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_34_pat_cur_offset_1 <= _source_stream_conv2d_16_source_34_pat_cur_offset_1 + _source_stream_conv2d_16_source_34_pat_stride_buf_1;
        _source_stream_conv2d_16_source_34_pat_count_1 <= _source_stream_conv2d_16_source_34_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_34_source_pat_fsm_17 == 1) && (_source_stream_conv2d_16_source_34_pat_count_0 == 0) && (_source_stream_conv2d_16_source_34_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_34_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_34_pat_count_1 <= _source_stream_conv2d_16_source_34_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_34_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_16_source_34_pat_count_0 == 0) && (_source_stream_conv2d_16_source_34_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_34_pat_cur_offset_2 <= _source_stream_conv2d_16_source_34_pat_cur_offset_2 + _source_stream_conv2d_16_source_34_pat_stride_buf_2;
        _source_stream_conv2d_16_source_34_pat_count_2 <= _source_stream_conv2d_16_source_34_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_34_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_16_source_34_pat_count_0 == 0) && (_source_stream_conv2d_16_source_34_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_34_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_34_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_34_pat_count_2 <= _source_stream_conv2d_16_source_34_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_34_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_16_source_34_pat_count_0 == 0) && (_source_stream_conv2d_16_source_34_pat_count_1 == 0) && (_source_stream_conv2d_16_source_34_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_34_pat_cur_offset_3 <= _source_stream_conv2d_16_source_34_pat_cur_offset_3 + _source_stream_conv2d_16_source_34_pat_stride_buf_3;
        _source_stream_conv2d_16_source_34_pat_count_3 <= _source_stream_conv2d_16_source_34_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_34_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_16_source_34_pat_count_0 == 0) && (_source_stream_conv2d_16_source_34_pat_count_1 == 0) && (_source_stream_conv2d_16_source_34_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_34_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_34_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_34_pat_count_3 <= _source_stream_conv2d_16_source_34_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_34_source_pat_fsm_17 == 2) begin
        _stream_conv2d_16_source_34_source_ram_renable <= 0;
        _stream_conv2d_16_source_34_idle <= 1;
      end 
      _set_flag_682 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_682 <= 1;
      end 
      if(_set_flag_682) begin
        _stream_conv2d_16_source_35_source_mode <= 3'b10;
        _stream_conv2d_16_source_35_source_offset <= conv2d_16_filter_page_comp_offset_buf;
      end 
      if(_set_flag_682) begin
        _source_stream_conv2d_16_source_35_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_35_pat_stride_0 <= 1;
      end 
      if(_set_flag_682) begin
        _source_stream_conv2d_16_source_35_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_35_pat_stride_1 <= cparam_conv2d_16_stream_aligned_reduce_size;
      end 
      if(_set_flag_682) begin
        _source_stream_conv2d_16_source_35_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_35_pat_stride_2 <= 0;
      end 
      if(_set_flag_682) begin
        _source_stream_conv2d_16_source_35_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_35_pat_stride_3 <= 0;
      end 
      if(_set_flag_682) begin
        _stream_conv2d_16_source_35_source_ram_sel <= 19;
      end 
      __tmp_695_1 <= _tmp_695;
      if(__tmp_695_1) begin
        _stream_conv2d_16_source_35_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_35_source_ram_rvalid) begin
        __variable_wdata_509 <= _stream_conv2d_16_source_35_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _stream_conv2d_16_source_35_idle <= 0;
        _stream_conv2d_16_source_35_source_offset_buf <= _stream_conv2d_16_source_35_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_count_0 <= _source_stream_conv2d_16_source_35_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_count_1 <= _source_stream_conv2d_16_source_35_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_count_2 <= _source_stream_conv2d_16_source_35_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_count_3 <= _source_stream_conv2d_16_source_35_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_size_buf_0 <= _source_stream_conv2d_16_source_35_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_size_buf_1 <= _source_stream_conv2d_16_source_35_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_size_buf_2 <= _source_stream_conv2d_16_source_35_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_size_buf_3 <= _source_stream_conv2d_16_source_35_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_stride_buf_0 <= _source_stream_conv2d_16_source_35_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_stride_buf_1 <= _source_stream_conv2d_16_source_35_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_stride_buf_2 <= _source_stream_conv2d_16_source_35_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_35_pat_stride_buf_3 <= _source_stream_conv2d_16_source_35_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_35_source_pat_fsm_18 == 1) begin
        _stream_conv2d_16_source_35_source_ram_raddr <= _stream_conv2d_16_source_35_source_pat_all_offset;
        _stream_conv2d_16_source_35_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_35_source_pat_fsm_18 == 1) begin
        _source_stream_conv2d_16_source_35_pat_cur_offset_0 <= _source_stream_conv2d_16_source_35_pat_cur_offset_0 + _source_stream_conv2d_16_source_35_pat_stride_buf_0;
        _source_stream_conv2d_16_source_35_pat_count_0 <= _source_stream_conv2d_16_source_35_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_35_source_pat_fsm_18 == 1) && (_source_stream_conv2d_16_source_35_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_35_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_35_pat_count_0 <= _source_stream_conv2d_16_source_35_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_35_source_pat_fsm_18 == 1) && (_source_stream_conv2d_16_source_35_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_35_pat_cur_offset_1 <= _source_stream_conv2d_16_source_35_pat_cur_offset_1 + _source_stream_conv2d_16_source_35_pat_stride_buf_1;
        _source_stream_conv2d_16_source_35_pat_count_1 <= _source_stream_conv2d_16_source_35_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_35_source_pat_fsm_18 == 1) && (_source_stream_conv2d_16_source_35_pat_count_0 == 0) && (_source_stream_conv2d_16_source_35_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_35_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_35_pat_count_1 <= _source_stream_conv2d_16_source_35_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_35_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_16_source_35_pat_count_0 == 0) && (_source_stream_conv2d_16_source_35_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_35_pat_cur_offset_2 <= _source_stream_conv2d_16_source_35_pat_cur_offset_2 + _source_stream_conv2d_16_source_35_pat_stride_buf_2;
        _source_stream_conv2d_16_source_35_pat_count_2 <= _source_stream_conv2d_16_source_35_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_35_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_16_source_35_pat_count_0 == 0) && (_source_stream_conv2d_16_source_35_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_35_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_35_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_35_pat_count_2 <= _source_stream_conv2d_16_source_35_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_35_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_16_source_35_pat_count_0 == 0) && (_source_stream_conv2d_16_source_35_pat_count_1 == 0) && (_source_stream_conv2d_16_source_35_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_35_pat_cur_offset_3 <= _source_stream_conv2d_16_source_35_pat_cur_offset_3 + _source_stream_conv2d_16_source_35_pat_stride_buf_3;
        _source_stream_conv2d_16_source_35_pat_count_3 <= _source_stream_conv2d_16_source_35_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_35_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_16_source_35_pat_count_0 == 0) && (_source_stream_conv2d_16_source_35_pat_count_1 == 0) && (_source_stream_conv2d_16_source_35_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_35_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_35_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_35_pat_count_3 <= _source_stream_conv2d_16_source_35_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_35_source_pat_fsm_18 == 2) begin
        _stream_conv2d_16_source_35_source_ram_renable <= 0;
        _stream_conv2d_16_source_35_idle <= 1;
      end 
      _set_flag_696 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_696 <= 1;
      end 
      if(_set_flag_696) begin
        _stream_conv2d_16_source_36_source_mode <= 3'b10;
        _stream_conv2d_16_source_36_source_offset <= conv2d_16_filter_page_comp_offset_buf;
      end 
      if(_set_flag_696) begin
        _source_stream_conv2d_16_source_36_pat_size_0 <= cparam_conv2d_16_stream_reduce_size;
        _source_stream_conv2d_16_source_36_pat_stride_0 <= 1;
      end 
      if(_set_flag_696) begin
        _source_stream_conv2d_16_source_36_pat_size_1 <= conv2d_16_next_stream_num_ops;
        _source_stream_conv2d_16_source_36_pat_stride_1 <= cparam_conv2d_16_stream_aligned_reduce_size;
      end 
      if(_set_flag_696) begin
        _source_stream_conv2d_16_source_36_pat_size_2 <= 1;
        _source_stream_conv2d_16_source_36_pat_stride_2 <= 0;
      end 
      if(_set_flag_696) begin
        _source_stream_conv2d_16_source_36_pat_size_3 <= 1;
        _source_stream_conv2d_16_source_36_pat_stride_3 <= 0;
      end 
      if(_set_flag_696) begin
        _stream_conv2d_16_source_36_source_ram_sel <= 20;
      end 
      __tmp_709_1 <= _tmp_709;
      if(__tmp_709_1) begin
        _stream_conv2d_16_source_36_source_ram_rvalid <= 1;
      end 
      if(_stream_conv2d_16_source_36_source_ram_rvalid) begin
        __variable_wdata_510 <= _stream_conv2d_16_source_36_source_ram_rdata;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _stream_conv2d_16_source_36_idle <= 0;
        _stream_conv2d_16_source_36_source_offset_buf <= _stream_conv2d_16_source_36_source_offset;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_count_0 <= _source_stream_conv2d_16_source_36_pat_size_0 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_count_1 <= _source_stream_conv2d_16_source_36_pat_size_1 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_count_2 <= _source_stream_conv2d_16_source_36_pat_size_2 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_count_3 <= _source_stream_conv2d_16_source_36_pat_size_3 - 1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_size_buf_0 <= _source_stream_conv2d_16_source_36_pat_size_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_size_buf_1 <= _source_stream_conv2d_16_source_36_pat_size_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_size_buf_2 <= _source_stream_conv2d_16_source_36_pat_size_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_size_buf_3 <= _source_stream_conv2d_16_source_36_pat_size_3;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_stride_buf_0 <= _source_stream_conv2d_16_source_36_pat_stride_0;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_stride_buf_1 <= _source_stream_conv2d_16_source_36_pat_stride_1;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_stride_buf_2 <= _source_stream_conv2d_16_source_36_pat_stride_2;
      end 
      if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
        _source_stream_conv2d_16_source_36_pat_stride_buf_3 <= _source_stream_conv2d_16_source_36_pat_stride_3;
      end 
      if(_stream_conv2d_16_source_36_source_pat_fsm_19 == 1) begin
        _stream_conv2d_16_source_36_source_ram_raddr <= _stream_conv2d_16_source_36_source_pat_all_offset;
        _stream_conv2d_16_source_36_source_ram_renable <= 1;
      end 
      if(_stream_conv2d_16_source_36_source_pat_fsm_19 == 1) begin
        _source_stream_conv2d_16_source_36_pat_cur_offset_0 <= _source_stream_conv2d_16_source_36_pat_cur_offset_0 + _source_stream_conv2d_16_source_36_pat_stride_buf_0;
        _source_stream_conv2d_16_source_36_pat_count_0 <= _source_stream_conv2d_16_source_36_pat_count_0 - 1;
      end 
      if((_stream_conv2d_16_source_36_source_pat_fsm_19 == 1) && (_source_stream_conv2d_16_source_36_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_36_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_16_source_36_pat_count_0 <= _source_stream_conv2d_16_source_36_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_16_source_36_source_pat_fsm_19 == 1) && (_source_stream_conv2d_16_source_36_pat_count_0 == 0)) begin
        _source_stream_conv2d_16_source_36_pat_cur_offset_1 <= _source_stream_conv2d_16_source_36_pat_cur_offset_1 + _source_stream_conv2d_16_source_36_pat_stride_buf_1;
        _source_stream_conv2d_16_source_36_pat_count_1 <= _source_stream_conv2d_16_source_36_pat_count_1 - 1;
      end 
      if((_stream_conv2d_16_source_36_source_pat_fsm_19 == 1) && (_source_stream_conv2d_16_source_36_pat_count_0 == 0) && (_source_stream_conv2d_16_source_36_pat_count_1 == 0)) begin
        _source_stream_conv2d_16_source_36_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_16_source_36_pat_count_1 <= _source_stream_conv2d_16_source_36_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_16_source_36_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_16_source_36_pat_count_0 == 0) && (_source_stream_conv2d_16_source_36_pat_count_1 == 0))) begin
        _source_stream_conv2d_16_source_36_pat_cur_offset_2 <= _source_stream_conv2d_16_source_36_pat_cur_offset_2 + _source_stream_conv2d_16_source_36_pat_stride_buf_2;
        _source_stream_conv2d_16_source_36_pat_count_2 <= _source_stream_conv2d_16_source_36_pat_count_2 - 1;
      end 
      if((_stream_conv2d_16_source_36_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_16_source_36_pat_count_0 == 0) && (_source_stream_conv2d_16_source_36_pat_count_1 == 0)) && (_source_stream_conv2d_16_source_36_pat_count_2 == 0)) begin
        _source_stream_conv2d_16_source_36_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_16_source_36_pat_count_2 <= _source_stream_conv2d_16_source_36_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_16_source_36_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_16_source_36_pat_count_0 == 0) && (_source_stream_conv2d_16_source_36_pat_count_1 == 0) && (_source_stream_conv2d_16_source_36_pat_count_2 == 0))) begin
        _source_stream_conv2d_16_source_36_pat_cur_offset_3 <= _source_stream_conv2d_16_source_36_pat_cur_offset_3 + _source_stream_conv2d_16_source_36_pat_stride_buf_3;
        _source_stream_conv2d_16_source_36_pat_count_3 <= _source_stream_conv2d_16_source_36_pat_count_3 - 1;
      end 
      if((_stream_conv2d_16_source_36_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_16_source_36_pat_count_0 == 0) && (_source_stream_conv2d_16_source_36_pat_count_1 == 0) && (_source_stream_conv2d_16_source_36_pat_count_2 == 0)) && (_source_stream_conv2d_16_source_36_pat_count_3 == 0)) begin
        _source_stream_conv2d_16_source_36_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_16_source_36_pat_count_3 <= _source_stream_conv2d_16_source_36_pat_size_buf_3 - 1;
      end 
      if(_stream_conv2d_16_source_36_source_pat_fsm_19 == 2) begin
        _stream_conv2d_16_source_36_source_ram_renable <= 0;
        _stream_conv2d_16_source_36_idle <= 1;
      end 
      _set_flag_710 <= 0;
      if(conv2d_16_comp_fsm == 3) begin
        _set_flag_710 <= 1;
      end 
      __stream_conv2d_16_sink_37_sink_offset_0_1 <= conv2d_16_stream_out_local + conv2d_16_out_page_comp_offset_buf;
      __stream_conv2d_16_sink_37_sink_size_1_1 <= conv2d_16_next_stream_num_ops;
      __stream_seq_14_cond_2_1 <= _set_flag_710;
      __set_flag_710_1 <= _set_flag_710;
      __set_flag_710_2 <= __set_flag_710_1;
      __set_flag_710_3 <= __set_flag_710_2;
      __set_flag_710_4 <= __set_flag_710_3;
      __set_flag_710_5 <= __set_flag_710_4;
      __set_flag_710_6 <= __set_flag_710_5;
      __set_flag_710_7 <= __set_flag_710_6;
      __set_flag_710_8 <= __set_flag_710_7;
      __set_flag_710_9 <= __set_flag_710_8;
      __set_flag_710_10 <= __set_flag_710_9;
      __set_flag_710_11 <= __set_flag_710_10;
      __set_flag_710_12 <= __set_flag_710_11;
      __set_flag_710_13 <= __set_flag_710_12;
      __set_flag_710_14 <= __set_flag_710_13;
      __set_flag_710_15 <= __set_flag_710_14;
      __set_flag_710_16 <= __set_flag_710_15;
      __set_flag_710_17 <= __set_flag_710_16;
      __set_flag_710_18 <= __set_flag_710_17;
      __set_flag_710_19 <= __set_flag_710_18;
      __set_flag_710_20 <= __set_flag_710_19;
      __set_flag_710_21 <= __set_flag_710_20;
      __set_flag_710_22 <= __set_flag_710_21;
      __set_flag_710_23 <= __set_flag_710_22;
      __set_flag_710_24 <= __set_flag_710_23;
      __set_flag_710_25 <= __set_flag_710_24;
      __set_flag_710_26 <= __set_flag_710_25;
      __set_flag_710_27 <= __set_flag_710_26;
      __set_flag_710_28 <= __set_flag_710_27;
      __set_flag_710_29 <= __set_flag_710_28;
      __set_flag_710_30 <= __set_flag_710_29;
      __set_flag_710_31 <= __set_flag_710_30;
      __set_flag_710_32 <= __set_flag_710_31;
      __set_flag_710_33 <= __set_flag_710_32;
      __set_flag_710_34 <= __set_flag_710_33;
      __set_flag_710_35 <= __set_flag_710_34;
      __set_flag_710_36 <= __set_flag_710_35;
      __set_flag_710_37 <= __set_flag_710_36;
      __set_flag_710_38 <= __set_flag_710_37;
      __set_flag_710_39 <= __set_flag_710_38;
      __set_flag_710_40 <= __set_flag_710_39;
      __set_flag_710_41 <= __set_flag_710_40;
      __set_flag_710_42 <= __set_flag_710_41;
      __set_flag_710_43 <= __set_flag_710_42;
      __set_flag_710_44 <= __set_flag_710_43;
      __set_flag_710_45 <= __set_flag_710_44;
      if(__set_flag_710_45) begin
        _stream_conv2d_16_sink_37_sink_ram_sel <= 21;
      end 
      __stream_conv2d_16_start_1 <= _stream_conv2d_16_start;
      __stream_conv2d_16_start_2 <= __stream_conv2d_16_start_1;
      __stream_conv2d_16_start_3 <= __stream_conv2d_16_start_2;
      __stream_conv2d_16_start_4 <= __stream_conv2d_16_start_3;
      __stream_conv2d_16_start_5 <= __stream_conv2d_16_start_4;
      __stream_conv2d_16_start_6 <= __stream_conv2d_16_start_5;
      __stream_conv2d_16_start_7 <= __stream_conv2d_16_start_6;
      __stream_conv2d_16_start_8 <= __stream_conv2d_16_start_7;
      __stream_conv2d_16_start_9 <= __stream_conv2d_16_start_8;
      __stream_conv2d_16_start_10 <= __stream_conv2d_16_start_9;
      __stream_conv2d_16_start_11 <= __stream_conv2d_16_start_10;
      __stream_conv2d_16_start_12 <= __stream_conv2d_16_start_11;
      __stream_conv2d_16_start_13 <= __stream_conv2d_16_start_12;
      __stream_conv2d_16_start_14 <= __stream_conv2d_16_start_13;
      __stream_conv2d_16_start_15 <= __stream_conv2d_16_start_14;
      __stream_conv2d_16_start_16 <= __stream_conv2d_16_start_15;
      __stream_conv2d_16_start_17 <= __stream_conv2d_16_start_16;
      __stream_conv2d_16_start_18 <= __stream_conv2d_16_start_17;
      __stream_conv2d_16_start_19 <= __stream_conv2d_16_start_18;
      __stream_conv2d_16_start_20 <= __stream_conv2d_16_start_19;
      __stream_conv2d_16_start_21 <= __stream_conv2d_16_start_20;
      __stream_conv2d_16_start_22 <= __stream_conv2d_16_start_21;
      __stream_conv2d_16_start_23 <= __stream_conv2d_16_start_22;
      __stream_conv2d_16_start_24 <= __stream_conv2d_16_start_23;
      __stream_conv2d_16_start_25 <= __stream_conv2d_16_start_24;
      __stream_conv2d_16_start_26 <= __stream_conv2d_16_start_25;
      __stream_conv2d_16_start_27 <= __stream_conv2d_16_start_26;
      __stream_conv2d_16_start_28 <= __stream_conv2d_16_start_27;
      __stream_conv2d_16_start_29 <= __stream_conv2d_16_start_28;
      __stream_conv2d_16_start_30 <= __stream_conv2d_16_start_29;
      __stream_conv2d_16_start_31 <= __stream_conv2d_16_start_30;
      __stream_conv2d_16_start_32 <= __stream_conv2d_16_start_31;
      __stream_conv2d_16_start_33 <= __stream_conv2d_16_start_32;
      __stream_conv2d_16_start_34 <= __stream_conv2d_16_start_33;
      __stream_conv2d_16_start_35 <= __stream_conv2d_16_start_34;
      __stream_conv2d_16_start_36 <= __stream_conv2d_16_start_35;
      __stream_conv2d_16_start_37 <= __stream_conv2d_16_start_36;
      __stream_conv2d_16_start_38 <= __stream_conv2d_16_start_37;
      __stream_conv2d_16_start_39 <= __stream_conv2d_16_start_38;
      __stream_conv2d_16_start_40 <= __stream_conv2d_16_start_39;
      __stream_conv2d_16_start_41 <= __stream_conv2d_16_start_40;
      __stream_conv2d_16_start_42 <= __stream_conv2d_16_start_41;
      __stream_conv2d_16_start_43 <= __stream_conv2d_16_start_42;
      __stream_conv2d_16_start_44 <= __stream_conv2d_16_start_43;
      __stream_conv2d_16_start_45 <= __stream_conv2d_16_start_44;
      __stream_conv2d_16_start_46 <= __stream_conv2d_16_start_45;
      if(__stream_conv2d_16_start_46 && _stream_conv2d_16_sink_37_sink_mode & 3'b1) begin
        _stream_conv2d_16_sink_37_sink_waddr <= _stream_conv2d_16_sink_37_sink_offset - _stream_conv2d_16_sink_37_sink_stride;
        _stream_conv2d_16_sink_37_sink_count <= _stream_conv2d_16_sink_37_sink_size;
        _stream_conv2d_16_sink_37_sink_offset_buf <= _stream_conv2d_16_sink_37_sink_offset;
        _stream_conv2d_16_sink_37_sink_stride_buf <= _stream_conv2d_16_sink_37_sink_stride;
      end 
      if((_stream_conv2d_16_sink_37_sink_fsm_20 == 1) && stream_conv2d_16_sink_38_data) begin
        _stream_conv2d_16_sink_37_sink_waddr <= _stream_conv2d_16_sink_37_sink_waddr + _stream_conv2d_16_sink_37_sink_stride_buf;
        _stream_conv2d_16_sink_37_sink_wdata <= stream_conv2d_16_sink_37_data;
        _stream_conv2d_16_sink_37_sink_wenable <= 1;
        _stream_conv2d_16_sink_37_sink_count <= _stream_conv2d_16_sink_37_sink_count - 1;
      end 
      __tmp_713_1 <= _tmp_713;
      __tmp_713_2 <= __tmp_713_1;
      __tmp_713_3 <= __tmp_713_2;
      __tmp_713_4 <= __tmp_713_3;
      __tmp_713_5 <= __tmp_713_4;
      __tmp_715_1 <= _tmp_715;
      __tmp_715_2 <= __tmp_715_1;
      __tmp_715_3 <= __tmp_715_2;
      __tmp_715_4 <= __tmp_715_3;
      __tmp_715_5 <= __tmp_715_4;
      __tmp_715_6 <= __tmp_715_5;
      __tmp_715_7 <= __tmp_715_6;
      __tmp_715_8 <= __tmp_715_7;
      __tmp_715_9 <= __tmp_715_8;
      __tmp_715_10 <= __tmp_715_9;
      __tmp_715_11 <= __tmp_715_10;
      __tmp_715_12 <= __tmp_715_11;
      __tmp_717_1 <= _tmp_717;
      __tmp_717_2 <= __tmp_717_1;
      __tmp_717_3 <= __tmp_717_2;
      __tmp_717_4 <= __tmp_717_3;
      __tmp_717_5 <= __tmp_717_4;
      __tmp_717_6 <= __tmp_717_5;
      __tmp_717_7 <= __tmp_717_6;
      __tmp_717_8 <= __tmp_717_7;
      __tmp_717_9 <= __tmp_717_8;
      __tmp_717_10 <= __tmp_717_9;
      __tmp_717_11 <= __tmp_717_10;
      __tmp_717_12 <= __tmp_717_11;
      __tmp_719_1 <= _tmp_719;
      __tmp_719_2 <= __tmp_719_1;
      __tmp_719_3 <= __tmp_719_2;
      __tmp_719_4 <= __tmp_719_3;
      __tmp_719_5 <= __tmp_719_4;
      __tmp_719_6 <= __tmp_719_5;
      __tmp_719_7 <= __tmp_719_6;
      __tmp_719_8 <= __tmp_719_7;
      __tmp_719_9 <= __tmp_719_8;
      __tmp_719_10 <= __tmp_719_9;
      __tmp_719_11 <= __tmp_719_10;
      __tmp_719_12 <= __tmp_719_11;
      __tmp_721_1 <= _tmp_721;
      __tmp_721_2 <= __tmp_721_1;
      __tmp_721_3 <= __tmp_721_2;
      __tmp_721_4 <= __tmp_721_3;
      __tmp_721_5 <= __tmp_721_4;
      __tmp_721_6 <= __tmp_721_5;
      __tmp_721_7 <= __tmp_721_6;
      __tmp_721_8 <= __tmp_721_7;
      __tmp_721_9 <= __tmp_721_8;
      __tmp_721_10 <= __tmp_721_9;
      __tmp_721_11 <= __tmp_721_10;
      __tmp_721_12 <= __tmp_721_11;
      __tmp_723_1 <= _tmp_723;
      __tmp_723_2 <= __tmp_723_1;
      __tmp_723_3 <= __tmp_723_2;
      __tmp_723_4 <= __tmp_723_3;
      __tmp_723_5 <= __tmp_723_4;
      __tmp_723_6 <= __tmp_723_5;
      __tmp_723_7 <= __tmp_723_6;
      __tmp_723_8 <= __tmp_723_7;
      __tmp_723_9 <= __tmp_723_8;
      __tmp_723_10 <= __tmp_723_9;
      __tmp_723_11 <= __tmp_723_10;
      __tmp_723_12 <= __tmp_723_11;
      __tmp_725_1 <= _tmp_725;
      __tmp_725_2 <= __tmp_725_1;
      __tmp_725_3 <= __tmp_725_2;
      __tmp_725_4 <= __tmp_725_3;
      __tmp_725_5 <= __tmp_725_4;
      __tmp_725_6 <= __tmp_725_5;
      __tmp_725_7 <= __tmp_725_6;
      __tmp_725_8 <= __tmp_725_7;
      __tmp_725_9 <= __tmp_725_8;
      __tmp_725_10 <= __tmp_725_9;
      __tmp_725_11 <= __tmp_725_10;
      __tmp_725_12 <= __tmp_725_11;
      __tmp_727_1 <= _tmp_727;
      __tmp_727_2 <= __tmp_727_1;
      __tmp_727_3 <= __tmp_727_2;
      __tmp_727_4 <= __tmp_727_3;
      __tmp_727_5 <= __tmp_727_4;
      __tmp_727_6 <= __tmp_727_5;
      __tmp_727_7 <= __tmp_727_6;
      __tmp_727_8 <= __tmp_727_7;
      __tmp_727_9 <= __tmp_727_8;
      __tmp_727_10 <= __tmp_727_9;
      __tmp_727_11 <= __tmp_727_10;
      __tmp_727_12 <= __tmp_727_11;
      __tmp_729_1 <= _tmp_729;
      __tmp_729_2 <= __tmp_729_1;
      __tmp_729_3 <= __tmp_729_2;
      __tmp_729_4 <= __tmp_729_3;
      __tmp_729_5 <= __tmp_729_4;
      __tmp_729_6 <= __tmp_729_5;
      __tmp_729_7 <= __tmp_729_6;
      __tmp_729_8 <= __tmp_729_7;
      __tmp_729_9 <= __tmp_729_8;
      __tmp_729_10 <= __tmp_729_9;
      __tmp_729_11 <= __tmp_729_10;
      __tmp_729_12 <= __tmp_729_11;
      __tmp_731_1 <= _tmp_731;
      __tmp_731_2 <= __tmp_731_1;
      __tmp_731_3 <= __tmp_731_2;
      __tmp_731_4 <= __tmp_731_3;
      __tmp_731_5 <= __tmp_731_4;
      __tmp_731_6 <= __tmp_731_5;
      __tmp_731_7 <= __tmp_731_6;
      __tmp_731_8 <= __tmp_731_7;
      __tmp_731_9 <= __tmp_731_8;
      __tmp_731_10 <= __tmp_731_9;
      __tmp_731_11 <= __tmp_731_10;
      __tmp_731_12 <= __tmp_731_11;
      __tmp_733_1 <= _tmp_733;
      __tmp_733_2 <= __tmp_733_1;
      __tmp_733_3 <= __tmp_733_2;
      __tmp_733_4 <= __tmp_733_3;
      __tmp_733_5 <= __tmp_733_4;
      __tmp_733_6 <= __tmp_733_5;
      __tmp_733_7 <= __tmp_733_6;
      __tmp_733_8 <= __tmp_733_7;
      __tmp_733_9 <= __tmp_733_8;
      __tmp_733_10 <= __tmp_733_9;
      __tmp_733_11 <= __tmp_733_10;
      __tmp_733_12 <= __tmp_733_11;
      __tmp_735_1 <= _tmp_735;
      __tmp_735_2 <= __tmp_735_1;
      __tmp_735_3 <= __tmp_735_2;
      __tmp_735_4 <= __tmp_735_3;
      __tmp_735_5 <= __tmp_735_4;
      __tmp_735_6 <= __tmp_735_5;
      __tmp_735_7 <= __tmp_735_6;
      __tmp_735_8 <= __tmp_735_7;
      __tmp_735_9 <= __tmp_735_8;
      __tmp_735_10 <= __tmp_735_9;
      __tmp_735_11 <= __tmp_735_10;
      __tmp_735_12 <= __tmp_735_11;
      __tmp_737_1 <= _tmp_737;
      __tmp_737_2 <= __tmp_737_1;
      __tmp_737_3 <= __tmp_737_2;
      __tmp_737_4 <= __tmp_737_3;
      __tmp_737_5 <= __tmp_737_4;
      __tmp_737_6 <= __tmp_737_5;
      __tmp_737_7 <= __tmp_737_6;
      __tmp_737_8 <= __tmp_737_7;
      __tmp_737_9 <= __tmp_737_8;
      __tmp_737_10 <= __tmp_737_9;
      __tmp_737_11 <= __tmp_737_10;
      __tmp_737_12 <= __tmp_737_11;
      __tmp_739_1 <= _tmp_739;
      __tmp_739_2 <= __tmp_739_1;
      __tmp_739_3 <= __tmp_739_2;
      __tmp_739_4 <= __tmp_739_3;
      __tmp_739_5 <= __tmp_739_4;
      __tmp_739_6 <= __tmp_739_5;
      __tmp_739_7 <= __tmp_739_6;
      __tmp_739_8 <= __tmp_739_7;
      __tmp_739_9 <= __tmp_739_8;
      __tmp_739_10 <= __tmp_739_9;
      __tmp_739_11 <= __tmp_739_10;
      __tmp_739_12 <= __tmp_739_11;
      __tmp_741_1 <= _tmp_741;
      __tmp_741_2 <= __tmp_741_1;
      __tmp_741_3 <= __tmp_741_2;
      __tmp_741_4 <= __tmp_741_3;
      __tmp_741_5 <= __tmp_741_4;
      __tmp_741_6 <= __tmp_741_5;
      __tmp_741_7 <= __tmp_741_6;
      __tmp_741_8 <= __tmp_741_7;
      __tmp_741_9 <= __tmp_741_8;
      __tmp_741_10 <= __tmp_741_9;
      __tmp_741_11 <= __tmp_741_10;
      __tmp_741_12 <= __tmp_741_11;
      __tmp_743_1 <= _tmp_743;
      __tmp_743_2 <= __tmp_743_1;
      __tmp_743_3 <= __tmp_743_2;
      __tmp_743_4 <= __tmp_743_3;
      __tmp_743_5 <= __tmp_743_4;
      __tmp_743_6 <= __tmp_743_5;
      __tmp_743_7 <= __tmp_743_6;
      __tmp_743_8 <= __tmp_743_7;
      __tmp_743_9 <= __tmp_743_8;
      __tmp_743_10 <= __tmp_743_9;
      __tmp_743_11 <= __tmp_743_10;
      __tmp_743_12 <= __tmp_743_11;
      __tmp_745_1 <= _tmp_745;
      __tmp_745_2 <= __tmp_745_1;
      __tmp_745_3 <= __tmp_745_2;
      __tmp_745_4 <= __tmp_745_3;
      __tmp_745_5 <= __tmp_745_4;
      __tmp_745_6 <= __tmp_745_5;
      __tmp_745_7 <= __tmp_745_6;
      __tmp_745_8 <= __tmp_745_7;
      __tmp_745_9 <= __tmp_745_8;
      __tmp_745_10 <= __tmp_745_9;
      __tmp_745_11 <= __tmp_745_10;
      __tmp_745_12 <= __tmp_745_11;
      __tmp_747_1 <= _tmp_747;
      __tmp_747_2 <= __tmp_747_1;
      __tmp_747_3 <= __tmp_747_2;
      __tmp_747_4 <= __tmp_747_3;
      __tmp_747_5 <= __tmp_747_4;
      __tmp_747_6 <= __tmp_747_5;
      __tmp_747_7 <= __tmp_747_6;
      __tmp_747_8 <= __tmp_747_7;
      __tmp_747_9 <= __tmp_747_8;
      __tmp_747_10 <= __tmp_747_9;
      __tmp_747_11 <= __tmp_747_10;
      __tmp_747_12 <= __tmp_747_11;
      __tmp_749_1 <= _tmp_749;
      __tmp_749_2 <= __tmp_749_1;
      __tmp_749_3 <= __tmp_749_2;
      __tmp_749_4 <= __tmp_749_3;
      __tmp_749_5 <= __tmp_749_4;
      __tmp_749_6 <= __tmp_749_5;
      __tmp_749_7 <= __tmp_749_6;
      __tmp_749_8 <= __tmp_749_7;
      __tmp_749_9 <= __tmp_749_8;
      __tmp_749_10 <= __tmp_749_9;
      __tmp_749_11 <= __tmp_749_10;
      __tmp_749_12 <= __tmp_749_11;
      __tmp_751_1 <= _tmp_751;
      __tmp_751_2 <= __tmp_751_1;
      __tmp_751_3 <= __tmp_751_2;
      __tmp_751_4 <= __tmp_751_3;
      __tmp_751_5 <= __tmp_751_4;
      __tmp_751_6 <= __tmp_751_5;
      __tmp_751_7 <= __tmp_751_6;
      __tmp_751_8 <= __tmp_751_7;
      __tmp_751_9 <= __tmp_751_8;
      __tmp_751_10 <= __tmp_751_9;
      __tmp_751_11 <= __tmp_751_10;
      __tmp_751_12 <= __tmp_751_11;
      __tmp_753_1 <= _tmp_753;
      __tmp_753_2 <= __tmp_753_1;
      __tmp_753_3 <= __tmp_753_2;
      __tmp_753_4 <= __tmp_753_3;
      __tmp_753_5 <= __tmp_753_4;
      __tmp_753_6 <= __tmp_753_5;
      __tmp_753_7 <= __tmp_753_6;
      __tmp_753_8 <= __tmp_753_7;
      __tmp_753_9 <= __tmp_753_8;
      __tmp_753_10 <= __tmp_753_9;
      __tmp_753_11 <= __tmp_753_10;
      __tmp_753_12 <= __tmp_753_11;
      __tmp_755_1 <= _tmp_755;
      __tmp_755_2 <= __tmp_755_1;
      __tmp_755_3 <= __tmp_755_2;
      __tmp_755_4 <= __tmp_755_3;
      __tmp_755_5 <= __tmp_755_4;
      __tmp_755_6 <= __tmp_755_5;
      __tmp_755_7 <= __tmp_755_6;
      __tmp_755_8 <= __tmp_755_7;
      __tmp_755_9 <= __tmp_755_8;
      __tmp_755_10 <= __tmp_755_9;
      __tmp_755_11 <= __tmp_755_10;
      __tmp_755_12 <= __tmp_755_11;
      __tmp_757_1 <= _tmp_757;
      __tmp_757_2 <= __tmp_757_1;
      __tmp_757_3 <= __tmp_757_2;
      __tmp_757_4 <= __tmp_757_3;
      __tmp_757_5 <= __tmp_757_4;
      __tmp_757_6 <= __tmp_757_5;
      __tmp_757_7 <= __tmp_757_6;
      __tmp_757_8 <= __tmp_757_7;
      __tmp_757_9 <= __tmp_757_8;
      __tmp_757_10 <= __tmp_757_9;
      __tmp_757_11 <= __tmp_757_10;
      __tmp_757_12 <= __tmp_757_11;
      __tmp_759_1 <= _tmp_759;
      __tmp_759_2 <= __tmp_759_1;
      __tmp_759_3 <= __tmp_759_2;
      __tmp_759_4 <= __tmp_759_3;
      __tmp_759_5 <= __tmp_759_4;
      __tmp_759_6 <= __tmp_759_5;
      __tmp_759_7 <= __tmp_759_6;
      __tmp_759_8 <= __tmp_759_7;
      __tmp_759_9 <= __tmp_759_8;
      __tmp_759_10 <= __tmp_759_9;
      __tmp_759_11 <= __tmp_759_10;
      __tmp_759_12 <= __tmp_759_11;
      __tmp_761_1 <= _tmp_761;
      __tmp_761_2 <= __tmp_761_1;
      __tmp_761_3 <= __tmp_761_2;
      __tmp_761_4 <= __tmp_761_3;
      __tmp_761_5 <= __tmp_761_4;
      __tmp_761_6 <= __tmp_761_5;
      __tmp_761_7 <= __tmp_761_6;
      __tmp_761_8 <= __tmp_761_7;
      __tmp_761_9 <= __tmp_761_8;
      __tmp_761_10 <= __tmp_761_9;
      __tmp_761_11 <= __tmp_761_10;
      __tmp_761_12 <= __tmp_761_11;
      __tmp_763_1 <= _tmp_763;
      __tmp_763_2 <= __tmp_763_1;
      __tmp_763_3 <= __tmp_763_2;
      __tmp_763_4 <= __tmp_763_3;
      __tmp_763_5 <= __tmp_763_4;
      __tmp_763_6 <= __tmp_763_5;
      __tmp_763_7 <= __tmp_763_6;
      __tmp_763_8 <= __tmp_763_7;
      __tmp_763_9 <= __tmp_763_8;
      __tmp_763_10 <= __tmp_763_9;
      __tmp_763_11 <= __tmp_763_10;
      __tmp_763_12 <= __tmp_763_11;
      __tmp_765_1 <= _tmp_765;
      __tmp_765_2 <= __tmp_765_1;
      __tmp_765_3 <= __tmp_765_2;
      __tmp_765_4 <= __tmp_765_3;
      __tmp_765_5 <= __tmp_765_4;
      __tmp_765_6 <= __tmp_765_5;
      __tmp_765_7 <= __tmp_765_6;
      __tmp_765_8 <= __tmp_765_7;
      __tmp_765_9 <= __tmp_765_8;
      __tmp_765_10 <= __tmp_765_9;
      __tmp_765_11 <= __tmp_765_10;
      __tmp_765_12 <= __tmp_765_11;
      __tmp_767_1 <= _tmp_767;
      __tmp_767_2 <= __tmp_767_1;
      __tmp_767_3 <= __tmp_767_2;
      __tmp_767_4 <= __tmp_767_3;
      __tmp_767_5 <= __tmp_767_4;
      __tmp_767_6 <= __tmp_767_5;
      __tmp_767_7 <= __tmp_767_6;
      __tmp_767_8 <= __tmp_767_7;
      __tmp_767_9 <= __tmp_767_8;
      __tmp_767_10 <= __tmp_767_9;
      __tmp_767_11 <= __tmp_767_10;
      __tmp_767_12 <= __tmp_767_11;
      __tmp_769_1 <= _tmp_769;
      __tmp_769_2 <= __tmp_769_1;
      __tmp_769_3 <= __tmp_769_2;
      __tmp_769_4 <= __tmp_769_3;
      __tmp_769_5 <= __tmp_769_4;
      __tmp_769_6 <= __tmp_769_5;
      __tmp_769_7 <= __tmp_769_6;
      __tmp_769_8 <= __tmp_769_7;
      __tmp_769_9 <= __tmp_769_8;
      __tmp_769_10 <= __tmp_769_9;
      __tmp_769_11 <= __tmp_769_10;
      __tmp_769_12 <= __tmp_769_11;
      __tmp_769_13 <= __tmp_769_12;
      __tmp_769_14 <= __tmp_769_13;
      __tmp_769_15 <= __tmp_769_14;
      __tmp_769_16 <= __tmp_769_15;
      __tmp_769_17 <= __tmp_769_16;
      __tmp_769_18 <= __tmp_769_17;
      __tmp_769_19 <= __tmp_769_18;
      __tmp_769_20 <= __tmp_769_19;
      __tmp_769_21 <= __tmp_769_20;
      __tmp_769_22 <= __tmp_769_21;
      __tmp_771_1 <= _tmp_771;
      __tmp_771_2 <= __tmp_771_1;
      __tmp_771_3 <= __tmp_771_2;
      __tmp_771_4 <= __tmp_771_3;
      __tmp_771_5 <= __tmp_771_4;
      __tmp_771_6 <= __tmp_771_5;
      __tmp_771_7 <= __tmp_771_6;
      __tmp_771_8 <= __tmp_771_7;
      __tmp_771_9 <= __tmp_771_8;
      __tmp_771_10 <= __tmp_771_9;
      __tmp_771_11 <= __tmp_771_10;
      __tmp_771_12 <= __tmp_771_11;
      __tmp_771_13 <= __tmp_771_12;
      __tmp_771_14 <= __tmp_771_13;
      __tmp_771_15 <= __tmp_771_14;
      __tmp_771_16 <= __tmp_771_15;
      __tmp_771_17 <= __tmp_771_16;
      __tmp_771_18 <= __tmp_771_17;
      __tmp_771_19 <= __tmp_771_18;
      __tmp_771_20 <= __tmp_771_19;
      __tmp_771_21 <= __tmp_771_20;
      __tmp_771_22 <= __tmp_771_21;
      __tmp_773_1 <= _tmp_773;
      __tmp_773_2 <= __tmp_773_1;
      __tmp_773_3 <= __tmp_773_2;
      __tmp_773_4 <= __tmp_773_3;
      __tmp_773_5 <= __tmp_773_4;
      __tmp_773_6 <= __tmp_773_5;
      __tmp_773_7 <= __tmp_773_6;
      __tmp_773_8 <= __tmp_773_7;
      __tmp_773_9 <= __tmp_773_8;
      __tmp_773_10 <= __tmp_773_9;
      __tmp_773_11 <= __tmp_773_10;
      __tmp_773_12 <= __tmp_773_11;
      __tmp_773_13 <= __tmp_773_12;
      __tmp_773_14 <= __tmp_773_13;
      __tmp_773_15 <= __tmp_773_14;
      __tmp_773_16 <= __tmp_773_15;
      __tmp_773_17 <= __tmp_773_16;
      __tmp_773_18 <= __tmp_773_17;
      __tmp_773_19 <= __tmp_773_18;
      __tmp_773_20 <= __tmp_773_19;
      __tmp_773_21 <= __tmp_773_20;
      __tmp_773_22 <= __tmp_773_21;
      __tmp_775_1 <= _tmp_775;
      __tmp_775_2 <= __tmp_775_1;
      __tmp_775_3 <= __tmp_775_2;
      __tmp_775_4 <= __tmp_775_3;
      __tmp_775_5 <= __tmp_775_4;
      __tmp_775_6 <= __tmp_775_5;
      __tmp_775_7 <= __tmp_775_6;
      __tmp_775_8 <= __tmp_775_7;
      __tmp_775_9 <= __tmp_775_8;
      __tmp_775_10 <= __tmp_775_9;
      __tmp_775_11 <= __tmp_775_10;
      __tmp_775_12 <= __tmp_775_11;
      __tmp_775_13 <= __tmp_775_12;
      __tmp_775_14 <= __tmp_775_13;
      __tmp_775_15 <= __tmp_775_14;
      __tmp_775_16 <= __tmp_775_15;
      __tmp_775_17 <= __tmp_775_16;
      __tmp_775_18 <= __tmp_775_17;
      __tmp_775_19 <= __tmp_775_18;
      __tmp_775_20 <= __tmp_775_19;
      __tmp_775_21 <= __tmp_775_20;
      __tmp_775_22 <= __tmp_775_21;
      __tmp_777_1 <= _tmp_777;
      __tmp_777_2 <= __tmp_777_1;
      __tmp_777_3 <= __tmp_777_2;
      __tmp_777_4 <= __tmp_777_3;
      __tmp_777_5 <= __tmp_777_4;
      __tmp_777_6 <= __tmp_777_5;
      __tmp_777_7 <= __tmp_777_6;
      __tmp_777_8 <= __tmp_777_7;
      __tmp_777_9 <= __tmp_777_8;
      __tmp_777_10 <= __tmp_777_9;
      __tmp_777_11 <= __tmp_777_10;
      __tmp_777_12 <= __tmp_777_11;
      __tmp_777_13 <= __tmp_777_12;
      __tmp_777_14 <= __tmp_777_13;
      __tmp_777_15 <= __tmp_777_14;
      __tmp_777_16 <= __tmp_777_15;
      __tmp_777_17 <= __tmp_777_16;
      __tmp_777_18 <= __tmp_777_17;
      __tmp_777_19 <= __tmp_777_18;
      __tmp_777_20 <= __tmp_777_19;
      __tmp_777_21 <= __tmp_777_20;
      __tmp_777_22 <= __tmp_777_21;
      __tmp_779_1 <= _tmp_779;
      __tmp_779_2 <= __tmp_779_1;
      __tmp_779_3 <= __tmp_779_2;
      __tmp_779_4 <= __tmp_779_3;
      __tmp_779_5 <= __tmp_779_4;
      __tmp_779_6 <= __tmp_779_5;
      __tmp_779_7 <= __tmp_779_6;
      __tmp_779_8 <= __tmp_779_7;
      __tmp_779_9 <= __tmp_779_8;
      __tmp_779_10 <= __tmp_779_9;
      __tmp_779_11 <= __tmp_779_10;
      __tmp_779_12 <= __tmp_779_11;
      __tmp_779_13 <= __tmp_779_12;
      __tmp_779_14 <= __tmp_779_13;
      __tmp_779_15 <= __tmp_779_14;
      __tmp_779_16 <= __tmp_779_15;
      __tmp_779_17 <= __tmp_779_16;
      __tmp_779_18 <= __tmp_779_17;
      __tmp_779_19 <= __tmp_779_18;
      __tmp_779_20 <= __tmp_779_19;
      __tmp_779_21 <= __tmp_779_20;
      __tmp_779_22 <= __tmp_779_21;
      __tmp_781_1 <= _tmp_781;
      __tmp_781_2 <= __tmp_781_1;
      __tmp_781_3 <= __tmp_781_2;
      __tmp_781_4 <= __tmp_781_3;
      __tmp_781_5 <= __tmp_781_4;
      __tmp_781_6 <= __tmp_781_5;
      __tmp_781_7 <= __tmp_781_6;
      __tmp_781_8 <= __tmp_781_7;
      __tmp_781_9 <= __tmp_781_8;
      __tmp_781_10 <= __tmp_781_9;
      __tmp_781_11 <= __tmp_781_10;
      __tmp_781_12 <= __tmp_781_11;
      __tmp_781_13 <= __tmp_781_12;
      __tmp_781_14 <= __tmp_781_13;
      __tmp_781_15 <= __tmp_781_14;
      __tmp_781_16 <= __tmp_781_15;
      __tmp_781_17 <= __tmp_781_16;
      __tmp_781_18 <= __tmp_781_17;
      __tmp_781_19 <= __tmp_781_18;
      __tmp_781_20 <= __tmp_781_19;
      __tmp_781_21 <= __tmp_781_20;
      __tmp_781_22 <= __tmp_781_21;
      __tmp_783_1 <= _tmp_783;
      __tmp_783_2 <= __tmp_783_1;
      __tmp_783_3 <= __tmp_783_2;
      __tmp_783_4 <= __tmp_783_3;
      __tmp_783_5 <= __tmp_783_4;
      __tmp_783_6 <= __tmp_783_5;
      __tmp_783_7 <= __tmp_783_6;
      __tmp_783_8 <= __tmp_783_7;
      __tmp_783_9 <= __tmp_783_8;
      __tmp_783_10 <= __tmp_783_9;
      __tmp_783_11 <= __tmp_783_10;
      __tmp_783_12 <= __tmp_783_11;
      __tmp_783_13 <= __tmp_783_12;
      __tmp_783_14 <= __tmp_783_13;
      __tmp_783_15 <= __tmp_783_14;
      __tmp_783_16 <= __tmp_783_15;
      __tmp_783_17 <= __tmp_783_16;
      __tmp_783_18 <= __tmp_783_17;
      __tmp_783_19 <= __tmp_783_18;
      __tmp_783_20 <= __tmp_783_19;
      __tmp_783_21 <= __tmp_783_20;
      __tmp_783_22 <= __tmp_783_21;
      __tmp_785_1 <= _tmp_785;
      __tmp_785_2 <= __tmp_785_1;
      __tmp_785_3 <= __tmp_785_2;
      __tmp_785_4 <= __tmp_785_3;
      __tmp_785_5 <= __tmp_785_4;
      __tmp_785_6 <= __tmp_785_5;
      __tmp_785_7 <= __tmp_785_6;
      __tmp_785_8 <= __tmp_785_7;
      __tmp_785_9 <= __tmp_785_8;
      __tmp_785_10 <= __tmp_785_9;
      __tmp_785_11 <= __tmp_785_10;
      __tmp_785_12 <= __tmp_785_11;
      __tmp_785_13 <= __tmp_785_12;
      __tmp_785_14 <= __tmp_785_13;
      __tmp_785_15 <= __tmp_785_14;
      __tmp_785_16 <= __tmp_785_15;
      __tmp_785_17 <= __tmp_785_16;
      __tmp_785_18 <= __tmp_785_17;
      __tmp_785_19 <= __tmp_785_18;
      __tmp_785_20 <= __tmp_785_19;
      __tmp_785_21 <= __tmp_785_20;
      __tmp_785_22 <= __tmp_785_21;
      __tmp_787_1 <= _tmp_787;
      __tmp_787_2 <= __tmp_787_1;
      __tmp_787_3 <= __tmp_787_2;
      __tmp_787_4 <= __tmp_787_3;
      __tmp_787_5 <= __tmp_787_4;
      __tmp_787_6 <= __tmp_787_5;
      __tmp_787_7 <= __tmp_787_6;
      __tmp_787_8 <= __tmp_787_7;
      __tmp_787_9 <= __tmp_787_8;
      __tmp_787_10 <= __tmp_787_9;
      __tmp_787_11 <= __tmp_787_10;
      __tmp_787_12 <= __tmp_787_11;
      __tmp_787_13 <= __tmp_787_12;
      __tmp_787_14 <= __tmp_787_13;
      __tmp_787_15 <= __tmp_787_14;
      __tmp_787_16 <= __tmp_787_15;
      __tmp_787_17 <= __tmp_787_16;
      __tmp_787_18 <= __tmp_787_17;
      __tmp_787_19 <= __tmp_787_18;
      __tmp_787_20 <= __tmp_787_19;
      __tmp_787_21 <= __tmp_787_20;
      __tmp_787_22 <= __tmp_787_21;
      __tmp_787_23 <= __tmp_787_22;
      __tmp_787_24 <= __tmp_787_23;
      __tmp_787_25 <= __tmp_787_24;
      __tmp_787_26 <= __tmp_787_25;
      __tmp_787_27 <= __tmp_787_26;
      __tmp_787_28 <= __tmp_787_27;
      __tmp_789_1 <= _tmp_789;
      __tmp_789_2 <= __tmp_789_1;
      __tmp_789_3 <= __tmp_789_2;
      __tmp_789_4 <= __tmp_789_3;
      __tmp_789_5 <= __tmp_789_4;
      __tmp_789_6 <= __tmp_789_5;
      __tmp_789_7 <= __tmp_789_6;
      __tmp_789_8 <= __tmp_789_7;
      __tmp_789_9 <= __tmp_789_8;
      __tmp_789_10 <= __tmp_789_9;
      __tmp_789_11 <= __tmp_789_10;
      __tmp_789_12 <= __tmp_789_11;
      __tmp_789_13 <= __tmp_789_12;
      __tmp_789_14 <= __tmp_789_13;
      __tmp_789_15 <= __tmp_789_14;
      __tmp_789_16 <= __tmp_789_15;
      __tmp_789_17 <= __tmp_789_16;
      __tmp_789_18 <= __tmp_789_17;
      __tmp_789_19 <= __tmp_789_18;
      __tmp_789_20 <= __tmp_789_19;
      __tmp_789_21 <= __tmp_789_20;
      __tmp_789_22 <= __tmp_789_21;
      __tmp_789_23 <= __tmp_789_22;
      __tmp_789_24 <= __tmp_789_23;
      __tmp_789_25 <= __tmp_789_24;
      __tmp_789_26 <= __tmp_789_25;
      __tmp_791_1 <= _tmp_791;
      __tmp_791_2 <= __tmp_791_1;
      __tmp_791_3 <= __tmp_791_2;
      __tmp_791_4 <= __tmp_791_3;
      __tmp_791_5 <= __tmp_791_4;
      __tmp_791_6 <= __tmp_791_5;
      __tmp_791_7 <= __tmp_791_6;
      __tmp_791_8 <= __tmp_791_7;
      __tmp_791_9 <= __tmp_791_8;
      __tmp_791_10 <= __tmp_791_9;
      __tmp_791_11 <= __tmp_791_10;
      __tmp_791_12 <= __tmp_791_11;
      __tmp_791_13 <= __tmp_791_12;
      __tmp_791_14 <= __tmp_791_13;
      __tmp_791_15 <= __tmp_791_14;
      __tmp_791_16 <= __tmp_791_15;
      __tmp_791_17 <= __tmp_791_16;
      __tmp_791_18 <= __tmp_791_17;
      __tmp_791_19 <= __tmp_791_18;
      __tmp_791_20 <= __tmp_791_19;
      __tmp_791_21 <= __tmp_791_20;
      __tmp_791_22 <= __tmp_791_21;
      __tmp_791_23 <= __tmp_791_22;
      __tmp_791_24 <= __tmp_791_23;
      __tmp_791_25 <= __tmp_791_24;
      __tmp_791_26 <= __tmp_791_25;
      __tmp_793_1 <= _tmp_793;
      __tmp_793_2 <= __tmp_793_1;
      __tmp_793_3 <= __tmp_793_2;
      __tmp_793_4 <= __tmp_793_3;
      __tmp_793_5 <= __tmp_793_4;
      __tmp_793_6 <= __tmp_793_5;
      __tmp_793_7 <= __tmp_793_6;
      __tmp_793_8 <= __tmp_793_7;
      __tmp_793_9 <= __tmp_793_8;
      __tmp_793_10 <= __tmp_793_9;
      __tmp_793_11 <= __tmp_793_10;
      __tmp_793_12 <= __tmp_793_11;
      __tmp_793_13 <= __tmp_793_12;
      __tmp_793_14 <= __tmp_793_13;
      __tmp_793_15 <= __tmp_793_14;
      __tmp_793_16 <= __tmp_793_15;
      __tmp_793_17 <= __tmp_793_16;
      __tmp_793_18 <= __tmp_793_17;
      __tmp_793_19 <= __tmp_793_18;
      __tmp_793_20 <= __tmp_793_19;
      __tmp_793_21 <= __tmp_793_20;
      __tmp_793_22 <= __tmp_793_21;
      __tmp_793_23 <= __tmp_793_22;
      __tmp_793_24 <= __tmp_793_23;
      __tmp_793_25 <= __tmp_793_24;
      __tmp_793_26 <= __tmp_793_25;
      __tmp_795_1 <= _tmp_795;
      __tmp_795_2 <= __tmp_795_1;
      __tmp_795_3 <= __tmp_795_2;
      __tmp_795_4 <= __tmp_795_3;
      __tmp_795_5 <= __tmp_795_4;
      __tmp_795_6 <= __tmp_795_5;
      __tmp_795_7 <= __tmp_795_6;
      __tmp_795_8 <= __tmp_795_7;
      __tmp_795_9 <= __tmp_795_8;
      __tmp_795_10 <= __tmp_795_9;
      __tmp_795_11 <= __tmp_795_10;
      __tmp_795_12 <= __tmp_795_11;
      __tmp_795_13 <= __tmp_795_12;
      __tmp_795_14 <= __tmp_795_13;
      __tmp_795_15 <= __tmp_795_14;
      __tmp_795_16 <= __tmp_795_15;
      __tmp_795_17 <= __tmp_795_16;
      __tmp_795_18 <= __tmp_795_17;
      __tmp_795_19 <= __tmp_795_18;
      __tmp_795_20 <= __tmp_795_19;
      __tmp_795_21 <= __tmp_795_20;
      __tmp_795_22 <= __tmp_795_21;
      __tmp_795_23 <= __tmp_795_22;
      __tmp_795_24 <= __tmp_795_23;
      __tmp_795_25 <= __tmp_795_24;
      __tmp_795_26 <= __tmp_795_25;
      __tmp_795_27 <= __tmp_795_26;
      __tmp_795_28 <= __tmp_795_27;
      __tmp_795_29 <= __tmp_795_28;
      __tmp_795_30 <= __tmp_795_29;
      __tmp_795_31 <= __tmp_795_30;
      __tmp_795_32 <= __tmp_795_31;
      __tmp_795_33 <= __tmp_795_32;
      __tmp_795_34 <= __tmp_795_33;
      __tmp_797_1 <= _tmp_797;
      __tmp_797_2 <= __tmp_797_1;
      __tmp_797_3 <= __tmp_797_2;
      __tmp_797_4 <= __tmp_797_3;
      __tmp_797_5 <= __tmp_797_4;
      __tmp_797_6 <= __tmp_797_5;
      __tmp_797_7 <= __tmp_797_6;
      __tmp_797_8 <= __tmp_797_7;
      __tmp_797_9 <= __tmp_797_8;
      __tmp_797_10 <= __tmp_797_9;
      __tmp_797_11 <= __tmp_797_10;
      __tmp_797_12 <= __tmp_797_11;
      __tmp_797_13 <= __tmp_797_12;
      __tmp_797_14 <= __tmp_797_13;
      __tmp_797_15 <= __tmp_797_14;
      __tmp_797_16 <= __tmp_797_15;
      __tmp_797_17 <= __tmp_797_16;
      __tmp_797_18 <= __tmp_797_17;
      __tmp_797_19 <= __tmp_797_18;
      __tmp_797_20 <= __tmp_797_19;
      __tmp_797_21 <= __tmp_797_20;
      __tmp_797_22 <= __tmp_797_21;
      __tmp_797_23 <= __tmp_797_22;
      __tmp_797_24 <= __tmp_797_23;
      __tmp_797_25 <= __tmp_797_24;
      __tmp_797_26 <= __tmp_797_25;
      __tmp_797_27 <= __tmp_797_26;
      __tmp_797_28 <= __tmp_797_27;
      __tmp_797_29 <= __tmp_797_28;
      __tmp_797_30 <= __tmp_797_29;
      __tmp_797_31 <= __tmp_797_30;
      __tmp_797_32 <= __tmp_797_31;
      __tmp_797_33 <= __tmp_797_32;
      __tmp_797_34 <= __tmp_797_33;
      __tmp_799_1 <= _tmp_799;
      __tmp_799_2 <= __tmp_799_1;
      __tmp_799_3 <= __tmp_799_2;
      __tmp_799_4 <= __tmp_799_3;
      __tmp_799_5 <= __tmp_799_4;
      __tmp_799_6 <= __tmp_799_5;
      __tmp_799_7 <= __tmp_799_6;
      __tmp_799_8 <= __tmp_799_7;
      __tmp_799_9 <= __tmp_799_8;
      __tmp_799_10 <= __tmp_799_9;
      __tmp_799_11 <= __tmp_799_10;
      __tmp_799_12 <= __tmp_799_11;
      __tmp_799_13 <= __tmp_799_12;
      __tmp_799_14 <= __tmp_799_13;
      __tmp_799_15 <= __tmp_799_14;
      __tmp_799_16 <= __tmp_799_15;
      __tmp_799_17 <= __tmp_799_16;
      __tmp_799_18 <= __tmp_799_17;
      __tmp_799_19 <= __tmp_799_18;
      __tmp_799_20 <= __tmp_799_19;
      __tmp_799_21 <= __tmp_799_20;
      __tmp_799_22 <= __tmp_799_21;
      __tmp_799_23 <= __tmp_799_22;
      __tmp_799_24 <= __tmp_799_23;
      __tmp_799_25 <= __tmp_799_24;
      __tmp_799_26 <= __tmp_799_25;
      __tmp_799_27 <= __tmp_799_26;
      __tmp_799_28 <= __tmp_799_27;
      __tmp_799_29 <= __tmp_799_28;
      __tmp_799_30 <= __tmp_799_29;
      __tmp_799_31 <= __tmp_799_30;
      __tmp_799_32 <= __tmp_799_31;
      __tmp_799_33 <= __tmp_799_32;
      __tmp_799_34 <= __tmp_799_33;
      __tmp_801_1 <= _tmp_801;
      __tmp_803_1 <= _tmp_803;
      __tmp_803_2 <= __tmp_803_1;
      __tmp_803_3 <= __tmp_803_2;
      __tmp_803_4 <= __tmp_803_3;
      __tmp_803_5 <= __tmp_803_4;
      __tmp_803_6 <= __tmp_803_5;
      __tmp_803_7 <= __tmp_803_6;
      __tmp_803_8 <= __tmp_803_7;
      __tmp_803_9 <= __tmp_803_8;
      __tmp_805_1 <= _tmp_805;
      __tmp_805_2 <= __tmp_805_1;
      __tmp_805_3 <= __tmp_805_2;
      __tmp_805_4 <= __tmp_805_3;
      __tmp_805_5 <= __tmp_805_4;
      __tmp_805_6 <= __tmp_805_5;
      __tmp_805_7 <= __tmp_805_6;
      __tmp_805_8 <= __tmp_805_7;
      __tmp_805_9 <= __tmp_805_8;
      __tmp_807_1 <= _tmp_807;
      __tmp_807_2 <= __tmp_807_1;
      __tmp_807_3 <= __tmp_807_2;
      __tmp_807_4 <= __tmp_807_3;
      __tmp_807_5 <= __tmp_807_4;
      __tmp_807_6 <= __tmp_807_5;
      __tmp_807_7 <= __tmp_807_6;
      __tmp_807_8 <= __tmp_807_7;
      __tmp_807_9 <= __tmp_807_8;
      __tmp_815_1 <= _tmp_815;
      __tmp_815_2 <= __tmp_815_1;
      __tmp_815_3 <= __tmp_815_2;
      __tmp_815_4 <= __tmp_815_3;
      __tmp_815_5 <= __tmp_815_4;
      __tmp_815_6 <= __tmp_815_5;
      __tmp_815_7 <= __tmp_815_6;
      __tmp_815_8 <= __tmp_815_7;
      __tmp_815_9 <= __tmp_815_8;
      __tmp_817_1 <= _tmp_817;
      __tmp_817_2 <= __tmp_817_1;
      __tmp_817_3 <= __tmp_817_2;
      __tmp_817_4 <= __tmp_817_3;
      __tmp_817_5 <= __tmp_817_4;
      __tmp_817_6 <= __tmp_817_5;
      __tmp_817_7 <= __tmp_817_6;
      __tmp_817_8 <= __tmp_817_7;
      __tmp_817_9 <= __tmp_817_8;
      __tmp_819_1 <= _tmp_819;
      __tmp_819_2 <= __tmp_819_1;
      __tmp_819_3 <= __tmp_819_2;
      __tmp_819_4 <= __tmp_819_3;
      __tmp_819_5 <= __tmp_819_4;
      __tmp_819_6 <= __tmp_819_5;
      __tmp_819_7 <= __tmp_819_6;
      __tmp_819_8 <= __tmp_819_7;
      __tmp_819_9 <= __tmp_819_8;
      __tmp_827_1 <= _tmp_827;
      __tmp_827_2 <= __tmp_827_1;
      __tmp_827_3 <= __tmp_827_2;
      __tmp_827_4 <= __tmp_827_3;
      __tmp_827_5 <= __tmp_827_4;
      __tmp_827_6 <= __tmp_827_5;
      __tmp_827_7 <= __tmp_827_6;
      __tmp_827_8 <= __tmp_827_7;
      __tmp_827_9 <= __tmp_827_8;
      __tmp_829_1 <= _tmp_829;
      __tmp_829_2 <= __tmp_829_1;
      __tmp_829_3 <= __tmp_829_2;
      __tmp_829_4 <= __tmp_829_3;
      __tmp_829_5 <= __tmp_829_4;
      __tmp_829_6 <= __tmp_829_5;
      __tmp_829_7 <= __tmp_829_6;
      __tmp_829_8 <= __tmp_829_7;
      __tmp_829_9 <= __tmp_829_8;
      __tmp_831_1 <= _tmp_831;
      __tmp_831_2 <= __tmp_831_1;
      __tmp_831_3 <= __tmp_831_2;
      __tmp_831_4 <= __tmp_831_3;
      __tmp_831_5 <= __tmp_831_4;
      __tmp_831_6 <= __tmp_831_5;
      __tmp_831_7 <= __tmp_831_6;
      __tmp_831_8 <= __tmp_831_7;
      __tmp_831_9 <= __tmp_831_8;
      __tmp_839_1 <= _tmp_839;
      __tmp_839_2 <= __tmp_839_1;
      __tmp_839_3 <= __tmp_839_2;
      __tmp_839_4 <= __tmp_839_3;
      __tmp_839_5 <= __tmp_839_4;
      __tmp_839_6 <= __tmp_839_5;
      __tmp_839_7 <= __tmp_839_6;
      __tmp_839_8 <= __tmp_839_7;
      __tmp_839_9 <= __tmp_839_8;
      __tmp_841_1 <= _tmp_841;
      __tmp_841_2 <= __tmp_841_1;
      __tmp_841_3 <= __tmp_841_2;
      __tmp_841_4 <= __tmp_841_3;
      __tmp_841_5 <= __tmp_841_4;
      __tmp_841_6 <= __tmp_841_5;
      __tmp_841_7 <= __tmp_841_6;
      __tmp_841_8 <= __tmp_841_7;
      __tmp_841_9 <= __tmp_841_8;
      __tmp_843_1 <= _tmp_843;
      __tmp_843_2 <= __tmp_843_1;
      __tmp_843_3 <= __tmp_843_2;
      __tmp_843_4 <= __tmp_843_3;
      __tmp_843_5 <= __tmp_843_4;
      __tmp_843_6 <= __tmp_843_5;
      __tmp_843_7 <= __tmp_843_6;
      __tmp_843_8 <= __tmp_843_7;
      __tmp_843_9 <= __tmp_843_8;
      __tmp_851_1 <= _tmp_851;
      __tmp_851_2 <= __tmp_851_1;
      __tmp_851_3 <= __tmp_851_2;
      __tmp_851_4 <= __tmp_851_3;
      __tmp_851_5 <= __tmp_851_4;
      __tmp_851_6 <= __tmp_851_5;
      __tmp_851_7 <= __tmp_851_6;
      __tmp_851_8 <= __tmp_851_7;
      __tmp_851_9 <= __tmp_851_8;
      __tmp_853_1 <= _tmp_853;
      __tmp_853_2 <= __tmp_853_1;
      __tmp_853_3 <= __tmp_853_2;
      __tmp_853_4 <= __tmp_853_3;
      __tmp_853_5 <= __tmp_853_4;
      __tmp_853_6 <= __tmp_853_5;
      __tmp_853_7 <= __tmp_853_6;
      __tmp_853_8 <= __tmp_853_7;
      __tmp_853_9 <= __tmp_853_8;
      __tmp_855_1 <= _tmp_855;
      __tmp_855_2 <= __tmp_855_1;
      __tmp_855_3 <= __tmp_855_2;
      __tmp_855_4 <= __tmp_855_3;
      __tmp_855_5 <= __tmp_855_4;
      __tmp_855_6 <= __tmp_855_5;
      __tmp_855_7 <= __tmp_855_6;
      __tmp_855_8 <= __tmp_855_7;
      __tmp_855_9 <= __tmp_855_8;
      __tmp_863_1 <= _tmp_863;
      __tmp_863_2 <= __tmp_863_1;
      __tmp_863_3 <= __tmp_863_2;
      __tmp_863_4 <= __tmp_863_3;
      __tmp_863_5 <= __tmp_863_4;
      __tmp_863_6 <= __tmp_863_5;
      __tmp_863_7 <= __tmp_863_6;
      __tmp_863_8 <= __tmp_863_7;
      __tmp_863_9 <= __tmp_863_8;
      __tmp_865_1 <= _tmp_865;
      __tmp_865_2 <= __tmp_865_1;
      __tmp_865_3 <= __tmp_865_2;
      __tmp_865_4 <= __tmp_865_3;
      __tmp_865_5 <= __tmp_865_4;
      __tmp_865_6 <= __tmp_865_5;
      __tmp_865_7 <= __tmp_865_6;
      __tmp_865_8 <= __tmp_865_7;
      __tmp_865_9 <= __tmp_865_8;
      __tmp_867_1 <= _tmp_867;
      __tmp_867_2 <= __tmp_867_1;
      __tmp_867_3 <= __tmp_867_2;
      __tmp_867_4 <= __tmp_867_3;
      __tmp_867_5 <= __tmp_867_4;
      __tmp_867_6 <= __tmp_867_5;
      __tmp_867_7 <= __tmp_867_6;
      __tmp_867_8 <= __tmp_867_7;
      __tmp_867_9 <= __tmp_867_8;
      __tmp_875_1 <= _tmp_875;
      __tmp_875_2 <= __tmp_875_1;
      __tmp_875_3 <= __tmp_875_2;
      __tmp_875_4 <= __tmp_875_3;
      __tmp_875_5 <= __tmp_875_4;
      __tmp_875_6 <= __tmp_875_5;
      __tmp_875_7 <= __tmp_875_6;
      __tmp_875_8 <= __tmp_875_7;
      __tmp_875_9 <= __tmp_875_8;
      __tmp_877_1 <= _tmp_877;
      __tmp_877_2 <= __tmp_877_1;
      __tmp_877_3 <= __tmp_877_2;
      __tmp_877_4 <= __tmp_877_3;
      __tmp_877_5 <= __tmp_877_4;
      __tmp_877_6 <= __tmp_877_5;
      __tmp_877_7 <= __tmp_877_6;
      __tmp_877_8 <= __tmp_877_7;
      __tmp_877_9 <= __tmp_877_8;
      __tmp_879_1 <= _tmp_879;
      __tmp_879_2 <= __tmp_879_1;
      __tmp_879_3 <= __tmp_879_2;
      __tmp_879_4 <= __tmp_879_3;
      __tmp_879_5 <= __tmp_879_4;
      __tmp_879_6 <= __tmp_879_5;
      __tmp_879_7 <= __tmp_879_6;
      __tmp_879_8 <= __tmp_879_7;
      __tmp_879_9 <= __tmp_879_8;
      __tmp_887_1 <= _tmp_887;
      __tmp_887_2 <= __tmp_887_1;
      __tmp_887_3 <= __tmp_887_2;
      __tmp_887_4 <= __tmp_887_3;
      __tmp_887_5 <= __tmp_887_4;
      __tmp_887_6 <= __tmp_887_5;
      __tmp_887_7 <= __tmp_887_6;
      __tmp_887_8 <= __tmp_887_7;
      __tmp_887_9 <= __tmp_887_8;
      __tmp_889_1 <= _tmp_889;
      __tmp_889_2 <= __tmp_889_1;
      __tmp_889_3 <= __tmp_889_2;
      __tmp_889_4 <= __tmp_889_3;
      __tmp_889_5 <= __tmp_889_4;
      __tmp_889_6 <= __tmp_889_5;
      __tmp_889_7 <= __tmp_889_6;
      __tmp_889_8 <= __tmp_889_7;
      __tmp_889_9 <= __tmp_889_8;
      __tmp_891_1 <= _tmp_891;
      __tmp_891_2 <= __tmp_891_1;
      __tmp_891_3 <= __tmp_891_2;
      __tmp_891_4 <= __tmp_891_3;
      __tmp_891_5 <= __tmp_891_4;
      __tmp_891_6 <= __tmp_891_5;
      __tmp_891_7 <= __tmp_891_6;
      __tmp_891_8 <= __tmp_891_7;
      __tmp_891_9 <= __tmp_891_8;
      __tmp_899_1 <= _tmp_899;
      __tmp_899_2 <= __tmp_899_1;
      __tmp_899_3 <= __tmp_899_2;
      __tmp_899_4 <= __tmp_899_3;
      __tmp_899_5 <= __tmp_899_4;
      __tmp_899_6 <= __tmp_899_5;
      __tmp_899_7 <= __tmp_899_6;
      __tmp_899_8 <= __tmp_899_7;
      __tmp_899_9 <= __tmp_899_8;
      __tmp_901_1 <= _tmp_901;
      __tmp_901_2 <= __tmp_901_1;
      __tmp_901_3 <= __tmp_901_2;
      __tmp_901_4 <= __tmp_901_3;
      __tmp_901_5 <= __tmp_901_4;
      __tmp_901_6 <= __tmp_901_5;
      __tmp_901_7 <= __tmp_901_6;
      __tmp_901_8 <= __tmp_901_7;
      __tmp_901_9 <= __tmp_901_8;
      __tmp_903_1 <= _tmp_903;
      __tmp_903_2 <= __tmp_903_1;
      __tmp_903_3 <= __tmp_903_2;
      __tmp_903_4 <= __tmp_903_3;
      __tmp_903_5 <= __tmp_903_4;
      __tmp_903_6 <= __tmp_903_5;
      __tmp_903_7 <= __tmp_903_6;
      __tmp_903_8 <= __tmp_903_7;
      __tmp_903_9 <= __tmp_903_8;
      __tmp_911_1 <= _tmp_911;
      __tmp_911_2 <= __tmp_911_1;
      __tmp_911_3 <= __tmp_911_2;
      __tmp_911_4 <= __tmp_911_3;
      __tmp_911_5 <= __tmp_911_4;
      __tmp_911_6 <= __tmp_911_5;
      __tmp_911_7 <= __tmp_911_6;
      __tmp_911_8 <= __tmp_911_7;
      __tmp_911_9 <= __tmp_911_8;
      __tmp_911_10 <= __tmp_911_9;
      __tmp_911_11 <= __tmp_911_10;
      __tmp_911_12 <= __tmp_911_11;
      __tmp_911_13 <= __tmp_911_12;
      __tmp_911_14 <= __tmp_911_13;
      __tmp_911_15 <= __tmp_911_14;
      __tmp_911_16 <= __tmp_911_15;
      __tmp_911_17 <= __tmp_911_16;
      __tmp_911_18 <= __tmp_911_17;
      __tmp_911_19 <= __tmp_911_18;
      __tmp_913_1 <= _tmp_913;
      __tmp_913_2 <= __tmp_913_1;
      __tmp_913_3 <= __tmp_913_2;
      __tmp_913_4 <= __tmp_913_3;
      __tmp_913_5 <= __tmp_913_4;
      __tmp_913_6 <= __tmp_913_5;
      __tmp_913_7 <= __tmp_913_6;
      __tmp_913_8 <= __tmp_913_7;
      __tmp_913_9 <= __tmp_913_8;
      __tmp_913_10 <= __tmp_913_9;
      __tmp_913_11 <= __tmp_913_10;
      __tmp_913_12 <= __tmp_913_11;
      __tmp_913_13 <= __tmp_913_12;
      __tmp_913_14 <= __tmp_913_13;
      __tmp_913_15 <= __tmp_913_14;
      __tmp_913_16 <= __tmp_913_15;
      __tmp_913_17 <= __tmp_913_16;
      __tmp_913_18 <= __tmp_913_17;
      __tmp_913_19 <= __tmp_913_18;
      __tmp_915_1 <= _tmp_915;
      __tmp_915_2 <= __tmp_915_1;
      __tmp_915_3 <= __tmp_915_2;
      __tmp_915_4 <= __tmp_915_3;
      __tmp_915_5 <= __tmp_915_4;
      __tmp_915_6 <= __tmp_915_5;
      __tmp_915_7 <= __tmp_915_6;
      __tmp_915_8 <= __tmp_915_7;
      __tmp_915_9 <= __tmp_915_8;
      __tmp_915_10 <= __tmp_915_9;
      __tmp_915_11 <= __tmp_915_10;
      __tmp_915_12 <= __tmp_915_11;
      __tmp_915_13 <= __tmp_915_12;
      __tmp_915_14 <= __tmp_915_13;
      __tmp_915_15 <= __tmp_915_14;
      __tmp_915_16 <= __tmp_915_15;
      __tmp_915_17 <= __tmp_915_16;
      __tmp_915_18 <= __tmp_915_17;
      __tmp_915_19 <= __tmp_915_18;
      __tmp_917_1 <= _tmp_917;
      __tmp_917_2 <= __tmp_917_1;
      __tmp_917_3 <= __tmp_917_2;
      __tmp_917_4 <= __tmp_917_3;
      __tmp_917_5 <= __tmp_917_4;
      __tmp_917_6 <= __tmp_917_5;
      __tmp_917_7 <= __tmp_917_6;
      __tmp_917_8 <= __tmp_917_7;
      __tmp_917_9 <= __tmp_917_8;
      __tmp_917_10 <= __tmp_917_9;
      __tmp_917_11 <= __tmp_917_10;
      __tmp_917_12 <= __tmp_917_11;
      __tmp_917_13 <= __tmp_917_12;
      __tmp_917_14 <= __tmp_917_13;
      __tmp_917_15 <= __tmp_917_14;
      __tmp_917_16 <= __tmp_917_15;
      __tmp_917_17 <= __tmp_917_16;
      __tmp_917_18 <= __tmp_917_17;
      __tmp_917_19 <= __tmp_917_18;
      __tmp_919_1 <= _tmp_919;
      __tmp_919_2 <= __tmp_919_1;
      __tmp_919_3 <= __tmp_919_2;
      __tmp_919_4 <= __tmp_919_3;
      __tmp_919_5 <= __tmp_919_4;
      __tmp_919_6 <= __tmp_919_5;
      __tmp_919_7 <= __tmp_919_6;
      __tmp_919_8 <= __tmp_919_7;
      __tmp_919_9 <= __tmp_919_8;
      __tmp_919_10 <= __tmp_919_9;
      __tmp_919_11 <= __tmp_919_10;
      __tmp_919_12 <= __tmp_919_11;
      __tmp_919_13 <= __tmp_919_12;
      __tmp_919_14 <= __tmp_919_13;
      __tmp_919_15 <= __tmp_919_14;
      __tmp_919_16 <= __tmp_919_15;
      __tmp_919_17 <= __tmp_919_16;
      __tmp_919_18 <= __tmp_919_17;
      __tmp_919_19 <= __tmp_919_18;
      __tmp_921_1 <= _tmp_921;
      __tmp_921_2 <= __tmp_921_1;
      __tmp_921_3 <= __tmp_921_2;
      __tmp_921_4 <= __tmp_921_3;
      __tmp_921_5 <= __tmp_921_4;
      __tmp_921_6 <= __tmp_921_5;
      __tmp_921_7 <= __tmp_921_6;
      __tmp_921_8 <= __tmp_921_7;
      __tmp_921_9 <= __tmp_921_8;
      __tmp_921_10 <= __tmp_921_9;
      __tmp_921_11 <= __tmp_921_10;
      __tmp_921_12 <= __tmp_921_11;
      __tmp_921_13 <= __tmp_921_12;
      __tmp_921_14 <= __tmp_921_13;
      __tmp_921_15 <= __tmp_921_14;
      __tmp_921_16 <= __tmp_921_15;
      __tmp_921_17 <= __tmp_921_16;
      __tmp_921_18 <= __tmp_921_17;
      __tmp_921_19 <= __tmp_921_18;
      __tmp_923_1 <= _tmp_923;
      __tmp_923_2 <= __tmp_923_1;
      __tmp_923_3 <= __tmp_923_2;
      __tmp_923_4 <= __tmp_923_3;
      __tmp_923_5 <= __tmp_923_4;
      __tmp_923_6 <= __tmp_923_5;
      __tmp_923_7 <= __tmp_923_6;
      __tmp_923_8 <= __tmp_923_7;
      __tmp_923_9 <= __tmp_923_8;
      __tmp_923_10 <= __tmp_923_9;
      __tmp_923_11 <= __tmp_923_10;
      __tmp_923_12 <= __tmp_923_11;
      __tmp_923_13 <= __tmp_923_12;
      __tmp_923_14 <= __tmp_923_13;
      __tmp_923_15 <= __tmp_923_14;
      __tmp_923_16 <= __tmp_923_15;
      __tmp_923_17 <= __tmp_923_16;
      __tmp_923_18 <= __tmp_923_17;
      __tmp_923_19 <= __tmp_923_18;
      __tmp_925_1 <= _tmp_925;
      __tmp_925_2 <= __tmp_925_1;
      __tmp_925_3 <= __tmp_925_2;
      __tmp_925_4 <= __tmp_925_3;
      __tmp_925_5 <= __tmp_925_4;
      __tmp_925_6 <= __tmp_925_5;
      __tmp_925_7 <= __tmp_925_6;
      __tmp_925_8 <= __tmp_925_7;
      __tmp_925_9 <= __tmp_925_8;
      __tmp_925_10 <= __tmp_925_9;
      __tmp_925_11 <= __tmp_925_10;
      __tmp_925_12 <= __tmp_925_11;
      __tmp_925_13 <= __tmp_925_12;
      __tmp_925_14 <= __tmp_925_13;
      __tmp_925_15 <= __tmp_925_14;
      __tmp_925_16 <= __tmp_925_15;
      __tmp_925_17 <= __tmp_925_16;
      __tmp_925_18 <= __tmp_925_17;
      __tmp_925_19 <= __tmp_925_18;
      __tmp_927_1 <= _tmp_927;
      __tmp_927_2 <= __tmp_927_1;
      __tmp_927_3 <= __tmp_927_2;
      __tmp_927_4 <= __tmp_927_3;
      __tmp_927_5 <= __tmp_927_4;
      __tmp_927_6 <= __tmp_927_5;
      __tmp_927_7 <= __tmp_927_6;
      __tmp_927_8 <= __tmp_927_7;
      __tmp_927_9 <= __tmp_927_8;
      __tmp_927_10 <= __tmp_927_9;
      __tmp_927_11 <= __tmp_927_10;
      __tmp_927_12 <= __tmp_927_11;
      __tmp_927_13 <= __tmp_927_12;
      __tmp_927_14 <= __tmp_927_13;
      __tmp_927_15 <= __tmp_927_14;
      __tmp_927_16 <= __tmp_927_15;
      __tmp_927_17 <= __tmp_927_16;
      __tmp_927_18 <= __tmp_927_17;
      __tmp_927_19 <= __tmp_927_18;
      __tmp_935_1 <= _tmp_935;
      __tmp_935_2 <= __tmp_935_1;
      __tmp_935_3 <= __tmp_935_2;
      __tmp_935_4 <= __tmp_935_3;
      __tmp_935_5 <= __tmp_935_4;
      __tmp_935_6 <= __tmp_935_5;
      __tmp_935_7 <= __tmp_935_6;
      __tmp_935_8 <= __tmp_935_7;
      __tmp_935_9 <= __tmp_935_8;
      __tmp_935_10 <= __tmp_935_9;
      __tmp_935_11 <= __tmp_935_10;
      __tmp_935_12 <= __tmp_935_11;
      __tmp_935_13 <= __tmp_935_12;
      __tmp_935_14 <= __tmp_935_13;
      __tmp_935_15 <= __tmp_935_14;
      __tmp_935_16 <= __tmp_935_15;
      __tmp_935_17 <= __tmp_935_16;
      __tmp_935_18 <= __tmp_935_17;
      __tmp_935_19 <= __tmp_935_18;
      __tmp_935_20 <= __tmp_935_19;
      __tmp_935_21 <= __tmp_935_20;
      __tmp_935_22 <= __tmp_935_21;
      __tmp_935_23 <= __tmp_935_22;
      __tmp_935_24 <= __tmp_935_23;
      __tmp_937_1 <= _tmp_937;
      __tmp_937_2 <= __tmp_937_1;
      __tmp_937_3 <= __tmp_937_2;
      __tmp_937_4 <= __tmp_937_3;
      __tmp_937_5 <= __tmp_937_4;
      __tmp_937_6 <= __tmp_937_5;
      __tmp_937_7 <= __tmp_937_6;
      __tmp_937_8 <= __tmp_937_7;
      __tmp_937_9 <= __tmp_937_8;
      __tmp_937_10 <= __tmp_937_9;
      __tmp_937_11 <= __tmp_937_10;
      __tmp_937_12 <= __tmp_937_11;
      __tmp_937_13 <= __tmp_937_12;
      __tmp_937_14 <= __tmp_937_13;
      __tmp_937_15 <= __tmp_937_14;
      __tmp_937_16 <= __tmp_937_15;
      __tmp_937_17 <= __tmp_937_16;
      __tmp_937_18 <= __tmp_937_17;
      __tmp_937_19 <= __tmp_937_18;
      __tmp_937_20 <= __tmp_937_19;
      __tmp_937_21 <= __tmp_937_20;
      __tmp_937_22 <= __tmp_937_21;
      __tmp_937_23 <= __tmp_937_22;
      __tmp_939_1 <= _tmp_939;
      __tmp_939_2 <= __tmp_939_1;
      __tmp_939_3 <= __tmp_939_2;
      __tmp_939_4 <= __tmp_939_3;
      __tmp_939_5 <= __tmp_939_4;
      __tmp_939_6 <= __tmp_939_5;
      __tmp_939_7 <= __tmp_939_6;
      __tmp_939_8 <= __tmp_939_7;
      __tmp_939_9 <= __tmp_939_8;
      __tmp_939_10 <= __tmp_939_9;
      __tmp_939_11 <= __tmp_939_10;
      __tmp_939_12 <= __tmp_939_11;
      __tmp_939_13 <= __tmp_939_12;
      __tmp_939_14 <= __tmp_939_13;
      __tmp_939_15 <= __tmp_939_14;
      __tmp_939_16 <= __tmp_939_15;
      __tmp_939_17 <= __tmp_939_16;
      __tmp_939_18 <= __tmp_939_17;
      __tmp_939_19 <= __tmp_939_18;
      __tmp_939_20 <= __tmp_939_19;
      __tmp_939_21 <= __tmp_939_20;
      __tmp_939_22 <= __tmp_939_21;
      __tmp_939_23 <= __tmp_939_22;
      __tmp_941_1 <= _tmp_941;
      __tmp_941_2 <= __tmp_941_1;
      __tmp_941_3 <= __tmp_941_2;
      __tmp_941_4 <= __tmp_941_3;
      __tmp_941_5 <= __tmp_941_4;
      __tmp_941_6 <= __tmp_941_5;
      __tmp_941_7 <= __tmp_941_6;
      __tmp_941_8 <= __tmp_941_7;
      __tmp_941_9 <= __tmp_941_8;
      __tmp_941_10 <= __tmp_941_9;
      __tmp_941_11 <= __tmp_941_10;
      __tmp_941_12 <= __tmp_941_11;
      __tmp_941_13 <= __tmp_941_12;
      __tmp_941_14 <= __tmp_941_13;
      __tmp_941_15 <= __tmp_941_14;
      __tmp_941_16 <= __tmp_941_15;
      __tmp_941_17 <= __tmp_941_16;
      __tmp_941_18 <= __tmp_941_17;
      __tmp_941_19 <= __tmp_941_18;
      __tmp_941_20 <= __tmp_941_19;
      __tmp_941_21 <= __tmp_941_20;
      __tmp_941_22 <= __tmp_941_21;
      __tmp_941_23 <= __tmp_941_22;
      __tmp_949_1 <= _tmp_949;
      __tmp_949_2 <= __tmp_949_1;
      __tmp_949_3 <= __tmp_949_2;
      __tmp_949_4 <= __tmp_949_3;
      __tmp_949_5 <= __tmp_949_4;
      __tmp_949_6 <= __tmp_949_5;
      __tmp_949_7 <= __tmp_949_6;
      __tmp_949_8 <= __tmp_949_7;
      __tmp_949_9 <= __tmp_949_8;
      __tmp_949_10 <= __tmp_949_9;
      __tmp_949_11 <= __tmp_949_10;
      __tmp_949_12 <= __tmp_949_11;
      __tmp_949_13 <= __tmp_949_12;
      __tmp_949_14 <= __tmp_949_13;
      __tmp_949_15 <= __tmp_949_14;
      __tmp_949_16 <= __tmp_949_15;
      __tmp_949_17 <= __tmp_949_16;
      __tmp_949_18 <= __tmp_949_17;
      __tmp_949_19 <= __tmp_949_18;
      __tmp_949_20 <= __tmp_949_19;
      __tmp_949_21 <= __tmp_949_20;
      __tmp_949_22 <= __tmp_949_21;
      __tmp_949_23 <= __tmp_949_22;
      __tmp_949_24 <= __tmp_949_23;
      __tmp_949_25 <= __tmp_949_24;
      __tmp_949_26 <= __tmp_949_25;
      __tmp_949_27 <= __tmp_949_26;
      __tmp_949_28 <= __tmp_949_27;
      __tmp_949_29 <= __tmp_949_28;
      __tmp_949_30 <= __tmp_949_29;
      __tmp_949_31 <= __tmp_949_30;
      __tmp_951_1 <= _tmp_951;
      __tmp_951_2 <= __tmp_951_1;
      __tmp_951_3 <= __tmp_951_2;
      __tmp_951_4 <= __tmp_951_3;
      __tmp_951_5 <= __tmp_951_4;
      __tmp_951_6 <= __tmp_951_5;
      __tmp_951_7 <= __tmp_951_6;
      __tmp_951_8 <= __tmp_951_7;
      __tmp_951_9 <= __tmp_951_8;
      __tmp_951_10 <= __tmp_951_9;
      __tmp_951_11 <= __tmp_951_10;
      __tmp_951_12 <= __tmp_951_11;
      __tmp_951_13 <= __tmp_951_12;
      __tmp_951_14 <= __tmp_951_13;
      __tmp_951_15 <= __tmp_951_14;
      __tmp_951_16 <= __tmp_951_15;
      __tmp_951_17 <= __tmp_951_16;
      __tmp_951_18 <= __tmp_951_17;
      __tmp_951_19 <= __tmp_951_18;
      __tmp_951_20 <= __tmp_951_19;
      __tmp_951_21 <= __tmp_951_20;
      __tmp_951_22 <= __tmp_951_21;
      __tmp_951_23 <= __tmp_951_22;
      __tmp_951_24 <= __tmp_951_23;
      __tmp_951_25 <= __tmp_951_24;
      __tmp_951_26 <= __tmp_951_25;
      __tmp_951_27 <= __tmp_951_26;
      __tmp_951_28 <= __tmp_951_27;
      __tmp_951_29 <= __tmp_951_28;
      __tmp_951_30 <= __tmp_951_29;
      __tmp_951_31 <= __tmp_951_30;
      __tmp_953_1 <= _tmp_953;
      __tmp_953_2 <= __tmp_953_1;
      __tmp_953_3 <= __tmp_953_2;
      __tmp_953_4 <= __tmp_953_3;
      __tmp_953_5 <= __tmp_953_4;
      __tmp_953_6 <= __tmp_953_5;
      __tmp_953_7 <= __tmp_953_6;
      __tmp_953_8 <= __tmp_953_7;
      __tmp_953_9 <= __tmp_953_8;
      __tmp_953_10 <= __tmp_953_9;
      __tmp_953_11 <= __tmp_953_10;
      __tmp_953_12 <= __tmp_953_11;
      __tmp_953_13 <= __tmp_953_12;
      __tmp_953_14 <= __tmp_953_13;
      __tmp_953_15 <= __tmp_953_14;
      __tmp_953_16 <= __tmp_953_15;
      __tmp_953_17 <= __tmp_953_16;
      __tmp_953_18 <= __tmp_953_17;
      __tmp_953_19 <= __tmp_953_18;
      __tmp_953_20 <= __tmp_953_19;
      __tmp_953_21 <= __tmp_953_20;
      __tmp_953_22 <= __tmp_953_21;
      __tmp_953_23 <= __tmp_953_22;
      __tmp_953_24 <= __tmp_953_23;
      __tmp_953_25 <= __tmp_953_24;
      __tmp_953_26 <= __tmp_953_25;
      __tmp_953_27 <= __tmp_953_26;
      __tmp_953_28 <= __tmp_953_27;
      __tmp_953_29 <= __tmp_953_28;
      __tmp_953_30 <= __tmp_953_29;
      __tmp_953_31 <= __tmp_953_30;
      __tmp_961_1 <= _tmp_961;
      __tmp_961_2 <= __tmp_961_1;
      __tmp_961_3 <= __tmp_961_2;
      __tmp_961_4 <= __tmp_961_3;
      __tmp_961_5 <= __tmp_961_4;
      __tmp_961_6 <= __tmp_961_5;
      __tmp_961_7 <= __tmp_961_6;
      __tmp_961_8 <= __tmp_961_7;
      __tmp_961_9 <= __tmp_961_8;
      __tmp_961_10 <= __tmp_961_9;
      __tmp_961_11 <= __tmp_961_10;
      __tmp_961_12 <= __tmp_961_11;
      __tmp_961_13 <= __tmp_961_12;
      __tmp_961_14 <= __tmp_961_13;
      __tmp_961_15 <= __tmp_961_14;
      __tmp_961_16 <= __tmp_961_15;
      __tmp_961_17 <= __tmp_961_16;
      __tmp_961_18 <= __tmp_961_17;
      __tmp_961_19 <= __tmp_961_18;
      __tmp_961_20 <= __tmp_961_19;
      __tmp_961_21 <= __tmp_961_20;
      __tmp_961_22 <= __tmp_961_21;
      __tmp_961_23 <= __tmp_961_22;
      __tmp_961_24 <= __tmp_961_23;
      __tmp_961_25 <= __tmp_961_24;
      __tmp_961_26 <= __tmp_961_25;
      __tmp_961_27 <= __tmp_961_26;
      __tmp_961_28 <= __tmp_961_27;
      __tmp_961_29 <= __tmp_961_28;
      __tmp_961_30 <= __tmp_961_29;
      __tmp_961_31 <= __tmp_961_30;
      __tmp_961_32 <= __tmp_961_31;
      __tmp_961_33 <= __tmp_961_32;
      __tmp_961_34 <= __tmp_961_33;
      __tmp_961_35 <= __tmp_961_34;
      __tmp_961_36 <= __tmp_961_35;
      __tmp_961_37 <= __tmp_961_36;
      __tmp_961_38 <= __tmp_961_37;
      __tmp_961_39 <= __tmp_961_38;
      __tmp_961_40 <= __tmp_961_39;
      __tmp_961_41 <= __tmp_961_40;
      __tmp_961_42 <= __tmp_961_41;
      __tmp_961_43 <= __tmp_961_42;
      __tmp_961_44 <= __tmp_961_43;
      __tmp_961_45 <= __tmp_961_44;
      __tmp_961_46 <= __tmp_961_45;
      __tmp_963_1 <= _tmp_963;
      __tmp_963_2 <= __tmp_963_1;
      __tmp_963_3 <= __tmp_963_2;
      __tmp_963_4 <= __tmp_963_3;
      __tmp_963_5 <= __tmp_963_4;
      __tmp_963_6 <= __tmp_963_5;
      __tmp_963_7 <= __tmp_963_6;
      __tmp_963_8 <= __tmp_963_7;
      __tmp_963_9 <= __tmp_963_8;
      __tmp_963_10 <= __tmp_963_9;
      __tmp_963_11 <= __tmp_963_10;
      __tmp_963_12 <= __tmp_963_11;
      __tmp_963_13 <= __tmp_963_12;
      __tmp_963_14 <= __tmp_963_13;
      __tmp_963_15 <= __tmp_963_14;
      __tmp_963_16 <= __tmp_963_15;
      __tmp_963_17 <= __tmp_963_16;
      __tmp_963_18 <= __tmp_963_17;
      __tmp_963_19 <= __tmp_963_18;
      __tmp_963_20 <= __tmp_963_19;
      __tmp_963_21 <= __tmp_963_20;
      __tmp_963_22 <= __tmp_963_21;
      __tmp_963_23 <= __tmp_963_22;
      __tmp_963_24 <= __tmp_963_23;
      __tmp_963_25 <= __tmp_963_24;
      __tmp_963_26 <= __tmp_963_25;
      __tmp_963_27 <= __tmp_963_26;
      __tmp_963_28 <= __tmp_963_27;
      __tmp_963_29 <= __tmp_963_28;
      __tmp_963_30 <= __tmp_963_29;
      __tmp_963_31 <= __tmp_963_30;
      __tmp_963_32 <= __tmp_963_31;
      __tmp_963_33 <= __tmp_963_32;
      __tmp_963_34 <= __tmp_963_33;
      __tmp_963_35 <= __tmp_963_34;
      __tmp_963_36 <= __tmp_963_35;
      __tmp_963_37 <= __tmp_963_36;
      __tmp_963_38 <= __tmp_963_37;
      __tmp_963_39 <= __tmp_963_38;
      __tmp_963_40 <= __tmp_963_39;
      __tmp_963_41 <= __tmp_963_40;
      __tmp_963_42 <= __tmp_963_41;
      __tmp_963_43 <= __tmp_963_42;
      __tmp_963_44 <= __tmp_963_43;
      __tmp_963_45 <= __tmp_963_44;
      __tmp_963_46 <= __tmp_963_45;
      __tmp_965_1 <= _tmp_965;
      __tmp_965_2 <= __tmp_965_1;
      __tmp_965_3 <= __tmp_965_2;
      __tmp_965_4 <= __tmp_965_3;
      __tmp_965_5 <= __tmp_965_4;
      __tmp_965_6 <= __tmp_965_5;
      __tmp_965_7 <= __tmp_965_6;
      __tmp_965_8 <= __tmp_965_7;
      __tmp_965_9 <= __tmp_965_8;
      __tmp_965_10 <= __tmp_965_9;
      __tmp_965_11 <= __tmp_965_10;
      __tmp_965_12 <= __tmp_965_11;
      __tmp_965_13 <= __tmp_965_12;
      __tmp_965_14 <= __tmp_965_13;
      __tmp_965_15 <= __tmp_965_14;
      __tmp_965_16 <= __tmp_965_15;
      __tmp_965_17 <= __tmp_965_16;
      __tmp_965_18 <= __tmp_965_17;
      __tmp_965_19 <= __tmp_965_18;
      __tmp_965_20 <= __tmp_965_19;
      __tmp_965_21 <= __tmp_965_20;
      __tmp_965_22 <= __tmp_965_21;
      __tmp_965_23 <= __tmp_965_22;
      __tmp_965_24 <= __tmp_965_23;
      __tmp_965_25 <= __tmp_965_24;
      __tmp_965_26 <= __tmp_965_25;
      __tmp_965_27 <= __tmp_965_26;
      __tmp_965_28 <= __tmp_965_27;
      __tmp_965_29 <= __tmp_965_28;
      __tmp_965_30 <= __tmp_965_29;
      __tmp_965_31 <= __tmp_965_30;
      __tmp_965_32 <= __tmp_965_31;
      __tmp_965_33 <= __tmp_965_32;
      __tmp_965_34 <= __tmp_965_33;
      __tmp_965_35 <= __tmp_965_34;
      __tmp_965_36 <= __tmp_965_35;
      __tmp_965_37 <= __tmp_965_36;
      __tmp_965_38 <= __tmp_965_37;
      __tmp_965_39 <= __tmp_965_38;
      __tmp_965_40 <= __tmp_965_39;
      __tmp_965_41 <= __tmp_965_40;
      __tmp_965_42 <= __tmp_965_41;
      __tmp_965_43 <= __tmp_965_42;
      __tmp_965_44 <= __tmp_965_43;
      __tmp_965_45 <= __tmp_965_44;
      __tmp_965_46 <= __tmp_965_45;
      __tmp_967_1 <= _tmp_967;
      __tmp_967_2 <= __tmp_967_1;
      __tmp_967_3 <= __tmp_967_2;
      __tmp_967_4 <= __tmp_967_3;
      __tmp_967_5 <= __tmp_967_4;
      __tmp_967_6 <= __tmp_967_5;
      __tmp_967_7 <= __tmp_967_6;
      __tmp_967_8 <= __tmp_967_7;
      __tmp_967_9 <= __tmp_967_8;
      __tmp_967_10 <= __tmp_967_9;
      __tmp_967_11 <= __tmp_967_10;
      __tmp_967_12 <= __tmp_967_11;
      __tmp_967_13 <= __tmp_967_12;
      __tmp_967_14 <= __tmp_967_13;
      __tmp_967_15 <= __tmp_967_14;
      __tmp_967_16 <= __tmp_967_15;
      __tmp_967_17 <= __tmp_967_16;
      __tmp_967_18 <= __tmp_967_17;
      __tmp_967_19 <= __tmp_967_18;
      __tmp_967_20 <= __tmp_967_19;
      __tmp_967_21 <= __tmp_967_20;
      __tmp_967_22 <= __tmp_967_21;
      __tmp_967_23 <= __tmp_967_22;
      __tmp_967_24 <= __tmp_967_23;
      __tmp_967_25 <= __tmp_967_24;
      __tmp_967_26 <= __tmp_967_25;
      __tmp_967_27 <= __tmp_967_26;
      __tmp_967_28 <= __tmp_967_27;
      __tmp_967_29 <= __tmp_967_28;
      __tmp_967_30 <= __tmp_967_29;
      __tmp_967_31 <= __tmp_967_30;
      __tmp_967_32 <= __tmp_967_31;
      __tmp_967_33 <= __tmp_967_32;
      __tmp_967_34 <= __tmp_967_33;
      __tmp_967_35 <= __tmp_967_34;
      __tmp_967_36 <= __tmp_967_35;
      __tmp_967_37 <= __tmp_967_36;
      __tmp_967_38 <= __tmp_967_37;
      __tmp_967_39 <= __tmp_967_38;
      __tmp_967_40 <= __tmp_967_39;
      __tmp_967_41 <= __tmp_967_40;
      __tmp_967_42 <= __tmp_967_41;
      __tmp_967_43 <= __tmp_967_42;
      __tmp_967_44 <= __tmp_967_43;
      __tmp_967_45 <= __tmp_967_44;
      __tmp_967_46 <= __tmp_967_45;
      __tmp_969_1 <= _tmp_969;
      __tmp_969_2 <= __tmp_969_1;
      __tmp_969_3 <= __tmp_969_2;
      __tmp_969_4 <= __tmp_969_3;
      __tmp_969_5 <= __tmp_969_4;
      __tmp_969_6 <= __tmp_969_5;
      __tmp_969_7 <= __tmp_969_6;
      __tmp_969_8 <= __tmp_969_7;
      __tmp_969_9 <= __tmp_969_8;
      __tmp_969_10 <= __tmp_969_9;
      __tmp_969_11 <= __tmp_969_10;
      __tmp_969_12 <= __tmp_969_11;
      __tmp_969_13 <= __tmp_969_12;
      __tmp_969_14 <= __tmp_969_13;
      __tmp_969_15 <= __tmp_969_14;
      __tmp_969_16 <= __tmp_969_15;
      __tmp_969_17 <= __tmp_969_16;
      __tmp_969_18 <= __tmp_969_17;
      __tmp_969_19 <= __tmp_969_18;
      __tmp_969_20 <= __tmp_969_19;
      __tmp_969_21 <= __tmp_969_20;
      __tmp_969_22 <= __tmp_969_21;
      __tmp_969_23 <= __tmp_969_22;
      __tmp_969_24 <= __tmp_969_23;
      __tmp_969_25 <= __tmp_969_24;
      __tmp_969_26 <= __tmp_969_25;
      __tmp_969_27 <= __tmp_969_26;
      __tmp_969_28 <= __tmp_969_27;
      __tmp_969_29 <= __tmp_969_28;
      __tmp_969_30 <= __tmp_969_29;
      __tmp_969_31 <= __tmp_969_30;
      __tmp_969_32 <= __tmp_969_31;
      __tmp_969_33 <= __tmp_969_32;
      __tmp_969_34 <= __tmp_969_33;
      __tmp_969_35 <= __tmp_969_34;
      __tmp_969_36 <= __tmp_969_35;
      __tmp_969_37 <= __tmp_969_36;
      __tmp_969_38 <= __tmp_969_37;
      __tmp_969_39 <= __tmp_969_38;
      __tmp_969_40 <= __tmp_969_39;
      __tmp_969_41 <= __tmp_969_40;
      __tmp_969_42 <= __tmp_969_41;
    end
  end

  localparam _stream_conv2d_16_fsm_1 = 1;
  localparam _stream_conv2d_16_fsm_2 = 2;
  localparam _stream_conv2d_16_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_fsm <= _stream_conv2d_16_fsm_init;
      _stream_conv2d_16_start <= 0;
      _stream_conv2d_16_source_busy <= 0;
      _stream_conv2d_16_reduce_reset <= 1;
      _stream_conv2d_16_sink_busy <= 0;
      _stream_conv2d_16_sink_wait_count <= 0;
      _stream_conv2d_16_end_flag <= 0;
      _stream_conv2d_16_term_sink <= 0;
    end else begin
      _stream_conv2d_16_start <= 0;
      if(__tmp_713_5) begin
        _stream_conv2d_16_reduce_reset <= 0;
      end 
      if(__tmp_801_1) begin
        _stream_conv2d_16_reduce_reset <= 1;
      end 
      if((_stream_conv2d_16_sink_wait_count == 1) && !((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_961_46) begin
        _stream_conv2d_16_sink_busy <= 0;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) begin
        _stream_conv2d_16_sink_busy <= 1;
      end 
      if(!((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag) && __tmp_963_46) begin
        _stream_conv2d_16_sink_wait_count <= _stream_conv2d_16_sink_wait_count - 1;
      end 
      if((_stream_conv2d_16_fsm == 0) && _stream_conv2d_16_start_flag && !__tmp_965_46) begin
        _stream_conv2d_16_sink_wait_count <= _stream_conv2d_16_sink_wait_count + 1;
      end 
      _stream_conv2d_16_end_flag <= 0;
      if(__tmp_967_46) begin
        _stream_conv2d_16_end_flag <= 1;
      end 
      _stream_conv2d_16_term_sink <= 0;
      if(__tmp_969_42) begin
        _stream_conv2d_16_term_sink <= 1;
      end 
      case(_stream_conv2d_16_fsm)
        _stream_conv2d_16_fsm_init: begin
          if(_stream_conv2d_16_start_flag) begin
            _stream_conv2d_16_start <= 1;
            _stream_conv2d_16_source_busy <= 1;
          end 
          if(_stream_conv2d_16_start_flag) begin
            _stream_conv2d_16_fsm <= _stream_conv2d_16_fsm_1;
          end 
        end
        _stream_conv2d_16_fsm_1: begin
          _stream_conv2d_16_fsm <= _stream_conv2d_16_fsm_2;
        end
        _stream_conv2d_16_fsm_2: begin
          if(_stream_conv2d_16_done) begin
            _stream_conv2d_16_fsm <= _stream_conv2d_16_fsm_3;
          end 
        end
        _stream_conv2d_16_fsm_3: begin
          _stream_conv2d_16_source_busy <= 0;
          _stream_conv2d_16_fsm <= _stream_conv2d_16_fsm_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_18_source_1_idle <= 1;
      _stream_max_pool_serial_18_source_1_source_ram_rvalid <= 0;
      _stream_max_pool_serial_18_sink_3_sink_wenable <= 0;
      _stream_max_pool_serial_18_sink_4_sink_wenable <= 0;
      _counter_count_782 <= 1'sd0;
      _counter_data_782 <= 1'sd0;
      __delay_data_1411 <= 0;
      __delay_data_1412 <= 0;
      __delay_data_1414 <= 0;
      _pointer_data_784 <= 0;
      __delay_data_1413 <= 0;
      __delay_data_1415 <= 0;
      _cond_data_791 <= 0;
      __delay_data_1416 <= 0;
      __substreamoutput_data_793 <= 0;
      __substreamoutput_data_794 <= 0;
      _set_flag_1024 <= 0;
      _stream_max_pool_serial_18_constant_0_next_constant_data <= 0;
      __variable_wdata_777 <= 0;
      _set_flag_1025 <= 0;
      _stream_max_pool_serial_18_constant_2_next_constant_data <= 0;
      __variable_wdata_779 <= 0;
      _set_flag_1026 <= 0;
      _stream_max_pool_serial_18_source_1_source_mode <= 3'b0;
      _stream_max_pool_serial_18_source_1_source_offset <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_size_0 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_stride_0 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_size_1 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_stride_1 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_size_2 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_stride_2 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_size_3 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_stride_3 <= 0;
      _stream_max_pool_serial_18_source_1_source_ram_sel <= 0;
      __tmp_1035_1 <= 0;
      __variable_wdata_778 <= 0;
      _stream_max_pool_serial_18_source_1_source_offset_buf <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_cur_offset_0 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_cur_offset_1 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_cur_offset_2 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_cur_offset_3 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_count_0 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_count_1 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_count_2 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_count_3 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_size_buf_0 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_size_buf_1 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_size_buf_2 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_size_buf_3 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_stride_buf_0 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_stride_buf_1 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_stride_buf_2 <= 0;
      _source_stream_max_pool_serial_18_source_1_pat_stride_buf_3 <= 0;
      _stream_max_pool_serial_18_source_1_source_ram_raddr <= 0;
      _stream_max_pool_serial_18_source_1_source_ram_renable <= 0;
      _set_flag_1036 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_1 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_2 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_3 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_4 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_5 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_6 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_7 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_8 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_9 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_size_1_1 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_size_1_2 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_size_1_3 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_size_1_4 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_size_1_5 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_size_1_6 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_size_1_7 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_size_1_8 <= 0;
      __stream_max_pool_serial_18_sink_3_sink_size_1_9 <= 0;
      __stream_seq_15_cond_2_1 <= 0;
      __stream_seq_15_cond_2_2 <= 0;
      __stream_seq_15_cond_2_3 <= 0;
      __stream_seq_15_cond_2_4 <= 0;
      __stream_seq_15_cond_2_5 <= 0;
      __stream_seq_15_cond_2_6 <= 0;
      __stream_seq_15_cond_2_7 <= 0;
      __stream_seq_15_cond_2_8 <= 0;
      __stream_seq_15_cond_2_9 <= 0;
      _stream_max_pool_serial_18_sink_3_sink_mode <= 3'b0;
      _stream_max_pool_serial_18_sink_3_sink_offset <= 0;
      _stream_max_pool_serial_18_sink_3_sink_size <= 0;
      _stream_max_pool_serial_18_sink_3_sink_stride <= 0;
      __set_flag_1036_1 <= 0;
      __set_flag_1036_2 <= 0;
      __set_flag_1036_3 <= 0;
      __set_flag_1036_4 <= 0;
      __set_flag_1036_5 <= 0;
      __set_flag_1036_6 <= 0;
      __set_flag_1036_7 <= 0;
      __set_flag_1036_8 <= 0;
      __set_flag_1036_9 <= 0;
      _stream_max_pool_serial_18_sink_3_sink_ram_sel <= 0;
      __stream_max_pool_serial_18_start_1 <= 0;
      __stream_max_pool_serial_18_start_2 <= 0;
      __stream_max_pool_serial_18_start_3 <= 0;
      __stream_max_pool_serial_18_start_4 <= 0;
      __stream_max_pool_serial_18_start_5 <= 0;
      __stream_max_pool_serial_18_start_6 <= 0;
      __stream_max_pool_serial_18_start_7 <= 0;
      __stream_max_pool_serial_18_start_8 <= 0;
      __stream_max_pool_serial_18_start_9 <= 0;
      __stream_max_pool_serial_18_start_10 <= 0;
      _stream_max_pool_serial_18_sink_3_sink_waddr <= 0;
      _stream_max_pool_serial_18_sink_3_sink_count <= 0;
      _stream_max_pool_serial_18_sink_3_sink_offset_buf <= 0;
      _stream_max_pool_serial_18_sink_3_sink_stride_buf <= 0;
      _stream_max_pool_serial_18_sink_3_sink_wdata <= 0;
      _set_flag_1038 <= 0;
      __tmp_1040_1 <= 0;
      __tmp_1040_2 <= 0;
      __tmp_1040_3 <= 0;
      __tmp_1040_4 <= 0;
      __tmp_1040_5 <= 0;
      __tmp_1042_1 <= 0;
      __tmp_1042_2 <= 0;
      __tmp_1042_3 <= 0;
      __tmp_1042_4 <= 0;
      __tmp_1042_5 <= 0;
      __tmp_1042_6 <= 0;
      __tmp_1042_7 <= 0;
      __tmp_1042_8 <= 0;
      __tmp_1042_9 <= 0;
      __tmp_1044_1 <= 0;
      __tmp_1044_2 <= 0;
      __tmp_1044_3 <= 0;
      __tmp_1044_4 <= 0;
      __tmp_1044_5 <= 0;
      __tmp_1044_6 <= 0;
      __tmp_1044_7 <= 0;
      __tmp_1046_1 <= 0;
      __tmp_1046_2 <= 0;
      __tmp_1046_3 <= 0;
      __tmp_1046_4 <= 0;
      __tmp_1046_5 <= 0;
      __tmp_1046_6 <= 0;
      __tmp_1046_7 <= 0;
      __tmp_1048_1 <= 0;
      __tmp_1050_1 <= 0;
      __tmp_1050_2 <= 0;
      __tmp_1050_3 <= 0;
      __tmp_1050_4 <= 0;
      __tmp_1050_5 <= 0;
      __tmp_1052_1 <= 0;
      __tmp_1052_2 <= 0;
      __tmp_1052_3 <= 0;
      __tmp_1052_4 <= 0;
      __tmp_1054_1 <= 0;
      __tmp_1054_2 <= 0;
      __tmp_1054_3 <= 0;
      __tmp_1054_4 <= 0;
      __tmp_1062_1 <= 0;
      __tmp_1062_2 <= 0;
      __tmp_1062_3 <= 0;
      __tmp_1062_4 <= 0;
      __tmp_1062_5 <= 0;
      __tmp_1062_6 <= 0;
      __tmp_1062_7 <= 0;
      __tmp_1062_8 <= 0;
      __tmp_1062_9 <= 0;
      __tmp_1062_10 <= 0;
      __tmp_1064_1 <= 0;
      __tmp_1064_2 <= 0;
      __tmp_1064_3 <= 0;
      __tmp_1064_4 <= 0;
      __tmp_1064_5 <= 0;
      __tmp_1064_6 <= 0;
      __tmp_1064_7 <= 0;
      __tmp_1064_8 <= 0;
      __tmp_1064_9 <= 0;
      __tmp_1064_10 <= 0;
      __tmp_1066_1 <= 0;
      __tmp_1066_2 <= 0;
      __tmp_1066_3 <= 0;
      __tmp_1066_4 <= 0;
      __tmp_1066_5 <= 0;
      __tmp_1066_6 <= 0;
      __tmp_1066_7 <= 0;
      __tmp_1066_8 <= 0;
      __tmp_1066_9 <= 0;
      __tmp_1066_10 <= 0;
      __tmp_1068_1 <= 0;
      __tmp_1068_2 <= 0;
      __tmp_1068_3 <= 0;
      __tmp_1068_4 <= 0;
      __tmp_1068_5 <= 0;
      __tmp_1068_6 <= 0;
      __tmp_1068_7 <= 0;
      __tmp_1068_8 <= 0;
      __tmp_1068_9 <= 0;
      __tmp_1068_10 <= 0;
      __tmp_1070_1 <= 0;
      __tmp_1070_2 <= 0;
      __tmp_1070_3 <= 0;
      __tmp_1070_4 <= 0;
      __tmp_1070_5 <= 0;
      __tmp_1070_6 <= 0;
    end else begin
      if(__stream_seq_15_cond_2_9) begin
        _stream_max_pool_serial_18_sink_3_sink_mode <= 3'b1;
        _stream_max_pool_serial_18_sink_3_sink_offset <= __stream_max_pool_serial_18_sink_3_sink_offset_0_9;
        _stream_max_pool_serial_18_sink_3_sink_size <= __stream_max_pool_serial_18_sink_3_sink_size_1_9;
        _stream_max_pool_serial_18_sink_3_sink_stride <= 1;
      end 
      __stream_max_pool_serial_18_sink_3_sink_offset_0_9 <= __stream_max_pool_serial_18_sink_3_sink_offset_0_8;
      __stream_max_pool_serial_18_sink_3_sink_size_1_9 <= __stream_max_pool_serial_18_sink_3_sink_size_1_8;
      __stream_seq_15_cond_2_9 <= __stream_seq_15_cond_2_8;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_8 <= __stream_max_pool_serial_18_sink_3_sink_offset_0_7;
      __stream_max_pool_serial_18_sink_3_sink_size_1_8 <= __stream_max_pool_serial_18_sink_3_sink_size_1_7;
      __stream_seq_15_cond_2_8 <= __stream_seq_15_cond_2_7;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_7 <= __stream_max_pool_serial_18_sink_3_sink_offset_0_6;
      __stream_max_pool_serial_18_sink_3_sink_size_1_7 <= __stream_max_pool_serial_18_sink_3_sink_size_1_6;
      __stream_seq_15_cond_2_7 <= __stream_seq_15_cond_2_6;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_6 <= __stream_max_pool_serial_18_sink_3_sink_offset_0_5;
      __stream_max_pool_serial_18_sink_3_sink_size_1_6 <= __stream_max_pool_serial_18_sink_3_sink_size_1_5;
      __stream_seq_15_cond_2_6 <= __stream_seq_15_cond_2_5;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_5 <= __stream_max_pool_serial_18_sink_3_sink_offset_0_4;
      __stream_max_pool_serial_18_sink_3_sink_size_1_5 <= __stream_max_pool_serial_18_sink_3_sink_size_1_4;
      __stream_seq_15_cond_2_5 <= __stream_seq_15_cond_2_4;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_4 <= __stream_max_pool_serial_18_sink_3_sink_offset_0_3;
      __stream_max_pool_serial_18_sink_3_sink_size_1_4 <= __stream_max_pool_serial_18_sink_3_sink_size_1_3;
      __stream_seq_15_cond_2_4 <= __stream_seq_15_cond_2_3;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_3 <= __stream_max_pool_serial_18_sink_3_sink_offset_0_2;
      __stream_max_pool_serial_18_sink_3_sink_size_1_3 <= __stream_max_pool_serial_18_sink_3_sink_size_1_2;
      __stream_seq_15_cond_2_3 <= __stream_seq_15_cond_2_2;
      __stream_max_pool_serial_18_sink_3_sink_offset_0_2 <= __stream_max_pool_serial_18_sink_3_sink_offset_0_1;
      __stream_max_pool_serial_18_sink_3_sink_size_1_2 <= __stream_max_pool_serial_18_sink_3_sink_size_1_1;
      __stream_seq_15_cond_2_2 <= __stream_seq_15_cond_2_1;
      _stream_max_pool_serial_18_source_1_idle <= _stream_max_pool_serial_18_source_1_idle;
      _stream_max_pool_serial_18_source_1_source_ram_rvalid <= 0;
      _stream_max_pool_serial_18_sink_3_sink_wenable <= 0;
      _stream_max_pool_serial_18_sink_4_sink_wenable <= 0;
      _counter_count_782 <= (_counter_count_782 >= stream_max_pool_serial_18_constant_0_data - 2'sd1)? _counter_count_782 + 2'sd1 - stream_max_pool_serial_18_constant_0_data : _counter_count_782 + 2'sd1;
      _counter_data_782 <= _counter_count_782;
      if(_stream_max_pool_serial_18_reduce_reset) begin
        _counter_count_782 <= 1'sd0;
      end 
      if(_stream_max_pool_serial_18_reduce_reset) begin
        _counter_data_782 <= 1'sd0;
      end 
      __delay_data_1411 <= stream_max_pool_serial_18_constant_2_data;
      __delay_data_1412 <= _reinterpretcast_data_789;
      __delay_data_1414 <= stream_max_pool_serial_18_constant_0_data;
      _pointer_data_784 <= __delay_data_1411[_counter_data_782];
      __delay_data_1413 <= __delay_data_1412;
      __delay_data_1415 <= __delay_data_1414;
      _cond_data_791 <= (_pointer_data_784)? -9'sd128 : __delay_data_1413;
      __delay_data_1416 <= __delay_data_1415;
      __substreamoutput_data_793 <= _reduce_max_13_data_data;
      __substreamoutput_data_794 <= _reduce_max_13_valid_data;
      _set_flag_1024 <= 0;
      if(max_pool_serial_18_comp_fsm == 4) begin
        _set_flag_1024 <= 1;
      end 
      if(_set_flag_1024) begin
        _stream_max_pool_serial_18_constant_0_next_constant_data <= 4;
      end 
      if(_stream_max_pool_serial_18_start) begin
        __variable_wdata_777 <= _stream_max_pool_serial_18_constant_0_next_constant_data;
      end 
      _set_flag_1025 <= 0;
      if(max_pool_serial_18_comp_fsm == 4) begin
        _set_flag_1025 <= 1;
      end 
      if(_set_flag_1025) begin
        _stream_max_pool_serial_18_constant_2_next_constant_data <= max_pool_serial_18_stream_pad_masks;
      end 
      if(_stream_max_pool_serial_18_start) begin
        __variable_wdata_779 <= _stream_max_pool_serial_18_constant_2_next_constant_data;
      end 
      _set_flag_1026 <= 0;
      if(max_pool_serial_18_comp_fsm == 4) begin
        _set_flag_1026 <= 1;
      end 
      if(_set_flag_1026) begin
        _stream_max_pool_serial_18_source_1_source_mode <= 3'b10;
        _stream_max_pool_serial_18_source_1_source_offset <= max_pool_serial_18_stream_act_local + max_pool_serial_18_act_page_comp_offset_buf;
      end 
      if(_set_flag_1026) begin
        _source_stream_max_pool_serial_18_source_1_pat_size_0 <= 2;
        _source_stream_max_pool_serial_18_source_1_pat_stride_0 <= cparam_max_pool_serial_18_act_read_block;
      end 
      if(_set_flag_1026) begin
        _source_stream_max_pool_serial_18_source_1_pat_size_1 <= 2;
        _source_stream_max_pool_serial_18_source_1_pat_stride_1 <= cparam_max_pool_serial_18_act_read_size;
      end 
      if(_set_flag_1026) begin
        _source_stream_max_pool_serial_18_source_1_pat_size_2 <= cparam_max_pool_serial_18_stream_size;
        _source_stream_max_pool_serial_18_source_1_pat_stride_2 <= 1;
      end 
      if(_set_flag_1026) begin
        _source_stream_max_pool_serial_18_source_1_pat_size_3 <= 1;
        _source_stream_max_pool_serial_18_source_1_pat_stride_3 <= 0;
      end 
      if(_set_flag_1026) begin
        _stream_max_pool_serial_18_source_1_source_ram_sel <= 1;
      end 
      __tmp_1035_1 <= _tmp_1035;
      if(__tmp_1035_1) begin
        _stream_max_pool_serial_18_source_1_source_ram_rvalid <= 1;
      end 
      if(_stream_max_pool_serial_18_source_1_source_ram_rvalid) begin
        __variable_wdata_778 <= _stream_max_pool_serial_18_source_1_source_ram_rdata;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _stream_max_pool_serial_18_source_1_idle <= 0;
        _stream_max_pool_serial_18_source_1_source_offset_buf <= _stream_max_pool_serial_18_source_1_source_offset;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_cur_offset_0 <= 0;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_cur_offset_1 <= 0;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_cur_offset_2 <= 0;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_cur_offset_3 <= 0;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_count_0 <= _source_stream_max_pool_serial_18_source_1_pat_size_0 - 1;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_count_1 <= _source_stream_max_pool_serial_18_source_1_pat_size_1 - 1;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_count_2 <= _source_stream_max_pool_serial_18_source_1_pat_size_2 - 1;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_count_3 <= _source_stream_max_pool_serial_18_source_1_pat_size_3 - 1;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_size_buf_0 <= _source_stream_max_pool_serial_18_source_1_pat_size_0;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_size_buf_1 <= _source_stream_max_pool_serial_18_source_1_pat_size_1;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_size_buf_2 <= _source_stream_max_pool_serial_18_source_1_pat_size_2;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_size_buf_3 <= _source_stream_max_pool_serial_18_source_1_pat_size_3;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_stride_buf_0 <= _source_stream_max_pool_serial_18_source_1_pat_stride_0;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_stride_buf_1 <= _source_stream_max_pool_serial_18_source_1_pat_stride_1;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_stride_buf_2 <= _source_stream_max_pool_serial_18_source_1_pat_stride_2;
      end 
      if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
        _source_stream_max_pool_serial_18_source_1_pat_stride_buf_3 <= _source_stream_max_pool_serial_18_source_1_pat_stride_3;
      end 
      if(_stream_max_pool_serial_18_source_1_source_pat_fsm_0 == 1) begin
        _stream_max_pool_serial_18_source_1_source_ram_raddr <= _stream_max_pool_serial_18_source_1_source_pat_all_offset;
        _stream_max_pool_serial_18_source_1_source_ram_renable <= 1;
      end 
      if(_stream_max_pool_serial_18_source_1_source_pat_fsm_0 == 1) begin
        _source_stream_max_pool_serial_18_source_1_pat_cur_offset_0 <= _source_stream_max_pool_serial_18_source_1_pat_cur_offset_0 + _source_stream_max_pool_serial_18_source_1_pat_stride_buf_0;
        _source_stream_max_pool_serial_18_source_1_pat_count_0 <= _source_stream_max_pool_serial_18_source_1_pat_count_0 - 1;
      end 
      if((_stream_max_pool_serial_18_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_18_source_1_pat_count_0 == 0)) begin
        _source_stream_max_pool_serial_18_source_1_pat_cur_offset_0 <= 0;
        _source_stream_max_pool_serial_18_source_1_pat_count_0 <= _source_stream_max_pool_serial_18_source_1_pat_size_buf_0 - 1;
      end 
      if((_stream_max_pool_serial_18_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_18_source_1_pat_count_0 == 0)) begin
        _source_stream_max_pool_serial_18_source_1_pat_cur_offset_1 <= _source_stream_max_pool_serial_18_source_1_pat_cur_offset_1 + _source_stream_max_pool_serial_18_source_1_pat_stride_buf_1;
        _source_stream_max_pool_serial_18_source_1_pat_count_1 <= _source_stream_max_pool_serial_18_source_1_pat_count_1 - 1;
      end 
      if((_stream_max_pool_serial_18_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_18_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_18_source_1_pat_count_1 == 0)) begin
        _source_stream_max_pool_serial_18_source_1_pat_cur_offset_1 <= 0;
        _source_stream_max_pool_serial_18_source_1_pat_count_1 <= _source_stream_max_pool_serial_18_source_1_pat_size_buf_1 - 1;
      end 
      if((_stream_max_pool_serial_18_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_18_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_18_source_1_pat_count_1 == 0))) begin
        _source_stream_max_pool_serial_18_source_1_pat_cur_offset_2 <= _source_stream_max_pool_serial_18_source_1_pat_cur_offset_2 + _source_stream_max_pool_serial_18_source_1_pat_stride_buf_2;
        _source_stream_max_pool_serial_18_source_1_pat_count_2 <= _source_stream_max_pool_serial_18_source_1_pat_count_2 - 1;
      end 
      if((_stream_max_pool_serial_18_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_18_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_18_source_1_pat_count_1 == 0)) && (_source_stream_max_pool_serial_18_source_1_pat_count_2 == 0)) begin
        _source_stream_max_pool_serial_18_source_1_pat_cur_offset_2 <= 0;
        _source_stream_max_pool_serial_18_source_1_pat_count_2 <= _source_stream_max_pool_serial_18_source_1_pat_size_buf_2 - 1;
      end 
      if((_stream_max_pool_serial_18_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_18_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_18_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_18_source_1_pat_count_2 == 0))) begin
        _source_stream_max_pool_serial_18_source_1_pat_cur_offset_3 <= _source_stream_max_pool_serial_18_source_1_pat_cur_offset_3 + _source_stream_max_pool_serial_18_source_1_pat_stride_buf_3;
        _source_stream_max_pool_serial_18_source_1_pat_count_3 <= _source_stream_max_pool_serial_18_source_1_pat_count_3 - 1;
      end 
      if((_stream_max_pool_serial_18_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_18_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_18_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_18_source_1_pat_count_2 == 0)) && (_source_stream_max_pool_serial_18_source_1_pat_count_3 == 0)) begin
        _source_stream_max_pool_serial_18_source_1_pat_cur_offset_3 <= 0;
        _source_stream_max_pool_serial_18_source_1_pat_count_3 <= _source_stream_max_pool_serial_18_source_1_pat_size_buf_3 - 1;
      end 
      if(_stream_max_pool_serial_18_source_1_source_pat_fsm_0 == 2) begin
        _stream_max_pool_serial_18_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_18_source_1_idle <= 1;
      end 
      _set_flag_1036 <= 0;
      if(max_pool_serial_18_comp_fsm == 4) begin
        _set_flag_1036 <= 1;
      end 
      __stream_max_pool_serial_18_sink_3_sink_offset_0_1 <= max_pool_serial_18_stream_out_local + max_pool_serial_18_out_page_comp_offset_buf;
      __stream_max_pool_serial_18_sink_3_sink_size_1_1 <= cparam_max_pool_serial_18_stream_size;
      __stream_seq_15_cond_2_1 <= _set_flag_1036;
      __set_flag_1036_1 <= _set_flag_1036;
      __set_flag_1036_2 <= __set_flag_1036_1;
      __set_flag_1036_3 <= __set_flag_1036_2;
      __set_flag_1036_4 <= __set_flag_1036_3;
      __set_flag_1036_5 <= __set_flag_1036_4;
      __set_flag_1036_6 <= __set_flag_1036_5;
      __set_flag_1036_7 <= __set_flag_1036_6;
      __set_flag_1036_8 <= __set_flag_1036_7;
      __set_flag_1036_9 <= __set_flag_1036_8;
      if(__set_flag_1036_9) begin
        _stream_max_pool_serial_18_sink_3_sink_ram_sel <= 2;
      end 
      __stream_max_pool_serial_18_start_1 <= _stream_max_pool_serial_18_start;
      __stream_max_pool_serial_18_start_2 <= __stream_max_pool_serial_18_start_1;
      __stream_max_pool_serial_18_start_3 <= __stream_max_pool_serial_18_start_2;
      __stream_max_pool_serial_18_start_4 <= __stream_max_pool_serial_18_start_3;
      __stream_max_pool_serial_18_start_5 <= __stream_max_pool_serial_18_start_4;
      __stream_max_pool_serial_18_start_6 <= __stream_max_pool_serial_18_start_5;
      __stream_max_pool_serial_18_start_7 <= __stream_max_pool_serial_18_start_6;
      __stream_max_pool_serial_18_start_8 <= __stream_max_pool_serial_18_start_7;
      __stream_max_pool_serial_18_start_9 <= __stream_max_pool_serial_18_start_8;
      __stream_max_pool_serial_18_start_10 <= __stream_max_pool_serial_18_start_9;
      if(__stream_max_pool_serial_18_start_10 && _stream_max_pool_serial_18_sink_3_sink_mode & 3'b1) begin
        _stream_max_pool_serial_18_sink_3_sink_waddr <= _stream_max_pool_serial_18_sink_3_sink_offset - _stream_max_pool_serial_18_sink_3_sink_stride;
        _stream_max_pool_serial_18_sink_3_sink_count <= _stream_max_pool_serial_18_sink_3_sink_size;
        _stream_max_pool_serial_18_sink_3_sink_offset_buf <= _stream_max_pool_serial_18_sink_3_sink_offset;
        _stream_max_pool_serial_18_sink_3_sink_stride_buf <= _stream_max_pool_serial_18_sink_3_sink_stride;
      end 
      if((_stream_max_pool_serial_18_sink_3_sink_fsm_1 == 1) && stream_max_pool_serial_18_sink_4_data) begin
        _stream_max_pool_serial_18_sink_3_sink_waddr <= _stream_max_pool_serial_18_sink_3_sink_waddr + _stream_max_pool_serial_18_sink_3_sink_stride_buf;
        _stream_max_pool_serial_18_sink_3_sink_wdata <= stream_max_pool_serial_18_sink_3_data;
        _stream_max_pool_serial_18_sink_3_sink_wenable <= 1;
        _stream_max_pool_serial_18_sink_3_sink_count <= _stream_max_pool_serial_18_sink_3_sink_count - 1;
      end 
      _set_flag_1038 <= 0;
      if(max_pool_serial_18_comp_fsm == 5) begin
        _set_flag_1038 <= 1;
      end 
      __tmp_1040_1 <= _tmp_1040;
      __tmp_1040_2 <= __tmp_1040_1;
      __tmp_1040_3 <= __tmp_1040_2;
      __tmp_1040_4 <= __tmp_1040_3;
      __tmp_1040_5 <= __tmp_1040_4;
      __tmp_1042_1 <= _tmp_1042;
      __tmp_1042_2 <= __tmp_1042_1;
      __tmp_1042_3 <= __tmp_1042_2;
      __tmp_1042_4 <= __tmp_1042_3;
      __tmp_1042_5 <= __tmp_1042_4;
      __tmp_1042_6 <= __tmp_1042_5;
      __tmp_1042_7 <= __tmp_1042_6;
      __tmp_1042_8 <= __tmp_1042_7;
      __tmp_1042_9 <= __tmp_1042_8;
      __tmp_1044_1 <= _tmp_1044;
      __tmp_1044_2 <= __tmp_1044_1;
      __tmp_1044_3 <= __tmp_1044_2;
      __tmp_1044_4 <= __tmp_1044_3;
      __tmp_1044_5 <= __tmp_1044_4;
      __tmp_1044_6 <= __tmp_1044_5;
      __tmp_1044_7 <= __tmp_1044_6;
      __tmp_1046_1 <= _tmp_1046;
      __tmp_1046_2 <= __tmp_1046_1;
      __tmp_1046_3 <= __tmp_1046_2;
      __tmp_1046_4 <= __tmp_1046_3;
      __tmp_1046_5 <= __tmp_1046_4;
      __tmp_1046_6 <= __tmp_1046_5;
      __tmp_1046_7 <= __tmp_1046_6;
      __tmp_1048_1 <= _tmp_1048;
      __tmp_1050_1 <= _tmp_1050;
      __tmp_1050_2 <= __tmp_1050_1;
      __tmp_1050_3 <= __tmp_1050_2;
      __tmp_1050_4 <= __tmp_1050_3;
      __tmp_1050_5 <= __tmp_1050_4;
      __tmp_1052_1 <= _tmp_1052;
      __tmp_1052_2 <= __tmp_1052_1;
      __tmp_1052_3 <= __tmp_1052_2;
      __tmp_1052_4 <= __tmp_1052_3;
      __tmp_1054_1 <= _tmp_1054;
      __tmp_1054_2 <= __tmp_1054_1;
      __tmp_1054_3 <= __tmp_1054_2;
      __tmp_1054_4 <= __tmp_1054_3;
      __tmp_1062_1 <= _tmp_1062;
      __tmp_1062_2 <= __tmp_1062_1;
      __tmp_1062_3 <= __tmp_1062_2;
      __tmp_1062_4 <= __tmp_1062_3;
      __tmp_1062_5 <= __tmp_1062_4;
      __tmp_1062_6 <= __tmp_1062_5;
      __tmp_1062_7 <= __tmp_1062_6;
      __tmp_1062_8 <= __tmp_1062_7;
      __tmp_1062_9 <= __tmp_1062_8;
      __tmp_1062_10 <= __tmp_1062_9;
      __tmp_1064_1 <= _tmp_1064;
      __tmp_1064_2 <= __tmp_1064_1;
      __tmp_1064_3 <= __tmp_1064_2;
      __tmp_1064_4 <= __tmp_1064_3;
      __tmp_1064_5 <= __tmp_1064_4;
      __tmp_1064_6 <= __tmp_1064_5;
      __tmp_1064_7 <= __tmp_1064_6;
      __tmp_1064_8 <= __tmp_1064_7;
      __tmp_1064_9 <= __tmp_1064_8;
      __tmp_1064_10 <= __tmp_1064_9;
      __tmp_1066_1 <= _tmp_1066;
      __tmp_1066_2 <= __tmp_1066_1;
      __tmp_1066_3 <= __tmp_1066_2;
      __tmp_1066_4 <= __tmp_1066_3;
      __tmp_1066_5 <= __tmp_1066_4;
      __tmp_1066_6 <= __tmp_1066_5;
      __tmp_1066_7 <= __tmp_1066_6;
      __tmp_1066_8 <= __tmp_1066_7;
      __tmp_1066_9 <= __tmp_1066_8;
      __tmp_1066_10 <= __tmp_1066_9;
      __tmp_1068_1 <= _tmp_1068;
      __tmp_1068_2 <= __tmp_1068_1;
      __tmp_1068_3 <= __tmp_1068_2;
      __tmp_1068_4 <= __tmp_1068_3;
      __tmp_1068_5 <= __tmp_1068_4;
      __tmp_1068_6 <= __tmp_1068_5;
      __tmp_1068_7 <= __tmp_1068_6;
      __tmp_1068_8 <= __tmp_1068_7;
      __tmp_1068_9 <= __tmp_1068_8;
      __tmp_1068_10 <= __tmp_1068_9;
      __tmp_1070_1 <= _tmp_1070;
      __tmp_1070_2 <= __tmp_1070_1;
      __tmp_1070_3 <= __tmp_1070_2;
      __tmp_1070_4 <= __tmp_1070_3;
      __tmp_1070_5 <= __tmp_1070_4;
      __tmp_1070_6 <= __tmp_1070_5;
    end
  end

  localparam _stream_max_pool_serial_18_fsm_1 = 1;
  localparam _stream_max_pool_serial_18_fsm_2 = 2;
  localparam _stream_max_pool_serial_18_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_18_fsm <= _stream_max_pool_serial_18_fsm_init;
      _stream_max_pool_serial_18_start <= 0;
      _stream_max_pool_serial_18_source_busy <= 0;
      _stream_max_pool_serial_18_reduce_reset <= 1;
      _stream_max_pool_serial_18_sink_busy <= 0;
      _stream_max_pool_serial_18_sink_wait_count <= 0;
      _stream_max_pool_serial_18_end_flag <= 0;
      _stream_max_pool_serial_18_term_sink <= 0;
    end else begin
      _stream_max_pool_serial_18_start <= 0;
      if(__tmp_1040_5) begin
        _stream_max_pool_serial_18_reduce_reset <= 0;
      end 
      if(__tmp_1048_1) begin
        _stream_max_pool_serial_18_reduce_reset <= 1;
      end 
      if((_stream_max_pool_serial_18_sink_wait_count == 1) && !((_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag) && __tmp_1062_10) begin
        _stream_max_pool_serial_18_sink_busy <= 0;
      end 
      if((_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag) begin
        _stream_max_pool_serial_18_sink_busy <= 1;
      end 
      if(!((_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag) && __tmp_1064_10) begin
        _stream_max_pool_serial_18_sink_wait_count <= _stream_max_pool_serial_18_sink_wait_count - 1;
      end 
      if((_stream_max_pool_serial_18_fsm == 0) && _stream_max_pool_serial_18_start_flag && !__tmp_1066_10) begin
        _stream_max_pool_serial_18_sink_wait_count <= _stream_max_pool_serial_18_sink_wait_count + 1;
      end 
      _stream_max_pool_serial_18_end_flag <= 0;
      if(__tmp_1068_10) begin
        _stream_max_pool_serial_18_end_flag <= 1;
      end 
      _stream_max_pool_serial_18_term_sink <= 0;
      if(__tmp_1070_6) begin
        _stream_max_pool_serial_18_term_sink <= 1;
      end 
      case(_stream_max_pool_serial_18_fsm)
        _stream_max_pool_serial_18_fsm_init: begin
          if(_stream_max_pool_serial_18_start_flag) begin
            _stream_max_pool_serial_18_start <= 1;
            _stream_max_pool_serial_18_source_busy <= 1;
          end 
          if(_stream_max_pool_serial_18_start_flag) begin
            _stream_max_pool_serial_18_fsm <= _stream_max_pool_serial_18_fsm_1;
          end 
        end
        _stream_max_pool_serial_18_fsm_1: begin
          _stream_max_pool_serial_18_fsm <= _stream_max_pool_serial_18_fsm_2;
        end
        _stream_max_pool_serial_18_fsm_2: begin
          if(_stream_max_pool_serial_18_done) begin
            _stream_max_pool_serial_18_fsm <= _stream_max_pool_serial_18_fsm_3;
          end 
        end
        _stream_max_pool_serial_18_fsm_3: begin
          _stream_max_pool_serial_18_source_busy <= 0;
          _stream_max_pool_serial_18_fsm <= _stream_max_pool_serial_18_fsm_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_29_source_6_idle <= 1;
      _stream_matmul_29_source_6_source_ram_rvalid <= 0;
      _stream_matmul_29_source_8_idle <= 1;
      _stream_matmul_29_source_8_source_ram_rvalid <= 0;
      _stream_matmul_29_source_10_idle <= 1;
      _stream_matmul_29_source_10_source_ram_rvalid <= 0;
      _stream_matmul_29_source_12_idle <= 1;
      _stream_matmul_29_source_12_source_ram_rvalid <= 0;
      _stream_matmul_29_source_14_idle <= 1;
      _stream_matmul_29_source_14_source_ram_rvalid <= 0;
      _stream_matmul_29_source_19_idle <= 1;
      _stream_matmul_29_source_19_source_ram_rvalid <= 0;
      _stream_matmul_29_source_20_idle <= 1;
      _stream_matmul_29_source_20_source_ram_rvalid <= 0;
      _stream_matmul_29_sink_21_sink_wenable <= 0;
      _stream_matmul_29_sink_22_sink_wenable <= 0;
      _cond_data_817 <= 0;
      _cond_data_824 <= 0;
      _cond_data_831 <= 0;
      _cond_data_838 <= 0;
      _cond_data_845 <= 0;
      _eq_data_851 <= 0;
      _eq_data_855 <= 0;
      _eq_data_891 <= 0;
      _eq_data_894 <= 0;
      __delay_data_1417 <= 0;
      __delay_data_1419 <= 0;
      __delay_data_1422 <= 0;
      __delay_data_1423 <= 0;
      __delay_data_1429 <= 0;
      __delay_data_1444 <= 0;
      __delay_data_1482 <= 0;
      _cond_data_853 <= 0;
      _plus_data_875 <= 0;
      _plus_data_880 <= 0;
      _plus_data_885 <= 0;
      __delay_data_1418 <= 0;
      __delay_data_1420 <= 0;
      __delay_data_1424 <= 0;
      __delay_data_1445 <= 0;
      __delay_data_1460 <= 0;
      __delay_data_1483 <= 0;
      __delay_data_1529 <= 0;
      __delay_data_1565 <= 0;
      _cond_data_857 <= 0;
      __delay_data_1421 <= 0;
      __delay_data_1425 <= 0;
      __delay_data_1427 <= 0;
      __delay_data_1430 <= 0;
      __delay_data_1446 <= 0;
      __delay_data_1461 <= 0;
      __delay_data_1484 <= 0;
      __delay_data_1506 <= 0;
      __delay_data_1530 <= 0;
      __delay_data_1566 <= 0;
      _cond_data_873 <= 0;
      __delay_data_1426 <= 0;
      __delay_data_1428 <= 0;
      __delay_data_1431 <= 0;
      __delay_data_1447 <= 0;
      __delay_data_1462 <= 0;
      __delay_data_1485 <= 0;
      __delay_data_1507 <= 0;
      __delay_data_1531 <= 0;
      __delay_data_1567 <= 0;
      __delay_data_1432 <= 0;
      __delay_data_1448 <= 0;
      __delay_data_1463 <= 0;
      __delay_data_1486 <= 0;
      __delay_data_1508 <= 0;
      __delay_data_1532 <= 0;
      __delay_data_1568 <= 0;
      __delay_data_1433 <= 0;
      __delay_data_1449 <= 0;
      __delay_data_1464 <= 0;
      __delay_data_1487 <= 0;
      __delay_data_1509 <= 0;
      __delay_data_1533 <= 0;
      __delay_data_1569 <= 0;
      __delay_data_1434 <= 0;
      __delay_data_1450 <= 0;
      __delay_data_1465 <= 0;
      __delay_data_1488 <= 0;
      __delay_data_1510 <= 0;
      __delay_data_1534 <= 0;
      __delay_data_1570 <= 0;
      __delay_data_1435 <= 0;
      __delay_data_1451 <= 0;
      __delay_data_1466 <= 0;
      __delay_data_1489 <= 0;
      __delay_data_1511 <= 0;
      __delay_data_1535 <= 0;
      __delay_data_1571 <= 0;
      __delay_data_1436 <= 0;
      __delay_data_1452 <= 0;
      __delay_data_1467 <= 0;
      __delay_data_1490 <= 0;
      __delay_data_1512 <= 0;
      __delay_data_1536 <= 0;
      __delay_data_1572 <= 0;
      __delay_data_1437 <= 0;
      __delay_data_1453 <= 0;
      __delay_data_1468 <= 0;
      __delay_data_1491 <= 0;
      __delay_data_1513 <= 0;
      __delay_data_1537 <= 0;
      __delay_data_1573 <= 0;
      __delay_data_1438 <= 0;
      __delay_data_1454 <= 0;
      __delay_data_1469 <= 0;
      __delay_data_1492 <= 0;
      __delay_data_1514 <= 0;
      __delay_data_1538 <= 0;
      __delay_data_1574 <= 0;
      __delay_data_1439 <= 0;
      __delay_data_1455 <= 0;
      __delay_data_1470 <= 0;
      __delay_data_1493 <= 0;
      __delay_data_1515 <= 0;
      __delay_data_1539 <= 0;
      __delay_data_1575 <= 0;
      __delay_data_1440 <= 0;
      __delay_data_1456 <= 0;
      __delay_data_1471 <= 0;
      __delay_data_1494 <= 0;
      __delay_data_1516 <= 0;
      __delay_data_1540 <= 0;
      __delay_data_1576 <= 0;
      __substreamoutput_data_876 <= 0;
      __delay_data_1441 <= 0;
      __delay_data_1457 <= 0;
      __delay_data_1472 <= 0;
      __delay_data_1495 <= 0;
      __delay_data_1517 <= 0;
      __delay_data_1541 <= 0;
      __delay_data_1577 <= 0;
      __delay_data_1442 <= 0;
      __delay_data_1458 <= 0;
      __delay_data_1473 <= 0;
      __delay_data_1496 <= 0;
      __delay_data_1518 <= 0;
      __delay_data_1542 <= 0;
      __delay_data_1578 <= 0;
      __substreamoutput_data_878 <= 0;
      __delay_data_1443 <= 0;
      __delay_data_1459 <= 0;
      __delay_data_1474 <= 0;
      __delay_data_1497 <= 0;
      __delay_data_1519 <= 0;
      __delay_data_1543 <= 0;
      __delay_data_1579 <= 0;
      __delay_data_1475 <= 0;
      __delay_data_1498 <= 0;
      __delay_data_1520 <= 0;
      __delay_data_1544 <= 0;
      __delay_data_1580 <= 0;
      __delay_data_1476 <= 0;
      __delay_data_1499 <= 0;
      __delay_data_1521 <= 0;
      __delay_data_1545 <= 0;
      __delay_data_1581 <= 0;
      __delay_data_1477 <= 0;
      __delay_data_1500 <= 0;
      __delay_data_1522 <= 0;
      __delay_data_1546 <= 0;
      __delay_data_1582 <= 0;
      __delay_data_1478 <= 0;
      __delay_data_1501 <= 0;
      __delay_data_1523 <= 0;
      __delay_data_1547 <= 0;
      __delay_data_1583 <= 0;
      __delay_data_1479 <= 0;
      __delay_data_1502 <= 0;
      __delay_data_1524 <= 0;
      __delay_data_1548 <= 0;
      __delay_data_1584 <= 0;
      __delay_data_1480 <= 0;
      __delay_data_1503 <= 0;
      __delay_data_1525 <= 0;
      __delay_data_1549 <= 0;
      __delay_data_1585 <= 0;
      __substreamoutput_data_881 <= 0;
      __substreamoutput_data_882 <= 0;
      __delay_data_1481 <= 0;
      __delay_data_1504 <= 0;
      __delay_data_1526 <= 0;
      __delay_data_1550 <= 0;
      __delay_data_1586 <= 0;
      _plus_data_883 <= 0;
      __delay_data_1505 <= 0;
      __delay_data_1527 <= 0;
      __delay_data_1551 <= 0;
      __delay_data_1587 <= 0;
      __delay_data_1602 <= 0;
      __delay_data_1552 <= 0;
      __delay_data_1588 <= 0;
      __delay_data_1603 <= 0;
      __delay_data_1553 <= 0;
      __delay_data_1589 <= 0;
      __delay_data_1604 <= 0;
      __delay_data_1554 <= 0;
      __delay_data_1590 <= 0;
      __delay_data_1605 <= 0;
      __delay_data_1555 <= 0;
      __delay_data_1591 <= 0;
      __delay_data_1606 <= 0;
      __delay_data_1556 <= 0;
      __delay_data_1592 <= 0;
      __delay_data_1607 <= 0;
      __delay_data_1557 <= 0;
      __delay_data_1593 <= 0;
      __delay_data_1608 <= 0;
      __delay_data_1558 <= 0;
      __delay_data_1594 <= 0;
      __delay_data_1609 <= 0;
      __delay_data_1559 <= 0;
      __delay_data_1595 <= 0;
      __delay_data_1610 <= 0;
      __delay_data_1560 <= 0;
      __delay_data_1596 <= 0;
      __delay_data_1611 <= 0;
      __substreamoutput_data_886 <= 0;
      __delay_data_1561 <= 0;
      __delay_data_1597 <= 0;
      __delay_data_1612 <= 0;
      _greaterthan_data_888 <= 0;
      __delay_data_1528 <= 0;
      __delay_data_1562 <= 0;
      __delay_data_1598 <= 0;
      __delay_data_1613 <= 0;
      _cond_data_890 <= 0;
      __delay_data_1563 <= 0;
      __delay_data_1564 <= 0;
      __delay_data_1599 <= 0;
      __delay_data_1614 <= 0;
      _cond_data_893 <= 0;
      __delay_data_1600 <= 0;
      __delay_data_1601 <= 0;
      __delay_data_1615 <= 0;
      _cond_data_896 <= 0;
      __delay_data_1616 <= 0;
      _set_flag_1163 <= 0;
      _stream_matmul_29_constant_0_next_constant_data <= 0;
      __variable_wdata_796 <= 0;
      _set_flag_1164 <= 0;
      _stream_matmul_29_constant_1_next_constant_data <= 0;
      __variable_wdata_797 <= 0;
      _set_flag_1165 <= 0;
      _stream_matmul_29_constant_2_next_constant_data <= 0;
      __variable_wdata_798 <= 0;
      _set_flag_1166 <= 0;
      _stream_matmul_29_constant_3_next_constant_data <= 0;
      __variable_wdata_799 <= 0;
      _set_flag_1167 <= 0;
      _stream_matmul_29_constant_4_next_constant_data <= 0;
      __variable_wdata_800 <= 0;
      _set_flag_1168 <= 0;
      _stream_matmul_29_constant_5_next_constant_data <= 0;
      __variable_wdata_811 <= 0;
      _set_flag_1169 <= 0;
      _stream_matmul_29_source_6_source_mode <= 3'b0;
      _stream_matmul_29_source_6_source_offset <= 0;
      _source_stream_matmul_29_source_6_pat_size_0 <= 0;
      _source_stream_matmul_29_source_6_pat_stride_0 <= 0;
      _source_stream_matmul_29_source_6_pat_size_1 <= 0;
      _source_stream_matmul_29_source_6_pat_stride_1 <= 0;
      _source_stream_matmul_29_source_6_pat_size_2 <= 0;
      _source_stream_matmul_29_source_6_pat_stride_2 <= 0;
      _source_stream_matmul_29_source_6_pat_size_3 <= 0;
      _source_stream_matmul_29_source_6_pat_stride_3 <= 0;
      _stream_matmul_29_source_6_source_ram_sel <= 0;
      __tmp_1178_1 <= 0;
      __variable_wdata_812 <= 0;
      _stream_matmul_29_source_6_source_offset_buf <= 0;
      _source_stream_matmul_29_source_6_pat_cur_offset_0 <= 0;
      _source_stream_matmul_29_source_6_pat_cur_offset_1 <= 0;
      _source_stream_matmul_29_source_6_pat_cur_offset_2 <= 0;
      _source_stream_matmul_29_source_6_pat_cur_offset_3 <= 0;
      _source_stream_matmul_29_source_6_pat_count_0 <= 0;
      _source_stream_matmul_29_source_6_pat_count_1 <= 0;
      _source_stream_matmul_29_source_6_pat_count_2 <= 0;
      _source_stream_matmul_29_source_6_pat_count_3 <= 0;
      _source_stream_matmul_29_source_6_pat_size_buf_0 <= 0;
      _source_stream_matmul_29_source_6_pat_size_buf_1 <= 0;
      _source_stream_matmul_29_source_6_pat_size_buf_2 <= 0;
      _source_stream_matmul_29_source_6_pat_size_buf_3 <= 0;
      _source_stream_matmul_29_source_6_pat_stride_buf_0 <= 0;
      _source_stream_matmul_29_source_6_pat_stride_buf_1 <= 0;
      _source_stream_matmul_29_source_6_pat_stride_buf_2 <= 0;
      _source_stream_matmul_29_source_6_pat_stride_buf_3 <= 0;
      _stream_matmul_29_source_6_source_ram_raddr <= 0;
      _stream_matmul_29_source_6_source_ram_renable <= 0;
      _set_flag_1179 <= 0;
      _stream_matmul_29_constant_7_next_constant_data <= 0;
      __variable_wdata_818 <= 0;
      _set_flag_1180 <= 0;
      _stream_matmul_29_source_8_source_mode <= 3'b0;
      _stream_matmul_29_source_8_source_offset <= 0;
      _source_stream_matmul_29_source_8_pat_size_0 <= 0;
      _source_stream_matmul_29_source_8_pat_stride_0 <= 0;
      _source_stream_matmul_29_source_8_pat_size_1 <= 0;
      _source_stream_matmul_29_source_8_pat_stride_1 <= 0;
      _source_stream_matmul_29_source_8_pat_size_2 <= 0;
      _source_stream_matmul_29_source_8_pat_stride_2 <= 0;
      _source_stream_matmul_29_source_8_pat_size_3 <= 0;
      _source_stream_matmul_29_source_8_pat_stride_3 <= 0;
      _stream_matmul_29_source_8_source_ram_sel <= 0;
      __tmp_1189_1 <= 0;
      __variable_wdata_819 <= 0;
      _stream_matmul_29_source_8_source_offset_buf <= 0;
      _source_stream_matmul_29_source_8_pat_cur_offset_0 <= 0;
      _source_stream_matmul_29_source_8_pat_cur_offset_1 <= 0;
      _source_stream_matmul_29_source_8_pat_cur_offset_2 <= 0;
      _source_stream_matmul_29_source_8_pat_cur_offset_3 <= 0;
      _source_stream_matmul_29_source_8_pat_count_0 <= 0;
      _source_stream_matmul_29_source_8_pat_count_1 <= 0;
      _source_stream_matmul_29_source_8_pat_count_2 <= 0;
      _source_stream_matmul_29_source_8_pat_count_3 <= 0;
      _source_stream_matmul_29_source_8_pat_size_buf_0 <= 0;
      _source_stream_matmul_29_source_8_pat_size_buf_1 <= 0;
      _source_stream_matmul_29_source_8_pat_size_buf_2 <= 0;
      _source_stream_matmul_29_source_8_pat_size_buf_3 <= 0;
      _source_stream_matmul_29_source_8_pat_stride_buf_0 <= 0;
      _source_stream_matmul_29_source_8_pat_stride_buf_1 <= 0;
      _source_stream_matmul_29_source_8_pat_stride_buf_2 <= 0;
      _source_stream_matmul_29_source_8_pat_stride_buf_3 <= 0;
      _stream_matmul_29_source_8_source_ram_raddr <= 0;
      _stream_matmul_29_source_8_source_ram_renable <= 0;
      _set_flag_1190 <= 0;
      _stream_matmul_29_constant_9_next_constant_data <= 0;
      __variable_wdata_825 <= 0;
      _set_flag_1191 <= 0;
      _stream_matmul_29_source_10_source_mode <= 3'b0;
      _stream_matmul_29_source_10_source_empty_data <= 0;
      __variable_wdata_826 <= 0;
      _set_flag_1192 <= 0;
      _stream_matmul_29_constant_11_next_constant_data <= 0;
      __variable_wdata_832 <= 0;
      _set_flag_1193 <= 0;
      _stream_matmul_29_source_12_source_mode <= 3'b0;
      _stream_matmul_29_source_12_source_empty_data <= 0;
      __variable_wdata_833 <= 0;
      _set_flag_1194 <= 0;
      _stream_matmul_29_constant_13_next_constant_data <= 0;
      __variable_wdata_839 <= 0;
      _set_flag_1195 <= 0;
      _stream_matmul_29_source_14_source_mode <= 3'b0;
      _stream_matmul_29_source_14_source_empty_data <= 0;
      __variable_wdata_840 <= 0;
      _set_flag_1196 <= 0;
      _stream_matmul_29_constant_15_next_constant_data <= 0;
      __variable_wdata_846 <= 0;
      _set_flag_1197 <= 0;
      _stream_matmul_29_constant_16_next_constant_data <= 0;
      __variable_wdata_847 <= 0;
      _set_flag_1198 <= 0;
      _stream_matmul_29_constant_17_next_constant_data <= 0;
      __variable_wdata_848 <= 0;
      _set_flag_1199 <= 0;
      _stream_matmul_29_constant_18_next_constant_data <= 0;
      __variable_wdata_849 <= 0;
      _set_flag_1200 <= 0;
      _stream_matmul_29_source_19_source_mode <= 3'b0;
      _stream_matmul_29_source_19_source_offset <= 0;
      _source_stream_matmul_29_source_19_pat_size_0 <= 0;
      _source_stream_matmul_29_source_19_pat_stride_0 <= 0;
      _source_stream_matmul_29_source_19_pat_size_1 <= 0;
      _source_stream_matmul_29_source_19_pat_stride_1 <= 0;
      _source_stream_matmul_29_source_19_pat_size_2 <= 0;
      _source_stream_matmul_29_source_19_pat_stride_2 <= 0;
      _source_stream_matmul_29_source_19_pat_size_3 <= 0;
      _source_stream_matmul_29_source_19_pat_stride_3 <= 0;
      _stream_matmul_29_source_19_source_ram_sel <= 0;
      __tmp_1209_1 <= 0;
      __variable_wdata_850 <= 0;
      _stream_matmul_29_source_19_source_offset_buf <= 0;
      _source_stream_matmul_29_source_19_pat_cur_offset_0 <= 0;
      _source_stream_matmul_29_source_19_pat_cur_offset_1 <= 0;
      _source_stream_matmul_29_source_19_pat_cur_offset_2 <= 0;
      _source_stream_matmul_29_source_19_pat_cur_offset_3 <= 0;
      _source_stream_matmul_29_source_19_pat_count_0 <= 0;
      _source_stream_matmul_29_source_19_pat_count_1 <= 0;
      _source_stream_matmul_29_source_19_pat_count_2 <= 0;
      _source_stream_matmul_29_source_19_pat_count_3 <= 0;
      _source_stream_matmul_29_source_19_pat_size_buf_0 <= 0;
      _source_stream_matmul_29_source_19_pat_size_buf_1 <= 0;
      _source_stream_matmul_29_source_19_pat_size_buf_2 <= 0;
      _source_stream_matmul_29_source_19_pat_size_buf_3 <= 0;
      _source_stream_matmul_29_source_19_pat_stride_buf_0 <= 0;
      _source_stream_matmul_29_source_19_pat_stride_buf_1 <= 0;
      _source_stream_matmul_29_source_19_pat_stride_buf_2 <= 0;
      _source_stream_matmul_29_source_19_pat_stride_buf_3 <= 0;
      _stream_matmul_29_source_19_source_ram_raddr <= 0;
      _stream_matmul_29_source_19_source_ram_renable <= 0;
      _set_flag_1210 <= 0;
      _stream_matmul_29_source_20_source_mode <= 3'b0;
      _stream_matmul_29_source_20_source_offset <= 0;
      _source_stream_matmul_29_source_20_pat_size_0 <= 0;
      _source_stream_matmul_29_source_20_pat_stride_0 <= 0;
      _source_stream_matmul_29_source_20_pat_size_1 <= 0;
      _source_stream_matmul_29_source_20_pat_stride_1 <= 0;
      _source_stream_matmul_29_source_20_pat_size_2 <= 0;
      _source_stream_matmul_29_source_20_pat_stride_2 <= 0;
      _source_stream_matmul_29_source_20_pat_size_3 <= 0;
      _source_stream_matmul_29_source_20_pat_stride_3 <= 0;
      _stream_matmul_29_source_20_source_ram_sel <= 0;
      __tmp_1223_1 <= 0;
      __variable_wdata_864 <= 0;
      _stream_matmul_29_source_20_source_offset_buf <= 0;
      _source_stream_matmul_29_source_20_pat_cur_offset_0 <= 0;
      _source_stream_matmul_29_source_20_pat_cur_offset_1 <= 0;
      _source_stream_matmul_29_source_20_pat_cur_offset_2 <= 0;
      _source_stream_matmul_29_source_20_pat_cur_offset_3 <= 0;
      _source_stream_matmul_29_source_20_pat_count_0 <= 0;
      _source_stream_matmul_29_source_20_pat_count_1 <= 0;
      _source_stream_matmul_29_source_20_pat_count_2 <= 0;
      _source_stream_matmul_29_source_20_pat_count_3 <= 0;
      _source_stream_matmul_29_source_20_pat_size_buf_0 <= 0;
      _source_stream_matmul_29_source_20_pat_size_buf_1 <= 0;
      _source_stream_matmul_29_source_20_pat_size_buf_2 <= 0;
      _source_stream_matmul_29_source_20_pat_size_buf_3 <= 0;
      _source_stream_matmul_29_source_20_pat_stride_buf_0 <= 0;
      _source_stream_matmul_29_source_20_pat_stride_buf_1 <= 0;
      _source_stream_matmul_29_source_20_pat_stride_buf_2 <= 0;
      _source_stream_matmul_29_source_20_pat_stride_buf_3 <= 0;
      _stream_matmul_29_source_20_source_ram_raddr <= 0;
      _stream_matmul_29_source_20_source_ram_renable <= 0;
      _set_flag_1224 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_1 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_2 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_3 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_4 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_5 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_6 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_7 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_8 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_9 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_10 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_11 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_12 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_13 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_14 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_15 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_16 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_17 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_18 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_19 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_20 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_21 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_22 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_23 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_24 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_25 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_26 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_27 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_28 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_29 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_30 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_31 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_32 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_33 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_34 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_35 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_36 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_37 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_38 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_39 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_40 <= 0;
      __stream_matmul_29_sink_21_sink_offset_0_41 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_1 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_2 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_3 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_4 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_5 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_6 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_7 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_8 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_9 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_10 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_11 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_12 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_13 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_14 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_15 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_16 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_17 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_18 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_19 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_20 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_21 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_22 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_23 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_24 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_25 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_26 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_27 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_28 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_29 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_30 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_31 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_32 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_33 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_34 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_35 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_36 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_37 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_38 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_39 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_40 <= 0;
      __stream_matmul_29_sink_21_sink_size_1_41 <= 0;
      __stream_seq_16_cond_2_1 <= 0;
      __stream_seq_16_cond_2_2 <= 0;
      __stream_seq_16_cond_2_3 <= 0;
      __stream_seq_16_cond_2_4 <= 0;
      __stream_seq_16_cond_2_5 <= 0;
      __stream_seq_16_cond_2_6 <= 0;
      __stream_seq_16_cond_2_7 <= 0;
      __stream_seq_16_cond_2_8 <= 0;
      __stream_seq_16_cond_2_9 <= 0;
      __stream_seq_16_cond_2_10 <= 0;
      __stream_seq_16_cond_2_11 <= 0;
      __stream_seq_16_cond_2_12 <= 0;
      __stream_seq_16_cond_2_13 <= 0;
      __stream_seq_16_cond_2_14 <= 0;
      __stream_seq_16_cond_2_15 <= 0;
      __stream_seq_16_cond_2_16 <= 0;
      __stream_seq_16_cond_2_17 <= 0;
      __stream_seq_16_cond_2_18 <= 0;
      __stream_seq_16_cond_2_19 <= 0;
      __stream_seq_16_cond_2_20 <= 0;
      __stream_seq_16_cond_2_21 <= 0;
      __stream_seq_16_cond_2_22 <= 0;
      __stream_seq_16_cond_2_23 <= 0;
      __stream_seq_16_cond_2_24 <= 0;
      __stream_seq_16_cond_2_25 <= 0;
      __stream_seq_16_cond_2_26 <= 0;
      __stream_seq_16_cond_2_27 <= 0;
      __stream_seq_16_cond_2_28 <= 0;
      __stream_seq_16_cond_2_29 <= 0;
      __stream_seq_16_cond_2_30 <= 0;
      __stream_seq_16_cond_2_31 <= 0;
      __stream_seq_16_cond_2_32 <= 0;
      __stream_seq_16_cond_2_33 <= 0;
      __stream_seq_16_cond_2_34 <= 0;
      __stream_seq_16_cond_2_35 <= 0;
      __stream_seq_16_cond_2_36 <= 0;
      __stream_seq_16_cond_2_37 <= 0;
      __stream_seq_16_cond_2_38 <= 0;
      __stream_seq_16_cond_2_39 <= 0;
      __stream_seq_16_cond_2_40 <= 0;
      __stream_seq_16_cond_2_41 <= 0;
      _stream_matmul_29_sink_21_sink_mode <= 3'b0;
      _stream_matmul_29_sink_21_sink_offset <= 0;
      _stream_matmul_29_sink_21_sink_size <= 0;
      _stream_matmul_29_sink_21_sink_stride <= 0;
      __set_flag_1224_1 <= 0;
      __set_flag_1224_2 <= 0;
      __set_flag_1224_3 <= 0;
      __set_flag_1224_4 <= 0;
      __set_flag_1224_5 <= 0;
      __set_flag_1224_6 <= 0;
      __set_flag_1224_7 <= 0;
      __set_flag_1224_8 <= 0;
      __set_flag_1224_9 <= 0;
      __set_flag_1224_10 <= 0;
      __set_flag_1224_11 <= 0;
      __set_flag_1224_12 <= 0;
      __set_flag_1224_13 <= 0;
      __set_flag_1224_14 <= 0;
      __set_flag_1224_15 <= 0;
      __set_flag_1224_16 <= 0;
      __set_flag_1224_17 <= 0;
      __set_flag_1224_18 <= 0;
      __set_flag_1224_19 <= 0;
      __set_flag_1224_20 <= 0;
      __set_flag_1224_21 <= 0;
      __set_flag_1224_22 <= 0;
      __set_flag_1224_23 <= 0;
      __set_flag_1224_24 <= 0;
      __set_flag_1224_25 <= 0;
      __set_flag_1224_26 <= 0;
      __set_flag_1224_27 <= 0;
      __set_flag_1224_28 <= 0;
      __set_flag_1224_29 <= 0;
      __set_flag_1224_30 <= 0;
      __set_flag_1224_31 <= 0;
      __set_flag_1224_32 <= 0;
      __set_flag_1224_33 <= 0;
      __set_flag_1224_34 <= 0;
      __set_flag_1224_35 <= 0;
      __set_flag_1224_36 <= 0;
      __set_flag_1224_37 <= 0;
      __set_flag_1224_38 <= 0;
      __set_flag_1224_39 <= 0;
      __set_flag_1224_40 <= 0;
      __set_flag_1224_41 <= 0;
      _stream_matmul_29_sink_21_sink_ram_sel <= 0;
      __stream_matmul_29_start_1 <= 0;
      __stream_matmul_29_start_2 <= 0;
      __stream_matmul_29_start_3 <= 0;
      __stream_matmul_29_start_4 <= 0;
      __stream_matmul_29_start_5 <= 0;
      __stream_matmul_29_start_6 <= 0;
      __stream_matmul_29_start_7 <= 0;
      __stream_matmul_29_start_8 <= 0;
      __stream_matmul_29_start_9 <= 0;
      __stream_matmul_29_start_10 <= 0;
      __stream_matmul_29_start_11 <= 0;
      __stream_matmul_29_start_12 <= 0;
      __stream_matmul_29_start_13 <= 0;
      __stream_matmul_29_start_14 <= 0;
      __stream_matmul_29_start_15 <= 0;
      __stream_matmul_29_start_16 <= 0;
      __stream_matmul_29_start_17 <= 0;
      __stream_matmul_29_start_18 <= 0;
      __stream_matmul_29_start_19 <= 0;
      __stream_matmul_29_start_20 <= 0;
      __stream_matmul_29_start_21 <= 0;
      __stream_matmul_29_start_22 <= 0;
      __stream_matmul_29_start_23 <= 0;
      __stream_matmul_29_start_24 <= 0;
      __stream_matmul_29_start_25 <= 0;
      __stream_matmul_29_start_26 <= 0;
      __stream_matmul_29_start_27 <= 0;
      __stream_matmul_29_start_28 <= 0;
      __stream_matmul_29_start_29 <= 0;
      __stream_matmul_29_start_30 <= 0;
      __stream_matmul_29_start_31 <= 0;
      __stream_matmul_29_start_32 <= 0;
      __stream_matmul_29_start_33 <= 0;
      __stream_matmul_29_start_34 <= 0;
      __stream_matmul_29_start_35 <= 0;
      __stream_matmul_29_start_36 <= 0;
      __stream_matmul_29_start_37 <= 0;
      __stream_matmul_29_start_38 <= 0;
      __stream_matmul_29_start_39 <= 0;
      __stream_matmul_29_start_40 <= 0;
      __stream_matmul_29_start_41 <= 0;
      __stream_matmul_29_start_42 <= 0;
      _stream_matmul_29_sink_21_sink_waddr <= 0;
      _stream_matmul_29_sink_21_sink_count <= 0;
      _stream_matmul_29_sink_21_sink_offset_buf <= 0;
      _stream_matmul_29_sink_21_sink_stride_buf <= 0;
      _stream_matmul_29_sink_21_sink_wdata <= 0;
      __tmp_1227_1 <= 0;
      __tmp_1227_2 <= 0;
      __tmp_1227_3 <= 0;
      __tmp_1227_4 <= 0;
      __tmp_1227_5 <= 0;
      __tmp_1229_1 <= 0;
      __tmp_1229_2 <= 0;
      __tmp_1229_3 <= 0;
      __tmp_1229_4 <= 0;
      __tmp_1229_5 <= 0;
      __tmp_1229_6 <= 0;
      __tmp_1229_7 <= 0;
      __tmp_1229_8 <= 0;
      __tmp_1231_1 <= 0;
      __tmp_1231_2 <= 0;
      __tmp_1231_3 <= 0;
      __tmp_1231_4 <= 0;
      __tmp_1231_5 <= 0;
      __tmp_1231_6 <= 0;
      __tmp_1231_7 <= 0;
      __tmp_1231_8 <= 0;
      __tmp_1233_1 <= 0;
      __tmp_1233_2 <= 0;
      __tmp_1233_3 <= 0;
      __tmp_1233_4 <= 0;
      __tmp_1233_5 <= 0;
      __tmp_1233_6 <= 0;
      __tmp_1233_7 <= 0;
      __tmp_1233_8 <= 0;
      __tmp_1235_1 <= 0;
      __tmp_1235_2 <= 0;
      __tmp_1235_3 <= 0;
      __tmp_1235_4 <= 0;
      __tmp_1235_5 <= 0;
      __tmp_1235_6 <= 0;
      __tmp_1235_7 <= 0;
      __tmp_1235_8 <= 0;
      __tmp_1235_9 <= 0;
      __tmp_1235_10 <= 0;
      __tmp_1235_11 <= 0;
      __tmp_1235_12 <= 0;
      __tmp_1235_13 <= 0;
      __tmp_1235_14 <= 0;
      __tmp_1235_15 <= 0;
      __tmp_1235_16 <= 0;
      __tmp_1235_17 <= 0;
      __tmp_1235_18 <= 0;
      __tmp_1237_1 <= 0;
      __tmp_1237_2 <= 0;
      __tmp_1237_3 <= 0;
      __tmp_1237_4 <= 0;
      __tmp_1237_5 <= 0;
      __tmp_1237_6 <= 0;
      __tmp_1237_7 <= 0;
      __tmp_1237_8 <= 0;
      __tmp_1237_9 <= 0;
      __tmp_1237_10 <= 0;
      __tmp_1237_11 <= 0;
      __tmp_1237_12 <= 0;
      __tmp_1237_13 <= 0;
      __tmp_1237_14 <= 0;
      __tmp_1237_15 <= 0;
      __tmp_1237_16 <= 0;
      __tmp_1237_17 <= 0;
      __tmp_1237_18 <= 0;
      __tmp_1237_19 <= 0;
      __tmp_1237_20 <= 0;
      __tmp_1237_21 <= 0;
      __tmp_1237_22 <= 0;
      __tmp_1239_1 <= 0;
      __tmp_1239_2 <= 0;
      __tmp_1239_3 <= 0;
      __tmp_1239_4 <= 0;
      __tmp_1239_5 <= 0;
      __tmp_1239_6 <= 0;
      __tmp_1239_7 <= 0;
      __tmp_1239_8 <= 0;
      __tmp_1239_9 <= 0;
      __tmp_1239_10 <= 0;
      __tmp_1239_11 <= 0;
      __tmp_1239_12 <= 0;
      __tmp_1239_13 <= 0;
      __tmp_1239_14 <= 0;
      __tmp_1239_15 <= 0;
      __tmp_1239_16 <= 0;
      __tmp_1239_17 <= 0;
      __tmp_1239_18 <= 0;
      __tmp_1239_19 <= 0;
      __tmp_1239_20 <= 0;
      __tmp_1241_1 <= 0;
      __tmp_1241_2 <= 0;
      __tmp_1241_3 <= 0;
      __tmp_1241_4 <= 0;
      __tmp_1241_5 <= 0;
      __tmp_1241_6 <= 0;
      __tmp_1241_7 <= 0;
      __tmp_1241_8 <= 0;
      __tmp_1241_9 <= 0;
      __tmp_1241_10 <= 0;
      __tmp_1241_11 <= 0;
      __tmp_1241_12 <= 0;
      __tmp_1241_13 <= 0;
      __tmp_1241_14 <= 0;
      __tmp_1241_15 <= 0;
      __tmp_1241_16 <= 0;
      __tmp_1241_17 <= 0;
      __tmp_1241_18 <= 0;
      __tmp_1241_19 <= 0;
      __tmp_1241_20 <= 0;
      __tmp_1243_1 <= 0;
      __tmp_1243_2 <= 0;
      __tmp_1243_3 <= 0;
      __tmp_1243_4 <= 0;
      __tmp_1243_5 <= 0;
      __tmp_1243_6 <= 0;
      __tmp_1243_7 <= 0;
      __tmp_1243_8 <= 0;
      __tmp_1243_9 <= 0;
      __tmp_1243_10 <= 0;
      __tmp_1243_11 <= 0;
      __tmp_1243_12 <= 0;
      __tmp_1243_13 <= 0;
      __tmp_1243_14 <= 0;
      __tmp_1243_15 <= 0;
      __tmp_1243_16 <= 0;
      __tmp_1243_17 <= 0;
      __tmp_1243_18 <= 0;
      __tmp_1243_19 <= 0;
      __tmp_1243_20 <= 0;
      __tmp_1245_1 <= 0;
      __tmp_1245_2 <= 0;
      __tmp_1245_3 <= 0;
      __tmp_1245_4 <= 0;
      __tmp_1245_5 <= 0;
      __tmp_1245_6 <= 0;
      __tmp_1245_7 <= 0;
      __tmp_1245_8 <= 0;
      __tmp_1245_9 <= 0;
      __tmp_1245_10 <= 0;
      __tmp_1245_11 <= 0;
      __tmp_1245_12 <= 0;
      __tmp_1245_13 <= 0;
      __tmp_1245_14 <= 0;
      __tmp_1245_15 <= 0;
      __tmp_1245_16 <= 0;
      __tmp_1245_17 <= 0;
      __tmp_1245_18 <= 0;
      __tmp_1245_19 <= 0;
      __tmp_1245_20 <= 0;
      __tmp_1245_21 <= 0;
      __tmp_1245_22 <= 0;
      __tmp_1245_23 <= 0;
      __tmp_1245_24 <= 0;
      __tmp_1245_25 <= 0;
      __tmp_1245_26 <= 0;
      __tmp_1245_27 <= 0;
      __tmp_1245_28 <= 0;
      __tmp_1247_1 <= 0;
      __tmp_1247_2 <= 0;
      __tmp_1247_3 <= 0;
      __tmp_1247_4 <= 0;
      __tmp_1247_5 <= 0;
      __tmp_1247_6 <= 0;
      __tmp_1247_7 <= 0;
      __tmp_1247_8 <= 0;
      __tmp_1247_9 <= 0;
      __tmp_1247_10 <= 0;
      __tmp_1247_11 <= 0;
      __tmp_1247_12 <= 0;
      __tmp_1247_13 <= 0;
      __tmp_1247_14 <= 0;
      __tmp_1247_15 <= 0;
      __tmp_1247_16 <= 0;
      __tmp_1247_17 <= 0;
      __tmp_1247_18 <= 0;
      __tmp_1247_19 <= 0;
      __tmp_1247_20 <= 0;
      __tmp_1247_21 <= 0;
      __tmp_1247_22 <= 0;
      __tmp_1247_23 <= 0;
      __tmp_1247_24 <= 0;
      __tmp_1247_25 <= 0;
      __tmp_1247_26 <= 0;
      __tmp_1247_27 <= 0;
      __tmp_1247_28 <= 0;
      __tmp_1249_1 <= 0;
      __tmp_1249_2 <= 0;
      __tmp_1249_3 <= 0;
      __tmp_1249_4 <= 0;
      __tmp_1249_5 <= 0;
      __tmp_1249_6 <= 0;
      __tmp_1249_7 <= 0;
      __tmp_1249_8 <= 0;
      __tmp_1249_9 <= 0;
      __tmp_1249_10 <= 0;
      __tmp_1249_11 <= 0;
      __tmp_1249_12 <= 0;
      __tmp_1249_13 <= 0;
      __tmp_1249_14 <= 0;
      __tmp_1249_15 <= 0;
      __tmp_1249_16 <= 0;
      __tmp_1249_17 <= 0;
      __tmp_1249_18 <= 0;
      __tmp_1249_19 <= 0;
      __tmp_1249_20 <= 0;
      __tmp_1249_21 <= 0;
      __tmp_1249_22 <= 0;
      __tmp_1249_23 <= 0;
      __tmp_1249_24 <= 0;
      __tmp_1249_25 <= 0;
      __tmp_1249_26 <= 0;
      __tmp_1249_27 <= 0;
      __tmp_1249_28 <= 0;
      __tmp_1251_1 <= 0;
      __tmp_1253_1 <= 0;
      __tmp_1253_2 <= 0;
      __tmp_1253_3 <= 0;
      __tmp_1253_4 <= 0;
      __tmp_1253_5 <= 0;
      __tmp_1255_1 <= 0;
      __tmp_1255_2 <= 0;
      __tmp_1255_3 <= 0;
      __tmp_1255_4 <= 0;
      __tmp_1255_5 <= 0;
      __tmp_1257_1 <= 0;
      __tmp_1257_2 <= 0;
      __tmp_1257_3 <= 0;
      __tmp_1257_4 <= 0;
      __tmp_1257_5 <= 0;
      __tmp_1265_1 <= 0;
      __tmp_1265_2 <= 0;
      __tmp_1265_3 <= 0;
      __tmp_1265_4 <= 0;
      __tmp_1265_5 <= 0;
      __tmp_1265_6 <= 0;
      __tmp_1265_7 <= 0;
      __tmp_1265_8 <= 0;
      __tmp_1265_9 <= 0;
      __tmp_1265_10 <= 0;
      __tmp_1265_11 <= 0;
      __tmp_1265_12 <= 0;
      __tmp_1265_13 <= 0;
      __tmp_1265_14 <= 0;
      __tmp_1265_15 <= 0;
      __tmp_1273_1 <= 0;
      __tmp_1273_2 <= 0;
      __tmp_1273_3 <= 0;
      __tmp_1273_4 <= 0;
      __tmp_1273_5 <= 0;
      __tmp_1273_6 <= 0;
      __tmp_1273_7 <= 0;
      __tmp_1273_8 <= 0;
      __tmp_1273_9 <= 0;
      __tmp_1273_10 <= 0;
      __tmp_1273_11 <= 0;
      __tmp_1273_12 <= 0;
      __tmp_1273_13 <= 0;
      __tmp_1273_14 <= 0;
      __tmp_1273_15 <= 0;
      __tmp_1273_16 <= 0;
      __tmp_1273_17 <= 0;
      __tmp_1273_18 <= 0;
      __tmp_1275_1 <= 0;
      __tmp_1275_2 <= 0;
      __tmp_1275_3 <= 0;
      __tmp_1275_4 <= 0;
      __tmp_1275_5 <= 0;
      __tmp_1275_6 <= 0;
      __tmp_1275_7 <= 0;
      __tmp_1275_8 <= 0;
      __tmp_1275_9 <= 0;
      __tmp_1275_10 <= 0;
      __tmp_1275_11 <= 0;
      __tmp_1275_12 <= 0;
      __tmp_1275_13 <= 0;
      __tmp_1275_14 <= 0;
      __tmp_1275_15 <= 0;
      __tmp_1275_16 <= 0;
      __tmp_1275_17 <= 0;
      __tmp_1277_1 <= 0;
      __tmp_1277_2 <= 0;
      __tmp_1277_3 <= 0;
      __tmp_1277_4 <= 0;
      __tmp_1277_5 <= 0;
      __tmp_1277_6 <= 0;
      __tmp_1277_7 <= 0;
      __tmp_1277_8 <= 0;
      __tmp_1277_9 <= 0;
      __tmp_1277_10 <= 0;
      __tmp_1277_11 <= 0;
      __tmp_1277_12 <= 0;
      __tmp_1277_13 <= 0;
      __tmp_1277_14 <= 0;
      __tmp_1277_15 <= 0;
      __tmp_1277_16 <= 0;
      __tmp_1277_17 <= 0;
      __tmp_1279_1 <= 0;
      __tmp_1279_2 <= 0;
      __tmp_1279_3 <= 0;
      __tmp_1279_4 <= 0;
      __tmp_1279_5 <= 0;
      __tmp_1279_6 <= 0;
      __tmp_1279_7 <= 0;
      __tmp_1279_8 <= 0;
      __tmp_1279_9 <= 0;
      __tmp_1279_10 <= 0;
      __tmp_1279_11 <= 0;
      __tmp_1279_12 <= 0;
      __tmp_1279_13 <= 0;
      __tmp_1279_14 <= 0;
      __tmp_1279_15 <= 0;
      __tmp_1279_16 <= 0;
      __tmp_1279_17 <= 0;
      __tmp_1287_1 <= 0;
      __tmp_1287_2 <= 0;
      __tmp_1287_3 <= 0;
      __tmp_1287_4 <= 0;
      __tmp_1287_5 <= 0;
      __tmp_1287_6 <= 0;
      __tmp_1287_7 <= 0;
      __tmp_1287_8 <= 0;
      __tmp_1287_9 <= 0;
      __tmp_1287_10 <= 0;
      __tmp_1287_11 <= 0;
      __tmp_1287_12 <= 0;
      __tmp_1287_13 <= 0;
      __tmp_1287_14 <= 0;
      __tmp_1287_15 <= 0;
      __tmp_1287_16 <= 0;
      __tmp_1287_17 <= 0;
      __tmp_1287_18 <= 0;
      __tmp_1287_19 <= 0;
      __tmp_1287_20 <= 0;
      __tmp_1287_21 <= 0;
      __tmp_1287_22 <= 0;
      __tmp_1287_23 <= 0;
      __tmp_1287_24 <= 0;
      __tmp_1287_25 <= 0;
      __tmp_1289_1 <= 0;
      __tmp_1289_2 <= 0;
      __tmp_1289_3 <= 0;
      __tmp_1289_4 <= 0;
      __tmp_1289_5 <= 0;
      __tmp_1289_6 <= 0;
      __tmp_1289_7 <= 0;
      __tmp_1289_8 <= 0;
      __tmp_1289_9 <= 0;
      __tmp_1289_10 <= 0;
      __tmp_1289_11 <= 0;
      __tmp_1289_12 <= 0;
      __tmp_1289_13 <= 0;
      __tmp_1289_14 <= 0;
      __tmp_1289_15 <= 0;
      __tmp_1289_16 <= 0;
      __tmp_1289_17 <= 0;
      __tmp_1289_18 <= 0;
      __tmp_1289_19 <= 0;
      __tmp_1289_20 <= 0;
      __tmp_1289_21 <= 0;
      __tmp_1289_22 <= 0;
      __tmp_1289_23 <= 0;
      __tmp_1289_24 <= 0;
      __tmp_1289_25 <= 0;
      __tmp_1291_1 <= 0;
      __tmp_1291_2 <= 0;
      __tmp_1291_3 <= 0;
      __tmp_1291_4 <= 0;
      __tmp_1291_5 <= 0;
      __tmp_1291_6 <= 0;
      __tmp_1291_7 <= 0;
      __tmp_1291_8 <= 0;
      __tmp_1291_9 <= 0;
      __tmp_1291_10 <= 0;
      __tmp_1291_11 <= 0;
      __tmp_1291_12 <= 0;
      __tmp_1291_13 <= 0;
      __tmp_1291_14 <= 0;
      __tmp_1291_15 <= 0;
      __tmp_1291_16 <= 0;
      __tmp_1291_17 <= 0;
      __tmp_1291_18 <= 0;
      __tmp_1291_19 <= 0;
      __tmp_1291_20 <= 0;
      __tmp_1291_21 <= 0;
      __tmp_1291_22 <= 0;
      __tmp_1291_23 <= 0;
      __tmp_1291_24 <= 0;
      __tmp_1291_25 <= 0;
      __tmp_1299_1 <= 0;
      __tmp_1299_2 <= 0;
      __tmp_1299_3 <= 0;
      __tmp_1299_4 <= 0;
      __tmp_1299_5 <= 0;
      __tmp_1299_6 <= 0;
      __tmp_1299_7 <= 0;
      __tmp_1299_8 <= 0;
      __tmp_1299_9 <= 0;
      __tmp_1299_10 <= 0;
      __tmp_1299_11 <= 0;
      __tmp_1299_12 <= 0;
      __tmp_1299_13 <= 0;
      __tmp_1299_14 <= 0;
      __tmp_1299_15 <= 0;
      __tmp_1299_16 <= 0;
      __tmp_1299_17 <= 0;
      __tmp_1299_18 <= 0;
      __tmp_1299_19 <= 0;
      __tmp_1299_20 <= 0;
      __tmp_1299_21 <= 0;
      __tmp_1299_22 <= 0;
      __tmp_1299_23 <= 0;
      __tmp_1299_24 <= 0;
      __tmp_1299_25 <= 0;
      __tmp_1299_26 <= 0;
      __tmp_1299_27 <= 0;
      __tmp_1299_28 <= 0;
      __tmp_1299_29 <= 0;
      __tmp_1299_30 <= 0;
      __tmp_1299_31 <= 0;
      __tmp_1299_32 <= 0;
      __tmp_1299_33 <= 0;
      __tmp_1299_34 <= 0;
      __tmp_1299_35 <= 0;
      __tmp_1299_36 <= 0;
      __tmp_1299_37 <= 0;
      __tmp_1299_38 <= 0;
      __tmp_1299_39 <= 0;
      __tmp_1299_40 <= 0;
      __tmp_1299_41 <= 0;
      __tmp_1299_42 <= 0;
      __tmp_1301_1 <= 0;
      __tmp_1301_2 <= 0;
      __tmp_1301_3 <= 0;
      __tmp_1301_4 <= 0;
      __tmp_1301_5 <= 0;
      __tmp_1301_6 <= 0;
      __tmp_1301_7 <= 0;
      __tmp_1301_8 <= 0;
      __tmp_1301_9 <= 0;
      __tmp_1301_10 <= 0;
      __tmp_1301_11 <= 0;
      __tmp_1301_12 <= 0;
      __tmp_1301_13 <= 0;
      __tmp_1301_14 <= 0;
      __tmp_1301_15 <= 0;
      __tmp_1301_16 <= 0;
      __tmp_1301_17 <= 0;
      __tmp_1301_18 <= 0;
      __tmp_1301_19 <= 0;
      __tmp_1301_20 <= 0;
      __tmp_1301_21 <= 0;
      __tmp_1301_22 <= 0;
      __tmp_1301_23 <= 0;
      __tmp_1301_24 <= 0;
      __tmp_1301_25 <= 0;
      __tmp_1301_26 <= 0;
      __tmp_1301_27 <= 0;
      __tmp_1301_28 <= 0;
      __tmp_1301_29 <= 0;
      __tmp_1301_30 <= 0;
      __tmp_1301_31 <= 0;
      __tmp_1301_32 <= 0;
      __tmp_1301_33 <= 0;
      __tmp_1301_34 <= 0;
      __tmp_1301_35 <= 0;
      __tmp_1301_36 <= 0;
      __tmp_1301_37 <= 0;
      __tmp_1301_38 <= 0;
      __tmp_1301_39 <= 0;
      __tmp_1301_40 <= 0;
      __tmp_1301_41 <= 0;
      __tmp_1301_42 <= 0;
      __tmp_1303_1 <= 0;
      __tmp_1303_2 <= 0;
      __tmp_1303_3 <= 0;
      __tmp_1303_4 <= 0;
      __tmp_1303_5 <= 0;
      __tmp_1303_6 <= 0;
      __tmp_1303_7 <= 0;
      __tmp_1303_8 <= 0;
      __tmp_1303_9 <= 0;
      __tmp_1303_10 <= 0;
      __tmp_1303_11 <= 0;
      __tmp_1303_12 <= 0;
      __tmp_1303_13 <= 0;
      __tmp_1303_14 <= 0;
      __tmp_1303_15 <= 0;
      __tmp_1303_16 <= 0;
      __tmp_1303_17 <= 0;
      __tmp_1303_18 <= 0;
      __tmp_1303_19 <= 0;
      __tmp_1303_20 <= 0;
      __tmp_1303_21 <= 0;
      __tmp_1303_22 <= 0;
      __tmp_1303_23 <= 0;
      __tmp_1303_24 <= 0;
      __tmp_1303_25 <= 0;
      __tmp_1303_26 <= 0;
      __tmp_1303_27 <= 0;
      __tmp_1303_28 <= 0;
      __tmp_1303_29 <= 0;
      __tmp_1303_30 <= 0;
      __tmp_1303_31 <= 0;
      __tmp_1303_32 <= 0;
      __tmp_1303_33 <= 0;
      __tmp_1303_34 <= 0;
      __tmp_1303_35 <= 0;
      __tmp_1303_36 <= 0;
      __tmp_1303_37 <= 0;
      __tmp_1303_38 <= 0;
      __tmp_1303_39 <= 0;
      __tmp_1303_40 <= 0;
      __tmp_1303_41 <= 0;
      __tmp_1303_42 <= 0;
      __tmp_1305_1 <= 0;
      __tmp_1305_2 <= 0;
      __tmp_1305_3 <= 0;
      __tmp_1305_4 <= 0;
      __tmp_1305_5 <= 0;
      __tmp_1305_6 <= 0;
      __tmp_1305_7 <= 0;
      __tmp_1305_8 <= 0;
      __tmp_1305_9 <= 0;
      __tmp_1305_10 <= 0;
      __tmp_1305_11 <= 0;
      __tmp_1305_12 <= 0;
      __tmp_1305_13 <= 0;
      __tmp_1305_14 <= 0;
      __tmp_1305_15 <= 0;
      __tmp_1305_16 <= 0;
      __tmp_1305_17 <= 0;
      __tmp_1305_18 <= 0;
      __tmp_1305_19 <= 0;
      __tmp_1305_20 <= 0;
      __tmp_1305_21 <= 0;
      __tmp_1305_22 <= 0;
      __tmp_1305_23 <= 0;
      __tmp_1305_24 <= 0;
      __tmp_1305_25 <= 0;
      __tmp_1305_26 <= 0;
      __tmp_1305_27 <= 0;
      __tmp_1305_28 <= 0;
      __tmp_1305_29 <= 0;
      __tmp_1305_30 <= 0;
      __tmp_1305_31 <= 0;
      __tmp_1305_32 <= 0;
      __tmp_1305_33 <= 0;
      __tmp_1305_34 <= 0;
      __tmp_1305_35 <= 0;
      __tmp_1305_36 <= 0;
      __tmp_1305_37 <= 0;
      __tmp_1305_38 <= 0;
      __tmp_1305_39 <= 0;
      __tmp_1305_40 <= 0;
      __tmp_1305_41 <= 0;
      __tmp_1305_42 <= 0;
      __tmp_1307_1 <= 0;
      __tmp_1307_2 <= 0;
      __tmp_1307_3 <= 0;
      __tmp_1307_4 <= 0;
      __tmp_1307_5 <= 0;
      __tmp_1307_6 <= 0;
      __tmp_1307_7 <= 0;
      __tmp_1307_8 <= 0;
      __tmp_1307_9 <= 0;
      __tmp_1307_10 <= 0;
      __tmp_1307_11 <= 0;
      __tmp_1307_12 <= 0;
      __tmp_1307_13 <= 0;
      __tmp_1307_14 <= 0;
      __tmp_1307_15 <= 0;
      __tmp_1307_16 <= 0;
      __tmp_1307_17 <= 0;
      __tmp_1307_18 <= 0;
      __tmp_1307_19 <= 0;
      __tmp_1307_20 <= 0;
      __tmp_1307_21 <= 0;
      __tmp_1307_22 <= 0;
      __tmp_1307_23 <= 0;
      __tmp_1307_24 <= 0;
      __tmp_1307_25 <= 0;
      __tmp_1307_26 <= 0;
      __tmp_1307_27 <= 0;
      __tmp_1307_28 <= 0;
      __tmp_1307_29 <= 0;
      __tmp_1307_30 <= 0;
      __tmp_1307_31 <= 0;
      __tmp_1307_32 <= 0;
      __tmp_1307_33 <= 0;
      __tmp_1307_34 <= 0;
      __tmp_1307_35 <= 0;
      __tmp_1307_36 <= 0;
      __tmp_1307_37 <= 0;
      __tmp_1307_38 <= 0;
    end else begin
      if(__stream_seq_16_cond_2_41) begin
        _stream_matmul_29_sink_21_sink_mode <= 3'b1;
        _stream_matmul_29_sink_21_sink_offset <= __stream_matmul_29_sink_21_sink_offset_0_41;
        _stream_matmul_29_sink_21_sink_size <= __stream_matmul_29_sink_21_sink_size_1_41;
        _stream_matmul_29_sink_21_sink_stride <= 1;
      end 
      __stream_matmul_29_sink_21_sink_offset_0_41 <= __stream_matmul_29_sink_21_sink_offset_0_40;
      __stream_matmul_29_sink_21_sink_size_1_41 <= __stream_matmul_29_sink_21_sink_size_1_40;
      __stream_seq_16_cond_2_41 <= __stream_seq_16_cond_2_40;
      __stream_matmul_29_sink_21_sink_offset_0_40 <= __stream_matmul_29_sink_21_sink_offset_0_39;
      __stream_matmul_29_sink_21_sink_size_1_40 <= __stream_matmul_29_sink_21_sink_size_1_39;
      __stream_seq_16_cond_2_40 <= __stream_seq_16_cond_2_39;
      __stream_matmul_29_sink_21_sink_offset_0_39 <= __stream_matmul_29_sink_21_sink_offset_0_38;
      __stream_matmul_29_sink_21_sink_size_1_39 <= __stream_matmul_29_sink_21_sink_size_1_38;
      __stream_seq_16_cond_2_39 <= __stream_seq_16_cond_2_38;
      __stream_matmul_29_sink_21_sink_offset_0_38 <= __stream_matmul_29_sink_21_sink_offset_0_37;
      __stream_matmul_29_sink_21_sink_size_1_38 <= __stream_matmul_29_sink_21_sink_size_1_37;
      __stream_seq_16_cond_2_38 <= __stream_seq_16_cond_2_37;
      __stream_matmul_29_sink_21_sink_offset_0_37 <= __stream_matmul_29_sink_21_sink_offset_0_36;
      __stream_matmul_29_sink_21_sink_size_1_37 <= __stream_matmul_29_sink_21_sink_size_1_36;
      __stream_seq_16_cond_2_37 <= __stream_seq_16_cond_2_36;
      __stream_matmul_29_sink_21_sink_offset_0_36 <= __stream_matmul_29_sink_21_sink_offset_0_35;
      __stream_matmul_29_sink_21_sink_size_1_36 <= __stream_matmul_29_sink_21_sink_size_1_35;
      __stream_seq_16_cond_2_36 <= __stream_seq_16_cond_2_35;
      __stream_matmul_29_sink_21_sink_offset_0_35 <= __stream_matmul_29_sink_21_sink_offset_0_34;
      __stream_matmul_29_sink_21_sink_size_1_35 <= __stream_matmul_29_sink_21_sink_size_1_34;
      __stream_seq_16_cond_2_35 <= __stream_seq_16_cond_2_34;
      __stream_matmul_29_sink_21_sink_offset_0_34 <= __stream_matmul_29_sink_21_sink_offset_0_33;
      __stream_matmul_29_sink_21_sink_size_1_34 <= __stream_matmul_29_sink_21_sink_size_1_33;
      __stream_seq_16_cond_2_34 <= __stream_seq_16_cond_2_33;
      __stream_matmul_29_sink_21_sink_offset_0_33 <= __stream_matmul_29_sink_21_sink_offset_0_32;
      __stream_matmul_29_sink_21_sink_size_1_33 <= __stream_matmul_29_sink_21_sink_size_1_32;
      __stream_seq_16_cond_2_33 <= __stream_seq_16_cond_2_32;
      __stream_matmul_29_sink_21_sink_offset_0_32 <= __stream_matmul_29_sink_21_sink_offset_0_31;
      __stream_matmul_29_sink_21_sink_size_1_32 <= __stream_matmul_29_sink_21_sink_size_1_31;
      __stream_seq_16_cond_2_32 <= __stream_seq_16_cond_2_31;
      __stream_matmul_29_sink_21_sink_offset_0_31 <= __stream_matmul_29_sink_21_sink_offset_0_30;
      __stream_matmul_29_sink_21_sink_size_1_31 <= __stream_matmul_29_sink_21_sink_size_1_30;
      __stream_seq_16_cond_2_31 <= __stream_seq_16_cond_2_30;
      __stream_matmul_29_sink_21_sink_offset_0_30 <= __stream_matmul_29_sink_21_sink_offset_0_29;
      __stream_matmul_29_sink_21_sink_size_1_30 <= __stream_matmul_29_sink_21_sink_size_1_29;
      __stream_seq_16_cond_2_30 <= __stream_seq_16_cond_2_29;
      __stream_matmul_29_sink_21_sink_offset_0_29 <= __stream_matmul_29_sink_21_sink_offset_0_28;
      __stream_matmul_29_sink_21_sink_size_1_29 <= __stream_matmul_29_sink_21_sink_size_1_28;
      __stream_seq_16_cond_2_29 <= __stream_seq_16_cond_2_28;
      __stream_matmul_29_sink_21_sink_offset_0_28 <= __stream_matmul_29_sink_21_sink_offset_0_27;
      __stream_matmul_29_sink_21_sink_size_1_28 <= __stream_matmul_29_sink_21_sink_size_1_27;
      __stream_seq_16_cond_2_28 <= __stream_seq_16_cond_2_27;
      __stream_matmul_29_sink_21_sink_offset_0_27 <= __stream_matmul_29_sink_21_sink_offset_0_26;
      __stream_matmul_29_sink_21_sink_size_1_27 <= __stream_matmul_29_sink_21_sink_size_1_26;
      __stream_seq_16_cond_2_27 <= __stream_seq_16_cond_2_26;
      __stream_matmul_29_sink_21_sink_offset_0_26 <= __stream_matmul_29_sink_21_sink_offset_0_25;
      __stream_matmul_29_sink_21_sink_size_1_26 <= __stream_matmul_29_sink_21_sink_size_1_25;
      __stream_seq_16_cond_2_26 <= __stream_seq_16_cond_2_25;
      __stream_matmul_29_sink_21_sink_offset_0_25 <= __stream_matmul_29_sink_21_sink_offset_0_24;
      __stream_matmul_29_sink_21_sink_size_1_25 <= __stream_matmul_29_sink_21_sink_size_1_24;
      __stream_seq_16_cond_2_25 <= __stream_seq_16_cond_2_24;
      __stream_matmul_29_sink_21_sink_offset_0_24 <= __stream_matmul_29_sink_21_sink_offset_0_23;
      __stream_matmul_29_sink_21_sink_size_1_24 <= __stream_matmul_29_sink_21_sink_size_1_23;
      __stream_seq_16_cond_2_24 <= __stream_seq_16_cond_2_23;
      __stream_matmul_29_sink_21_sink_offset_0_23 <= __stream_matmul_29_sink_21_sink_offset_0_22;
      __stream_matmul_29_sink_21_sink_size_1_23 <= __stream_matmul_29_sink_21_sink_size_1_22;
      __stream_seq_16_cond_2_23 <= __stream_seq_16_cond_2_22;
      __stream_matmul_29_sink_21_sink_offset_0_22 <= __stream_matmul_29_sink_21_sink_offset_0_21;
      __stream_matmul_29_sink_21_sink_size_1_22 <= __stream_matmul_29_sink_21_sink_size_1_21;
      __stream_seq_16_cond_2_22 <= __stream_seq_16_cond_2_21;
      __stream_matmul_29_sink_21_sink_offset_0_21 <= __stream_matmul_29_sink_21_sink_offset_0_20;
      __stream_matmul_29_sink_21_sink_size_1_21 <= __stream_matmul_29_sink_21_sink_size_1_20;
      __stream_seq_16_cond_2_21 <= __stream_seq_16_cond_2_20;
      __stream_matmul_29_sink_21_sink_offset_0_20 <= __stream_matmul_29_sink_21_sink_offset_0_19;
      __stream_matmul_29_sink_21_sink_size_1_20 <= __stream_matmul_29_sink_21_sink_size_1_19;
      __stream_seq_16_cond_2_20 <= __stream_seq_16_cond_2_19;
      __stream_matmul_29_sink_21_sink_offset_0_19 <= __stream_matmul_29_sink_21_sink_offset_0_18;
      __stream_matmul_29_sink_21_sink_size_1_19 <= __stream_matmul_29_sink_21_sink_size_1_18;
      __stream_seq_16_cond_2_19 <= __stream_seq_16_cond_2_18;
      __stream_matmul_29_sink_21_sink_offset_0_18 <= __stream_matmul_29_sink_21_sink_offset_0_17;
      __stream_matmul_29_sink_21_sink_size_1_18 <= __stream_matmul_29_sink_21_sink_size_1_17;
      __stream_seq_16_cond_2_18 <= __stream_seq_16_cond_2_17;
      __stream_matmul_29_sink_21_sink_offset_0_17 <= __stream_matmul_29_sink_21_sink_offset_0_16;
      __stream_matmul_29_sink_21_sink_size_1_17 <= __stream_matmul_29_sink_21_sink_size_1_16;
      __stream_seq_16_cond_2_17 <= __stream_seq_16_cond_2_16;
      __stream_matmul_29_sink_21_sink_offset_0_16 <= __stream_matmul_29_sink_21_sink_offset_0_15;
      __stream_matmul_29_sink_21_sink_size_1_16 <= __stream_matmul_29_sink_21_sink_size_1_15;
      __stream_seq_16_cond_2_16 <= __stream_seq_16_cond_2_15;
      __stream_matmul_29_sink_21_sink_offset_0_15 <= __stream_matmul_29_sink_21_sink_offset_0_14;
      __stream_matmul_29_sink_21_sink_size_1_15 <= __stream_matmul_29_sink_21_sink_size_1_14;
      __stream_seq_16_cond_2_15 <= __stream_seq_16_cond_2_14;
      __stream_matmul_29_sink_21_sink_offset_0_14 <= __stream_matmul_29_sink_21_sink_offset_0_13;
      __stream_matmul_29_sink_21_sink_size_1_14 <= __stream_matmul_29_sink_21_sink_size_1_13;
      __stream_seq_16_cond_2_14 <= __stream_seq_16_cond_2_13;
      __stream_matmul_29_sink_21_sink_offset_0_13 <= __stream_matmul_29_sink_21_sink_offset_0_12;
      __stream_matmul_29_sink_21_sink_size_1_13 <= __stream_matmul_29_sink_21_sink_size_1_12;
      __stream_seq_16_cond_2_13 <= __stream_seq_16_cond_2_12;
      __stream_matmul_29_sink_21_sink_offset_0_12 <= __stream_matmul_29_sink_21_sink_offset_0_11;
      __stream_matmul_29_sink_21_sink_size_1_12 <= __stream_matmul_29_sink_21_sink_size_1_11;
      __stream_seq_16_cond_2_12 <= __stream_seq_16_cond_2_11;
      __stream_matmul_29_sink_21_sink_offset_0_11 <= __stream_matmul_29_sink_21_sink_offset_0_10;
      __stream_matmul_29_sink_21_sink_size_1_11 <= __stream_matmul_29_sink_21_sink_size_1_10;
      __stream_seq_16_cond_2_11 <= __stream_seq_16_cond_2_10;
      __stream_matmul_29_sink_21_sink_offset_0_10 <= __stream_matmul_29_sink_21_sink_offset_0_9;
      __stream_matmul_29_sink_21_sink_size_1_10 <= __stream_matmul_29_sink_21_sink_size_1_9;
      __stream_seq_16_cond_2_10 <= __stream_seq_16_cond_2_9;
      __stream_matmul_29_sink_21_sink_offset_0_9 <= __stream_matmul_29_sink_21_sink_offset_0_8;
      __stream_matmul_29_sink_21_sink_size_1_9 <= __stream_matmul_29_sink_21_sink_size_1_8;
      __stream_seq_16_cond_2_9 <= __stream_seq_16_cond_2_8;
      __stream_matmul_29_sink_21_sink_offset_0_8 <= __stream_matmul_29_sink_21_sink_offset_0_7;
      __stream_matmul_29_sink_21_sink_size_1_8 <= __stream_matmul_29_sink_21_sink_size_1_7;
      __stream_seq_16_cond_2_8 <= __stream_seq_16_cond_2_7;
      __stream_matmul_29_sink_21_sink_offset_0_7 <= __stream_matmul_29_sink_21_sink_offset_0_6;
      __stream_matmul_29_sink_21_sink_size_1_7 <= __stream_matmul_29_sink_21_sink_size_1_6;
      __stream_seq_16_cond_2_7 <= __stream_seq_16_cond_2_6;
      __stream_matmul_29_sink_21_sink_offset_0_6 <= __stream_matmul_29_sink_21_sink_offset_0_5;
      __stream_matmul_29_sink_21_sink_size_1_6 <= __stream_matmul_29_sink_21_sink_size_1_5;
      __stream_seq_16_cond_2_6 <= __stream_seq_16_cond_2_5;
      __stream_matmul_29_sink_21_sink_offset_0_5 <= __stream_matmul_29_sink_21_sink_offset_0_4;
      __stream_matmul_29_sink_21_sink_size_1_5 <= __stream_matmul_29_sink_21_sink_size_1_4;
      __stream_seq_16_cond_2_5 <= __stream_seq_16_cond_2_4;
      __stream_matmul_29_sink_21_sink_offset_0_4 <= __stream_matmul_29_sink_21_sink_offset_0_3;
      __stream_matmul_29_sink_21_sink_size_1_4 <= __stream_matmul_29_sink_21_sink_size_1_3;
      __stream_seq_16_cond_2_4 <= __stream_seq_16_cond_2_3;
      __stream_matmul_29_sink_21_sink_offset_0_3 <= __stream_matmul_29_sink_21_sink_offset_0_2;
      __stream_matmul_29_sink_21_sink_size_1_3 <= __stream_matmul_29_sink_21_sink_size_1_2;
      __stream_seq_16_cond_2_3 <= __stream_seq_16_cond_2_2;
      __stream_matmul_29_sink_21_sink_offset_0_2 <= __stream_matmul_29_sink_21_sink_offset_0_1;
      __stream_matmul_29_sink_21_sink_size_1_2 <= __stream_matmul_29_sink_21_sink_size_1_1;
      __stream_seq_16_cond_2_2 <= __stream_seq_16_cond_2_1;
      _stream_matmul_29_source_6_idle <= _stream_matmul_29_source_6_idle;
      _stream_matmul_29_source_6_source_ram_rvalid <= 0;
      _stream_matmul_29_source_8_idle <= _stream_matmul_29_source_8_idle;
      _stream_matmul_29_source_8_source_ram_rvalid <= 0;
      _stream_matmul_29_source_10_idle <= _stream_matmul_29_source_10_idle;
      _stream_matmul_29_source_10_source_ram_rvalid <= 0;
      _stream_matmul_29_source_12_idle <= _stream_matmul_29_source_12_idle;
      _stream_matmul_29_source_12_source_ram_rvalid <= 0;
      _stream_matmul_29_source_14_idle <= _stream_matmul_29_source_14_idle;
      _stream_matmul_29_source_14_source_ram_rvalid <= 0;
      _stream_matmul_29_source_19_idle <= _stream_matmul_29_source_19_idle;
      _stream_matmul_29_source_19_source_ram_rvalid <= 0;
      _stream_matmul_29_source_20_idle <= _stream_matmul_29_source_20_idle;
      _stream_matmul_29_source_20_source_ram_rvalid <= 0;
      _stream_matmul_29_sink_21_sink_wenable <= 0;
      _stream_matmul_29_sink_22_sink_wenable <= 0;
      _cond_data_817 <= (stream_matmul_29_constant_5_data)? _reinterpretcast_data_816 : _reinterpretcast_data_816;
      _cond_data_824 <= (stream_matmul_29_constant_7_data)? _reinterpretcast_data_823 : _reinterpretcast_data_823;
      _cond_data_831 <= (stream_matmul_29_constant_9_data)? _reinterpretcast_data_830 : _reinterpretcast_data_830;
      _cond_data_838 <= (stream_matmul_29_constant_11_data)? _reinterpretcast_data_837 : _reinterpretcast_data_837;
      _cond_data_845 <= (stream_matmul_29_constant_13_data)? _reinterpretcast_data_844 : _reinterpretcast_data_844;
      _eq_data_851 <= stream_matmul_29_constant_1_data == 1'sd0;
      _eq_data_855 <= stream_matmul_29_constant_2_data == 1'sd0;
      _eq_data_891 <= stream_matmul_29_constant_18_data == 1'sd0;
      _eq_data_894 <= stream_matmul_29_constant_18_data == 2'sd1;
      __delay_data_1417 <= stream_matmul_29_source_19_data;
      __delay_data_1419 <= _pointer_data_870;
      __delay_data_1422 <= stream_matmul_29_constant_15_data;
      __delay_data_1423 <= _reinterpretcast_data_869;
      __delay_data_1429 <= stream_matmul_29_constant_16_data;
      __delay_data_1444 <= stream_matmul_29_constant_0_data;
      __delay_data_1482 <= stream_matmul_29_constant_17_data;
      _cond_data_853 <= (_eq_data_851)? __delay_data_1417 : 1'sd0;
      _plus_data_875 <= _cond_data_831 + __delay_data_1422;
      _plus_data_880 <= _cond_data_838 + __delay_data_1429;
      _plus_data_885 <= _cond_data_845 + __delay_data_1482;
      __delay_data_1418 <= _eq_data_855;
      __delay_data_1420 <= __delay_data_1419;
      __delay_data_1424 <= __delay_data_1423;
      __delay_data_1445 <= __delay_data_1444;
      __delay_data_1460 <= _cond_data_817;
      __delay_data_1483 <= _cond_data_824;
      __delay_data_1529 <= _eq_data_891;
      __delay_data_1565 <= _eq_data_894;
      _cond_data_857 <= (__delay_data_1418)? _cond_data_853 : 1'sd0;
      __delay_data_1421 <= __delay_data_1420;
      __delay_data_1425 <= __delay_data_1424;
      __delay_data_1427 <= _plus_data_875;
      __delay_data_1430 <= _plus_data_880;
      __delay_data_1446 <= __delay_data_1445;
      __delay_data_1461 <= __delay_data_1460;
      __delay_data_1484 <= __delay_data_1483;
      __delay_data_1506 <= _plus_data_885;
      __delay_data_1530 <= __delay_data_1529;
      __delay_data_1566 <= __delay_data_1565;
      _cond_data_873 <= (__delay_data_1421)? 1'sd0 : _reinterpretcast_data_863;
      __delay_data_1426 <= __delay_data_1425;
      __delay_data_1428 <= __delay_data_1427;
      __delay_data_1431 <= __delay_data_1430;
      __delay_data_1447 <= __delay_data_1446;
      __delay_data_1462 <= __delay_data_1461;
      __delay_data_1485 <= __delay_data_1484;
      __delay_data_1507 <= __delay_data_1506;
      __delay_data_1531 <= __delay_data_1530;
      __delay_data_1567 <= __delay_data_1566;
      __delay_data_1432 <= __delay_data_1431;
      __delay_data_1448 <= __delay_data_1447;
      __delay_data_1463 <= __delay_data_1462;
      __delay_data_1486 <= __delay_data_1485;
      __delay_data_1508 <= __delay_data_1507;
      __delay_data_1532 <= __delay_data_1531;
      __delay_data_1568 <= __delay_data_1567;
      __delay_data_1433 <= __delay_data_1432;
      __delay_data_1449 <= __delay_data_1448;
      __delay_data_1464 <= __delay_data_1463;
      __delay_data_1487 <= __delay_data_1486;
      __delay_data_1509 <= __delay_data_1508;
      __delay_data_1533 <= __delay_data_1532;
      __delay_data_1569 <= __delay_data_1568;
      __delay_data_1434 <= __delay_data_1433;
      __delay_data_1450 <= __delay_data_1449;
      __delay_data_1465 <= __delay_data_1464;
      __delay_data_1488 <= __delay_data_1487;
      __delay_data_1510 <= __delay_data_1509;
      __delay_data_1534 <= __delay_data_1533;
      __delay_data_1570 <= __delay_data_1569;
      __delay_data_1435 <= __delay_data_1434;
      __delay_data_1451 <= __delay_data_1450;
      __delay_data_1466 <= __delay_data_1465;
      __delay_data_1489 <= __delay_data_1488;
      __delay_data_1511 <= __delay_data_1510;
      __delay_data_1535 <= __delay_data_1534;
      __delay_data_1571 <= __delay_data_1570;
      __delay_data_1436 <= __delay_data_1435;
      __delay_data_1452 <= __delay_data_1451;
      __delay_data_1467 <= __delay_data_1466;
      __delay_data_1490 <= __delay_data_1489;
      __delay_data_1512 <= __delay_data_1511;
      __delay_data_1536 <= __delay_data_1535;
      __delay_data_1572 <= __delay_data_1571;
      __delay_data_1437 <= __delay_data_1436;
      __delay_data_1453 <= __delay_data_1452;
      __delay_data_1468 <= __delay_data_1467;
      __delay_data_1491 <= __delay_data_1490;
      __delay_data_1513 <= __delay_data_1512;
      __delay_data_1537 <= __delay_data_1536;
      __delay_data_1573 <= __delay_data_1572;
      __delay_data_1438 <= __delay_data_1437;
      __delay_data_1454 <= __delay_data_1453;
      __delay_data_1469 <= __delay_data_1468;
      __delay_data_1492 <= __delay_data_1491;
      __delay_data_1514 <= __delay_data_1513;
      __delay_data_1538 <= __delay_data_1537;
      __delay_data_1574 <= __delay_data_1573;
      __delay_data_1439 <= __delay_data_1438;
      __delay_data_1455 <= __delay_data_1454;
      __delay_data_1470 <= __delay_data_1469;
      __delay_data_1493 <= __delay_data_1492;
      __delay_data_1515 <= __delay_data_1514;
      __delay_data_1539 <= __delay_data_1538;
      __delay_data_1575 <= __delay_data_1574;
      __delay_data_1440 <= __delay_data_1439;
      __delay_data_1456 <= __delay_data_1455;
      __delay_data_1471 <= __delay_data_1470;
      __delay_data_1494 <= __delay_data_1493;
      __delay_data_1516 <= __delay_data_1515;
      __delay_data_1540 <= __delay_data_1539;
      __delay_data_1576 <= __delay_data_1575;
      __substreamoutput_data_876 <= mul_4_z_data;
      __delay_data_1441 <= __delay_data_1440;
      __delay_data_1457 <= __delay_data_1456;
      __delay_data_1472 <= __delay_data_1471;
      __delay_data_1495 <= __delay_data_1494;
      __delay_data_1517 <= __delay_data_1516;
      __delay_data_1541 <= __delay_data_1540;
      __delay_data_1577 <= __delay_data_1576;
      __delay_data_1442 <= __delay_data_1441;
      __delay_data_1458 <= __delay_data_1457;
      __delay_data_1473 <= __delay_data_1472;
      __delay_data_1496 <= __delay_data_1495;
      __delay_data_1518 <= __delay_data_1517;
      __delay_data_1542 <= __delay_data_1541;
      __delay_data_1578 <= __delay_data_1577;
      __substreamoutput_data_878 <= add_tree_1_sum_data;
      __delay_data_1443 <= __delay_data_1442;
      __delay_data_1459 <= __delay_data_1458;
      __delay_data_1474 <= __delay_data_1473;
      __delay_data_1497 <= __delay_data_1496;
      __delay_data_1519 <= __delay_data_1518;
      __delay_data_1543 <= __delay_data_1542;
      __delay_data_1579 <= __delay_data_1578;
      __delay_data_1475 <= __delay_data_1474;
      __delay_data_1498 <= __delay_data_1497;
      __delay_data_1520 <= __delay_data_1519;
      __delay_data_1544 <= __delay_data_1543;
      __delay_data_1580 <= __delay_data_1579;
      __delay_data_1476 <= __delay_data_1475;
      __delay_data_1499 <= __delay_data_1498;
      __delay_data_1521 <= __delay_data_1520;
      __delay_data_1545 <= __delay_data_1544;
      __delay_data_1581 <= __delay_data_1580;
      __delay_data_1477 <= __delay_data_1476;
      __delay_data_1500 <= __delay_data_1499;
      __delay_data_1522 <= __delay_data_1521;
      __delay_data_1546 <= __delay_data_1545;
      __delay_data_1582 <= __delay_data_1581;
      __delay_data_1478 <= __delay_data_1477;
      __delay_data_1501 <= __delay_data_1500;
      __delay_data_1523 <= __delay_data_1522;
      __delay_data_1547 <= __delay_data_1546;
      __delay_data_1583 <= __delay_data_1582;
      __delay_data_1479 <= __delay_data_1478;
      __delay_data_1502 <= __delay_data_1501;
      __delay_data_1524 <= __delay_data_1523;
      __delay_data_1548 <= __delay_data_1547;
      __delay_data_1584 <= __delay_data_1583;
      __delay_data_1480 <= __delay_data_1479;
      __delay_data_1503 <= __delay_data_1502;
      __delay_data_1525 <= __delay_data_1524;
      __delay_data_1549 <= __delay_data_1548;
      __delay_data_1585 <= __delay_data_1584;
      __substreamoutput_data_881 <= acc_0_sum_data;
      __substreamoutput_data_882 <= acc_0_valid_data;
      __delay_data_1481 <= __delay_data_1480;
      __delay_data_1504 <= __delay_data_1503;
      __delay_data_1526 <= __delay_data_1525;
      __delay_data_1550 <= __delay_data_1549;
      __delay_data_1586 <= __delay_data_1585;
      _plus_data_883 <= __substreamoutput_data_881 + __delay_data_1481;
      __delay_data_1505 <= __delay_data_1504;
      __delay_data_1527 <= __delay_data_1526;
      __delay_data_1551 <= __delay_data_1550;
      __delay_data_1587 <= __delay_data_1586;
      __delay_data_1602 <= __substreamoutput_data_882;
      __delay_data_1552 <= __delay_data_1551;
      __delay_data_1588 <= __delay_data_1587;
      __delay_data_1603 <= __delay_data_1602;
      __delay_data_1553 <= __delay_data_1552;
      __delay_data_1589 <= __delay_data_1588;
      __delay_data_1604 <= __delay_data_1603;
      __delay_data_1554 <= __delay_data_1553;
      __delay_data_1590 <= __delay_data_1589;
      __delay_data_1605 <= __delay_data_1604;
      __delay_data_1555 <= __delay_data_1554;
      __delay_data_1591 <= __delay_data_1590;
      __delay_data_1606 <= __delay_data_1605;
      __delay_data_1556 <= __delay_data_1555;
      __delay_data_1592 <= __delay_data_1591;
      __delay_data_1607 <= __delay_data_1606;
      __delay_data_1557 <= __delay_data_1556;
      __delay_data_1593 <= __delay_data_1592;
      __delay_data_1608 <= __delay_data_1607;
      __delay_data_1558 <= __delay_data_1557;
      __delay_data_1594 <= __delay_data_1593;
      __delay_data_1609 <= __delay_data_1608;
      __delay_data_1559 <= __delay_data_1558;
      __delay_data_1595 <= __delay_data_1594;
      __delay_data_1610 <= __delay_data_1609;
      __delay_data_1560 <= __delay_data_1559;
      __delay_data_1596 <= __delay_data_1595;
      __delay_data_1611 <= __delay_data_1610;
      __substreamoutput_data_886 <= mul_rshift_clip_3_z_data;
      __delay_data_1561 <= __delay_data_1560;
      __delay_data_1597 <= __delay_data_1596;
      __delay_data_1612 <= __delay_data_1611;
      _greaterthan_data_888 <= __substreamoutput_data_886 > 1'sd0;
      __delay_data_1528 <= __substreamoutput_data_886;
      __delay_data_1562 <= __delay_data_1561;
      __delay_data_1598 <= __delay_data_1597;
      __delay_data_1613 <= __delay_data_1612;
      _cond_data_890 <= (_greaterthan_data_888)? __delay_data_1528 : 1'sd0;
      __delay_data_1563 <= __delay_data_1562;
      __delay_data_1564 <= __delay_data_1528;
      __delay_data_1599 <= __delay_data_1598;
      __delay_data_1614 <= __delay_data_1613;
      _cond_data_893 <= (__delay_data_1563)? _cond_data_890 : __delay_data_1564;
      __delay_data_1600 <= __delay_data_1599;
      __delay_data_1601 <= __delay_data_1564;
      __delay_data_1615 <= __delay_data_1614;
      _cond_data_896 <= (__delay_data_1600)? __delay_data_1601 : _cond_data_893;
      __delay_data_1616 <= __delay_data_1615;
      _set_flag_1163 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1163 <= 1;
      end 
      if(_set_flag_1163) begin
        _stream_matmul_29_constant_0_next_constant_data <= cparam_matmul_29_stream_reduce_size;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_796 <= _stream_matmul_29_constant_0_next_constant_data;
      end 
      _set_flag_1164 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1164 <= 1;
      end 
      if(_set_flag_1164) begin
        _stream_matmul_29_constant_1_next_constant_data <= matmul_29_col_select;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_797 <= _stream_matmul_29_constant_1_next_constant_data;
      end 
      _set_flag_1165 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1165 <= 1;
      end 
      if(_set_flag_1165) begin
        _stream_matmul_29_constant_2_next_constant_data <= matmul_29_row_select_buf;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_798 <= _stream_matmul_29_constant_2_next_constant_data;
      end 
      _set_flag_1166 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1166 <= 1;
      end 
      if(_set_flag_1166) begin
        _stream_matmul_29_constant_3_next_constant_data <= matmul_29_stream_pad_masks;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_799 <= _stream_matmul_29_constant_3_next_constant_data;
      end 
      _set_flag_1167 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1167 <= 1;
      end 
      if(_set_flag_1167) begin
        _stream_matmul_29_constant_4_next_constant_data <= cparam_matmul_29_stream_omit_mask;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_800 <= _stream_matmul_29_constant_4_next_constant_data;
      end 
      _set_flag_1168 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1168 <= 1;
      end 
      if(_set_flag_1168) begin
        _stream_matmul_29_constant_5_next_constant_data <= cparam_matmul_29_bias_scala;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_811 <= _stream_matmul_29_constant_5_next_constant_data;
      end 
      _set_flag_1169 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1169 <= 1;
      end 
      if(_set_flag_1169) begin
        _stream_matmul_29_source_6_source_mode <= 3'b10;
        _stream_matmul_29_source_6_source_offset <= (cparam_matmul_29_bias_num == 1)? 0 : matmul_29_och_count_buf;
      end 
      if(_set_flag_1169) begin
        _source_stream_matmul_29_source_6_pat_size_0 <= cparam_matmul_29_stream_reduce_size;
        _source_stream_matmul_29_source_6_pat_stride_0 <= 0;
      end 
      if(_set_flag_1169) begin
        _source_stream_matmul_29_source_6_pat_size_1 <= matmul_29_next_stream_num_ops;
        _source_stream_matmul_29_source_6_pat_stride_1 <= (cparam_matmul_29_bias_num == 1)? 0 : 1;
      end 
      if(_set_flag_1169) begin
        _source_stream_matmul_29_source_6_pat_size_2 <= 1;
        _source_stream_matmul_29_source_6_pat_stride_2 <= 0;
      end 
      if(_set_flag_1169) begin
        _source_stream_matmul_29_source_6_pat_size_3 <= 1;
        _source_stream_matmul_29_source_6_pat_stride_3 <= 0;
      end 
      if(_set_flag_1169) begin
        _stream_matmul_29_source_6_source_ram_sel <= 1;
      end 
      __tmp_1178_1 <= _tmp_1178;
      if(__tmp_1178_1) begin
        _stream_matmul_29_source_6_source_ram_rvalid <= 1;
      end 
      if(_stream_matmul_29_source_6_source_ram_rvalid) begin
        __variable_wdata_812 <= _stream_matmul_29_source_6_source_ram_rdata;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _stream_matmul_29_source_6_idle <= 0;
        _stream_matmul_29_source_6_source_offset_buf <= _stream_matmul_29_source_6_source_offset;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_count_0 <= _source_stream_matmul_29_source_6_pat_size_0 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_count_1 <= _source_stream_matmul_29_source_6_pat_size_1 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_count_2 <= _source_stream_matmul_29_source_6_pat_size_2 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_count_3 <= _source_stream_matmul_29_source_6_pat_size_3 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_size_buf_0 <= _source_stream_matmul_29_source_6_pat_size_0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_size_buf_1 <= _source_stream_matmul_29_source_6_pat_size_1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_size_buf_2 <= _source_stream_matmul_29_source_6_pat_size_2;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_size_buf_3 <= _source_stream_matmul_29_source_6_pat_size_3;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_stride_buf_0 <= _source_stream_matmul_29_source_6_pat_stride_0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_stride_buf_1 <= _source_stream_matmul_29_source_6_pat_stride_1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_stride_buf_2 <= _source_stream_matmul_29_source_6_pat_stride_2;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_6_pat_stride_buf_3 <= _source_stream_matmul_29_source_6_pat_stride_3;
      end 
      if(_stream_matmul_29_source_6_source_pat_fsm_0 == 1) begin
        _stream_matmul_29_source_6_source_ram_raddr <= _stream_matmul_29_source_6_source_pat_all_offset;
        _stream_matmul_29_source_6_source_ram_renable <= 1;
      end 
      if(_stream_matmul_29_source_6_source_pat_fsm_0 == 1) begin
        _source_stream_matmul_29_source_6_pat_cur_offset_0 <= _source_stream_matmul_29_source_6_pat_cur_offset_0 + _source_stream_matmul_29_source_6_pat_stride_buf_0;
        _source_stream_matmul_29_source_6_pat_count_0 <= _source_stream_matmul_29_source_6_pat_count_0 - 1;
      end 
      if((_stream_matmul_29_source_6_source_pat_fsm_0 == 1) && (_source_stream_matmul_29_source_6_pat_count_0 == 0)) begin
        _source_stream_matmul_29_source_6_pat_cur_offset_0 <= 0;
        _source_stream_matmul_29_source_6_pat_count_0 <= _source_stream_matmul_29_source_6_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_29_source_6_source_pat_fsm_0 == 1) && (_source_stream_matmul_29_source_6_pat_count_0 == 0)) begin
        _source_stream_matmul_29_source_6_pat_cur_offset_1 <= _source_stream_matmul_29_source_6_pat_cur_offset_1 + _source_stream_matmul_29_source_6_pat_stride_buf_1;
        _source_stream_matmul_29_source_6_pat_count_1 <= _source_stream_matmul_29_source_6_pat_count_1 - 1;
      end 
      if((_stream_matmul_29_source_6_source_pat_fsm_0 == 1) && (_source_stream_matmul_29_source_6_pat_count_0 == 0) && (_source_stream_matmul_29_source_6_pat_count_1 == 0)) begin
        _source_stream_matmul_29_source_6_pat_cur_offset_1 <= 0;
        _source_stream_matmul_29_source_6_pat_count_1 <= _source_stream_matmul_29_source_6_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_29_source_6_source_pat_fsm_0 == 1) && ((_source_stream_matmul_29_source_6_pat_count_0 == 0) && (_source_stream_matmul_29_source_6_pat_count_1 == 0))) begin
        _source_stream_matmul_29_source_6_pat_cur_offset_2 <= _source_stream_matmul_29_source_6_pat_cur_offset_2 + _source_stream_matmul_29_source_6_pat_stride_buf_2;
        _source_stream_matmul_29_source_6_pat_count_2 <= _source_stream_matmul_29_source_6_pat_count_2 - 1;
      end 
      if((_stream_matmul_29_source_6_source_pat_fsm_0 == 1) && ((_source_stream_matmul_29_source_6_pat_count_0 == 0) && (_source_stream_matmul_29_source_6_pat_count_1 == 0)) && (_source_stream_matmul_29_source_6_pat_count_2 == 0)) begin
        _source_stream_matmul_29_source_6_pat_cur_offset_2 <= 0;
        _source_stream_matmul_29_source_6_pat_count_2 <= _source_stream_matmul_29_source_6_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_29_source_6_source_pat_fsm_0 == 1) && ((_source_stream_matmul_29_source_6_pat_count_0 == 0) && (_source_stream_matmul_29_source_6_pat_count_1 == 0) && (_source_stream_matmul_29_source_6_pat_count_2 == 0))) begin
        _source_stream_matmul_29_source_6_pat_cur_offset_3 <= _source_stream_matmul_29_source_6_pat_cur_offset_3 + _source_stream_matmul_29_source_6_pat_stride_buf_3;
        _source_stream_matmul_29_source_6_pat_count_3 <= _source_stream_matmul_29_source_6_pat_count_3 - 1;
      end 
      if((_stream_matmul_29_source_6_source_pat_fsm_0 == 1) && ((_source_stream_matmul_29_source_6_pat_count_0 == 0) && (_source_stream_matmul_29_source_6_pat_count_1 == 0) && (_source_stream_matmul_29_source_6_pat_count_2 == 0)) && (_source_stream_matmul_29_source_6_pat_count_3 == 0)) begin
        _source_stream_matmul_29_source_6_pat_cur_offset_3 <= 0;
        _source_stream_matmul_29_source_6_pat_count_3 <= _source_stream_matmul_29_source_6_pat_size_buf_3 - 1;
      end 
      if(_stream_matmul_29_source_6_source_pat_fsm_0 == 2) begin
        _stream_matmul_29_source_6_source_ram_renable <= 0;
        _stream_matmul_29_source_6_idle <= 1;
      end 
      _set_flag_1179 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1179 <= 1;
      end 
      if(_set_flag_1179) begin
        _stream_matmul_29_constant_7_next_constant_data <= cparam_matmul_29_scale_scala;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_818 <= _stream_matmul_29_constant_7_next_constant_data;
      end 
      _set_flag_1180 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1180 <= 1;
      end 
      if(_set_flag_1180) begin
        _stream_matmul_29_source_8_source_mode <= 3'b10;
        _stream_matmul_29_source_8_source_offset <= (cparam_matmul_29_scale_num == 1)? 0 : matmul_29_och_count_buf;
      end 
      if(_set_flag_1180) begin
        _source_stream_matmul_29_source_8_pat_size_0 <= cparam_matmul_29_stream_reduce_size;
        _source_stream_matmul_29_source_8_pat_stride_0 <= 0;
      end 
      if(_set_flag_1180) begin
        _source_stream_matmul_29_source_8_pat_size_1 <= matmul_29_next_stream_num_ops;
        _source_stream_matmul_29_source_8_pat_stride_1 <= (cparam_matmul_29_scale_num == 1)? 0 : 1;
      end 
      if(_set_flag_1180) begin
        _source_stream_matmul_29_source_8_pat_size_2 <= 1;
        _source_stream_matmul_29_source_8_pat_stride_2 <= 0;
      end 
      if(_set_flag_1180) begin
        _source_stream_matmul_29_source_8_pat_size_3 <= 1;
        _source_stream_matmul_29_source_8_pat_stride_3 <= 0;
      end 
      if(_set_flag_1180) begin
        _stream_matmul_29_source_8_source_ram_sel <= 2;
      end 
      __tmp_1189_1 <= _tmp_1189;
      if(__tmp_1189_1) begin
        _stream_matmul_29_source_8_source_ram_rvalid <= 1;
      end 
      if(_stream_matmul_29_source_8_source_ram_rvalid) begin
        __variable_wdata_819 <= _stream_matmul_29_source_8_source_ram_rdata;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _stream_matmul_29_source_8_idle <= 0;
        _stream_matmul_29_source_8_source_offset_buf <= _stream_matmul_29_source_8_source_offset;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_count_0 <= _source_stream_matmul_29_source_8_pat_size_0 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_count_1 <= _source_stream_matmul_29_source_8_pat_size_1 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_count_2 <= _source_stream_matmul_29_source_8_pat_size_2 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_count_3 <= _source_stream_matmul_29_source_8_pat_size_3 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_size_buf_0 <= _source_stream_matmul_29_source_8_pat_size_0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_size_buf_1 <= _source_stream_matmul_29_source_8_pat_size_1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_size_buf_2 <= _source_stream_matmul_29_source_8_pat_size_2;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_size_buf_3 <= _source_stream_matmul_29_source_8_pat_size_3;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_stride_buf_0 <= _source_stream_matmul_29_source_8_pat_stride_0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_stride_buf_1 <= _source_stream_matmul_29_source_8_pat_stride_1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_stride_buf_2 <= _source_stream_matmul_29_source_8_pat_stride_2;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_8_pat_stride_buf_3 <= _source_stream_matmul_29_source_8_pat_stride_3;
      end 
      if(_stream_matmul_29_source_8_source_pat_fsm_1 == 1) begin
        _stream_matmul_29_source_8_source_ram_raddr <= _stream_matmul_29_source_8_source_pat_all_offset;
        _stream_matmul_29_source_8_source_ram_renable <= 1;
      end 
      if(_stream_matmul_29_source_8_source_pat_fsm_1 == 1) begin
        _source_stream_matmul_29_source_8_pat_cur_offset_0 <= _source_stream_matmul_29_source_8_pat_cur_offset_0 + _source_stream_matmul_29_source_8_pat_stride_buf_0;
        _source_stream_matmul_29_source_8_pat_count_0 <= _source_stream_matmul_29_source_8_pat_count_0 - 1;
      end 
      if((_stream_matmul_29_source_8_source_pat_fsm_1 == 1) && (_source_stream_matmul_29_source_8_pat_count_0 == 0)) begin
        _source_stream_matmul_29_source_8_pat_cur_offset_0 <= 0;
        _source_stream_matmul_29_source_8_pat_count_0 <= _source_stream_matmul_29_source_8_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_29_source_8_source_pat_fsm_1 == 1) && (_source_stream_matmul_29_source_8_pat_count_0 == 0)) begin
        _source_stream_matmul_29_source_8_pat_cur_offset_1 <= _source_stream_matmul_29_source_8_pat_cur_offset_1 + _source_stream_matmul_29_source_8_pat_stride_buf_1;
        _source_stream_matmul_29_source_8_pat_count_1 <= _source_stream_matmul_29_source_8_pat_count_1 - 1;
      end 
      if((_stream_matmul_29_source_8_source_pat_fsm_1 == 1) && (_source_stream_matmul_29_source_8_pat_count_0 == 0) && (_source_stream_matmul_29_source_8_pat_count_1 == 0)) begin
        _source_stream_matmul_29_source_8_pat_cur_offset_1 <= 0;
        _source_stream_matmul_29_source_8_pat_count_1 <= _source_stream_matmul_29_source_8_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_29_source_8_source_pat_fsm_1 == 1) && ((_source_stream_matmul_29_source_8_pat_count_0 == 0) && (_source_stream_matmul_29_source_8_pat_count_1 == 0))) begin
        _source_stream_matmul_29_source_8_pat_cur_offset_2 <= _source_stream_matmul_29_source_8_pat_cur_offset_2 + _source_stream_matmul_29_source_8_pat_stride_buf_2;
        _source_stream_matmul_29_source_8_pat_count_2 <= _source_stream_matmul_29_source_8_pat_count_2 - 1;
      end 
      if((_stream_matmul_29_source_8_source_pat_fsm_1 == 1) && ((_source_stream_matmul_29_source_8_pat_count_0 == 0) && (_source_stream_matmul_29_source_8_pat_count_1 == 0)) && (_source_stream_matmul_29_source_8_pat_count_2 == 0)) begin
        _source_stream_matmul_29_source_8_pat_cur_offset_2 <= 0;
        _source_stream_matmul_29_source_8_pat_count_2 <= _source_stream_matmul_29_source_8_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_29_source_8_source_pat_fsm_1 == 1) && ((_source_stream_matmul_29_source_8_pat_count_0 == 0) && (_source_stream_matmul_29_source_8_pat_count_1 == 0) && (_source_stream_matmul_29_source_8_pat_count_2 == 0))) begin
        _source_stream_matmul_29_source_8_pat_cur_offset_3 <= _source_stream_matmul_29_source_8_pat_cur_offset_3 + _source_stream_matmul_29_source_8_pat_stride_buf_3;
        _source_stream_matmul_29_source_8_pat_count_3 <= _source_stream_matmul_29_source_8_pat_count_3 - 1;
      end 
      if((_stream_matmul_29_source_8_source_pat_fsm_1 == 1) && ((_source_stream_matmul_29_source_8_pat_count_0 == 0) && (_source_stream_matmul_29_source_8_pat_count_1 == 0) && (_source_stream_matmul_29_source_8_pat_count_2 == 0)) && (_source_stream_matmul_29_source_8_pat_count_3 == 0)) begin
        _source_stream_matmul_29_source_8_pat_cur_offset_3 <= 0;
        _source_stream_matmul_29_source_8_pat_count_3 <= _source_stream_matmul_29_source_8_pat_size_buf_3 - 1;
      end 
      if(_stream_matmul_29_source_8_source_pat_fsm_1 == 2) begin
        _stream_matmul_29_source_8_source_ram_renable <= 0;
        _stream_matmul_29_source_8_idle <= 1;
      end 
      _set_flag_1190 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1190 <= 1;
      end 
      if(_set_flag_1190) begin
        _stream_matmul_29_constant_9_next_constant_data <= 1;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_825 <= _stream_matmul_29_constant_9_next_constant_data;
      end 
      _set_flag_1191 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1191 <= 1;
      end 
      if(_set_flag_1191) begin
        _stream_matmul_29_source_10_source_mode <= 3'b0;
        _stream_matmul_29_source_10_source_empty_data <= 0;
      end 
      if(_stream_matmul_29_start && !(|(_stream_matmul_29_source_10_source_mode & 3'b0))) begin
        _stream_matmul_29_source_10_idle <= 1;
      end 
      if(_stream_matmul_29_start && !(|(_stream_matmul_29_source_10_source_mode & 3'b0))) begin
        __variable_wdata_826 <= _stream_matmul_29_source_10_source_empty_data;
      end 
      _set_flag_1192 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1192 <= 1;
      end 
      if(_set_flag_1192) begin
        _stream_matmul_29_constant_11_next_constant_data <= 1;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_832 <= _stream_matmul_29_constant_11_next_constant_data;
      end 
      _set_flag_1193 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1193 <= 1;
      end 
      if(_set_flag_1193) begin
        _stream_matmul_29_source_12_source_mode <= 3'b0;
        _stream_matmul_29_source_12_source_empty_data <= 0;
      end 
      if(_stream_matmul_29_start && !(|(_stream_matmul_29_source_12_source_mode & 3'b0))) begin
        _stream_matmul_29_source_12_idle <= 1;
      end 
      if(_stream_matmul_29_start && !(|(_stream_matmul_29_source_12_source_mode & 3'b0))) begin
        __variable_wdata_833 <= _stream_matmul_29_source_12_source_empty_data;
      end 
      _set_flag_1194 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1194 <= 1;
      end 
      if(_set_flag_1194) begin
        _stream_matmul_29_constant_13_next_constant_data <= 1;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_839 <= _stream_matmul_29_constant_13_next_constant_data;
      end 
      _set_flag_1195 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1195 <= 1;
      end 
      if(_set_flag_1195) begin
        _stream_matmul_29_source_14_source_mode <= 3'b0;
        _stream_matmul_29_source_14_source_empty_data <= 0;
      end 
      if(_stream_matmul_29_start && !(|(_stream_matmul_29_source_14_source_mode & 3'b0))) begin
        _stream_matmul_29_source_14_idle <= 1;
      end 
      if(_stream_matmul_29_start && !(|(_stream_matmul_29_source_14_source_mode & 3'b0))) begin
        __variable_wdata_840 <= _stream_matmul_29_source_14_source_empty_data;
      end 
      _set_flag_1196 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1196 <= 1;
      end 
      if(_set_flag_1196) begin
        _stream_matmul_29_constant_15_next_constant_data <= cparam_matmul_29_cshamt_mul_value;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_846 <= _stream_matmul_29_constant_15_next_constant_data;
      end 
      _set_flag_1197 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1197 <= 1;
      end 
      if(_set_flag_1197) begin
        _stream_matmul_29_constant_16_next_constant_data <= cparam_matmul_29_cshamt_sum_value;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_847 <= _stream_matmul_29_constant_16_next_constant_data;
      end 
      _set_flag_1198 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1198 <= 1;
      end 
      if(_set_flag_1198) begin
        _stream_matmul_29_constant_17_next_constant_data <= cparam_matmul_29_cshamt_out_value;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_848 <= _stream_matmul_29_constant_17_next_constant_data;
      end 
      _set_flag_1199 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1199 <= 1;
      end 
      if(_set_flag_1199) begin
        _stream_matmul_29_constant_18_next_constant_data <= cparam_matmul_29_act_func_index;
      end 
      if(_stream_matmul_29_start) begin
        __variable_wdata_849 <= _stream_matmul_29_constant_18_next_constant_data;
      end 
      _set_flag_1200 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1200 <= 1;
      end 
      if(_set_flag_1200) begin
        _stream_matmul_29_source_19_source_mode <= 3'b10;
        _stream_matmul_29_source_19_source_offset <= matmul_29_stream_act_local_0 + matmul_29_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_1200) begin
        _source_stream_matmul_29_source_19_pat_size_0 <= cparam_matmul_29_stream_reduce_size;
        _source_stream_matmul_29_source_19_pat_stride_0 <= 1;
      end 
      if(_set_flag_1200) begin
        _source_stream_matmul_29_source_19_pat_size_1 <= matmul_29_next_stream_num_ops;
        _source_stream_matmul_29_source_19_pat_stride_1 <= 0;
      end 
      if(_set_flag_1200) begin
        _source_stream_matmul_29_source_19_pat_size_2 <= 1;
        _source_stream_matmul_29_source_19_pat_stride_2 <= 0;
      end 
      if(_set_flag_1200) begin
        _source_stream_matmul_29_source_19_pat_size_3 <= 1;
        _source_stream_matmul_29_source_19_pat_stride_3 <= 0;
      end 
      if(_set_flag_1200) begin
        _stream_matmul_29_source_19_source_ram_sel <= 3;
      end 
      __tmp_1209_1 <= _tmp_1209;
      if(__tmp_1209_1) begin
        _stream_matmul_29_source_19_source_ram_rvalid <= 1;
      end 
      if(_stream_matmul_29_source_19_source_ram_rvalid) begin
        __variable_wdata_850 <= _stream_matmul_29_source_19_source_ram_rdata;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _stream_matmul_29_source_19_idle <= 0;
        _stream_matmul_29_source_19_source_offset_buf <= _stream_matmul_29_source_19_source_offset;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_count_0 <= _source_stream_matmul_29_source_19_pat_size_0 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_count_1 <= _source_stream_matmul_29_source_19_pat_size_1 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_count_2 <= _source_stream_matmul_29_source_19_pat_size_2 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_count_3 <= _source_stream_matmul_29_source_19_pat_size_3 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_size_buf_0 <= _source_stream_matmul_29_source_19_pat_size_0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_size_buf_1 <= _source_stream_matmul_29_source_19_pat_size_1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_size_buf_2 <= _source_stream_matmul_29_source_19_pat_size_2;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_size_buf_3 <= _source_stream_matmul_29_source_19_pat_size_3;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_stride_buf_0 <= _source_stream_matmul_29_source_19_pat_stride_0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_stride_buf_1 <= _source_stream_matmul_29_source_19_pat_stride_1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_stride_buf_2 <= _source_stream_matmul_29_source_19_pat_stride_2;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_19_pat_stride_buf_3 <= _source_stream_matmul_29_source_19_pat_stride_3;
      end 
      if(_stream_matmul_29_source_19_source_pat_fsm_2 == 1) begin
        _stream_matmul_29_source_19_source_ram_raddr <= _stream_matmul_29_source_19_source_pat_all_offset;
        _stream_matmul_29_source_19_source_ram_renable <= 1;
      end 
      if(_stream_matmul_29_source_19_source_pat_fsm_2 == 1) begin
        _source_stream_matmul_29_source_19_pat_cur_offset_0 <= _source_stream_matmul_29_source_19_pat_cur_offset_0 + _source_stream_matmul_29_source_19_pat_stride_buf_0;
        _source_stream_matmul_29_source_19_pat_count_0 <= _source_stream_matmul_29_source_19_pat_count_0 - 1;
      end 
      if((_stream_matmul_29_source_19_source_pat_fsm_2 == 1) && (_source_stream_matmul_29_source_19_pat_count_0 == 0)) begin
        _source_stream_matmul_29_source_19_pat_cur_offset_0 <= 0;
        _source_stream_matmul_29_source_19_pat_count_0 <= _source_stream_matmul_29_source_19_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_29_source_19_source_pat_fsm_2 == 1) && (_source_stream_matmul_29_source_19_pat_count_0 == 0)) begin
        _source_stream_matmul_29_source_19_pat_cur_offset_1 <= _source_stream_matmul_29_source_19_pat_cur_offset_1 + _source_stream_matmul_29_source_19_pat_stride_buf_1;
        _source_stream_matmul_29_source_19_pat_count_1 <= _source_stream_matmul_29_source_19_pat_count_1 - 1;
      end 
      if((_stream_matmul_29_source_19_source_pat_fsm_2 == 1) && (_source_stream_matmul_29_source_19_pat_count_0 == 0) && (_source_stream_matmul_29_source_19_pat_count_1 == 0)) begin
        _source_stream_matmul_29_source_19_pat_cur_offset_1 <= 0;
        _source_stream_matmul_29_source_19_pat_count_1 <= _source_stream_matmul_29_source_19_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_29_source_19_source_pat_fsm_2 == 1) && ((_source_stream_matmul_29_source_19_pat_count_0 == 0) && (_source_stream_matmul_29_source_19_pat_count_1 == 0))) begin
        _source_stream_matmul_29_source_19_pat_cur_offset_2 <= _source_stream_matmul_29_source_19_pat_cur_offset_2 + _source_stream_matmul_29_source_19_pat_stride_buf_2;
        _source_stream_matmul_29_source_19_pat_count_2 <= _source_stream_matmul_29_source_19_pat_count_2 - 1;
      end 
      if((_stream_matmul_29_source_19_source_pat_fsm_2 == 1) && ((_source_stream_matmul_29_source_19_pat_count_0 == 0) && (_source_stream_matmul_29_source_19_pat_count_1 == 0)) && (_source_stream_matmul_29_source_19_pat_count_2 == 0)) begin
        _source_stream_matmul_29_source_19_pat_cur_offset_2 <= 0;
        _source_stream_matmul_29_source_19_pat_count_2 <= _source_stream_matmul_29_source_19_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_29_source_19_source_pat_fsm_2 == 1) && ((_source_stream_matmul_29_source_19_pat_count_0 == 0) && (_source_stream_matmul_29_source_19_pat_count_1 == 0) && (_source_stream_matmul_29_source_19_pat_count_2 == 0))) begin
        _source_stream_matmul_29_source_19_pat_cur_offset_3 <= _source_stream_matmul_29_source_19_pat_cur_offset_3 + _source_stream_matmul_29_source_19_pat_stride_buf_3;
        _source_stream_matmul_29_source_19_pat_count_3 <= _source_stream_matmul_29_source_19_pat_count_3 - 1;
      end 
      if((_stream_matmul_29_source_19_source_pat_fsm_2 == 1) && ((_source_stream_matmul_29_source_19_pat_count_0 == 0) && (_source_stream_matmul_29_source_19_pat_count_1 == 0) && (_source_stream_matmul_29_source_19_pat_count_2 == 0)) && (_source_stream_matmul_29_source_19_pat_count_3 == 0)) begin
        _source_stream_matmul_29_source_19_pat_cur_offset_3 <= 0;
        _source_stream_matmul_29_source_19_pat_count_3 <= _source_stream_matmul_29_source_19_pat_size_buf_3 - 1;
      end 
      if(_stream_matmul_29_source_19_source_pat_fsm_2 == 2) begin
        _stream_matmul_29_source_19_source_ram_renable <= 0;
        _stream_matmul_29_source_19_idle <= 1;
      end 
      _set_flag_1210 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1210 <= 1;
      end 
      if(_set_flag_1210) begin
        _stream_matmul_29_source_20_source_mode <= 3'b10;
        _stream_matmul_29_source_20_source_offset <= matmul_29_filter_page_comp_offset_buf;
      end 
      if(_set_flag_1210) begin
        _source_stream_matmul_29_source_20_pat_size_0 <= cparam_matmul_29_stream_reduce_size;
        _source_stream_matmul_29_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_1210) begin
        _source_stream_matmul_29_source_20_pat_size_1 <= matmul_29_next_stream_num_ops;
        _source_stream_matmul_29_source_20_pat_stride_1 <= cparam_matmul_29_stream_aligned_reduce_size;
      end 
      if(_set_flag_1210) begin
        _source_stream_matmul_29_source_20_pat_size_2 <= 1;
        _source_stream_matmul_29_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_1210) begin
        _source_stream_matmul_29_source_20_pat_size_3 <= 1;
        _source_stream_matmul_29_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_1210) begin
        _stream_matmul_29_source_20_source_ram_sel <= 4;
      end 
      __tmp_1223_1 <= _tmp_1223;
      if(__tmp_1223_1) begin
        _stream_matmul_29_source_20_source_ram_rvalid <= 1;
      end 
      if(_stream_matmul_29_source_20_source_ram_rvalid) begin
        __variable_wdata_864 <= _stream_matmul_29_source_20_source_ram_rdata;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _stream_matmul_29_source_20_idle <= 0;
        _stream_matmul_29_source_20_source_offset_buf <= _stream_matmul_29_source_20_source_offset;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_count_0 <= _source_stream_matmul_29_source_20_pat_size_0 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_count_1 <= _source_stream_matmul_29_source_20_pat_size_1 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_count_2 <= _source_stream_matmul_29_source_20_pat_size_2 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_count_3 <= _source_stream_matmul_29_source_20_pat_size_3 - 1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_size_buf_0 <= _source_stream_matmul_29_source_20_pat_size_0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_size_buf_1 <= _source_stream_matmul_29_source_20_pat_size_1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_size_buf_2 <= _source_stream_matmul_29_source_20_pat_size_2;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_size_buf_3 <= _source_stream_matmul_29_source_20_pat_size_3;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_stride_buf_0 <= _source_stream_matmul_29_source_20_pat_stride_0;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_stride_buf_1 <= _source_stream_matmul_29_source_20_pat_stride_1;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_stride_buf_2 <= _source_stream_matmul_29_source_20_pat_stride_2;
      end 
      if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
        _source_stream_matmul_29_source_20_pat_stride_buf_3 <= _source_stream_matmul_29_source_20_pat_stride_3;
      end 
      if(_stream_matmul_29_source_20_source_pat_fsm_3 == 1) begin
        _stream_matmul_29_source_20_source_ram_raddr <= _stream_matmul_29_source_20_source_pat_all_offset;
        _stream_matmul_29_source_20_source_ram_renable <= 1;
      end 
      if(_stream_matmul_29_source_20_source_pat_fsm_3 == 1) begin
        _source_stream_matmul_29_source_20_pat_cur_offset_0 <= _source_stream_matmul_29_source_20_pat_cur_offset_0 + _source_stream_matmul_29_source_20_pat_stride_buf_0;
        _source_stream_matmul_29_source_20_pat_count_0 <= _source_stream_matmul_29_source_20_pat_count_0 - 1;
      end 
      if((_stream_matmul_29_source_20_source_pat_fsm_3 == 1) && (_source_stream_matmul_29_source_20_pat_count_0 == 0)) begin
        _source_stream_matmul_29_source_20_pat_cur_offset_0 <= 0;
        _source_stream_matmul_29_source_20_pat_count_0 <= _source_stream_matmul_29_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_29_source_20_source_pat_fsm_3 == 1) && (_source_stream_matmul_29_source_20_pat_count_0 == 0)) begin
        _source_stream_matmul_29_source_20_pat_cur_offset_1 <= _source_stream_matmul_29_source_20_pat_cur_offset_1 + _source_stream_matmul_29_source_20_pat_stride_buf_1;
        _source_stream_matmul_29_source_20_pat_count_1 <= _source_stream_matmul_29_source_20_pat_count_1 - 1;
      end 
      if((_stream_matmul_29_source_20_source_pat_fsm_3 == 1) && (_source_stream_matmul_29_source_20_pat_count_0 == 0) && (_source_stream_matmul_29_source_20_pat_count_1 == 0)) begin
        _source_stream_matmul_29_source_20_pat_cur_offset_1 <= 0;
        _source_stream_matmul_29_source_20_pat_count_1 <= _source_stream_matmul_29_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_29_source_20_source_pat_fsm_3 == 1) && ((_source_stream_matmul_29_source_20_pat_count_0 == 0) && (_source_stream_matmul_29_source_20_pat_count_1 == 0))) begin
        _source_stream_matmul_29_source_20_pat_cur_offset_2 <= _source_stream_matmul_29_source_20_pat_cur_offset_2 + _source_stream_matmul_29_source_20_pat_stride_buf_2;
        _source_stream_matmul_29_source_20_pat_count_2 <= _source_stream_matmul_29_source_20_pat_count_2 - 1;
      end 
      if((_stream_matmul_29_source_20_source_pat_fsm_3 == 1) && ((_source_stream_matmul_29_source_20_pat_count_0 == 0) && (_source_stream_matmul_29_source_20_pat_count_1 == 0)) && (_source_stream_matmul_29_source_20_pat_count_2 == 0)) begin
        _source_stream_matmul_29_source_20_pat_cur_offset_2 <= 0;
        _source_stream_matmul_29_source_20_pat_count_2 <= _source_stream_matmul_29_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_29_source_20_source_pat_fsm_3 == 1) && ((_source_stream_matmul_29_source_20_pat_count_0 == 0) && (_source_stream_matmul_29_source_20_pat_count_1 == 0) && (_source_stream_matmul_29_source_20_pat_count_2 == 0))) begin
        _source_stream_matmul_29_source_20_pat_cur_offset_3 <= _source_stream_matmul_29_source_20_pat_cur_offset_3 + _source_stream_matmul_29_source_20_pat_stride_buf_3;
        _source_stream_matmul_29_source_20_pat_count_3 <= _source_stream_matmul_29_source_20_pat_count_3 - 1;
      end 
      if((_stream_matmul_29_source_20_source_pat_fsm_3 == 1) && ((_source_stream_matmul_29_source_20_pat_count_0 == 0) && (_source_stream_matmul_29_source_20_pat_count_1 == 0) && (_source_stream_matmul_29_source_20_pat_count_2 == 0)) && (_source_stream_matmul_29_source_20_pat_count_3 == 0)) begin
        _source_stream_matmul_29_source_20_pat_cur_offset_3 <= 0;
        _source_stream_matmul_29_source_20_pat_count_3 <= _source_stream_matmul_29_source_20_pat_size_buf_3 - 1;
      end 
      if(_stream_matmul_29_source_20_source_pat_fsm_3 == 2) begin
        _stream_matmul_29_source_20_source_ram_renable <= 0;
        _stream_matmul_29_source_20_idle <= 1;
      end 
      _set_flag_1224 <= 0;
      if(matmul_29_comp_fsm == 3) begin
        _set_flag_1224 <= 1;
      end 
      __stream_matmul_29_sink_21_sink_offset_0_1 <= matmul_29_stream_out_local + matmul_29_out_page_comp_offset_buf;
      __stream_matmul_29_sink_21_sink_size_1_1 <= matmul_29_next_stream_num_ops;
      __stream_seq_16_cond_2_1 <= _set_flag_1224;
      __set_flag_1224_1 <= _set_flag_1224;
      __set_flag_1224_2 <= __set_flag_1224_1;
      __set_flag_1224_3 <= __set_flag_1224_2;
      __set_flag_1224_4 <= __set_flag_1224_3;
      __set_flag_1224_5 <= __set_flag_1224_4;
      __set_flag_1224_6 <= __set_flag_1224_5;
      __set_flag_1224_7 <= __set_flag_1224_6;
      __set_flag_1224_8 <= __set_flag_1224_7;
      __set_flag_1224_9 <= __set_flag_1224_8;
      __set_flag_1224_10 <= __set_flag_1224_9;
      __set_flag_1224_11 <= __set_flag_1224_10;
      __set_flag_1224_12 <= __set_flag_1224_11;
      __set_flag_1224_13 <= __set_flag_1224_12;
      __set_flag_1224_14 <= __set_flag_1224_13;
      __set_flag_1224_15 <= __set_flag_1224_14;
      __set_flag_1224_16 <= __set_flag_1224_15;
      __set_flag_1224_17 <= __set_flag_1224_16;
      __set_flag_1224_18 <= __set_flag_1224_17;
      __set_flag_1224_19 <= __set_flag_1224_18;
      __set_flag_1224_20 <= __set_flag_1224_19;
      __set_flag_1224_21 <= __set_flag_1224_20;
      __set_flag_1224_22 <= __set_flag_1224_21;
      __set_flag_1224_23 <= __set_flag_1224_22;
      __set_flag_1224_24 <= __set_flag_1224_23;
      __set_flag_1224_25 <= __set_flag_1224_24;
      __set_flag_1224_26 <= __set_flag_1224_25;
      __set_flag_1224_27 <= __set_flag_1224_26;
      __set_flag_1224_28 <= __set_flag_1224_27;
      __set_flag_1224_29 <= __set_flag_1224_28;
      __set_flag_1224_30 <= __set_flag_1224_29;
      __set_flag_1224_31 <= __set_flag_1224_30;
      __set_flag_1224_32 <= __set_flag_1224_31;
      __set_flag_1224_33 <= __set_flag_1224_32;
      __set_flag_1224_34 <= __set_flag_1224_33;
      __set_flag_1224_35 <= __set_flag_1224_34;
      __set_flag_1224_36 <= __set_flag_1224_35;
      __set_flag_1224_37 <= __set_flag_1224_36;
      __set_flag_1224_38 <= __set_flag_1224_37;
      __set_flag_1224_39 <= __set_flag_1224_38;
      __set_flag_1224_40 <= __set_flag_1224_39;
      __set_flag_1224_41 <= __set_flag_1224_40;
      if(__set_flag_1224_41) begin
        _stream_matmul_29_sink_21_sink_ram_sel <= 5;
      end 
      __stream_matmul_29_start_1 <= _stream_matmul_29_start;
      __stream_matmul_29_start_2 <= __stream_matmul_29_start_1;
      __stream_matmul_29_start_3 <= __stream_matmul_29_start_2;
      __stream_matmul_29_start_4 <= __stream_matmul_29_start_3;
      __stream_matmul_29_start_5 <= __stream_matmul_29_start_4;
      __stream_matmul_29_start_6 <= __stream_matmul_29_start_5;
      __stream_matmul_29_start_7 <= __stream_matmul_29_start_6;
      __stream_matmul_29_start_8 <= __stream_matmul_29_start_7;
      __stream_matmul_29_start_9 <= __stream_matmul_29_start_8;
      __stream_matmul_29_start_10 <= __stream_matmul_29_start_9;
      __stream_matmul_29_start_11 <= __stream_matmul_29_start_10;
      __stream_matmul_29_start_12 <= __stream_matmul_29_start_11;
      __stream_matmul_29_start_13 <= __stream_matmul_29_start_12;
      __stream_matmul_29_start_14 <= __stream_matmul_29_start_13;
      __stream_matmul_29_start_15 <= __stream_matmul_29_start_14;
      __stream_matmul_29_start_16 <= __stream_matmul_29_start_15;
      __stream_matmul_29_start_17 <= __stream_matmul_29_start_16;
      __stream_matmul_29_start_18 <= __stream_matmul_29_start_17;
      __stream_matmul_29_start_19 <= __stream_matmul_29_start_18;
      __stream_matmul_29_start_20 <= __stream_matmul_29_start_19;
      __stream_matmul_29_start_21 <= __stream_matmul_29_start_20;
      __stream_matmul_29_start_22 <= __stream_matmul_29_start_21;
      __stream_matmul_29_start_23 <= __stream_matmul_29_start_22;
      __stream_matmul_29_start_24 <= __stream_matmul_29_start_23;
      __stream_matmul_29_start_25 <= __stream_matmul_29_start_24;
      __stream_matmul_29_start_26 <= __stream_matmul_29_start_25;
      __stream_matmul_29_start_27 <= __stream_matmul_29_start_26;
      __stream_matmul_29_start_28 <= __stream_matmul_29_start_27;
      __stream_matmul_29_start_29 <= __stream_matmul_29_start_28;
      __stream_matmul_29_start_30 <= __stream_matmul_29_start_29;
      __stream_matmul_29_start_31 <= __stream_matmul_29_start_30;
      __stream_matmul_29_start_32 <= __stream_matmul_29_start_31;
      __stream_matmul_29_start_33 <= __stream_matmul_29_start_32;
      __stream_matmul_29_start_34 <= __stream_matmul_29_start_33;
      __stream_matmul_29_start_35 <= __stream_matmul_29_start_34;
      __stream_matmul_29_start_36 <= __stream_matmul_29_start_35;
      __stream_matmul_29_start_37 <= __stream_matmul_29_start_36;
      __stream_matmul_29_start_38 <= __stream_matmul_29_start_37;
      __stream_matmul_29_start_39 <= __stream_matmul_29_start_38;
      __stream_matmul_29_start_40 <= __stream_matmul_29_start_39;
      __stream_matmul_29_start_41 <= __stream_matmul_29_start_40;
      __stream_matmul_29_start_42 <= __stream_matmul_29_start_41;
      if(__stream_matmul_29_start_42 && _stream_matmul_29_sink_21_sink_mode & 3'b1) begin
        _stream_matmul_29_sink_21_sink_waddr <= _stream_matmul_29_sink_21_sink_offset - _stream_matmul_29_sink_21_sink_stride;
        _stream_matmul_29_sink_21_sink_count <= _stream_matmul_29_sink_21_sink_size;
        _stream_matmul_29_sink_21_sink_offset_buf <= _stream_matmul_29_sink_21_sink_offset;
        _stream_matmul_29_sink_21_sink_stride_buf <= _stream_matmul_29_sink_21_sink_stride;
      end 
      if((_stream_matmul_29_sink_21_sink_fsm_4 == 1) && stream_matmul_29_sink_22_data) begin
        _stream_matmul_29_sink_21_sink_waddr <= _stream_matmul_29_sink_21_sink_waddr + _stream_matmul_29_sink_21_sink_stride_buf;
        _stream_matmul_29_sink_21_sink_wdata <= stream_matmul_29_sink_21_data;
        _stream_matmul_29_sink_21_sink_wenable <= 1;
        _stream_matmul_29_sink_21_sink_count <= _stream_matmul_29_sink_21_sink_count - 1;
      end 
      __tmp_1227_1 <= _tmp_1227;
      __tmp_1227_2 <= __tmp_1227_1;
      __tmp_1227_3 <= __tmp_1227_2;
      __tmp_1227_4 <= __tmp_1227_3;
      __tmp_1227_5 <= __tmp_1227_4;
      __tmp_1229_1 <= _tmp_1229;
      __tmp_1229_2 <= __tmp_1229_1;
      __tmp_1229_3 <= __tmp_1229_2;
      __tmp_1229_4 <= __tmp_1229_3;
      __tmp_1229_5 <= __tmp_1229_4;
      __tmp_1229_6 <= __tmp_1229_5;
      __tmp_1229_7 <= __tmp_1229_6;
      __tmp_1229_8 <= __tmp_1229_7;
      __tmp_1231_1 <= _tmp_1231;
      __tmp_1231_2 <= __tmp_1231_1;
      __tmp_1231_3 <= __tmp_1231_2;
      __tmp_1231_4 <= __tmp_1231_3;
      __tmp_1231_5 <= __tmp_1231_4;
      __tmp_1231_6 <= __tmp_1231_5;
      __tmp_1231_7 <= __tmp_1231_6;
      __tmp_1231_8 <= __tmp_1231_7;
      __tmp_1233_1 <= _tmp_1233;
      __tmp_1233_2 <= __tmp_1233_1;
      __tmp_1233_3 <= __tmp_1233_2;
      __tmp_1233_4 <= __tmp_1233_3;
      __tmp_1233_5 <= __tmp_1233_4;
      __tmp_1233_6 <= __tmp_1233_5;
      __tmp_1233_7 <= __tmp_1233_6;
      __tmp_1233_8 <= __tmp_1233_7;
      __tmp_1235_1 <= _tmp_1235;
      __tmp_1235_2 <= __tmp_1235_1;
      __tmp_1235_3 <= __tmp_1235_2;
      __tmp_1235_4 <= __tmp_1235_3;
      __tmp_1235_5 <= __tmp_1235_4;
      __tmp_1235_6 <= __tmp_1235_5;
      __tmp_1235_7 <= __tmp_1235_6;
      __tmp_1235_8 <= __tmp_1235_7;
      __tmp_1235_9 <= __tmp_1235_8;
      __tmp_1235_10 <= __tmp_1235_9;
      __tmp_1235_11 <= __tmp_1235_10;
      __tmp_1235_12 <= __tmp_1235_11;
      __tmp_1235_13 <= __tmp_1235_12;
      __tmp_1235_14 <= __tmp_1235_13;
      __tmp_1235_15 <= __tmp_1235_14;
      __tmp_1235_16 <= __tmp_1235_15;
      __tmp_1235_17 <= __tmp_1235_16;
      __tmp_1235_18 <= __tmp_1235_17;
      __tmp_1237_1 <= _tmp_1237;
      __tmp_1237_2 <= __tmp_1237_1;
      __tmp_1237_3 <= __tmp_1237_2;
      __tmp_1237_4 <= __tmp_1237_3;
      __tmp_1237_5 <= __tmp_1237_4;
      __tmp_1237_6 <= __tmp_1237_5;
      __tmp_1237_7 <= __tmp_1237_6;
      __tmp_1237_8 <= __tmp_1237_7;
      __tmp_1237_9 <= __tmp_1237_8;
      __tmp_1237_10 <= __tmp_1237_9;
      __tmp_1237_11 <= __tmp_1237_10;
      __tmp_1237_12 <= __tmp_1237_11;
      __tmp_1237_13 <= __tmp_1237_12;
      __tmp_1237_14 <= __tmp_1237_13;
      __tmp_1237_15 <= __tmp_1237_14;
      __tmp_1237_16 <= __tmp_1237_15;
      __tmp_1237_17 <= __tmp_1237_16;
      __tmp_1237_18 <= __tmp_1237_17;
      __tmp_1237_19 <= __tmp_1237_18;
      __tmp_1237_20 <= __tmp_1237_19;
      __tmp_1237_21 <= __tmp_1237_20;
      __tmp_1237_22 <= __tmp_1237_21;
      __tmp_1239_1 <= _tmp_1239;
      __tmp_1239_2 <= __tmp_1239_1;
      __tmp_1239_3 <= __tmp_1239_2;
      __tmp_1239_4 <= __tmp_1239_3;
      __tmp_1239_5 <= __tmp_1239_4;
      __tmp_1239_6 <= __tmp_1239_5;
      __tmp_1239_7 <= __tmp_1239_6;
      __tmp_1239_8 <= __tmp_1239_7;
      __tmp_1239_9 <= __tmp_1239_8;
      __tmp_1239_10 <= __tmp_1239_9;
      __tmp_1239_11 <= __tmp_1239_10;
      __tmp_1239_12 <= __tmp_1239_11;
      __tmp_1239_13 <= __tmp_1239_12;
      __tmp_1239_14 <= __tmp_1239_13;
      __tmp_1239_15 <= __tmp_1239_14;
      __tmp_1239_16 <= __tmp_1239_15;
      __tmp_1239_17 <= __tmp_1239_16;
      __tmp_1239_18 <= __tmp_1239_17;
      __tmp_1239_19 <= __tmp_1239_18;
      __tmp_1239_20 <= __tmp_1239_19;
      __tmp_1241_1 <= _tmp_1241;
      __tmp_1241_2 <= __tmp_1241_1;
      __tmp_1241_3 <= __tmp_1241_2;
      __tmp_1241_4 <= __tmp_1241_3;
      __tmp_1241_5 <= __tmp_1241_4;
      __tmp_1241_6 <= __tmp_1241_5;
      __tmp_1241_7 <= __tmp_1241_6;
      __tmp_1241_8 <= __tmp_1241_7;
      __tmp_1241_9 <= __tmp_1241_8;
      __tmp_1241_10 <= __tmp_1241_9;
      __tmp_1241_11 <= __tmp_1241_10;
      __tmp_1241_12 <= __tmp_1241_11;
      __tmp_1241_13 <= __tmp_1241_12;
      __tmp_1241_14 <= __tmp_1241_13;
      __tmp_1241_15 <= __tmp_1241_14;
      __tmp_1241_16 <= __tmp_1241_15;
      __tmp_1241_17 <= __tmp_1241_16;
      __tmp_1241_18 <= __tmp_1241_17;
      __tmp_1241_19 <= __tmp_1241_18;
      __tmp_1241_20 <= __tmp_1241_19;
      __tmp_1243_1 <= _tmp_1243;
      __tmp_1243_2 <= __tmp_1243_1;
      __tmp_1243_3 <= __tmp_1243_2;
      __tmp_1243_4 <= __tmp_1243_3;
      __tmp_1243_5 <= __tmp_1243_4;
      __tmp_1243_6 <= __tmp_1243_5;
      __tmp_1243_7 <= __tmp_1243_6;
      __tmp_1243_8 <= __tmp_1243_7;
      __tmp_1243_9 <= __tmp_1243_8;
      __tmp_1243_10 <= __tmp_1243_9;
      __tmp_1243_11 <= __tmp_1243_10;
      __tmp_1243_12 <= __tmp_1243_11;
      __tmp_1243_13 <= __tmp_1243_12;
      __tmp_1243_14 <= __tmp_1243_13;
      __tmp_1243_15 <= __tmp_1243_14;
      __tmp_1243_16 <= __tmp_1243_15;
      __tmp_1243_17 <= __tmp_1243_16;
      __tmp_1243_18 <= __tmp_1243_17;
      __tmp_1243_19 <= __tmp_1243_18;
      __tmp_1243_20 <= __tmp_1243_19;
      __tmp_1245_1 <= _tmp_1245;
      __tmp_1245_2 <= __tmp_1245_1;
      __tmp_1245_3 <= __tmp_1245_2;
      __tmp_1245_4 <= __tmp_1245_3;
      __tmp_1245_5 <= __tmp_1245_4;
      __tmp_1245_6 <= __tmp_1245_5;
      __tmp_1245_7 <= __tmp_1245_6;
      __tmp_1245_8 <= __tmp_1245_7;
      __tmp_1245_9 <= __tmp_1245_8;
      __tmp_1245_10 <= __tmp_1245_9;
      __tmp_1245_11 <= __tmp_1245_10;
      __tmp_1245_12 <= __tmp_1245_11;
      __tmp_1245_13 <= __tmp_1245_12;
      __tmp_1245_14 <= __tmp_1245_13;
      __tmp_1245_15 <= __tmp_1245_14;
      __tmp_1245_16 <= __tmp_1245_15;
      __tmp_1245_17 <= __tmp_1245_16;
      __tmp_1245_18 <= __tmp_1245_17;
      __tmp_1245_19 <= __tmp_1245_18;
      __tmp_1245_20 <= __tmp_1245_19;
      __tmp_1245_21 <= __tmp_1245_20;
      __tmp_1245_22 <= __tmp_1245_21;
      __tmp_1245_23 <= __tmp_1245_22;
      __tmp_1245_24 <= __tmp_1245_23;
      __tmp_1245_25 <= __tmp_1245_24;
      __tmp_1245_26 <= __tmp_1245_25;
      __tmp_1245_27 <= __tmp_1245_26;
      __tmp_1245_28 <= __tmp_1245_27;
      __tmp_1247_1 <= _tmp_1247;
      __tmp_1247_2 <= __tmp_1247_1;
      __tmp_1247_3 <= __tmp_1247_2;
      __tmp_1247_4 <= __tmp_1247_3;
      __tmp_1247_5 <= __tmp_1247_4;
      __tmp_1247_6 <= __tmp_1247_5;
      __tmp_1247_7 <= __tmp_1247_6;
      __tmp_1247_8 <= __tmp_1247_7;
      __tmp_1247_9 <= __tmp_1247_8;
      __tmp_1247_10 <= __tmp_1247_9;
      __tmp_1247_11 <= __tmp_1247_10;
      __tmp_1247_12 <= __tmp_1247_11;
      __tmp_1247_13 <= __tmp_1247_12;
      __tmp_1247_14 <= __tmp_1247_13;
      __tmp_1247_15 <= __tmp_1247_14;
      __tmp_1247_16 <= __tmp_1247_15;
      __tmp_1247_17 <= __tmp_1247_16;
      __tmp_1247_18 <= __tmp_1247_17;
      __tmp_1247_19 <= __tmp_1247_18;
      __tmp_1247_20 <= __tmp_1247_19;
      __tmp_1247_21 <= __tmp_1247_20;
      __tmp_1247_22 <= __tmp_1247_21;
      __tmp_1247_23 <= __tmp_1247_22;
      __tmp_1247_24 <= __tmp_1247_23;
      __tmp_1247_25 <= __tmp_1247_24;
      __tmp_1247_26 <= __tmp_1247_25;
      __tmp_1247_27 <= __tmp_1247_26;
      __tmp_1247_28 <= __tmp_1247_27;
      __tmp_1249_1 <= _tmp_1249;
      __tmp_1249_2 <= __tmp_1249_1;
      __tmp_1249_3 <= __tmp_1249_2;
      __tmp_1249_4 <= __tmp_1249_3;
      __tmp_1249_5 <= __tmp_1249_4;
      __tmp_1249_6 <= __tmp_1249_5;
      __tmp_1249_7 <= __tmp_1249_6;
      __tmp_1249_8 <= __tmp_1249_7;
      __tmp_1249_9 <= __tmp_1249_8;
      __tmp_1249_10 <= __tmp_1249_9;
      __tmp_1249_11 <= __tmp_1249_10;
      __tmp_1249_12 <= __tmp_1249_11;
      __tmp_1249_13 <= __tmp_1249_12;
      __tmp_1249_14 <= __tmp_1249_13;
      __tmp_1249_15 <= __tmp_1249_14;
      __tmp_1249_16 <= __tmp_1249_15;
      __tmp_1249_17 <= __tmp_1249_16;
      __tmp_1249_18 <= __tmp_1249_17;
      __tmp_1249_19 <= __tmp_1249_18;
      __tmp_1249_20 <= __tmp_1249_19;
      __tmp_1249_21 <= __tmp_1249_20;
      __tmp_1249_22 <= __tmp_1249_21;
      __tmp_1249_23 <= __tmp_1249_22;
      __tmp_1249_24 <= __tmp_1249_23;
      __tmp_1249_25 <= __tmp_1249_24;
      __tmp_1249_26 <= __tmp_1249_25;
      __tmp_1249_27 <= __tmp_1249_26;
      __tmp_1249_28 <= __tmp_1249_27;
      __tmp_1251_1 <= _tmp_1251;
      __tmp_1253_1 <= _tmp_1253;
      __tmp_1253_2 <= __tmp_1253_1;
      __tmp_1253_3 <= __tmp_1253_2;
      __tmp_1253_4 <= __tmp_1253_3;
      __tmp_1253_5 <= __tmp_1253_4;
      __tmp_1255_1 <= _tmp_1255;
      __tmp_1255_2 <= __tmp_1255_1;
      __tmp_1255_3 <= __tmp_1255_2;
      __tmp_1255_4 <= __tmp_1255_3;
      __tmp_1255_5 <= __tmp_1255_4;
      __tmp_1257_1 <= _tmp_1257;
      __tmp_1257_2 <= __tmp_1257_1;
      __tmp_1257_3 <= __tmp_1257_2;
      __tmp_1257_4 <= __tmp_1257_3;
      __tmp_1257_5 <= __tmp_1257_4;
      __tmp_1265_1 <= _tmp_1265;
      __tmp_1265_2 <= __tmp_1265_1;
      __tmp_1265_3 <= __tmp_1265_2;
      __tmp_1265_4 <= __tmp_1265_3;
      __tmp_1265_5 <= __tmp_1265_4;
      __tmp_1265_6 <= __tmp_1265_5;
      __tmp_1265_7 <= __tmp_1265_6;
      __tmp_1265_8 <= __tmp_1265_7;
      __tmp_1265_9 <= __tmp_1265_8;
      __tmp_1265_10 <= __tmp_1265_9;
      __tmp_1265_11 <= __tmp_1265_10;
      __tmp_1265_12 <= __tmp_1265_11;
      __tmp_1265_13 <= __tmp_1265_12;
      __tmp_1265_14 <= __tmp_1265_13;
      __tmp_1265_15 <= __tmp_1265_14;
      __tmp_1273_1 <= _tmp_1273;
      __tmp_1273_2 <= __tmp_1273_1;
      __tmp_1273_3 <= __tmp_1273_2;
      __tmp_1273_4 <= __tmp_1273_3;
      __tmp_1273_5 <= __tmp_1273_4;
      __tmp_1273_6 <= __tmp_1273_5;
      __tmp_1273_7 <= __tmp_1273_6;
      __tmp_1273_8 <= __tmp_1273_7;
      __tmp_1273_9 <= __tmp_1273_8;
      __tmp_1273_10 <= __tmp_1273_9;
      __tmp_1273_11 <= __tmp_1273_10;
      __tmp_1273_12 <= __tmp_1273_11;
      __tmp_1273_13 <= __tmp_1273_12;
      __tmp_1273_14 <= __tmp_1273_13;
      __tmp_1273_15 <= __tmp_1273_14;
      __tmp_1273_16 <= __tmp_1273_15;
      __tmp_1273_17 <= __tmp_1273_16;
      __tmp_1273_18 <= __tmp_1273_17;
      __tmp_1275_1 <= _tmp_1275;
      __tmp_1275_2 <= __tmp_1275_1;
      __tmp_1275_3 <= __tmp_1275_2;
      __tmp_1275_4 <= __tmp_1275_3;
      __tmp_1275_5 <= __tmp_1275_4;
      __tmp_1275_6 <= __tmp_1275_5;
      __tmp_1275_7 <= __tmp_1275_6;
      __tmp_1275_8 <= __tmp_1275_7;
      __tmp_1275_9 <= __tmp_1275_8;
      __tmp_1275_10 <= __tmp_1275_9;
      __tmp_1275_11 <= __tmp_1275_10;
      __tmp_1275_12 <= __tmp_1275_11;
      __tmp_1275_13 <= __tmp_1275_12;
      __tmp_1275_14 <= __tmp_1275_13;
      __tmp_1275_15 <= __tmp_1275_14;
      __tmp_1275_16 <= __tmp_1275_15;
      __tmp_1275_17 <= __tmp_1275_16;
      __tmp_1277_1 <= _tmp_1277;
      __tmp_1277_2 <= __tmp_1277_1;
      __tmp_1277_3 <= __tmp_1277_2;
      __tmp_1277_4 <= __tmp_1277_3;
      __tmp_1277_5 <= __tmp_1277_4;
      __tmp_1277_6 <= __tmp_1277_5;
      __tmp_1277_7 <= __tmp_1277_6;
      __tmp_1277_8 <= __tmp_1277_7;
      __tmp_1277_9 <= __tmp_1277_8;
      __tmp_1277_10 <= __tmp_1277_9;
      __tmp_1277_11 <= __tmp_1277_10;
      __tmp_1277_12 <= __tmp_1277_11;
      __tmp_1277_13 <= __tmp_1277_12;
      __tmp_1277_14 <= __tmp_1277_13;
      __tmp_1277_15 <= __tmp_1277_14;
      __tmp_1277_16 <= __tmp_1277_15;
      __tmp_1277_17 <= __tmp_1277_16;
      __tmp_1279_1 <= _tmp_1279;
      __tmp_1279_2 <= __tmp_1279_1;
      __tmp_1279_3 <= __tmp_1279_2;
      __tmp_1279_4 <= __tmp_1279_3;
      __tmp_1279_5 <= __tmp_1279_4;
      __tmp_1279_6 <= __tmp_1279_5;
      __tmp_1279_7 <= __tmp_1279_6;
      __tmp_1279_8 <= __tmp_1279_7;
      __tmp_1279_9 <= __tmp_1279_8;
      __tmp_1279_10 <= __tmp_1279_9;
      __tmp_1279_11 <= __tmp_1279_10;
      __tmp_1279_12 <= __tmp_1279_11;
      __tmp_1279_13 <= __tmp_1279_12;
      __tmp_1279_14 <= __tmp_1279_13;
      __tmp_1279_15 <= __tmp_1279_14;
      __tmp_1279_16 <= __tmp_1279_15;
      __tmp_1279_17 <= __tmp_1279_16;
      __tmp_1287_1 <= _tmp_1287;
      __tmp_1287_2 <= __tmp_1287_1;
      __tmp_1287_3 <= __tmp_1287_2;
      __tmp_1287_4 <= __tmp_1287_3;
      __tmp_1287_5 <= __tmp_1287_4;
      __tmp_1287_6 <= __tmp_1287_5;
      __tmp_1287_7 <= __tmp_1287_6;
      __tmp_1287_8 <= __tmp_1287_7;
      __tmp_1287_9 <= __tmp_1287_8;
      __tmp_1287_10 <= __tmp_1287_9;
      __tmp_1287_11 <= __tmp_1287_10;
      __tmp_1287_12 <= __tmp_1287_11;
      __tmp_1287_13 <= __tmp_1287_12;
      __tmp_1287_14 <= __tmp_1287_13;
      __tmp_1287_15 <= __tmp_1287_14;
      __tmp_1287_16 <= __tmp_1287_15;
      __tmp_1287_17 <= __tmp_1287_16;
      __tmp_1287_18 <= __tmp_1287_17;
      __tmp_1287_19 <= __tmp_1287_18;
      __tmp_1287_20 <= __tmp_1287_19;
      __tmp_1287_21 <= __tmp_1287_20;
      __tmp_1287_22 <= __tmp_1287_21;
      __tmp_1287_23 <= __tmp_1287_22;
      __tmp_1287_24 <= __tmp_1287_23;
      __tmp_1287_25 <= __tmp_1287_24;
      __tmp_1289_1 <= _tmp_1289;
      __tmp_1289_2 <= __tmp_1289_1;
      __tmp_1289_3 <= __tmp_1289_2;
      __tmp_1289_4 <= __tmp_1289_3;
      __tmp_1289_5 <= __tmp_1289_4;
      __tmp_1289_6 <= __tmp_1289_5;
      __tmp_1289_7 <= __tmp_1289_6;
      __tmp_1289_8 <= __tmp_1289_7;
      __tmp_1289_9 <= __tmp_1289_8;
      __tmp_1289_10 <= __tmp_1289_9;
      __tmp_1289_11 <= __tmp_1289_10;
      __tmp_1289_12 <= __tmp_1289_11;
      __tmp_1289_13 <= __tmp_1289_12;
      __tmp_1289_14 <= __tmp_1289_13;
      __tmp_1289_15 <= __tmp_1289_14;
      __tmp_1289_16 <= __tmp_1289_15;
      __tmp_1289_17 <= __tmp_1289_16;
      __tmp_1289_18 <= __tmp_1289_17;
      __tmp_1289_19 <= __tmp_1289_18;
      __tmp_1289_20 <= __tmp_1289_19;
      __tmp_1289_21 <= __tmp_1289_20;
      __tmp_1289_22 <= __tmp_1289_21;
      __tmp_1289_23 <= __tmp_1289_22;
      __tmp_1289_24 <= __tmp_1289_23;
      __tmp_1289_25 <= __tmp_1289_24;
      __tmp_1291_1 <= _tmp_1291;
      __tmp_1291_2 <= __tmp_1291_1;
      __tmp_1291_3 <= __tmp_1291_2;
      __tmp_1291_4 <= __tmp_1291_3;
      __tmp_1291_5 <= __tmp_1291_4;
      __tmp_1291_6 <= __tmp_1291_5;
      __tmp_1291_7 <= __tmp_1291_6;
      __tmp_1291_8 <= __tmp_1291_7;
      __tmp_1291_9 <= __tmp_1291_8;
      __tmp_1291_10 <= __tmp_1291_9;
      __tmp_1291_11 <= __tmp_1291_10;
      __tmp_1291_12 <= __tmp_1291_11;
      __tmp_1291_13 <= __tmp_1291_12;
      __tmp_1291_14 <= __tmp_1291_13;
      __tmp_1291_15 <= __tmp_1291_14;
      __tmp_1291_16 <= __tmp_1291_15;
      __tmp_1291_17 <= __tmp_1291_16;
      __tmp_1291_18 <= __tmp_1291_17;
      __tmp_1291_19 <= __tmp_1291_18;
      __tmp_1291_20 <= __tmp_1291_19;
      __tmp_1291_21 <= __tmp_1291_20;
      __tmp_1291_22 <= __tmp_1291_21;
      __tmp_1291_23 <= __tmp_1291_22;
      __tmp_1291_24 <= __tmp_1291_23;
      __tmp_1291_25 <= __tmp_1291_24;
      __tmp_1299_1 <= _tmp_1299;
      __tmp_1299_2 <= __tmp_1299_1;
      __tmp_1299_3 <= __tmp_1299_2;
      __tmp_1299_4 <= __tmp_1299_3;
      __tmp_1299_5 <= __tmp_1299_4;
      __tmp_1299_6 <= __tmp_1299_5;
      __tmp_1299_7 <= __tmp_1299_6;
      __tmp_1299_8 <= __tmp_1299_7;
      __tmp_1299_9 <= __tmp_1299_8;
      __tmp_1299_10 <= __tmp_1299_9;
      __tmp_1299_11 <= __tmp_1299_10;
      __tmp_1299_12 <= __tmp_1299_11;
      __tmp_1299_13 <= __tmp_1299_12;
      __tmp_1299_14 <= __tmp_1299_13;
      __tmp_1299_15 <= __tmp_1299_14;
      __tmp_1299_16 <= __tmp_1299_15;
      __tmp_1299_17 <= __tmp_1299_16;
      __tmp_1299_18 <= __tmp_1299_17;
      __tmp_1299_19 <= __tmp_1299_18;
      __tmp_1299_20 <= __tmp_1299_19;
      __tmp_1299_21 <= __tmp_1299_20;
      __tmp_1299_22 <= __tmp_1299_21;
      __tmp_1299_23 <= __tmp_1299_22;
      __tmp_1299_24 <= __tmp_1299_23;
      __tmp_1299_25 <= __tmp_1299_24;
      __tmp_1299_26 <= __tmp_1299_25;
      __tmp_1299_27 <= __tmp_1299_26;
      __tmp_1299_28 <= __tmp_1299_27;
      __tmp_1299_29 <= __tmp_1299_28;
      __tmp_1299_30 <= __tmp_1299_29;
      __tmp_1299_31 <= __tmp_1299_30;
      __tmp_1299_32 <= __tmp_1299_31;
      __tmp_1299_33 <= __tmp_1299_32;
      __tmp_1299_34 <= __tmp_1299_33;
      __tmp_1299_35 <= __tmp_1299_34;
      __tmp_1299_36 <= __tmp_1299_35;
      __tmp_1299_37 <= __tmp_1299_36;
      __tmp_1299_38 <= __tmp_1299_37;
      __tmp_1299_39 <= __tmp_1299_38;
      __tmp_1299_40 <= __tmp_1299_39;
      __tmp_1299_41 <= __tmp_1299_40;
      __tmp_1299_42 <= __tmp_1299_41;
      __tmp_1301_1 <= _tmp_1301;
      __tmp_1301_2 <= __tmp_1301_1;
      __tmp_1301_3 <= __tmp_1301_2;
      __tmp_1301_4 <= __tmp_1301_3;
      __tmp_1301_5 <= __tmp_1301_4;
      __tmp_1301_6 <= __tmp_1301_5;
      __tmp_1301_7 <= __tmp_1301_6;
      __tmp_1301_8 <= __tmp_1301_7;
      __tmp_1301_9 <= __tmp_1301_8;
      __tmp_1301_10 <= __tmp_1301_9;
      __tmp_1301_11 <= __tmp_1301_10;
      __tmp_1301_12 <= __tmp_1301_11;
      __tmp_1301_13 <= __tmp_1301_12;
      __tmp_1301_14 <= __tmp_1301_13;
      __tmp_1301_15 <= __tmp_1301_14;
      __tmp_1301_16 <= __tmp_1301_15;
      __tmp_1301_17 <= __tmp_1301_16;
      __tmp_1301_18 <= __tmp_1301_17;
      __tmp_1301_19 <= __tmp_1301_18;
      __tmp_1301_20 <= __tmp_1301_19;
      __tmp_1301_21 <= __tmp_1301_20;
      __tmp_1301_22 <= __tmp_1301_21;
      __tmp_1301_23 <= __tmp_1301_22;
      __tmp_1301_24 <= __tmp_1301_23;
      __tmp_1301_25 <= __tmp_1301_24;
      __tmp_1301_26 <= __tmp_1301_25;
      __tmp_1301_27 <= __tmp_1301_26;
      __tmp_1301_28 <= __tmp_1301_27;
      __tmp_1301_29 <= __tmp_1301_28;
      __tmp_1301_30 <= __tmp_1301_29;
      __tmp_1301_31 <= __tmp_1301_30;
      __tmp_1301_32 <= __tmp_1301_31;
      __tmp_1301_33 <= __tmp_1301_32;
      __tmp_1301_34 <= __tmp_1301_33;
      __tmp_1301_35 <= __tmp_1301_34;
      __tmp_1301_36 <= __tmp_1301_35;
      __tmp_1301_37 <= __tmp_1301_36;
      __tmp_1301_38 <= __tmp_1301_37;
      __tmp_1301_39 <= __tmp_1301_38;
      __tmp_1301_40 <= __tmp_1301_39;
      __tmp_1301_41 <= __tmp_1301_40;
      __tmp_1301_42 <= __tmp_1301_41;
      __tmp_1303_1 <= _tmp_1303;
      __tmp_1303_2 <= __tmp_1303_1;
      __tmp_1303_3 <= __tmp_1303_2;
      __tmp_1303_4 <= __tmp_1303_3;
      __tmp_1303_5 <= __tmp_1303_4;
      __tmp_1303_6 <= __tmp_1303_5;
      __tmp_1303_7 <= __tmp_1303_6;
      __tmp_1303_8 <= __tmp_1303_7;
      __tmp_1303_9 <= __tmp_1303_8;
      __tmp_1303_10 <= __tmp_1303_9;
      __tmp_1303_11 <= __tmp_1303_10;
      __tmp_1303_12 <= __tmp_1303_11;
      __tmp_1303_13 <= __tmp_1303_12;
      __tmp_1303_14 <= __tmp_1303_13;
      __tmp_1303_15 <= __tmp_1303_14;
      __tmp_1303_16 <= __tmp_1303_15;
      __tmp_1303_17 <= __tmp_1303_16;
      __tmp_1303_18 <= __tmp_1303_17;
      __tmp_1303_19 <= __tmp_1303_18;
      __tmp_1303_20 <= __tmp_1303_19;
      __tmp_1303_21 <= __tmp_1303_20;
      __tmp_1303_22 <= __tmp_1303_21;
      __tmp_1303_23 <= __tmp_1303_22;
      __tmp_1303_24 <= __tmp_1303_23;
      __tmp_1303_25 <= __tmp_1303_24;
      __tmp_1303_26 <= __tmp_1303_25;
      __tmp_1303_27 <= __tmp_1303_26;
      __tmp_1303_28 <= __tmp_1303_27;
      __tmp_1303_29 <= __tmp_1303_28;
      __tmp_1303_30 <= __tmp_1303_29;
      __tmp_1303_31 <= __tmp_1303_30;
      __tmp_1303_32 <= __tmp_1303_31;
      __tmp_1303_33 <= __tmp_1303_32;
      __tmp_1303_34 <= __tmp_1303_33;
      __tmp_1303_35 <= __tmp_1303_34;
      __tmp_1303_36 <= __tmp_1303_35;
      __tmp_1303_37 <= __tmp_1303_36;
      __tmp_1303_38 <= __tmp_1303_37;
      __tmp_1303_39 <= __tmp_1303_38;
      __tmp_1303_40 <= __tmp_1303_39;
      __tmp_1303_41 <= __tmp_1303_40;
      __tmp_1303_42 <= __tmp_1303_41;
      __tmp_1305_1 <= _tmp_1305;
      __tmp_1305_2 <= __tmp_1305_1;
      __tmp_1305_3 <= __tmp_1305_2;
      __tmp_1305_4 <= __tmp_1305_3;
      __tmp_1305_5 <= __tmp_1305_4;
      __tmp_1305_6 <= __tmp_1305_5;
      __tmp_1305_7 <= __tmp_1305_6;
      __tmp_1305_8 <= __tmp_1305_7;
      __tmp_1305_9 <= __tmp_1305_8;
      __tmp_1305_10 <= __tmp_1305_9;
      __tmp_1305_11 <= __tmp_1305_10;
      __tmp_1305_12 <= __tmp_1305_11;
      __tmp_1305_13 <= __tmp_1305_12;
      __tmp_1305_14 <= __tmp_1305_13;
      __tmp_1305_15 <= __tmp_1305_14;
      __tmp_1305_16 <= __tmp_1305_15;
      __tmp_1305_17 <= __tmp_1305_16;
      __tmp_1305_18 <= __tmp_1305_17;
      __tmp_1305_19 <= __tmp_1305_18;
      __tmp_1305_20 <= __tmp_1305_19;
      __tmp_1305_21 <= __tmp_1305_20;
      __tmp_1305_22 <= __tmp_1305_21;
      __tmp_1305_23 <= __tmp_1305_22;
      __tmp_1305_24 <= __tmp_1305_23;
      __tmp_1305_25 <= __tmp_1305_24;
      __tmp_1305_26 <= __tmp_1305_25;
      __tmp_1305_27 <= __tmp_1305_26;
      __tmp_1305_28 <= __tmp_1305_27;
      __tmp_1305_29 <= __tmp_1305_28;
      __tmp_1305_30 <= __tmp_1305_29;
      __tmp_1305_31 <= __tmp_1305_30;
      __tmp_1305_32 <= __tmp_1305_31;
      __tmp_1305_33 <= __tmp_1305_32;
      __tmp_1305_34 <= __tmp_1305_33;
      __tmp_1305_35 <= __tmp_1305_34;
      __tmp_1305_36 <= __tmp_1305_35;
      __tmp_1305_37 <= __tmp_1305_36;
      __tmp_1305_38 <= __tmp_1305_37;
      __tmp_1305_39 <= __tmp_1305_38;
      __tmp_1305_40 <= __tmp_1305_39;
      __tmp_1305_41 <= __tmp_1305_40;
      __tmp_1305_42 <= __tmp_1305_41;
      __tmp_1307_1 <= _tmp_1307;
      __tmp_1307_2 <= __tmp_1307_1;
      __tmp_1307_3 <= __tmp_1307_2;
      __tmp_1307_4 <= __tmp_1307_3;
      __tmp_1307_5 <= __tmp_1307_4;
      __tmp_1307_6 <= __tmp_1307_5;
      __tmp_1307_7 <= __tmp_1307_6;
      __tmp_1307_8 <= __tmp_1307_7;
      __tmp_1307_9 <= __tmp_1307_8;
      __tmp_1307_10 <= __tmp_1307_9;
      __tmp_1307_11 <= __tmp_1307_10;
      __tmp_1307_12 <= __tmp_1307_11;
      __tmp_1307_13 <= __tmp_1307_12;
      __tmp_1307_14 <= __tmp_1307_13;
      __tmp_1307_15 <= __tmp_1307_14;
      __tmp_1307_16 <= __tmp_1307_15;
      __tmp_1307_17 <= __tmp_1307_16;
      __tmp_1307_18 <= __tmp_1307_17;
      __tmp_1307_19 <= __tmp_1307_18;
      __tmp_1307_20 <= __tmp_1307_19;
      __tmp_1307_21 <= __tmp_1307_20;
      __tmp_1307_22 <= __tmp_1307_21;
      __tmp_1307_23 <= __tmp_1307_22;
      __tmp_1307_24 <= __tmp_1307_23;
      __tmp_1307_25 <= __tmp_1307_24;
      __tmp_1307_26 <= __tmp_1307_25;
      __tmp_1307_27 <= __tmp_1307_26;
      __tmp_1307_28 <= __tmp_1307_27;
      __tmp_1307_29 <= __tmp_1307_28;
      __tmp_1307_30 <= __tmp_1307_29;
      __tmp_1307_31 <= __tmp_1307_30;
      __tmp_1307_32 <= __tmp_1307_31;
      __tmp_1307_33 <= __tmp_1307_32;
      __tmp_1307_34 <= __tmp_1307_33;
      __tmp_1307_35 <= __tmp_1307_34;
      __tmp_1307_36 <= __tmp_1307_35;
      __tmp_1307_37 <= __tmp_1307_36;
      __tmp_1307_38 <= __tmp_1307_37;
    end
  end

  localparam _stream_matmul_29_fsm_1 = 1;
  localparam _stream_matmul_29_fsm_2 = 2;
  localparam _stream_matmul_29_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_29_fsm <= _stream_matmul_29_fsm_init;
      _stream_matmul_29_start <= 0;
      _stream_matmul_29_source_busy <= 0;
      _stream_matmul_29_reduce_reset <= 1;
      _stream_matmul_29_sink_busy <= 0;
      _stream_matmul_29_sink_wait_count <= 0;
      _stream_matmul_29_end_flag <= 0;
      _stream_matmul_29_term_sink <= 0;
    end else begin
      _stream_matmul_29_start <= 0;
      if(__tmp_1227_5) begin
        _stream_matmul_29_reduce_reset <= 0;
      end 
      if(__tmp_1251_1) begin
        _stream_matmul_29_reduce_reset <= 1;
      end 
      if((_stream_matmul_29_sink_wait_count == 1) && !((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) && __tmp_1299_42) begin
        _stream_matmul_29_sink_busy <= 0;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) begin
        _stream_matmul_29_sink_busy <= 1;
      end 
      if(!((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag) && __tmp_1301_42) begin
        _stream_matmul_29_sink_wait_count <= _stream_matmul_29_sink_wait_count - 1;
      end 
      if((_stream_matmul_29_fsm == 0) && _stream_matmul_29_start_flag && !__tmp_1303_42) begin
        _stream_matmul_29_sink_wait_count <= _stream_matmul_29_sink_wait_count + 1;
      end 
      _stream_matmul_29_end_flag <= 0;
      if(__tmp_1305_42) begin
        _stream_matmul_29_end_flag <= 1;
      end 
      _stream_matmul_29_term_sink <= 0;
      if(__tmp_1307_38) begin
        _stream_matmul_29_term_sink <= 1;
      end 
      case(_stream_matmul_29_fsm)
        _stream_matmul_29_fsm_init: begin
          if(_stream_matmul_29_start_flag) begin
            _stream_matmul_29_start <= 1;
            _stream_matmul_29_source_busy <= 1;
          end 
          if(_stream_matmul_29_start_flag) begin
            _stream_matmul_29_fsm <= _stream_matmul_29_fsm_1;
          end 
        end
        _stream_matmul_29_fsm_1: begin
          _stream_matmul_29_fsm <= _stream_matmul_29_fsm_2;
        end
        _stream_matmul_29_fsm_2: begin
          if(_stream_matmul_29_done) begin
            _stream_matmul_29_fsm <= _stream_matmul_29_fsm_3;
          end 
        end
        _stream_matmul_29_fsm_3: begin
          _stream_matmul_29_source_busy <= 0;
          _stream_matmul_29_fsm <= _stream_matmul_29_fsm_init;
        end
      endcase
    end
  end

  localparam main_fsm_1 = 1;
  localparam main_fsm_2 = 2;
  localparam main_fsm_3 = 3;
  localparam main_fsm_4 = 4;
  localparam main_fsm_5 = 5;
  localparam main_fsm_6 = 6;
  localparam main_fsm_7 = 7;
  localparam main_fsm_8 = 8;
  localparam main_fsm_9 = 9;
  localparam main_fsm_10 = 10;
  localparam main_fsm_11 = 11;
  localparam main_fsm_12 = 12;
  localparam main_fsm_13 = 13;
  localparam main_fsm_14 = 14;
  localparam main_fsm_15 = 15;
  localparam main_fsm_16 = 16;
  localparam main_fsm_17 = 17;
  localparam main_fsm_18 = 18;
  localparam main_fsm_19 = 19;
  localparam main_fsm_20 = 20;
  localparam main_fsm_21 = 21;
  localparam main_fsm_22 = 22;
  localparam main_fsm_23 = 23;
  localparam main_fsm_24 = 24;
  localparam main_fsm_25 = 25;
  localparam main_fsm_26 = 26;
  localparam main_fsm_27 = 27;
  localparam main_fsm_28 = 28;
  localparam main_fsm_29 = 29;
  localparam main_fsm_30 = 30;
  localparam main_fsm_31 = 31;
  localparam main_fsm_32 = 32;
  localparam main_fsm_33 = 33;
  localparam main_fsm_34 = 34;
  localparam main_fsm_35 = 35;
  localparam main_fsm_36 = 36;
  localparam main_fsm_37 = 37;
  localparam main_fsm_38 = 38;
  localparam main_fsm_39 = 39;
  localparam main_fsm_40 = 40;
  localparam main_fsm_41 = 41;
  localparam main_fsm_42 = 42;
  localparam main_fsm_43 = 43;
  localparam main_fsm_44 = 44;
  localparam main_fsm_45 = 45;
  localparam main_fsm_46 = 46;
  localparam main_fsm_47 = 47;
  localparam main_fsm_48 = 48;
  localparam main_fsm_49 = 49;
  localparam main_fsm_50 = 50;
  localparam main_fsm_51 = 51;
  localparam main_fsm_52 = 52;
  localparam main_fsm_53 = 53;
  localparam main_fsm_54 = 54;
  localparam main_fsm_55 = 55;
  localparam main_fsm_56 = 56;
  localparam main_fsm_57 = 57;
  localparam main_fsm_58 = 58;
  localparam main_fsm_59 = 59;
  localparam main_fsm_60 = 60;
  localparam main_fsm_61 = 61;
  localparam main_fsm_62 = 62;
  localparam main_fsm_63 = 63;
  localparam main_fsm_64 = 64;
  localparam main_fsm_65 = 65;
  localparam main_fsm_66 = 66;
  localparam main_fsm_67 = 67;
  localparam main_fsm_68 = 68;
  localparam main_fsm_69 = 69;
  localparam main_fsm_70 = 70;
  localparam main_fsm_71 = 71;
  localparam main_fsm_72 = 72;
  localparam main_fsm_73 = 73;
  localparam main_fsm_74 = 74;
  localparam main_fsm_75 = 75;
  localparam main_fsm_76 = 76;
  localparam main_fsm_77 = 77;
  localparam main_fsm_78 = 78;
  localparam main_fsm_79 = 79;
  localparam main_fsm_80 = 80;
  localparam main_fsm_81 = 81;
  localparam main_fsm_82 = 82;
  localparam main_fsm_83 = 83;
  localparam main_fsm_84 = 84;
  localparam main_fsm_85 = 85;
  localparam main_fsm_86 = 86;
  localparam main_fsm_87 = 87;
  localparam main_fsm_88 = 88;
  localparam main_fsm_89 = 89;
  localparam main_fsm_90 = 90;
  localparam main_fsm_91 = 91;
  localparam main_fsm_92 = 92;

  always @(posedge CLK) begin
    if(RST) begin
      main_fsm <= main_fsm_init;
      conv2d_16_objaddr <= 0;
      conv2d_16_arg_objaddr_0 <= 0;
      conv2d_16_arg_objaddr_1 <= 0;
      conv2d_16_arg_objaddr_2 <= 0;
      conv2d_16_arg_objaddr_3 <= 0;
      conv2d_16_control_param_index <= 0;
      max_pool_serial_18_objaddr <= 0;
      max_pool_serial_18_arg_objaddr_0 <= 0;
      max_pool_serial_18_control_param_index <= 0;
      matmul_29_objaddr <= 0;
      matmul_29_arg_objaddr_0 <= 0;
      matmul_29_arg_objaddr_1 <= 0;
      matmul_29_arg_objaddr_2 <= 0;
      matmul_29_arg_objaddr_3 <= 0;
      matmul_29_control_param_index <= 0;
    end else begin
      case(main_fsm)
        main_fsm_init: begin
          if(_saxi_register_4 != 0) begin
            main_fsm <= main_fsm_1;
          end 
        end
        main_fsm_1: begin
          main_fsm <= main_fsm_2;
        end
        main_fsm_2: begin
          main_fsm <= main_fsm_3;
        end
        main_fsm_3: begin
          main_fsm <= main_fsm_4;
        end
        main_fsm_4: begin
          main_fsm <= main_fsm_5;
        end
        main_fsm_5: begin
          conv2d_16_objaddr <= _saxi_register_10;
          main_fsm <= main_fsm_6;
        end
        main_fsm_6: begin
          conv2d_16_arg_objaddr_0 <= _saxi_register_12;
          main_fsm <= main_fsm_7;
        end
        main_fsm_7: begin
          conv2d_16_arg_objaddr_1 <= _saxi_register_13;
          main_fsm <= main_fsm_8;
        end
        main_fsm_8: begin
          conv2d_16_arg_objaddr_2 <= _saxi_register_13 + 576;
          main_fsm <= main_fsm_9;
        end
        main_fsm_9: begin
          conv2d_16_arg_objaddr_3 <= _saxi_register_13 + 640;
          main_fsm <= main_fsm_10;
        end
        main_fsm_10: begin
          conv2d_16_control_param_index <= 0;
          main_fsm <= main_fsm_11;
        end
        main_fsm_11: begin
          main_fsm <= main_fsm_12;
        end
        main_fsm_12: begin
          main_fsm <= main_fsm_13;
        end
        main_fsm_13: begin
          if(control_conv2d_16 == 55) begin
            main_fsm <= main_fsm_14;
          end 
        end
        main_fsm_14: begin
          main_fsm <= main_fsm_15;
        end
        main_fsm_15: begin
          max_pool_serial_18_objaddr <= _saxi_register_10 + 16384;
          main_fsm <= main_fsm_16;
        end
        main_fsm_16: begin
          max_pool_serial_18_arg_objaddr_0 <= _saxi_register_10;
          main_fsm <= main_fsm_17;
        end
        main_fsm_17: begin
          max_pool_serial_18_control_param_index <= 0;
          main_fsm <= main_fsm_18;
        end
        main_fsm_18: begin
          main_fsm <= main_fsm_19;
        end
        main_fsm_19: begin
          main_fsm <= main_fsm_20;
        end
        main_fsm_20: begin
          if(control_max_pool_serial_18 == 25) begin
            main_fsm <= main_fsm_21;
          end 
        end
        main_fsm_21: begin
          main_fsm <= main_fsm_22;
        end
        main_fsm_22: begin
          conv2d_16_objaddr <= _saxi_register_10 + 20480;
          main_fsm <= main_fsm_23;
        end
        main_fsm_23: begin
          conv2d_16_arg_objaddr_0 <= _saxi_register_10 + 16384;
          main_fsm <= main_fsm_24;
        end
        main_fsm_24: begin
          conv2d_16_arg_objaddr_1 <= _saxi_register_13 + 704;
          main_fsm <= main_fsm_25;
        end
        main_fsm_25: begin
          conv2d_16_arg_objaddr_2 <= _saxi_register_13 + 3008;
          main_fsm <= main_fsm_26;
        end
        main_fsm_26: begin
          conv2d_16_arg_objaddr_3 <= _saxi_register_13 + 3072;
          main_fsm <= main_fsm_27;
        end
        main_fsm_27: begin
          conv2d_16_control_param_index <= 1;
          main_fsm <= main_fsm_28;
        end
        main_fsm_28: begin
          main_fsm <= main_fsm_29;
        end
        main_fsm_29: begin
          main_fsm <= main_fsm_30;
        end
        main_fsm_30: begin
          if(control_conv2d_16 == 55) begin
            main_fsm <= main_fsm_31;
          end 
        end
        main_fsm_31: begin
          main_fsm <= main_fsm_32;
        end
        main_fsm_32: begin
          max_pool_serial_18_objaddr <= _saxi_register_10 + 28672;
          main_fsm <= main_fsm_33;
        end
        main_fsm_33: begin
          max_pool_serial_18_arg_objaddr_0 <= _saxi_register_10 + 20480;
          main_fsm <= main_fsm_34;
        end
        main_fsm_34: begin
          max_pool_serial_18_control_param_index <= 1;
          main_fsm <= main_fsm_35;
        end
        main_fsm_35: begin
          main_fsm <= main_fsm_36;
        end
        main_fsm_36: begin
          main_fsm <= main_fsm_37;
        end
        main_fsm_37: begin
          if(control_max_pool_serial_18 == 25) begin
            main_fsm <= main_fsm_38;
          end 
        end
        main_fsm_38: begin
          main_fsm <= main_fsm_39;
        end
        main_fsm_39: begin
          conv2d_16_objaddr <= _saxi_register_10 + 30720;
          main_fsm <= main_fsm_40;
        end
        main_fsm_40: begin
          conv2d_16_arg_objaddr_0 <= _saxi_register_10 + 28672;
          main_fsm <= main_fsm_41;
        end
        main_fsm_41: begin
          conv2d_16_arg_objaddr_1 <= _saxi_register_13 + 3136;
          main_fsm <= main_fsm_42;
        end
        main_fsm_42: begin
          conv2d_16_arg_objaddr_2 <= _saxi_register_13 + 12352;
          main_fsm <= main_fsm_43;
        end
        main_fsm_43: begin
          conv2d_16_arg_objaddr_3 <= _saxi_register_13 + 12416;
          main_fsm <= main_fsm_44;
        end
        main_fsm_44: begin
          conv2d_16_control_param_index <= 2;
          main_fsm <= main_fsm_45;
        end
        main_fsm_45: begin
          main_fsm <= main_fsm_46;
        end
        main_fsm_46: begin
          main_fsm <= main_fsm_47;
        end
        main_fsm_47: begin
          if(control_conv2d_16 == 55) begin
            main_fsm <= main_fsm_48;
          end 
        end
        main_fsm_48: begin
          main_fsm <= main_fsm_49;
        end
        main_fsm_49: begin
          max_pool_serial_18_objaddr <= _saxi_register_10 + 34816;
          main_fsm <= main_fsm_50;
        end
        main_fsm_50: begin
          max_pool_serial_18_arg_objaddr_0 <= _saxi_register_10 + 30720;
          main_fsm <= main_fsm_51;
        end
        main_fsm_51: begin
          max_pool_serial_18_control_param_index <= 2;
          main_fsm <= main_fsm_52;
        end
        main_fsm_52: begin
          main_fsm <= main_fsm_53;
        end
        main_fsm_53: begin
          main_fsm <= main_fsm_54;
        end
        main_fsm_54: begin
          if(control_max_pool_serial_18 == 25) begin
            main_fsm <= main_fsm_55;
          end 
        end
        main_fsm_55: begin
          main_fsm <= main_fsm_56;
        end
        main_fsm_56: begin
          main_fsm <= main_fsm_57;
        end
        main_fsm_57: begin
          main_fsm <= main_fsm_58;
        end
        main_fsm_58: begin
          matmul_29_objaddr <= _saxi_register_10 + 35840;
          main_fsm <= main_fsm_59;
        end
        main_fsm_59: begin
          matmul_29_arg_objaddr_0 <= _saxi_register_10 + 34816;
          main_fsm <= main_fsm_60;
        end
        main_fsm_60: begin
          matmul_29_arg_objaddr_1 <= _saxi_register_13 + 12480;
          main_fsm <= main_fsm_61;
        end
        main_fsm_61: begin
          matmul_29_arg_objaddr_2 <= _saxi_register_13 + 143552;
          main_fsm <= main_fsm_62;
        end
        main_fsm_62: begin
          matmul_29_arg_objaddr_3 <= _saxi_register_13 + 143808;
          main_fsm <= main_fsm_63;
        end
        main_fsm_63: begin
          matmul_29_control_param_index <= 0;
          main_fsm <= main_fsm_64;
        end
        main_fsm_64: begin
          main_fsm <= main_fsm_65;
        end
        main_fsm_65: begin
          main_fsm <= main_fsm_66;
        end
        main_fsm_66: begin
          if(control_matmul_29 == 39) begin
            main_fsm <= main_fsm_67;
          end 
        end
        main_fsm_67: begin
          main_fsm <= main_fsm_68;
        end
        main_fsm_68: begin
          matmul_29_objaddr <= _saxi_register_10 + 36096;
          main_fsm <= main_fsm_69;
        end
        main_fsm_69: begin
          matmul_29_arg_objaddr_0 <= _saxi_register_10 + 35840;
          main_fsm <= main_fsm_70;
        end
        main_fsm_70: begin
          matmul_29_arg_objaddr_1 <= _saxi_register_13 + 143872;
          main_fsm <= main_fsm_71;
        end
        main_fsm_71: begin
          matmul_29_arg_objaddr_2 <= _saxi_register_13 + 160256;
          main_fsm <= main_fsm_72;
        end
        main_fsm_72: begin
          matmul_29_arg_objaddr_3 <= _saxi_register_13 + 160384;
          main_fsm <= main_fsm_73;
        end
        main_fsm_73: begin
          matmul_29_control_param_index <= 1;
          main_fsm <= main_fsm_74;
        end
        main_fsm_74: begin
          main_fsm <= main_fsm_75;
        end
        main_fsm_75: begin
          main_fsm <= main_fsm_76;
        end
        main_fsm_76: begin
          if(control_matmul_29 == 39) begin
            main_fsm <= main_fsm_77;
          end 
        end
        main_fsm_77: begin
          main_fsm <= main_fsm_78;
        end
        main_fsm_78: begin
          matmul_29_objaddr <= _saxi_register_11;
          main_fsm <= main_fsm_79;
        end
        main_fsm_79: begin
          matmul_29_arg_objaddr_0 <= _saxi_register_10 + 36096;
          main_fsm <= main_fsm_80;
        end
        main_fsm_80: begin
          matmul_29_arg_objaddr_1 <= _saxi_register_13 + 160448;
          main_fsm <= main_fsm_81;
        end
        main_fsm_81: begin
          matmul_29_arg_objaddr_2 <= _saxi_register_13 + 161088;
          main_fsm <= main_fsm_82;
        end
        main_fsm_82: begin
          matmul_29_arg_objaddr_3 <= _saxi_register_13 + 161152;
          main_fsm <= main_fsm_83;
        end
        main_fsm_83: begin
          matmul_29_control_param_index <= 2;
          main_fsm <= main_fsm_84;
        end
        main_fsm_84: begin
          main_fsm <= main_fsm_85;
        end
        main_fsm_85: begin
          main_fsm <= main_fsm_86;
        end
        main_fsm_86: begin
          if(control_matmul_29 == 39) begin
            main_fsm <= main_fsm_87;
          end 
        end
        main_fsm_87: begin
          main_fsm <= main_fsm_88;
        end
        main_fsm_88: begin
          main_fsm <= main_fsm_89;
        end
        main_fsm_89: begin
          main_fsm <= main_fsm_90;
        end
        main_fsm_90: begin
          main_fsm <= main_fsm_91;
        end
        main_fsm_91: begin
          main_fsm <= main_fsm_92;
        end
        main_fsm_92: begin
          main_fsm <= main_fsm_init;
        end
      endcase
    end
  end

  localparam control_conv2d_16_1 = 1;
  localparam control_conv2d_16_2 = 2;
  localparam control_conv2d_16_3 = 3;
  localparam control_conv2d_16_4 = 4;
  localparam control_conv2d_16_5 = 5;
  localparam control_conv2d_16_6 = 6;
  localparam control_conv2d_16_7 = 7;
  localparam control_conv2d_16_8 = 8;
  localparam control_conv2d_16_9 = 9;
  localparam control_conv2d_16_10 = 10;
  localparam control_conv2d_16_11 = 11;
  localparam control_conv2d_16_12 = 12;
  localparam control_conv2d_16_13 = 13;
  localparam control_conv2d_16_14 = 14;
  localparam control_conv2d_16_15 = 15;
  localparam control_conv2d_16_16 = 16;
  localparam control_conv2d_16_17 = 17;
  localparam control_conv2d_16_18 = 18;
  localparam control_conv2d_16_19 = 19;
  localparam control_conv2d_16_20 = 20;
  localparam control_conv2d_16_21 = 21;
  localparam control_conv2d_16_22 = 22;
  localparam control_conv2d_16_23 = 23;
  localparam control_conv2d_16_24 = 24;
  localparam control_conv2d_16_25 = 25;
  localparam control_conv2d_16_26 = 26;
  localparam control_conv2d_16_27 = 27;
  localparam control_conv2d_16_28 = 28;
  localparam control_conv2d_16_29 = 29;
  localparam control_conv2d_16_30 = 30;
  localparam control_conv2d_16_31 = 31;
  localparam control_conv2d_16_32 = 32;
  localparam control_conv2d_16_33 = 33;
  localparam control_conv2d_16_34 = 34;
  localparam control_conv2d_16_35 = 35;
  localparam control_conv2d_16_36 = 36;
  localparam control_conv2d_16_37 = 37;
  localparam control_conv2d_16_38 = 38;
  localparam control_conv2d_16_39 = 39;
  localparam control_conv2d_16_40 = 40;
  localparam control_conv2d_16_41 = 41;
  localparam control_conv2d_16_42 = 42;
  localparam control_conv2d_16_43 = 43;
  localparam control_conv2d_16_44 = 44;
  localparam control_conv2d_16_45 = 45;
  localparam control_conv2d_16_46 = 46;
  localparam control_conv2d_16_47 = 47;
  localparam control_conv2d_16_48 = 48;
  localparam control_conv2d_16_49 = 49;
  localparam control_conv2d_16_50 = 50;
  localparam control_conv2d_16_51 = 51;
  localparam control_conv2d_16_52 = 52;
  localparam control_conv2d_16_53 = 53;
  localparam control_conv2d_16_54 = 54;
  localparam control_conv2d_16_55 = 55;

  always @(posedge CLK) begin
    if(RST) begin
      control_conv2d_16 <= control_conv2d_16_init;
      _d1_control_conv2d_16 <= control_conv2d_16_init;
      _control_conv2d_16_called <= 0;
      conv2d_16_filter_base_offset <= 0;
      conv2d_16_filter_page_comp_offset <= 0;
      conv2d_16_filter_page_dma_offset <= 0;
      conv2d_16_act_base_offset_row <= 0;
      conv2d_16_act_base_offset_bat <= 0;
      conv2d_16_dma_flag_0 <= 0;
      conv2d_16_dma_flag_1 <= 0;
      conv2d_16_dma_flag_2 <= 0;
      conv2d_16_act_page_comp_offset_0 <= 0;
      conv2d_16_act_page_comp_offset_1 <= 0;
      conv2d_16_act_page_comp_offset_2 <= 0;
      conv2d_16_act_page_dma_offset_0 <= 0;
      conv2d_16_act_page_dma_offset_1 <= 0;
      conv2d_16_act_page_dma_offset_2 <= 0;
      conv2d_16_out_base_offset_val <= 0;
      conv2d_16_out_base_offset_col <= 0;
      conv2d_16_out_base_offset_row <= 0;
      conv2d_16_out_base_offset_bat <= 0;
      conv2d_16_out_base_offset_och <= 0;
      conv2d_16_out_page <= 0;
      conv2d_16_out_page_comp_offset <= 0;
      conv2d_16_out_page_dma_offset <= 0;
      conv2d_16_out_laddr_offset <= 0;
      conv2d_16_sync_out_count <= 0;
      conv2d_16_write_count <= 0;
      conv2d_16_next_out_write_size <= 0;
      conv2d_16_row_count <= 0;
      conv2d_16_bat_count <= 0;
      conv2d_16_och_count <= 0;
      conv2d_16_row_select <= 0;
      conv2d_16_prev_row_count <= 0;
      conv2d_16_prev_bat_count <= 0;
      conv2d_16_prev_och_count <= 0;
      conv2d_16_prev_row_select <= 0;
      conv2d_16_out_col_count <= 0;
      conv2d_16_out_row_count <= 0;
      conv2d_16_out_ram_select <= 0;
      conv2d_16_skip_read_filter <= 0;
      conv2d_16_skip_read_act <= 0;
      conv2d_16_skip_comp <= 0;
      conv2d_16_skip_write_out <= 1;
      axim_flag_9 <= 0;
      _control_conv2d_16_cond_3_0_1 <= 0;
      axim_flag_22 <= 0;
      _control_conv2d_16_cond_8_1_1 <= 0;
      set_req_34 <= 0;
      _control_conv2d_16_cond_14_2_1 <= 0;
      axim_flag_35 <= 0;
      _control_conv2d_16_cond_15_3_1 <= 0;
      set_req_287 <= 0;
      _control_conv2d_16_cond_23_4_1 <= 0;
      axim_flag_288 <= 0;
      _control_conv2d_16_cond_24_5_1 <= 0;
      set_req_344 <= 0;
      _control_conv2d_16_cond_30_6_1 <= 0;
      axim_flag_345 <= 0;
      _control_conv2d_16_cond_31_7_1 <= 0;
      set_req_401 <= 0;
      _control_conv2d_16_cond_37_8_1 <= 0;
      axim_flag_402 <= 0;
      _control_conv2d_16_cond_38_9_1 <= 0;
      axim_flag_970 <= 0;
      _control_conv2d_16_cond_48_10_1 <= 0;
    end else begin
      _d1_control_conv2d_16 <= control_conv2d_16;
      case(_d1_control_conv2d_16)
        control_conv2d_16_3: begin
          if(_control_conv2d_16_cond_3_0_1) begin
            axim_flag_9 <= 0;
          end 
        end
        control_conv2d_16_8: begin
          if(_control_conv2d_16_cond_8_1_1) begin
            axim_flag_22 <= 0;
          end 
        end
        control_conv2d_16_14: begin
          if(_control_conv2d_16_cond_14_2_1) begin
            set_req_34 <= 0;
          end 
        end
        control_conv2d_16_15: begin
          if(_control_conv2d_16_cond_15_3_1) begin
            axim_flag_35 <= 0;
          end 
        end
        control_conv2d_16_23: begin
          if(_control_conv2d_16_cond_23_4_1) begin
            set_req_287 <= 0;
          end 
        end
        control_conv2d_16_24: begin
          if(_control_conv2d_16_cond_24_5_1) begin
            axim_flag_288 <= 0;
          end 
        end
        control_conv2d_16_30: begin
          if(_control_conv2d_16_cond_30_6_1) begin
            set_req_344 <= 0;
          end 
        end
        control_conv2d_16_31: begin
          if(_control_conv2d_16_cond_31_7_1) begin
            axim_flag_345 <= 0;
          end 
        end
        control_conv2d_16_37: begin
          if(_control_conv2d_16_cond_37_8_1) begin
            set_req_401 <= 0;
          end 
        end
        control_conv2d_16_38: begin
          if(_control_conv2d_16_cond_38_9_1) begin
            axim_flag_402 <= 0;
          end 
        end
        control_conv2d_16_48: begin
          if(_control_conv2d_16_cond_48_10_1) begin
            axim_flag_970 <= 0;
          end 
        end
      endcase
      case(control_conv2d_16)
        control_conv2d_16_init: begin
          if(main_fsm == 11) begin
            _control_conv2d_16_called <= 1;
          end 
          if(main_fsm == 28) begin
            _control_conv2d_16_called <= 1;
          end 
          if(main_fsm == 45) begin
            _control_conv2d_16_called <= 1;
          end 
          if(main_fsm == 11) begin
            control_conv2d_16 <= control_conv2d_16_1;
          end 
          if(main_fsm == 28) begin
            control_conv2d_16 <= control_conv2d_16_1;
          end 
          if(main_fsm == 45) begin
            control_conv2d_16 <= control_conv2d_16_1;
          end 
        end
        control_conv2d_16_1: begin
          control_conv2d_16 <= control_conv2d_16_2;
        end
        control_conv2d_16_2: begin
          conv2d_16_filter_base_offset <= 0;
          conv2d_16_filter_page_comp_offset <= 0;
          conv2d_16_filter_page_dma_offset <= 0;
          conv2d_16_act_base_offset_row <= 0;
          conv2d_16_act_base_offset_bat <= 0;
          conv2d_16_dma_flag_0 <= 1;
          conv2d_16_dma_flag_1 <= 1;
          conv2d_16_dma_flag_2 <= 1;
          conv2d_16_act_page_comp_offset_0 <= 0;
          conv2d_16_act_page_comp_offset_1 <= 0;
          conv2d_16_act_page_comp_offset_2 <= 0;
          conv2d_16_act_page_dma_offset_0 <= 0;
          conv2d_16_act_page_dma_offset_1 <= 0;
          conv2d_16_act_page_dma_offset_2 <= 0;
          conv2d_16_out_base_offset_val <= 0;
          conv2d_16_out_base_offset_col <= 0;
          conv2d_16_out_base_offset_row <= 0;
          conv2d_16_out_base_offset_bat <= 0;
          conv2d_16_out_base_offset_och <= 0;
          conv2d_16_out_page <= 0;
          conv2d_16_out_page_comp_offset <= 0;
          conv2d_16_out_page_dma_offset <= 0;
          conv2d_16_out_laddr_offset <= 0;
          conv2d_16_sync_out_count <= 0;
          conv2d_16_write_count <= 0;
          conv2d_16_next_out_write_size <= (cparam_conv2d_16_max_och_count == 0)? cparam_conv2d_16_out_write_size_res : cparam_conv2d_16_out_write_size;
          conv2d_16_row_count <= 0;
          conv2d_16_bat_count <= 0;
          conv2d_16_och_count <= 0;
          conv2d_16_row_select <= 0;
          conv2d_16_prev_row_count <= 0;
          conv2d_16_prev_bat_count <= 0;
          conv2d_16_prev_och_count <= 0;
          conv2d_16_prev_row_select <= 0;
          conv2d_16_out_col_count <= 0;
          conv2d_16_out_row_count <= 0;
          conv2d_16_out_ram_select <= 0;
          conv2d_16_skip_read_filter <= 0;
          conv2d_16_skip_read_act <= 0;
          conv2d_16_skip_comp <= 0;
          conv2d_16_skip_write_out <= 1;
          if(_maxi_read_idle) begin
            control_conv2d_16 <= control_conv2d_16_3;
          end 
        end
        control_conv2d_16_3: begin
          axim_flag_9 <= 1;
          _control_conv2d_16_cond_3_0_1 <= 1;
          control_conv2d_16 <= control_conv2d_16_4;
        end
        control_conv2d_16_4: begin
          control_conv2d_16 <= control_conv2d_16_5;
        end
        control_conv2d_16_5: begin
          control_conv2d_16 <= control_conv2d_16_6;
        end
        control_conv2d_16_6: begin
          if(_maxi_read_idle) begin
            control_conv2d_16 <= control_conv2d_16_7;
          end 
        end
        control_conv2d_16_7: begin
          if(_maxi_read_idle) begin
            control_conv2d_16 <= control_conv2d_16_8;
          end 
        end
        control_conv2d_16_8: begin
          axim_flag_22 <= 1;
          _control_conv2d_16_cond_8_1_1 <= 1;
          control_conv2d_16 <= control_conv2d_16_9;
        end
        control_conv2d_16_9: begin
          control_conv2d_16 <= control_conv2d_16_10;
        end
        control_conv2d_16_10: begin
          control_conv2d_16 <= control_conv2d_16_11;
        end
        control_conv2d_16_11: begin
          if(_maxi_read_idle) begin
            control_conv2d_16 <= control_conv2d_16_12;
          end 
        end
        control_conv2d_16_12: begin
          if(cparam_conv2d_16_data_stationary == 0) begin
            control_conv2d_16 <= control_conv2d_16_13;
          end 
          if(cparam_conv2d_16_data_stationary == 1) begin
            control_conv2d_16 <= control_conv2d_16_21;
          end 
        end
        control_conv2d_16_13: begin
          if(_maxi_read_idle) begin
            control_conv2d_16 <= control_conv2d_16_14;
          end 
          if(conv2d_16_skip_read_filter) begin
            control_conv2d_16 <= control_conv2d_16_20;
          end 
        end
        control_conv2d_16_14: begin
          set_req_34 <= 1;
          _control_conv2d_16_cond_14_2_1 <= 1;
          control_conv2d_16 <= control_conv2d_16_15;
        end
        control_conv2d_16_15: begin
          axim_flag_35 <= 1;
          _control_conv2d_16_cond_15_3_1 <= 1;
          control_conv2d_16 <= control_conv2d_16_16;
        end
        control_conv2d_16_16: begin
          control_conv2d_16 <= control_conv2d_16_17;
        end
        control_conv2d_16_17: begin
          control_conv2d_16 <= control_conv2d_16_18;
        end
        control_conv2d_16_18: begin
          if(_maxi_read_idle) begin
            control_conv2d_16 <= control_conv2d_16_19;
          end 
        end
        control_conv2d_16_19: begin
          control_conv2d_16 <= control_conv2d_16_20;
        end
        control_conv2d_16_20: begin
          if(cparam_conv2d_16_data_stationary == 0) begin
            control_conv2d_16 <= control_conv2d_16_21;
          end 
          if(cparam_conv2d_16_data_stationary == 1) begin
            control_conv2d_16 <= control_conv2d_16_44;
          end 
        end
        control_conv2d_16_21: begin
          control_conv2d_16 <= control_conv2d_16_22;
          if(conv2d_16_mux_dma_pad_mask_0 || !conv2d_16_mux_dma_flag_0) begin
            control_conv2d_16 <= control_conv2d_16_28;
          end 
          if(conv2d_16_skip_read_act) begin
            control_conv2d_16 <= control_conv2d_16_43;
          end 
        end
        control_conv2d_16_22: begin
          if(_maxi_read_idle) begin
            control_conv2d_16 <= control_conv2d_16_23;
          end 
        end
        control_conv2d_16_23: begin
          set_req_287 <= 1;
          _control_conv2d_16_cond_23_4_1 <= 1;
          control_conv2d_16 <= control_conv2d_16_24;
        end
        control_conv2d_16_24: begin
          axim_flag_288 <= 1;
          _control_conv2d_16_cond_24_5_1 <= 1;
          control_conv2d_16 <= control_conv2d_16_25;
        end
        control_conv2d_16_25: begin
          control_conv2d_16 <= control_conv2d_16_26;
        end
        control_conv2d_16_26: begin
          control_conv2d_16 <= control_conv2d_16_27;
        end
        control_conv2d_16_27: begin
          if(_maxi_read_idle) begin
            control_conv2d_16 <= control_conv2d_16_28;
          end 
        end
        control_conv2d_16_28: begin
          control_conv2d_16 <= control_conv2d_16_29;
          if(conv2d_16_mux_dma_pad_mask_1 || !conv2d_16_mux_dma_flag_1) begin
            control_conv2d_16 <= control_conv2d_16_35;
          end 
        end
        control_conv2d_16_29: begin
          if(_maxi_read_idle) begin
            control_conv2d_16 <= control_conv2d_16_30;
          end 
        end
        control_conv2d_16_30: begin
          set_req_344 <= 1;
          _control_conv2d_16_cond_30_6_1 <= 1;
          control_conv2d_16 <= control_conv2d_16_31;
        end
        control_conv2d_16_31: begin
          axim_flag_345 <= 1;
          _control_conv2d_16_cond_31_7_1 <= 1;
          control_conv2d_16 <= control_conv2d_16_32;
        end
        control_conv2d_16_32: begin
          control_conv2d_16 <= control_conv2d_16_33;
        end
        control_conv2d_16_33: begin
          control_conv2d_16 <= control_conv2d_16_34;
        end
        control_conv2d_16_34: begin
          if(_maxi_read_idle) begin
            control_conv2d_16 <= control_conv2d_16_35;
          end 
        end
        control_conv2d_16_35: begin
          control_conv2d_16 <= control_conv2d_16_36;
          if(conv2d_16_mux_dma_pad_mask_2 || !conv2d_16_mux_dma_flag_2) begin
            control_conv2d_16 <= control_conv2d_16_42;
          end 
        end
        control_conv2d_16_36: begin
          if(_maxi_read_idle) begin
            control_conv2d_16 <= control_conv2d_16_37;
          end 
        end
        control_conv2d_16_37: begin
          set_req_401 <= 1;
          _control_conv2d_16_cond_37_8_1 <= 1;
          control_conv2d_16 <= control_conv2d_16_38;
        end
        control_conv2d_16_38: begin
          axim_flag_402 <= 1;
          _control_conv2d_16_cond_38_9_1 <= 1;
          control_conv2d_16 <= control_conv2d_16_39;
        end
        control_conv2d_16_39: begin
          control_conv2d_16 <= control_conv2d_16_40;
        end
        control_conv2d_16_40: begin
          control_conv2d_16 <= control_conv2d_16_41;
        end
        control_conv2d_16_41: begin
          if(_maxi_read_idle) begin
            control_conv2d_16 <= control_conv2d_16_42;
          end 
        end
        control_conv2d_16_42: begin
          control_conv2d_16 <= control_conv2d_16_43;
        end
        control_conv2d_16_43: begin
          if(cparam_conv2d_16_data_stationary == 0) begin
            control_conv2d_16 <= control_conv2d_16_44;
          end 
          if(cparam_conv2d_16_data_stationary == 1) begin
            control_conv2d_16 <= control_conv2d_16_13;
          end 
        end
        control_conv2d_16_44: begin
          if(conv2d_16_comp_fsm == 0) begin
            control_conv2d_16 <= control_conv2d_16_45;
          end 
        end
        control_conv2d_16_45: begin
          if(conv2d_16_sync_comp_count >= conv2d_16_sync_out_count + cparam_conv2d_16_inc_sync_out) begin
            control_conv2d_16 <= control_conv2d_16_46;
          end 
          if(conv2d_16_skip_write_out) begin
            control_conv2d_16 <= control_conv2d_16_53;
          end 
          if((cparam_conv2d_16_data_stationary == 1) && (conv2d_16_prev_och_count < cparam_conv2d_16_max_och_count)) begin
            control_conv2d_16 <= control_conv2d_16_53;
          end 
        end
        control_conv2d_16_46: begin
          if(!conv2d_16_dma_out_mask_0) begin
            control_conv2d_16 <= control_conv2d_16_47;
          end 
          if(conv2d_16_dma_out_mask_0) begin
            control_conv2d_16 <= control_conv2d_16_51;
          end 
        end
        control_conv2d_16_47: begin
          if(_maxi_write_idle) begin
            control_conv2d_16 <= control_conv2d_16_48;
          end 
        end
        control_conv2d_16_48: begin
          axim_flag_970 <= 1;
          _control_conv2d_16_cond_48_10_1 <= 1;
          control_conv2d_16 <= control_conv2d_16_49;
        end
        control_conv2d_16_49: begin
          control_conv2d_16 <= control_conv2d_16_50;
        end
        control_conv2d_16_50: begin
          control_conv2d_16 <= control_conv2d_16_51;
        end
        control_conv2d_16_51: begin
          control_conv2d_16 <= control_conv2d_16_52;
        end
        control_conv2d_16_52: begin
          conv2d_16_write_count <= conv2d_16_write_count + 1;
          if(conv2d_16_out_ram_select == 0) begin
            conv2d_16_out_laddr_offset <= conv2d_16_out_laddr_offset + conv2d_16_next_out_write_size;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && !cparam_conv2d_16_keep_filter) begin
            conv2d_16_out_base_offset_col <= conv2d_16_out_base_offset_col + cparam_conv2d_16_out_col_step;
            conv2d_16_out_col_count <= conv2d_16_out_col_count + 1;
          end 
          conv2d_16_out_ram_select <= conv2d_16_out_ram_select + 1;
          if(conv2d_16_out_ram_select == 0) begin
            conv2d_16_out_ram_select <= 0;
          end 
          conv2d_16_sync_out_count <= conv2d_16_sync_out_count + cparam_conv2d_16_inc_sync_out;
          if((cparam_conv2d_16_data_stationary == 0) && !cparam_conv2d_16_keep_filter && (conv2d_16_write_count >= cparam_conv2d_16_out_num_col - 1) || (cparam_conv2d_16_data_stationary == 0) && cparam_conv2d_16_keep_filter || (cparam_conv2d_16_data_stationary == 1)) begin
            conv2d_16_sync_out_count <= conv2d_16_sync_out_count + (cparam_conv2d_16_inc_sync_out + cparam_conv2d_16_inc_sync_out_res);
          end 
          if((cparam_conv2d_16_data_stationary == 0) && !cparam_conv2d_16_keep_filter) begin
            control_conv2d_16 <= control_conv2d_16_45;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && !cparam_conv2d_16_keep_filter && (conv2d_16_write_count >= cparam_conv2d_16_out_num_col - 1) || (cparam_conv2d_16_data_stationary == 0) && cparam_conv2d_16_keep_filter || (cparam_conv2d_16_data_stationary == 1)) begin
            control_conv2d_16 <= control_conv2d_16_53;
          end 
        end
        control_conv2d_16_53: begin
          if(conv2d_16_update_filter) begin
            conv2d_16_filter_base_offset <= conv2d_16_filter_base_offset + cparam_conv2d_16_filter_base_step;
          end 
          if((cparam_conv2d_16_data_stationary == 1) && (conv2d_16_och_count >= cparam_conv2d_16_max_och_count)) begin
            conv2d_16_filter_base_offset <= 0;
          end 
          if(conv2d_16_update_filter) begin
            conv2d_16_och_count <= conv2d_16_och_count + cparam_conv2d_16_och_count_step;
          end 
          if((cparam_conv2d_16_data_stationary == 1) && (conv2d_16_och_count >= cparam_conv2d_16_max_och_count)) begin
            conv2d_16_och_count <= 0;
          end 
          if(conv2d_16_update_filter) begin
            conv2d_16_filter_page_comp_offset <= conv2d_16_filter_page_comp_offset + cparam_conv2d_16_filter_read_step;
            conv2d_16_filter_page_dma_offset <= conv2d_16_filter_page_dma_offset + cparam_conv2d_16_filter_read_step;
          end 
          if(conv2d_16_update_filter && (conv2d_16_filter_page_comp_offset + cparam_conv2d_16_filter_read_step + cparam_conv2d_16_filter_read_step > 8192)) begin
            conv2d_16_filter_page_comp_offset <= 0;
            conv2d_16_filter_page_dma_offset <= 0;
          end 
          if(conv2d_16_update_act) begin
            conv2d_16_act_base_offset_row <= conv2d_16_act_base_offset_row + cparam_conv2d_16_act_row_step;
          end 
          if(conv2d_16_update_act && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)) begin
            conv2d_16_act_base_offset_row <= 0;
            conv2d_16_act_base_offset_bat <= conv2d_16_act_base_offset_bat + cparam_conv2d_16_act_bat_step;
          end 
          if(conv2d_16_update_act && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_bat_count >= cparam_conv2d_16_max_bat_count)) begin
            conv2d_16_act_base_offset_bat <= 0;
          end 
          if(!conv2d_16_update_act) begin
            conv2d_16_dma_flag_0 <= 0;
          end 
          if(conv2d_16_update_act) begin
            conv2d_16_dma_flag_0 <= cparam_conv2d_16_dma_flag_conds_0;
          end 
          if(conv2d_16_update_act && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)) begin
            conv2d_16_dma_flag_0 <= 1;
          end 
          if(!conv2d_16_update_act) begin
            conv2d_16_dma_flag_1 <= 0;
          end 
          if(conv2d_16_update_act) begin
            conv2d_16_dma_flag_1 <= cparam_conv2d_16_dma_flag_conds_1;
          end 
          if(conv2d_16_update_act && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)) begin
            conv2d_16_dma_flag_1 <= 1;
          end 
          if(!conv2d_16_update_act) begin
            conv2d_16_dma_flag_2 <= 0;
          end 
          if(conv2d_16_update_act) begin
            conv2d_16_dma_flag_2 <= cparam_conv2d_16_dma_flag_conds_2;
          end 
          if(conv2d_16_update_act && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)) begin
            conv2d_16_dma_flag_2 <= 1;
          end 
          if(conv2d_16_update_act) begin
            conv2d_16_row_count <= conv2d_16_row_count + cparam_conv2d_16_stride_row_par_row;
          end 
          if(conv2d_16_update_act && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)) begin
            conv2d_16_row_count <= 0;
            conv2d_16_bat_count <= conv2d_16_bat_count + 1;
          end 
          if(conv2d_16_update_act && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_bat_count >= cparam_conv2d_16_max_bat_count)) begin
            conv2d_16_bat_count <= 0;
          end 
          if(conv2d_16_update_act && (cparam_conv2d_16_stride_row_par_row < 3)) begin
            conv2d_16_row_select <= conv2d_16_row_select + cparam_conv2d_16_stride_row_par_row;
            conv2d_16_prev_row_select <= conv2d_16_row_select;
          end 
          if(conv2d_16_update_act && (cparam_conv2d_16_stride_row_par_row < 3) && (conv2d_16_row_select + cparam_conv2d_16_stride_row_par_row >= 3)) begin
            conv2d_16_row_select <= conv2d_16_row_select - (3 - cparam_conv2d_16_stride_row_par_row);
            conv2d_16_prev_row_select <= conv2d_16_row_select;
          end 
          if(conv2d_16_update_act && !(cparam_conv2d_16_stride_row_par_row < 3)) begin
            conv2d_16_row_select <= 0;
            conv2d_16_prev_row_select <= 0;
          end 
          if(conv2d_16_update_act && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count)) begin
            conv2d_16_row_select <= 0;
            conv2d_16_prev_row_select <= 0;
          end 
          if(conv2d_16_update_act && conv2d_16_mux_next_dma_flag_0) begin
            conv2d_16_act_page_comp_offset_0 <= conv2d_16_act_page_comp_offset_0 + cparam_conv2d_16_act_read_step;
            conv2d_16_act_page_dma_offset_0 <= conv2d_16_act_page_dma_offset_0 + cparam_conv2d_16_act_read_step;
          end 
          if(conv2d_16_update_act && conv2d_16_mux_next_dma_flag_0 && (conv2d_16_act_page_comp_offset_0 + cparam_conv2d_16_act_read_step + cparam_conv2d_16_act_read_step > 2048)) begin
            conv2d_16_act_page_comp_offset_0 <= 0;
            conv2d_16_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_bat_count >= cparam_conv2d_16_max_bat_count) && cparam_conv2d_16_keep_input) begin
            conv2d_16_act_page_comp_offset_0 <= 0;
            conv2d_16_act_page_dma_offset_0 <= 0;
          end 
          if(conv2d_16_update_act && conv2d_16_mux_next_dma_flag_1) begin
            conv2d_16_act_page_comp_offset_1 <= conv2d_16_act_page_comp_offset_1 + cparam_conv2d_16_act_read_step;
            conv2d_16_act_page_dma_offset_1 <= conv2d_16_act_page_dma_offset_1 + cparam_conv2d_16_act_read_step;
          end 
          if(conv2d_16_update_act && conv2d_16_mux_next_dma_flag_1 && (conv2d_16_act_page_comp_offset_1 + cparam_conv2d_16_act_read_step + cparam_conv2d_16_act_read_step > 2048)) begin
            conv2d_16_act_page_comp_offset_1 <= 0;
            conv2d_16_act_page_dma_offset_1 <= 0;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_bat_count >= cparam_conv2d_16_max_bat_count) && cparam_conv2d_16_keep_input) begin
            conv2d_16_act_page_comp_offset_1 <= 0;
            conv2d_16_act_page_dma_offset_1 <= 0;
          end 
          if(conv2d_16_update_act && conv2d_16_mux_next_dma_flag_2) begin
            conv2d_16_act_page_comp_offset_2 <= conv2d_16_act_page_comp_offset_2 + cparam_conv2d_16_act_read_step;
            conv2d_16_act_page_dma_offset_2 <= conv2d_16_act_page_dma_offset_2 + cparam_conv2d_16_act_read_step;
          end 
          if(conv2d_16_update_act && conv2d_16_mux_next_dma_flag_2 && (conv2d_16_act_page_comp_offset_2 + cparam_conv2d_16_act_read_step + cparam_conv2d_16_act_read_step > 2048)) begin
            conv2d_16_act_page_comp_offset_2 <= 0;
            conv2d_16_act_page_dma_offset_2 <= 0;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_bat_count >= cparam_conv2d_16_max_bat_count) && cparam_conv2d_16_keep_input) begin
            conv2d_16_act_page_comp_offset_2 <= 0;
            conv2d_16_act_page_dma_offset_2 <= 0;
          end 
          conv2d_16_next_out_write_size <= (conv2d_16_och_count >= cparam_conv2d_16_max_och_count)? cparam_conv2d_16_out_write_size_res : cparam_conv2d_16_out_write_size;
          if(!conv2d_16_skip_write_out) begin
            conv2d_16_write_count <= 0;
            conv2d_16_out_laddr_offset <= 0;
            conv2d_16_out_ram_select <= 0;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && !conv2d_16_skip_write_out) begin
            conv2d_16_out_base_offset_col <= 0;
            conv2d_16_out_base_offset_row <= conv2d_16_out_base_offset_row + cparam_conv2d_16_out_row_step;
            conv2d_16_out_col_count <= 0;
            conv2d_16_out_row_count <= conv2d_16_out_row_count + 1;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && !conv2d_16_skip_write_out && (conv2d_16_prev_row_count >= cparam_conv2d_16_max_row_count)) begin
            conv2d_16_out_base_offset_row <= 0;
            conv2d_16_out_base_offset_bat <= conv2d_16_out_base_offset_bat + cparam_conv2d_16_out_bat_step;
            conv2d_16_out_row_count <= 0;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && !conv2d_16_skip_write_out && (conv2d_16_prev_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_prev_bat_count >= cparam_conv2d_16_max_bat_count)) begin
            conv2d_16_out_base_offset_bat <= 0;
            conv2d_16_out_base_offset_och <= conv2d_16_out_base_offset_och + cparam_conv2d_16_out_och_step;
          end 
          if((cparam_conv2d_16_data_stationary == 1) && (conv2d_16_prev_och_count >= cparam_conv2d_16_max_och_count) && !conv2d_16_skip_write_out) begin
            conv2d_16_out_base_offset_row <= conv2d_16_out_base_offset_row + cparam_conv2d_16_out_row_step;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && !conv2d_16_out_page) begin
            conv2d_16_out_page_comp_offset <= 1024;
            conv2d_16_out_page_dma_offset <= 0;
            conv2d_16_out_page <= 1;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && conv2d_16_out_page) begin
            conv2d_16_out_page_comp_offset <= 0;
            conv2d_16_out_page_dma_offset <= 1024;
            conv2d_16_out_page <= 0;
          end 
          if((cparam_conv2d_16_data_stationary == 1) && (conv2d_16_och_count >= cparam_conv2d_16_max_och_count) && !conv2d_16_out_page) begin
            conv2d_16_out_page_comp_offset <= 1024;
            conv2d_16_out_page_dma_offset <= 0;
            conv2d_16_out_page <= 1;
          end 
          if((cparam_conv2d_16_data_stationary == 1) && (conv2d_16_och_count >= cparam_conv2d_16_max_och_count) && conv2d_16_out_page) begin
            conv2d_16_out_page_comp_offset <= 0;
            conv2d_16_out_page_dma_offset <= 1024;
            conv2d_16_out_page <= 0;
          end 
          conv2d_16_prev_row_count <= conv2d_16_row_count;
          conv2d_16_prev_bat_count <= conv2d_16_bat_count;
          conv2d_16_prev_och_count <= conv2d_16_och_count;
          if((conv2d_16_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_bat_count >= cparam_conv2d_16_max_bat_count) && (conv2d_16_och_count >= cparam_conv2d_16_max_och_count)) begin
            conv2d_16_skip_read_filter <= 1;
          end 
          if((cparam_conv2d_16_data_stationary == 1) && cparam_conv2d_16_keep_filter) begin
            conv2d_16_skip_read_filter <= 1;
          end 
          if((conv2d_16_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_bat_count >= cparam_conv2d_16_max_bat_count) && (conv2d_16_och_count >= cparam_conv2d_16_max_och_count)) begin
            conv2d_16_skip_read_act <= 1;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_bat_count >= cparam_conv2d_16_max_bat_count) && cparam_conv2d_16_keep_input) begin
            conv2d_16_skip_read_act <= 1;
          end 
          if((conv2d_16_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_bat_count >= cparam_conv2d_16_max_bat_count) && (conv2d_16_och_count >= cparam_conv2d_16_max_och_count)) begin
            conv2d_16_skip_comp <= 1;
          end 
          if(conv2d_16_skip_write_out && (conv2d_16_prev_row_count == 0) && (conv2d_16_prev_bat_count == 0) && (conv2d_16_prev_och_count == 0)) begin
            conv2d_16_skip_write_out <= 0;
          end 
          if(cparam_conv2d_16_data_stationary == 0) begin
            control_conv2d_16 <= control_conv2d_16_21;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && (conv2d_16_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_bat_count >= cparam_conv2d_16_max_bat_count)) begin
            control_conv2d_16 <= control_conv2d_16_13;
          end 
          if(cparam_conv2d_16_data_stationary == 1) begin
            control_conv2d_16 <= control_conv2d_16_13;
          end 
          if((cparam_conv2d_16_data_stationary == 1) && (conv2d_16_och_count >= cparam_conv2d_16_max_och_count)) begin
            control_conv2d_16 <= control_conv2d_16_21;
          end 
          if(!conv2d_16_skip_write_out && (conv2d_16_prev_och_count >= cparam_conv2d_16_max_och_count) && (conv2d_16_prev_row_count >= cparam_conv2d_16_max_row_count) && (conv2d_16_prev_bat_count >= cparam_conv2d_16_max_bat_count)) begin
            control_conv2d_16 <= control_conv2d_16_54;
          end 
        end
        control_conv2d_16_54: begin
          if(_maxi_write_idle) begin
            control_conv2d_16 <= control_conv2d_16_55;
          end 
        end
        control_conv2d_16_55: begin
          if(main_fsm == 14) begin
            _control_conv2d_16_called <= 0;
          end 
          if(main_fsm == 31) begin
            _control_conv2d_16_called <= 0;
          end 
          if(main_fsm == 48) begin
            _control_conv2d_16_called <= 0;
          end 
          if(main_fsm == 14) begin
            control_conv2d_16 <= control_conv2d_16_init;
          end 
          if(main_fsm == 31) begin
            control_conv2d_16 <= control_conv2d_16_init;
          end 
          if(main_fsm == 48) begin
            control_conv2d_16 <= control_conv2d_16_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_fsm_1 = 1;
  localparam _maxi_read_fsm_2 = 2;
  localparam _maxi_read_fsm_3 = 3;
  localparam _maxi_read_fsm_4 = 4;
  localparam _maxi_read_fsm_5 = 5;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_fsm <= _maxi_read_fsm_init;
      _d1__maxi_read_fsm <= _maxi_read_fsm_init;
      _maxi_read_cur_global_addr <= 0;
      _maxi_read_rest_size <= 0;
      _maxi_read_cur_size <= 0;
      __maxi_read_fsm_cond_3_0_1 <= 0;
      _wvalid_11 <= 0;
      _wdata_10 <= 0;
      axim_flag_21 <= 0;
      __maxi_read_fsm_cond_4_1_1 <= 0;
      __maxi_read_fsm_cond_3_2_1 <= 0;
      _wvalid_24 <= 0;
      _wdata_23 <= 0;
      __maxi_read_fsm_cond_3_3_1 <= 0;
      _wvalid_37 <= 0;
      _wdata_36 <= 0;
      __maxi_read_fsm_cond_3_4_1 <= 0;
      _wvalid_290 <= 0;
      _wdata_289 <= 0;
      __maxi_read_fsm_cond_3_5_1 <= 0;
      _wvalid_347 <= 0;
      _wdata_346 <= 0;
      __maxi_read_fsm_cond_3_6_1 <= 0;
      _wvalid_404 <= 0;
      _wdata_403 <= 0;
      __maxi_read_fsm_cond_3_7_1 <= 0;
      _wvalid_1123 <= 0;
      _wdata_1122 <= 0;
      __maxi_read_fsm_cond_3_8_1 <= 0;
      _wvalid_1135 <= 0;
      _wdata_1134 <= 0;
      __maxi_read_fsm_cond_3_9_1 <= 0;
      _wvalid_1154 <= 0;
      _wdata_1153 <= 0;
    end else begin
      _d1__maxi_read_fsm <= _maxi_read_fsm;
      case(_d1__maxi_read_fsm)
        _maxi_read_fsm_3: begin
          if(__maxi_read_fsm_cond_3_0_1) begin
            _wvalid_11 <= 0;
          end 
          if(__maxi_read_fsm_cond_3_2_1) begin
            _wvalid_24 <= 0;
          end 
          if(__maxi_read_fsm_cond_3_3_1) begin
            _wvalid_37 <= 0;
          end 
          if(__maxi_read_fsm_cond_3_4_1) begin
            _wvalid_290 <= 0;
          end 
          if(__maxi_read_fsm_cond_3_5_1) begin
            _wvalid_347 <= 0;
          end 
          if(__maxi_read_fsm_cond_3_6_1) begin
            _wvalid_404 <= 0;
          end 
          if(__maxi_read_fsm_cond_3_7_1) begin
            _wvalid_1123 <= 0;
          end 
          if(__maxi_read_fsm_cond_3_8_1) begin
            _wvalid_1135 <= 0;
          end 
          if(__maxi_read_fsm_cond_3_9_1) begin
            _wvalid_1154 <= 0;
          end 
        end
        _maxi_read_fsm_4: begin
          if(__maxi_read_fsm_cond_4_1_1) begin
            axim_flag_21 <= 0;
          end 
        end
      endcase
      case(_maxi_read_fsm)
        _maxi_read_fsm_init: begin
          if(_maxi_read_start) begin
            _maxi_read_cur_global_addr <= (_maxi_read_global_addr + _maxi_global_base_addr >> 2) << 2;
            _maxi_read_rest_size <= _maxi_read_size;
          end 
          if(_maxi_read_start && (_maxi_read_op_sel == 1)) begin
            _maxi_read_fsm <= _maxi_read_fsm_1;
          end 
          if(_maxi_read_start && (_maxi_read_op_sel == 2)) begin
            _maxi_read_fsm <= _maxi_read_fsm_1;
          end 
          if(_maxi_read_start && (_maxi_read_op_sel == 3)) begin
            _maxi_read_fsm <= _maxi_read_fsm_1;
          end 
          if(_maxi_read_start && (_maxi_read_op_sel == 4)) begin
            _maxi_read_fsm <= _maxi_read_fsm_1;
          end 
          if(_maxi_read_start && (_maxi_read_op_sel == 5)) begin
            _maxi_read_fsm <= _maxi_read_fsm_1;
          end 
          if(_maxi_read_start && (_maxi_read_op_sel == 6)) begin
            _maxi_read_fsm <= _maxi_read_fsm_1;
          end 
          if(_maxi_read_start && (_maxi_read_op_sel == 7)) begin
            _maxi_read_fsm <= _maxi_read_fsm_1;
          end 
          if(_maxi_read_start && (_maxi_read_op_sel == 8)) begin
            _maxi_read_fsm <= _maxi_read_fsm_1;
          end 
          if(_maxi_read_start && (_maxi_read_op_sel == 9)) begin
            _maxi_read_fsm <= _maxi_read_fsm_1;
          end 
        end
        _maxi_read_fsm_1: begin
          if((_maxi_read_rest_size <= 256) && ((_maxi_read_cur_global_addr & 4095) + (_maxi_read_rest_size << 2) >= 4096)) begin
            _maxi_read_cur_size <= 4096 - (_maxi_read_cur_global_addr & 4095) >> 2;
            _maxi_read_rest_size <= _maxi_read_rest_size - (4096 - (_maxi_read_cur_global_addr & 4095) >> 2);
          end else if(_maxi_read_rest_size <= 256) begin
            _maxi_read_cur_size <= _maxi_read_rest_size;
            _maxi_read_rest_size <= 0;
          end else if((_maxi_read_cur_global_addr & 4095) + 1024 >= 4096) begin
            _maxi_read_cur_size <= 4096 - (_maxi_read_cur_global_addr & 4095) >> 2;
            _maxi_read_rest_size <= _maxi_read_rest_size - (4096 - (_maxi_read_cur_global_addr & 4095) >> 2);
          end else begin
            _maxi_read_cur_size <= 256;
            _maxi_read_rest_size <= _maxi_read_rest_size - 256;
          end
          _maxi_read_fsm <= _maxi_read_fsm_2;
        end
        _maxi_read_fsm_2: begin
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_fsm <= _maxi_read_fsm_3;
          end 
        end
        _maxi_read_fsm_3: begin
          __maxi_read_fsm_cond_3_0_1 <= 1;
          if(maxi_rready && maxi_rvalid && (_maxi_read_op_sel == 1)) begin
            _wdata_10 <= maxi_rdata;
            _wvalid_11 <= 1;
          end 
          if(maxi_rready && maxi_rvalid && maxi_rlast) begin
            _maxi_read_cur_global_addr <= _maxi_read_cur_global_addr + (_maxi_read_cur_size << 2);
          end 
          __maxi_read_fsm_cond_3_2_1 <= 1;
          if(maxi_rready && maxi_rvalid && (_maxi_read_op_sel == 2)) begin
            _wdata_23 <= maxi_rdata;
            _wvalid_24 <= 1;
          end 
          __maxi_read_fsm_cond_3_3_1 <= 1;
          if(maxi_rready && maxi_rvalid && (_maxi_read_op_sel == 3)) begin
            _wdata_36 <= maxi_rdata;
            _wvalid_37 <= 1;
          end 
          __maxi_read_fsm_cond_3_4_1 <= 1;
          if(maxi_rready && maxi_rvalid && (_maxi_read_op_sel == 4)) begin
            _wdata_289 <= maxi_rdata;
            _wvalid_290 <= 1;
          end 
          __maxi_read_fsm_cond_3_5_1 <= 1;
          if(maxi_rready && maxi_rvalid && (_maxi_read_op_sel == 5)) begin
            _wdata_346 <= maxi_rdata;
            _wvalid_347 <= 1;
          end 
          __maxi_read_fsm_cond_3_6_1 <= 1;
          if(maxi_rready && maxi_rvalid && (_maxi_read_op_sel == 6)) begin
            _wdata_403 <= maxi_rdata;
            _wvalid_404 <= 1;
          end 
          __maxi_read_fsm_cond_3_7_1 <= 1;
          if(maxi_rready && maxi_rvalid && (_maxi_read_op_sel == 7)) begin
            _wdata_1122 <= maxi_rdata;
            _wvalid_1123 <= 1;
          end 
          __maxi_read_fsm_cond_3_8_1 <= 1;
          if(maxi_rready && maxi_rvalid && (_maxi_read_op_sel == 8)) begin
            _wdata_1134 <= maxi_rdata;
            _wvalid_1135 <= 1;
          end 
          __maxi_read_fsm_cond_3_9_1 <= 1;
          if(maxi_rready && maxi_rvalid && (_maxi_read_op_sel == 9)) begin
            _wdata_1153 <= maxi_rdata;
            _wvalid_1154 <= 1;
          end 
          if(maxi_rready && maxi_rvalid && maxi_rlast && (_maxi_read_rest_size > 0)) begin
            _maxi_read_fsm <= _maxi_read_fsm_1;
          end 
          if(maxi_rready && maxi_rvalid && maxi_rlast && (_maxi_read_rest_size == 0)) begin
            _maxi_read_fsm <= _maxi_read_fsm_4;
          end 
        end
        _maxi_read_fsm_4: begin
          axim_flag_21 <= 1;
          __maxi_read_fsm_cond_4_1_1 <= 1;
          _maxi_read_fsm <= _maxi_read_fsm_5;
        end
        _maxi_read_fsm_5: begin
          _maxi_read_fsm <= _maxi_read_fsm_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      req_block_size_33 <= 0;
    end else begin
      if(set_req_34) begin
        req_block_size_33 <= cparam_conv2d_16_filter_read_block >> 3;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      req_block_size_286 <= 0;
    end else begin
      if(set_req_287) begin
        req_block_size_286 <= cparam_conv2d_16_act_read_block >> 2;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      req_block_size_343 <= 0;
    end else begin
      if(set_req_344) begin
        req_block_size_343 <= cparam_conv2d_16_act_read_block >> 2;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      req_block_size_400 <= 0;
    end else begin
      if(set_req_401) begin
        req_block_size_400 <= cparam_conv2d_16_act_read_block >> 2;
      end 
    end
  end

  localparam conv2d_16_comp_fsm_1 = 1;
  localparam conv2d_16_comp_fsm_2 = 2;
  localparam conv2d_16_comp_fsm_3 = 3;
  localparam conv2d_16_comp_fsm_4 = 4;
  localparam conv2d_16_comp_fsm_5 = 5;
  localparam conv2d_16_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      conv2d_16_comp_fsm <= conv2d_16_comp_fsm_init;
      conv2d_16_stream_act_local_0 <= 0;
      conv2d_16_stream_act_local_1 <= 0;
      conv2d_16_stream_act_local_2 <= 0;
      conv2d_16_stream_act_local_3 <= 0;
      conv2d_16_stream_act_local_4 <= 0;
      conv2d_16_stream_act_local_5 <= 0;
      conv2d_16_stream_act_local_6 <= 0;
      conv2d_16_stream_act_local_7 <= 0;
      conv2d_16_stream_act_local_8 <= 0;
      conv2d_16_stream_out_local_col <= 0;
      conv2d_16_stream_out_local_val <= 0;
      conv2d_16_col_count <= 0;
      conv2d_16_col_select <= 0;
      conv2d_16_filter_page_comp_offset_buf <= 0;
      conv2d_16_act_page_comp_offset_buf_0 <= 0;
      conv2d_16_act_page_comp_offset_buf_1 <= 0;
      conv2d_16_act_page_comp_offset_buf_2 <= 0;
      conv2d_16_out_page_comp_offset_buf <= 0;
      conv2d_16_row_count_buf <= 0;
      conv2d_16_row_select_buf <= 0;
      conv2d_16_och_count_buf <= 0;
      conv2d_16_next_stream_num_ops <= 0;
      conv2d_16_stream_pad_masks <= 0;
      conv2d_16_sync_comp_count <= 0;
    end else begin
      if(_stream_conv2d_16_end_flag) begin
        conv2d_16_sync_comp_count <= conv2d_16_sync_comp_count + 1;
      end 
      if(control_conv2d_16 == 12) begin
        conv2d_16_sync_comp_count <= 0;
      end 
      case(conv2d_16_comp_fsm)
        conv2d_16_comp_fsm_init: begin
          if((control_conv2d_16 == 44) && !conv2d_16_skip_comp) begin
            conv2d_16_comp_fsm <= conv2d_16_comp_fsm_1;
          end 
        end
        conv2d_16_comp_fsm_1: begin
          conv2d_16_stream_act_local_0 <= 0;
          if(cparam_conv2d_16_stream_act_local_small_flags_0) begin
            conv2d_16_stream_act_local_0 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_16_stream_act_local_large_flags_0) begin
            conv2d_16_stream_act_local_0 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          conv2d_16_stream_act_local_1 <= 0;
          if(cparam_conv2d_16_stream_act_local_small_flags_1) begin
            conv2d_16_stream_act_local_1 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_16_stream_act_local_large_flags_1) begin
            conv2d_16_stream_act_local_1 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          conv2d_16_stream_act_local_2 <= 0;
          if(cparam_conv2d_16_stream_act_local_small_flags_2) begin
            conv2d_16_stream_act_local_2 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_16_stream_act_local_large_flags_2) begin
            conv2d_16_stream_act_local_2 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          conv2d_16_stream_act_local_3 <= 0;
          if(cparam_conv2d_16_stream_act_local_small_flags_0) begin
            conv2d_16_stream_act_local_3 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_16_stream_act_local_large_flags_0) begin
            conv2d_16_stream_act_local_3 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          conv2d_16_stream_act_local_4 <= 0;
          if(cparam_conv2d_16_stream_act_local_small_flags_1) begin
            conv2d_16_stream_act_local_4 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_16_stream_act_local_large_flags_1) begin
            conv2d_16_stream_act_local_4 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          conv2d_16_stream_act_local_5 <= 0;
          if(cparam_conv2d_16_stream_act_local_small_flags_2) begin
            conv2d_16_stream_act_local_5 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_16_stream_act_local_large_flags_2) begin
            conv2d_16_stream_act_local_5 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          conv2d_16_stream_act_local_6 <= 0;
          if(cparam_conv2d_16_stream_act_local_small_flags_0) begin
            conv2d_16_stream_act_local_6 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_16_stream_act_local_large_flags_0) begin
            conv2d_16_stream_act_local_6 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          conv2d_16_stream_act_local_7 <= 0;
          if(cparam_conv2d_16_stream_act_local_small_flags_1) begin
            conv2d_16_stream_act_local_7 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_16_stream_act_local_large_flags_1) begin
            conv2d_16_stream_act_local_7 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          conv2d_16_stream_act_local_8 <= 0;
          if(cparam_conv2d_16_stream_act_local_small_flags_2) begin
            conv2d_16_stream_act_local_8 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_16_stream_act_local_large_flags_2) begin
            conv2d_16_stream_act_local_8 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          conv2d_16_stream_out_local_col <= 0;
          if((cparam_conv2d_16_data_stationary == 1) && (conv2d_16_och_count == 0)) begin
            conv2d_16_stream_out_local_val <= 0;
          end 
          conv2d_16_col_count <= 0;
          conv2d_16_col_select <= cparam_conv2d_16_col_select_initval;
          conv2d_16_filter_page_comp_offset_buf <= conv2d_16_filter_page_comp_offset;
          conv2d_16_act_page_comp_offset_buf_0 <= conv2d_16_act_page_comp_offset_0;
          conv2d_16_act_page_comp_offset_buf_1 <= conv2d_16_act_page_comp_offset_1;
          conv2d_16_act_page_comp_offset_buf_2 <= conv2d_16_act_page_comp_offset_2;
          conv2d_16_out_page_comp_offset_buf <= conv2d_16_out_page_comp_offset;
          conv2d_16_row_count_buf <= conv2d_16_row_count;
          conv2d_16_row_select_buf <= conv2d_16_row_select;
          conv2d_16_och_count_buf <= conv2d_16_och_count;
          conv2d_16_next_stream_num_ops <= (conv2d_16_och_count >= cparam_conv2d_16_max_och_count)? cparam_conv2d_16_stream_num_ops_res : cparam_conv2d_16_stream_num_ops;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_2;
        end
        conv2d_16_comp_fsm_2: begin
          conv2d_16_stream_pad_masks <= { conv2d_16_stream_pad_mask_2_2, conv2d_16_stream_pad_mask_2_1, conv2d_16_stream_pad_mask_2_0, conv2d_16_stream_pad_mask_1_2, conv2d_16_stream_pad_mask_1_1, conv2d_16_stream_pad_mask_1_0, conv2d_16_stream_pad_mask_0_2, conv2d_16_stream_pad_mask_0_1, conv2d_16_stream_pad_mask_0_0 };
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_3;
        end
        conv2d_16_comp_fsm_3: begin
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_4;
        end
        conv2d_16_comp_fsm_4: begin
          if(!_stream_conv2d_16_source_busy) begin
            conv2d_16_comp_fsm <= conv2d_16_comp_fsm_5;
          end 
        end
        conv2d_16_comp_fsm_5: begin
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_6;
        end
        conv2d_16_comp_fsm_6: begin
          if(!((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_0 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_1 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_2 : 0)) begin
            conv2d_16_stream_act_local_0 <= conv2d_16_stream_act_local_0 + cparam_conv2d_16_inc_act_laddr_small;
          end 
          if((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_0 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_1 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_2 : 0) begin
            conv2d_16_stream_act_local_0 <= conv2d_16_stream_act_local_0 + cparam_conv2d_16_inc_act_laddr_large;
          end 
          if(conv2d_16_col_count >= cparam_conv2d_16_max_col_count) begin
            conv2d_16_stream_act_local_0 <= 0;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_small_flags_0) begin
            conv2d_16_stream_act_local_0 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_large_flags_0) begin
            conv2d_16_stream_act_local_0 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          if(!((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_3 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_4 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_5 : 0)) begin
            conv2d_16_stream_act_local_1 <= conv2d_16_stream_act_local_1 + cparam_conv2d_16_inc_act_laddr_small;
          end 
          if((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_3 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_4 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_5 : 0) begin
            conv2d_16_stream_act_local_1 <= conv2d_16_stream_act_local_1 + cparam_conv2d_16_inc_act_laddr_large;
          end 
          if(conv2d_16_col_count >= cparam_conv2d_16_max_col_count) begin
            conv2d_16_stream_act_local_1 <= 0;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_small_flags_1) begin
            conv2d_16_stream_act_local_1 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_large_flags_1) begin
            conv2d_16_stream_act_local_1 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          if(!((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_6 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_7 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_8 : 0)) begin
            conv2d_16_stream_act_local_2 <= conv2d_16_stream_act_local_2 + cparam_conv2d_16_inc_act_laddr_small;
          end 
          if((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_6 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_7 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_8 : 0) begin
            conv2d_16_stream_act_local_2 <= conv2d_16_stream_act_local_2 + cparam_conv2d_16_inc_act_laddr_large;
          end 
          if(conv2d_16_col_count >= cparam_conv2d_16_max_col_count) begin
            conv2d_16_stream_act_local_2 <= 0;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_small_flags_2) begin
            conv2d_16_stream_act_local_2 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_large_flags_2) begin
            conv2d_16_stream_act_local_2 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          if(!((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_9 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_10 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_11 : 0)) begin
            conv2d_16_stream_act_local_3 <= conv2d_16_stream_act_local_3 + cparam_conv2d_16_inc_act_laddr_small;
          end 
          if((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_9 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_10 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_11 : 0) begin
            conv2d_16_stream_act_local_3 <= conv2d_16_stream_act_local_3 + cparam_conv2d_16_inc_act_laddr_large;
          end 
          if(conv2d_16_col_count >= cparam_conv2d_16_max_col_count) begin
            conv2d_16_stream_act_local_3 <= 0;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_small_flags_0) begin
            conv2d_16_stream_act_local_3 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_large_flags_0) begin
            conv2d_16_stream_act_local_3 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          if(!((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_12 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_13 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_14 : 0)) begin
            conv2d_16_stream_act_local_4 <= conv2d_16_stream_act_local_4 + cparam_conv2d_16_inc_act_laddr_small;
          end 
          if((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_12 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_13 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_14 : 0) begin
            conv2d_16_stream_act_local_4 <= conv2d_16_stream_act_local_4 + cparam_conv2d_16_inc_act_laddr_large;
          end 
          if(conv2d_16_col_count >= cparam_conv2d_16_max_col_count) begin
            conv2d_16_stream_act_local_4 <= 0;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_small_flags_1) begin
            conv2d_16_stream_act_local_4 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_large_flags_1) begin
            conv2d_16_stream_act_local_4 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          if(!((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_15 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_16 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_17 : 0)) begin
            conv2d_16_stream_act_local_5 <= conv2d_16_stream_act_local_5 + cparam_conv2d_16_inc_act_laddr_small;
          end 
          if((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_15 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_16 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_17 : 0) begin
            conv2d_16_stream_act_local_5 <= conv2d_16_stream_act_local_5 + cparam_conv2d_16_inc_act_laddr_large;
          end 
          if(conv2d_16_col_count >= cparam_conv2d_16_max_col_count) begin
            conv2d_16_stream_act_local_5 <= 0;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_small_flags_2) begin
            conv2d_16_stream_act_local_5 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_large_flags_2) begin
            conv2d_16_stream_act_local_5 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          if(!((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_18 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_19 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_20 : 0)) begin
            conv2d_16_stream_act_local_6 <= conv2d_16_stream_act_local_6 + cparam_conv2d_16_inc_act_laddr_small;
          end 
          if((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_18 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_19 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_20 : 0) begin
            conv2d_16_stream_act_local_6 <= conv2d_16_stream_act_local_6 + cparam_conv2d_16_inc_act_laddr_large;
          end 
          if(conv2d_16_col_count >= cparam_conv2d_16_max_col_count) begin
            conv2d_16_stream_act_local_6 <= 0;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_small_flags_0) begin
            conv2d_16_stream_act_local_6 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_large_flags_0) begin
            conv2d_16_stream_act_local_6 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          if(!((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_21 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_22 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_23 : 0)) begin
            conv2d_16_stream_act_local_7 <= conv2d_16_stream_act_local_7 + cparam_conv2d_16_inc_act_laddr_small;
          end 
          if((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_21 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_22 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_23 : 0) begin
            conv2d_16_stream_act_local_7 <= conv2d_16_stream_act_local_7 + cparam_conv2d_16_inc_act_laddr_large;
          end 
          if(conv2d_16_col_count >= cparam_conv2d_16_max_col_count) begin
            conv2d_16_stream_act_local_7 <= 0;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_small_flags_1) begin
            conv2d_16_stream_act_local_7 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_large_flags_1) begin
            conv2d_16_stream_act_local_7 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          if(!((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_24 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_25 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_26 : 0)) begin
            conv2d_16_stream_act_local_8 <= conv2d_16_stream_act_local_8 + cparam_conv2d_16_inc_act_laddr_small;
          end 
          if((conv2d_16_col_select == 0)? cparam_conv2d_16_inc_act_laddr_conds_24 : 
          (conv2d_16_col_select == 1)? cparam_conv2d_16_inc_act_laddr_conds_25 : 
          (conv2d_16_col_select == 2)? cparam_conv2d_16_inc_act_laddr_conds_26 : 0) begin
            conv2d_16_stream_act_local_8 <= conv2d_16_stream_act_local_8 + cparam_conv2d_16_inc_act_laddr_large;
          end 
          if(conv2d_16_col_count >= cparam_conv2d_16_max_col_count) begin
            conv2d_16_stream_act_local_8 <= 0;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_small_flags_2) begin
            conv2d_16_stream_act_local_8 <= cparam_conv2d_16_stream_act_local_small_offset;
          end 
          if((conv2d_16_col_count >= cparam_conv2d_16_max_col_count) && cparam_conv2d_16_stream_act_local_large_flags_2) begin
            conv2d_16_stream_act_local_8 <= cparam_conv2d_16_stream_act_local_large_offset;
          end 
          if(cparam_conv2d_16_data_stationary == 0) begin
            conv2d_16_stream_out_local_col <= conv2d_16_stream_out_local_col + conv2d_16_next_stream_num_ops;
          end 
          if((cparam_conv2d_16_data_stationary == 0) && (conv2d_16_col_count >= cparam_conv2d_16_max_col_count)) begin
            conv2d_16_stream_out_local_col <= 0;
          end 
          if(cparam_conv2d_16_data_stationary == 1) begin
            conv2d_16_stream_out_local_col <= conv2d_16_stream_out_local_col + cparam_conv2d_16_inc_out_laddr_col;
          end 
          if((cparam_conv2d_16_data_stationary == 1) && (conv2d_16_col_count >= cparam_conv2d_16_max_col_count)) begin
            conv2d_16_stream_out_local_val <= conv2d_16_stream_out_local_val + conv2d_16_next_stream_num_ops;
            conv2d_16_stream_out_local_col <= 0;
          end 
          conv2d_16_col_count <= conv2d_16_col_count + cparam_conv2d_16_stride_col_par_col;
          if(conv2d_16_col_count >= cparam_conv2d_16_max_col_count) begin
            conv2d_16_col_count <= 0;
          end 
          conv2d_16_col_select <= conv2d_16_col_select + cparam_conv2d_16_stride_col_mod_filter_num;
          if(conv2d_16_col_select + cparam_conv2d_16_stride_col_mod_filter_num >= 3) begin
            conv2d_16_col_select <= conv2d_16_col_select - cparam_conv2d_16_filter_num_col_minus_stride_col_mod;
          end 
          if(conv2d_16_col_count >= cparam_conv2d_16_max_col_count) begin
            conv2d_16_col_select <= cparam_conv2d_16_col_select_initval;
          end 
          conv2d_16_comp_fsm <= conv2d_16_comp_fsm_2;
          if(conv2d_16_col_count >= cparam_conv2d_16_max_col_count) begin
            conv2d_16_comp_fsm <= conv2d_16_comp_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_464_1 <= 0;
      __tmp_464_2 <= 0;
      __tmp_1027_1 <= 0;
      __tmp_1027_2 <= 0;
    end else begin
      __tmp_464_1 <= _tmp_464;
      __tmp_464_2 <= __tmp_464_1;
      __tmp_1027_1 <= _tmp_1027;
      __tmp_1027_2 <= __tmp_1027_1;
    end
  end

  localparam _stream_conv2d_16_source_6_source_pat_fsm_0_1 = 1;
  localparam _stream_conv2d_16_source_6_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_6_source_pat_fsm_0 <= _stream_conv2d_16_source_6_source_pat_fsm_0_init;
    end else begin
      case(_stream_conv2d_16_source_6_source_pat_fsm_0)
        _stream_conv2d_16_source_6_source_pat_fsm_0_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_6_source_mode & 3'b10) begin
            _stream_conv2d_16_source_6_source_pat_fsm_0 <= _stream_conv2d_16_source_6_source_pat_fsm_0_1;
          end 
        end
        _stream_conv2d_16_source_6_source_pat_fsm_0_1: begin
          if((_source_stream_conv2d_16_source_6_pat_count_0 == 0) && (_source_stream_conv2d_16_source_6_pat_count_1 == 0) && (_source_stream_conv2d_16_source_6_pat_count_2 == 0) && (_source_stream_conv2d_16_source_6_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_6_source_pat_fsm_0 <= _stream_conv2d_16_source_6_source_pat_fsm_0_2;
          end 
        end
        _stream_conv2d_16_source_6_source_pat_fsm_0_2: begin
          _stream_conv2d_16_source_6_source_pat_fsm_0 <= _stream_conv2d_16_source_6_source_pat_fsm_0_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_475_1 <= 0;
      __tmp_475_2 <= 0;
      __tmp_1181_1 <= 0;
      __tmp_1181_2 <= 0;
    end else begin
      __tmp_475_1 <= _tmp_475;
      __tmp_475_2 <= __tmp_475_1;
      __tmp_1181_1 <= _tmp_1181;
      __tmp_1181_2 <= __tmp_1181_1;
    end
  end

  localparam _stream_conv2d_16_source_8_source_pat_fsm_1_1 = 1;
  localparam _stream_conv2d_16_source_8_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_8_source_pat_fsm_1 <= _stream_conv2d_16_source_8_source_pat_fsm_1_init;
    end else begin
      case(_stream_conv2d_16_source_8_source_pat_fsm_1)
        _stream_conv2d_16_source_8_source_pat_fsm_1_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_8_source_mode & 3'b10) begin
            _stream_conv2d_16_source_8_source_pat_fsm_1 <= _stream_conv2d_16_source_8_source_pat_fsm_1_1;
          end 
        end
        _stream_conv2d_16_source_8_source_pat_fsm_1_1: begin
          if((_source_stream_conv2d_16_source_8_pat_count_0 == 0) && (_source_stream_conv2d_16_source_8_pat_count_1 == 0) && (_source_stream_conv2d_16_source_8_pat_count_2 == 0) && (_source_stream_conv2d_16_source_8_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_8_source_pat_fsm_1 <= _stream_conv2d_16_source_8_source_pat_fsm_1_2;
          end 
        end
        _stream_conv2d_16_source_8_source_pat_fsm_1_2: begin
          _stream_conv2d_16_source_8_source_pat_fsm_1 <= _stream_conv2d_16_source_8_source_pat_fsm_1_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_495_1 <= 0;
      __tmp_495_2 <= 0;
      __tmp_1170_1 <= 0;
      __tmp_1170_2 <= 0;
    end else begin
      __tmp_495_1 <= _tmp_495;
      __tmp_495_2 <= __tmp_495_1;
      __tmp_1170_1 <= _tmp_1170;
      __tmp_1170_2 <= __tmp_1170_1;
    end
  end

  localparam _stream_conv2d_16_source_19_source_pat_fsm_2_1 = 1;
  localparam _stream_conv2d_16_source_19_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_19_source_pat_fsm_2 <= _stream_conv2d_16_source_19_source_pat_fsm_2_init;
    end else begin
      case(_stream_conv2d_16_source_19_source_pat_fsm_2)
        _stream_conv2d_16_source_19_source_pat_fsm_2_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_19_source_mode & 3'b10) begin
            _stream_conv2d_16_source_19_source_pat_fsm_2 <= _stream_conv2d_16_source_19_source_pat_fsm_2_1;
          end 
        end
        _stream_conv2d_16_source_19_source_pat_fsm_2_1: begin
          if((_source_stream_conv2d_16_source_19_pat_count_0 == 0) && (_source_stream_conv2d_16_source_19_pat_count_1 == 0) && (_source_stream_conv2d_16_source_19_pat_count_2 == 0) && (_source_stream_conv2d_16_source_19_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_19_source_pat_fsm_2 <= _stream_conv2d_16_source_19_source_pat_fsm_2_2;
          end 
        end
        _stream_conv2d_16_source_19_source_pat_fsm_2_2: begin
          _stream_conv2d_16_source_19_source_pat_fsm_2 <= _stream_conv2d_16_source_19_source_pat_fsm_2_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_505_1 <= 0;
      __tmp_505_2 <= 0;
      __tmp_1201_1 <= 0;
      __tmp_1201_2 <= 0;
    end else begin
      __tmp_505_1 <= _tmp_505;
      __tmp_505_2 <= __tmp_505_1;
      __tmp_1201_1 <= _tmp_1201;
      __tmp_1201_2 <= __tmp_1201_1;
    end
  end

  localparam _stream_conv2d_16_source_20_source_pat_fsm_3_1 = 1;
  localparam _stream_conv2d_16_source_20_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_20_source_pat_fsm_3 <= _stream_conv2d_16_source_20_source_pat_fsm_3_init;
    end else begin
      case(_stream_conv2d_16_source_20_source_pat_fsm_3)
        _stream_conv2d_16_source_20_source_pat_fsm_3_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_20_source_mode & 3'b10) begin
            _stream_conv2d_16_source_20_source_pat_fsm_3 <= _stream_conv2d_16_source_20_source_pat_fsm_3_1;
          end 
        end
        _stream_conv2d_16_source_20_source_pat_fsm_3_1: begin
          if((_source_stream_conv2d_16_source_20_pat_count_0 == 0) && (_source_stream_conv2d_16_source_20_pat_count_1 == 0) && (_source_stream_conv2d_16_source_20_pat_count_2 == 0) && (_source_stream_conv2d_16_source_20_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_20_source_pat_fsm_3 <= _stream_conv2d_16_source_20_source_pat_fsm_3_2;
          end 
        end
        _stream_conv2d_16_source_20_source_pat_fsm_3_2: begin
          _stream_conv2d_16_source_20_source_pat_fsm_3 <= _stream_conv2d_16_source_20_source_pat_fsm_3_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_515_1 <= 0;
      __tmp_515_2 <= 0;
    end else begin
      __tmp_515_1 <= _tmp_515;
      __tmp_515_2 <= __tmp_515_1;
    end
  end

  localparam _stream_conv2d_16_source_21_source_pat_fsm_4_1 = 1;
  localparam _stream_conv2d_16_source_21_source_pat_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_21_source_pat_fsm_4 <= _stream_conv2d_16_source_21_source_pat_fsm_4_init;
    end else begin
      case(_stream_conv2d_16_source_21_source_pat_fsm_4)
        _stream_conv2d_16_source_21_source_pat_fsm_4_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_21_source_mode & 3'b10) begin
            _stream_conv2d_16_source_21_source_pat_fsm_4 <= _stream_conv2d_16_source_21_source_pat_fsm_4_1;
          end 
        end
        _stream_conv2d_16_source_21_source_pat_fsm_4_1: begin
          if((_source_stream_conv2d_16_source_21_pat_count_0 == 0) && (_source_stream_conv2d_16_source_21_pat_count_1 == 0) && (_source_stream_conv2d_16_source_21_pat_count_2 == 0) && (_source_stream_conv2d_16_source_21_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_21_source_pat_fsm_4 <= _stream_conv2d_16_source_21_source_pat_fsm_4_2;
          end 
        end
        _stream_conv2d_16_source_21_source_pat_fsm_4_2: begin
          _stream_conv2d_16_source_21_source_pat_fsm_4 <= _stream_conv2d_16_source_21_source_pat_fsm_4_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_525_1 <= 0;
      __tmp_525_2 <= 0;
    end else begin
      __tmp_525_1 <= _tmp_525;
      __tmp_525_2 <= __tmp_525_1;
    end
  end

  localparam _stream_conv2d_16_source_22_source_pat_fsm_5_1 = 1;
  localparam _stream_conv2d_16_source_22_source_pat_fsm_5_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_22_source_pat_fsm_5 <= _stream_conv2d_16_source_22_source_pat_fsm_5_init;
    end else begin
      case(_stream_conv2d_16_source_22_source_pat_fsm_5)
        _stream_conv2d_16_source_22_source_pat_fsm_5_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_22_source_mode & 3'b10) begin
            _stream_conv2d_16_source_22_source_pat_fsm_5 <= _stream_conv2d_16_source_22_source_pat_fsm_5_1;
          end 
        end
        _stream_conv2d_16_source_22_source_pat_fsm_5_1: begin
          if((_source_stream_conv2d_16_source_22_pat_count_0 == 0) && (_source_stream_conv2d_16_source_22_pat_count_1 == 0) && (_source_stream_conv2d_16_source_22_pat_count_2 == 0) && (_source_stream_conv2d_16_source_22_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_22_source_pat_fsm_5 <= _stream_conv2d_16_source_22_source_pat_fsm_5_2;
          end 
        end
        _stream_conv2d_16_source_22_source_pat_fsm_5_2: begin
          _stream_conv2d_16_source_22_source_pat_fsm_5 <= _stream_conv2d_16_source_22_source_pat_fsm_5_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_535_1 <= 0;
      __tmp_535_2 <= 0;
    end else begin
      __tmp_535_1 <= _tmp_535;
      __tmp_535_2 <= __tmp_535_1;
    end
  end

  localparam _stream_conv2d_16_source_23_source_pat_fsm_6_1 = 1;
  localparam _stream_conv2d_16_source_23_source_pat_fsm_6_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_23_source_pat_fsm_6 <= _stream_conv2d_16_source_23_source_pat_fsm_6_init;
    end else begin
      case(_stream_conv2d_16_source_23_source_pat_fsm_6)
        _stream_conv2d_16_source_23_source_pat_fsm_6_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_23_source_mode & 3'b10) begin
            _stream_conv2d_16_source_23_source_pat_fsm_6 <= _stream_conv2d_16_source_23_source_pat_fsm_6_1;
          end 
        end
        _stream_conv2d_16_source_23_source_pat_fsm_6_1: begin
          if((_source_stream_conv2d_16_source_23_pat_count_0 == 0) && (_source_stream_conv2d_16_source_23_pat_count_1 == 0) && (_source_stream_conv2d_16_source_23_pat_count_2 == 0) && (_source_stream_conv2d_16_source_23_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_23_source_pat_fsm_6 <= _stream_conv2d_16_source_23_source_pat_fsm_6_2;
          end 
        end
        _stream_conv2d_16_source_23_source_pat_fsm_6_2: begin
          _stream_conv2d_16_source_23_source_pat_fsm_6 <= _stream_conv2d_16_source_23_source_pat_fsm_6_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_545_1 <= 0;
      __tmp_545_2 <= 0;
    end else begin
      __tmp_545_1 <= _tmp_545;
      __tmp_545_2 <= __tmp_545_1;
    end
  end

  localparam _stream_conv2d_16_source_24_source_pat_fsm_7_1 = 1;
  localparam _stream_conv2d_16_source_24_source_pat_fsm_7_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_24_source_pat_fsm_7 <= _stream_conv2d_16_source_24_source_pat_fsm_7_init;
    end else begin
      case(_stream_conv2d_16_source_24_source_pat_fsm_7)
        _stream_conv2d_16_source_24_source_pat_fsm_7_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_24_source_mode & 3'b10) begin
            _stream_conv2d_16_source_24_source_pat_fsm_7 <= _stream_conv2d_16_source_24_source_pat_fsm_7_1;
          end 
        end
        _stream_conv2d_16_source_24_source_pat_fsm_7_1: begin
          if((_source_stream_conv2d_16_source_24_pat_count_0 == 0) && (_source_stream_conv2d_16_source_24_pat_count_1 == 0) && (_source_stream_conv2d_16_source_24_pat_count_2 == 0) && (_source_stream_conv2d_16_source_24_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_24_source_pat_fsm_7 <= _stream_conv2d_16_source_24_source_pat_fsm_7_2;
          end 
        end
        _stream_conv2d_16_source_24_source_pat_fsm_7_2: begin
          _stream_conv2d_16_source_24_source_pat_fsm_7 <= _stream_conv2d_16_source_24_source_pat_fsm_7_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_555_1 <= 0;
      __tmp_555_2 <= 0;
    end else begin
      __tmp_555_1 <= _tmp_555;
      __tmp_555_2 <= __tmp_555_1;
    end
  end

  localparam _stream_conv2d_16_source_25_source_pat_fsm_8_1 = 1;
  localparam _stream_conv2d_16_source_25_source_pat_fsm_8_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_25_source_pat_fsm_8 <= _stream_conv2d_16_source_25_source_pat_fsm_8_init;
    end else begin
      case(_stream_conv2d_16_source_25_source_pat_fsm_8)
        _stream_conv2d_16_source_25_source_pat_fsm_8_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_25_source_mode & 3'b10) begin
            _stream_conv2d_16_source_25_source_pat_fsm_8 <= _stream_conv2d_16_source_25_source_pat_fsm_8_1;
          end 
        end
        _stream_conv2d_16_source_25_source_pat_fsm_8_1: begin
          if((_source_stream_conv2d_16_source_25_pat_count_0 == 0) && (_source_stream_conv2d_16_source_25_pat_count_1 == 0) && (_source_stream_conv2d_16_source_25_pat_count_2 == 0) && (_source_stream_conv2d_16_source_25_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_25_source_pat_fsm_8 <= _stream_conv2d_16_source_25_source_pat_fsm_8_2;
          end 
        end
        _stream_conv2d_16_source_25_source_pat_fsm_8_2: begin
          _stream_conv2d_16_source_25_source_pat_fsm_8 <= _stream_conv2d_16_source_25_source_pat_fsm_8_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_565_1 <= 0;
      __tmp_565_2 <= 0;
    end else begin
      __tmp_565_1 <= _tmp_565;
      __tmp_565_2 <= __tmp_565_1;
    end
  end

  localparam _stream_conv2d_16_source_26_source_pat_fsm_9_1 = 1;
  localparam _stream_conv2d_16_source_26_source_pat_fsm_9_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_26_source_pat_fsm_9 <= _stream_conv2d_16_source_26_source_pat_fsm_9_init;
    end else begin
      case(_stream_conv2d_16_source_26_source_pat_fsm_9)
        _stream_conv2d_16_source_26_source_pat_fsm_9_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_26_source_mode & 3'b10) begin
            _stream_conv2d_16_source_26_source_pat_fsm_9 <= _stream_conv2d_16_source_26_source_pat_fsm_9_1;
          end 
        end
        _stream_conv2d_16_source_26_source_pat_fsm_9_1: begin
          if((_source_stream_conv2d_16_source_26_pat_count_0 == 0) && (_source_stream_conv2d_16_source_26_pat_count_1 == 0) && (_source_stream_conv2d_16_source_26_pat_count_2 == 0) && (_source_stream_conv2d_16_source_26_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_26_source_pat_fsm_9 <= _stream_conv2d_16_source_26_source_pat_fsm_9_2;
          end 
        end
        _stream_conv2d_16_source_26_source_pat_fsm_9_2: begin
          _stream_conv2d_16_source_26_source_pat_fsm_9 <= _stream_conv2d_16_source_26_source_pat_fsm_9_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_575_1 <= 0;
      __tmp_575_2 <= 0;
    end else begin
      __tmp_575_1 <= _tmp_575;
      __tmp_575_2 <= __tmp_575_1;
    end
  end

  localparam _stream_conv2d_16_source_27_source_pat_fsm_10_1 = 1;
  localparam _stream_conv2d_16_source_27_source_pat_fsm_10_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_27_source_pat_fsm_10 <= _stream_conv2d_16_source_27_source_pat_fsm_10_init;
    end else begin
      case(_stream_conv2d_16_source_27_source_pat_fsm_10)
        _stream_conv2d_16_source_27_source_pat_fsm_10_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_27_source_mode & 3'b10) begin
            _stream_conv2d_16_source_27_source_pat_fsm_10 <= _stream_conv2d_16_source_27_source_pat_fsm_10_1;
          end 
        end
        _stream_conv2d_16_source_27_source_pat_fsm_10_1: begin
          if((_source_stream_conv2d_16_source_27_pat_count_0 == 0) && (_source_stream_conv2d_16_source_27_pat_count_1 == 0) && (_source_stream_conv2d_16_source_27_pat_count_2 == 0) && (_source_stream_conv2d_16_source_27_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_27_source_pat_fsm_10 <= _stream_conv2d_16_source_27_source_pat_fsm_10_2;
          end 
        end
        _stream_conv2d_16_source_27_source_pat_fsm_10_2: begin
          _stream_conv2d_16_source_27_source_pat_fsm_10 <= _stream_conv2d_16_source_27_source_pat_fsm_10_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_585_1 <= 0;
      __tmp_585_2 <= 0;
      __tmp_1211_1 <= 0;
      __tmp_1211_2 <= 0;
    end else begin
      __tmp_585_1 <= _tmp_585;
      __tmp_585_2 <= __tmp_585_1;
      __tmp_1211_1 <= _tmp_1211;
      __tmp_1211_2 <= __tmp_1211_1;
    end
  end

  localparam _stream_conv2d_16_source_28_source_pat_fsm_11_1 = 1;
  localparam _stream_conv2d_16_source_28_source_pat_fsm_11_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_28_source_pat_fsm_11 <= _stream_conv2d_16_source_28_source_pat_fsm_11_init;
    end else begin
      case(_stream_conv2d_16_source_28_source_pat_fsm_11)
        _stream_conv2d_16_source_28_source_pat_fsm_11_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_28_source_mode & 3'b10) begin
            _stream_conv2d_16_source_28_source_pat_fsm_11 <= _stream_conv2d_16_source_28_source_pat_fsm_11_1;
          end 
        end
        _stream_conv2d_16_source_28_source_pat_fsm_11_1: begin
          if((_source_stream_conv2d_16_source_28_pat_count_0 == 0) && (_source_stream_conv2d_16_source_28_pat_count_1 == 0) && (_source_stream_conv2d_16_source_28_pat_count_2 == 0) && (_source_stream_conv2d_16_source_28_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_28_source_pat_fsm_11 <= _stream_conv2d_16_source_28_source_pat_fsm_11_2;
          end 
        end
        _stream_conv2d_16_source_28_source_pat_fsm_11_2: begin
          _stream_conv2d_16_source_28_source_pat_fsm_11 <= _stream_conv2d_16_source_28_source_pat_fsm_11_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_599_1 <= 0;
      __tmp_599_2 <= 0;
    end else begin
      __tmp_599_1 <= _tmp_599;
      __tmp_599_2 <= __tmp_599_1;
    end
  end

  localparam _stream_conv2d_16_source_29_source_pat_fsm_12_1 = 1;
  localparam _stream_conv2d_16_source_29_source_pat_fsm_12_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_29_source_pat_fsm_12 <= _stream_conv2d_16_source_29_source_pat_fsm_12_init;
    end else begin
      case(_stream_conv2d_16_source_29_source_pat_fsm_12)
        _stream_conv2d_16_source_29_source_pat_fsm_12_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_29_source_mode & 3'b10) begin
            _stream_conv2d_16_source_29_source_pat_fsm_12 <= _stream_conv2d_16_source_29_source_pat_fsm_12_1;
          end 
        end
        _stream_conv2d_16_source_29_source_pat_fsm_12_1: begin
          if((_source_stream_conv2d_16_source_29_pat_count_0 == 0) && (_source_stream_conv2d_16_source_29_pat_count_1 == 0) && (_source_stream_conv2d_16_source_29_pat_count_2 == 0) && (_source_stream_conv2d_16_source_29_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_29_source_pat_fsm_12 <= _stream_conv2d_16_source_29_source_pat_fsm_12_2;
          end 
        end
        _stream_conv2d_16_source_29_source_pat_fsm_12_2: begin
          _stream_conv2d_16_source_29_source_pat_fsm_12 <= _stream_conv2d_16_source_29_source_pat_fsm_12_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_613_1 <= 0;
      __tmp_613_2 <= 0;
    end else begin
      __tmp_613_1 <= _tmp_613;
      __tmp_613_2 <= __tmp_613_1;
    end
  end

  localparam _stream_conv2d_16_source_30_source_pat_fsm_13_1 = 1;
  localparam _stream_conv2d_16_source_30_source_pat_fsm_13_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_30_source_pat_fsm_13 <= _stream_conv2d_16_source_30_source_pat_fsm_13_init;
    end else begin
      case(_stream_conv2d_16_source_30_source_pat_fsm_13)
        _stream_conv2d_16_source_30_source_pat_fsm_13_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_30_source_mode & 3'b10) begin
            _stream_conv2d_16_source_30_source_pat_fsm_13 <= _stream_conv2d_16_source_30_source_pat_fsm_13_1;
          end 
        end
        _stream_conv2d_16_source_30_source_pat_fsm_13_1: begin
          if((_source_stream_conv2d_16_source_30_pat_count_0 == 0) && (_source_stream_conv2d_16_source_30_pat_count_1 == 0) && (_source_stream_conv2d_16_source_30_pat_count_2 == 0) && (_source_stream_conv2d_16_source_30_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_30_source_pat_fsm_13 <= _stream_conv2d_16_source_30_source_pat_fsm_13_2;
          end 
        end
        _stream_conv2d_16_source_30_source_pat_fsm_13_2: begin
          _stream_conv2d_16_source_30_source_pat_fsm_13 <= _stream_conv2d_16_source_30_source_pat_fsm_13_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_627_1 <= 0;
      __tmp_627_2 <= 0;
    end else begin
      __tmp_627_1 <= _tmp_627;
      __tmp_627_2 <= __tmp_627_1;
    end
  end

  localparam _stream_conv2d_16_source_31_source_pat_fsm_14_1 = 1;
  localparam _stream_conv2d_16_source_31_source_pat_fsm_14_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_31_source_pat_fsm_14 <= _stream_conv2d_16_source_31_source_pat_fsm_14_init;
    end else begin
      case(_stream_conv2d_16_source_31_source_pat_fsm_14)
        _stream_conv2d_16_source_31_source_pat_fsm_14_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_31_source_mode & 3'b10) begin
            _stream_conv2d_16_source_31_source_pat_fsm_14 <= _stream_conv2d_16_source_31_source_pat_fsm_14_1;
          end 
        end
        _stream_conv2d_16_source_31_source_pat_fsm_14_1: begin
          if((_source_stream_conv2d_16_source_31_pat_count_0 == 0) && (_source_stream_conv2d_16_source_31_pat_count_1 == 0) && (_source_stream_conv2d_16_source_31_pat_count_2 == 0) && (_source_stream_conv2d_16_source_31_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_31_source_pat_fsm_14 <= _stream_conv2d_16_source_31_source_pat_fsm_14_2;
          end 
        end
        _stream_conv2d_16_source_31_source_pat_fsm_14_2: begin
          _stream_conv2d_16_source_31_source_pat_fsm_14 <= _stream_conv2d_16_source_31_source_pat_fsm_14_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_641_1 <= 0;
      __tmp_641_2 <= 0;
    end else begin
      __tmp_641_1 <= _tmp_641;
      __tmp_641_2 <= __tmp_641_1;
    end
  end

  localparam _stream_conv2d_16_source_32_source_pat_fsm_15_1 = 1;
  localparam _stream_conv2d_16_source_32_source_pat_fsm_15_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_32_source_pat_fsm_15 <= _stream_conv2d_16_source_32_source_pat_fsm_15_init;
    end else begin
      case(_stream_conv2d_16_source_32_source_pat_fsm_15)
        _stream_conv2d_16_source_32_source_pat_fsm_15_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_32_source_mode & 3'b10) begin
            _stream_conv2d_16_source_32_source_pat_fsm_15 <= _stream_conv2d_16_source_32_source_pat_fsm_15_1;
          end 
        end
        _stream_conv2d_16_source_32_source_pat_fsm_15_1: begin
          if((_source_stream_conv2d_16_source_32_pat_count_0 == 0) && (_source_stream_conv2d_16_source_32_pat_count_1 == 0) && (_source_stream_conv2d_16_source_32_pat_count_2 == 0) && (_source_stream_conv2d_16_source_32_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_32_source_pat_fsm_15 <= _stream_conv2d_16_source_32_source_pat_fsm_15_2;
          end 
        end
        _stream_conv2d_16_source_32_source_pat_fsm_15_2: begin
          _stream_conv2d_16_source_32_source_pat_fsm_15 <= _stream_conv2d_16_source_32_source_pat_fsm_15_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_655_1 <= 0;
      __tmp_655_2 <= 0;
    end else begin
      __tmp_655_1 <= _tmp_655;
      __tmp_655_2 <= __tmp_655_1;
    end
  end

  localparam _stream_conv2d_16_source_33_source_pat_fsm_16_1 = 1;
  localparam _stream_conv2d_16_source_33_source_pat_fsm_16_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_33_source_pat_fsm_16 <= _stream_conv2d_16_source_33_source_pat_fsm_16_init;
    end else begin
      case(_stream_conv2d_16_source_33_source_pat_fsm_16)
        _stream_conv2d_16_source_33_source_pat_fsm_16_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_33_source_mode & 3'b10) begin
            _stream_conv2d_16_source_33_source_pat_fsm_16 <= _stream_conv2d_16_source_33_source_pat_fsm_16_1;
          end 
        end
        _stream_conv2d_16_source_33_source_pat_fsm_16_1: begin
          if((_source_stream_conv2d_16_source_33_pat_count_0 == 0) && (_source_stream_conv2d_16_source_33_pat_count_1 == 0) && (_source_stream_conv2d_16_source_33_pat_count_2 == 0) && (_source_stream_conv2d_16_source_33_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_33_source_pat_fsm_16 <= _stream_conv2d_16_source_33_source_pat_fsm_16_2;
          end 
        end
        _stream_conv2d_16_source_33_source_pat_fsm_16_2: begin
          _stream_conv2d_16_source_33_source_pat_fsm_16 <= _stream_conv2d_16_source_33_source_pat_fsm_16_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_669_1 <= 0;
      __tmp_669_2 <= 0;
    end else begin
      __tmp_669_1 <= _tmp_669;
      __tmp_669_2 <= __tmp_669_1;
    end
  end

  localparam _stream_conv2d_16_source_34_source_pat_fsm_17_1 = 1;
  localparam _stream_conv2d_16_source_34_source_pat_fsm_17_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_34_source_pat_fsm_17 <= _stream_conv2d_16_source_34_source_pat_fsm_17_init;
    end else begin
      case(_stream_conv2d_16_source_34_source_pat_fsm_17)
        _stream_conv2d_16_source_34_source_pat_fsm_17_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_34_source_mode & 3'b10) begin
            _stream_conv2d_16_source_34_source_pat_fsm_17 <= _stream_conv2d_16_source_34_source_pat_fsm_17_1;
          end 
        end
        _stream_conv2d_16_source_34_source_pat_fsm_17_1: begin
          if((_source_stream_conv2d_16_source_34_pat_count_0 == 0) && (_source_stream_conv2d_16_source_34_pat_count_1 == 0) && (_source_stream_conv2d_16_source_34_pat_count_2 == 0) && (_source_stream_conv2d_16_source_34_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_34_source_pat_fsm_17 <= _stream_conv2d_16_source_34_source_pat_fsm_17_2;
          end 
        end
        _stream_conv2d_16_source_34_source_pat_fsm_17_2: begin
          _stream_conv2d_16_source_34_source_pat_fsm_17 <= _stream_conv2d_16_source_34_source_pat_fsm_17_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_683_1 <= 0;
      __tmp_683_2 <= 0;
    end else begin
      __tmp_683_1 <= _tmp_683;
      __tmp_683_2 <= __tmp_683_1;
    end
  end

  localparam _stream_conv2d_16_source_35_source_pat_fsm_18_1 = 1;
  localparam _stream_conv2d_16_source_35_source_pat_fsm_18_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_35_source_pat_fsm_18 <= _stream_conv2d_16_source_35_source_pat_fsm_18_init;
    end else begin
      case(_stream_conv2d_16_source_35_source_pat_fsm_18)
        _stream_conv2d_16_source_35_source_pat_fsm_18_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_35_source_mode & 3'b10) begin
            _stream_conv2d_16_source_35_source_pat_fsm_18 <= _stream_conv2d_16_source_35_source_pat_fsm_18_1;
          end 
        end
        _stream_conv2d_16_source_35_source_pat_fsm_18_1: begin
          if((_source_stream_conv2d_16_source_35_pat_count_0 == 0) && (_source_stream_conv2d_16_source_35_pat_count_1 == 0) && (_source_stream_conv2d_16_source_35_pat_count_2 == 0) && (_source_stream_conv2d_16_source_35_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_35_source_pat_fsm_18 <= _stream_conv2d_16_source_35_source_pat_fsm_18_2;
          end 
        end
        _stream_conv2d_16_source_35_source_pat_fsm_18_2: begin
          _stream_conv2d_16_source_35_source_pat_fsm_18 <= _stream_conv2d_16_source_35_source_pat_fsm_18_init;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_697_1 <= 0;
      __tmp_697_2 <= 0;
    end else begin
      __tmp_697_1 <= _tmp_697;
      __tmp_697_2 <= __tmp_697_1;
    end
  end

  localparam _stream_conv2d_16_source_36_source_pat_fsm_19_1 = 1;
  localparam _stream_conv2d_16_source_36_source_pat_fsm_19_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_source_36_source_pat_fsm_19 <= _stream_conv2d_16_source_36_source_pat_fsm_19_init;
    end else begin
      case(_stream_conv2d_16_source_36_source_pat_fsm_19)
        _stream_conv2d_16_source_36_source_pat_fsm_19_init: begin
          if(_stream_conv2d_16_start && _stream_conv2d_16_source_36_source_mode & 3'b10) begin
            _stream_conv2d_16_source_36_source_pat_fsm_19 <= _stream_conv2d_16_source_36_source_pat_fsm_19_1;
          end 
        end
        _stream_conv2d_16_source_36_source_pat_fsm_19_1: begin
          if((_source_stream_conv2d_16_source_36_pat_count_0 == 0) && (_source_stream_conv2d_16_source_36_pat_count_1 == 0) && (_source_stream_conv2d_16_source_36_pat_count_2 == 0) && (_source_stream_conv2d_16_source_36_pat_count_3 == 0)) begin
            _stream_conv2d_16_source_36_source_pat_fsm_19 <= _stream_conv2d_16_source_36_source_pat_fsm_19_2;
          end 
        end
        _stream_conv2d_16_source_36_source_pat_fsm_19_2: begin
          _stream_conv2d_16_source_36_source_pat_fsm_19 <= _stream_conv2d_16_source_36_source_pat_fsm_19_init;
        end
      endcase
    end
  end

  localparam _stream_conv2d_16_sink_37_sink_fsm_20_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_16_sink_37_sink_fsm_20 <= _stream_conv2d_16_sink_37_sink_fsm_20_init;
    end else begin
      case(_stream_conv2d_16_sink_37_sink_fsm_20)
        _stream_conv2d_16_sink_37_sink_fsm_20_init: begin
          if(__stream_conv2d_16_start_46 && _stream_conv2d_16_sink_37_sink_mode & 3'b1) begin
            _stream_conv2d_16_sink_37_sink_fsm_20 <= _stream_conv2d_16_sink_37_sink_fsm_20_1;
          end 
        end
        _stream_conv2d_16_sink_37_sink_fsm_20_1: begin
          if(stream_conv2d_16_sink_38_data && (_stream_conv2d_16_sink_37_sink_count == 1)) begin
            _stream_conv2d_16_sink_37_sink_fsm_20 <= _stream_conv2d_16_sink_37_sink_fsm_20_init;
          end 
          if(_stream_conv2d_16_term_sink) begin
            _stream_conv2d_16_sink_37_sink_fsm_20 <= _stream_conv2d_16_sink_37_sink_fsm_20_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_fsm_1 = 1;
  localparam _maxi_write_fsm_2 = 2;
  localparam _maxi_write_fsm_3 = 3;
  localparam _maxi_write_fsm_4 = 4;
  localparam _maxi_write_fsm_5 = 5;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_fsm <= _maxi_write_fsm_init;
      _d1__maxi_write_fsm <= _maxi_write_fsm_init;
      _maxi_write_cur_global_addr <= 0;
      _maxi_write_rest_size <= 0;
      _maxi_write_cur_size <= 0;
      axim_flag_1021 <= 0;
      __maxi_write_fsm_cond_4_0_1 <= 0;
    end else begin
      _d1__maxi_write_fsm <= _maxi_write_fsm;
      case(_d1__maxi_write_fsm)
        _maxi_write_fsm_4: begin
          if(__maxi_write_fsm_cond_4_0_1) begin
            axim_flag_1021 <= 0;
          end 
        end
      endcase
      case(_maxi_write_fsm)
        _maxi_write_fsm_init: begin
          if(_maxi_write_start) begin
            _maxi_write_cur_global_addr <= (_maxi_write_global_addr + _maxi_global_base_addr >> 2) << 2;
            _maxi_write_rest_size <= _maxi_write_size;
          end 
          if(_maxi_write_start && (_maxi_write_op_sel == 1)) begin
            _maxi_write_fsm <= _maxi_write_fsm_1;
          end 
          if(_maxi_write_start && (_maxi_write_op_sel == 2)) begin
            _maxi_write_fsm <= _maxi_write_fsm_1;
          end 
          if(_maxi_write_start && (_maxi_write_op_sel == 3)) begin
            _maxi_write_fsm <= _maxi_write_fsm_1;
          end 
        end
        _maxi_write_fsm_1: begin
          if((_maxi_write_rest_size <= 256) && ((_maxi_write_cur_global_addr & 4095) + (_maxi_write_rest_size << 2) >= 4096)) begin
            _maxi_write_cur_size <= 4096 - (_maxi_write_cur_global_addr & 4095) >> 2;
            _maxi_write_rest_size <= _maxi_write_rest_size - (4096 - (_maxi_write_cur_global_addr & 4095) >> 2);
          end else if(_maxi_write_rest_size <= 256) begin
            _maxi_write_cur_size <= _maxi_write_rest_size;
            _maxi_write_rest_size <= 0;
          end else if((_maxi_write_cur_global_addr & 4095) + 1024 >= 4096) begin
            _maxi_write_cur_size <= 4096 - (_maxi_write_cur_global_addr & 4095) >> 2;
            _maxi_write_rest_size <= _maxi_write_rest_size - (4096 - (_maxi_write_cur_global_addr & 4095) >> 2);
          end else begin
            _maxi_write_cur_size <= 256;
            _maxi_write_rest_size <= _maxi_write_rest_size - 256;
          end
          _maxi_write_fsm <= _maxi_write_fsm_2;
        end
        _maxi_write_fsm_2: begin
          if(maxi_awready || !maxi_awvalid) begin
            _maxi_write_fsm <= _maxi_write_fsm_3;
          end 
        end
        _maxi_write_fsm_3: begin
          if(_maxi_write_data_done) begin
            _maxi_write_cur_global_addr <= _maxi_write_cur_global_addr + (_maxi_write_cur_size << 2);
          end 
          if(_maxi_write_data_done && (_maxi_write_rest_size > 0)) begin
            _maxi_write_fsm <= _maxi_write_fsm_1;
          end 
          if(_maxi_write_data_done && (_maxi_write_rest_size == 0)) begin
            _maxi_write_fsm <= _maxi_write_fsm_4;
          end 
        end
        _maxi_write_fsm_4: begin
          axim_flag_1021 <= 1;
          __maxi_write_fsm_cond_4_0_1 <= 1;
          _maxi_write_fsm <= _maxi_write_fsm_5;
        end
        _maxi_write_fsm_5: begin
          _maxi_write_fsm <= _maxi_write_fsm_init;
        end
      endcase
    end
  end

  localparam control_max_pool_serial_18_1 = 1;
  localparam control_max_pool_serial_18_2 = 2;
  localparam control_max_pool_serial_18_3 = 3;
  localparam control_max_pool_serial_18_4 = 4;
  localparam control_max_pool_serial_18_5 = 5;
  localparam control_max_pool_serial_18_6 = 6;
  localparam control_max_pool_serial_18_7 = 7;
  localparam control_max_pool_serial_18_8 = 8;
  localparam control_max_pool_serial_18_9 = 9;
  localparam control_max_pool_serial_18_10 = 10;
  localparam control_max_pool_serial_18_11 = 11;
  localparam control_max_pool_serial_18_12 = 12;
  localparam control_max_pool_serial_18_13 = 13;
  localparam control_max_pool_serial_18_14 = 14;
  localparam control_max_pool_serial_18_15 = 15;
  localparam control_max_pool_serial_18_16 = 16;
  localparam control_max_pool_serial_18_17 = 17;
  localparam control_max_pool_serial_18_18 = 18;
  localparam control_max_pool_serial_18_19 = 19;
  localparam control_max_pool_serial_18_20 = 20;
  localparam control_max_pool_serial_18_21 = 21;
  localparam control_max_pool_serial_18_22 = 22;
  localparam control_max_pool_serial_18_23 = 23;
  localparam control_max_pool_serial_18_24 = 24;
  localparam control_max_pool_serial_18_25 = 25;

  always @(posedge CLK) begin
    if(RST) begin
      control_max_pool_serial_18 <= control_max_pool_serial_18_init;
      _d1_control_max_pool_serial_18 <= control_max_pool_serial_18_init;
      _control_max_pool_serial_18_called <= 0;
      max_pool_serial_18_act_base_offset_row <= 0;
      max_pool_serial_18_act_base_offset_bat <= 0;
      max_pool_serial_18_act_page <= 0;
      max_pool_serial_18_act_page_comp_offset <= 0;
      max_pool_serial_18_act_page_dma_offset <= 0;
      max_pool_serial_18_out_base_offset_row <= 0;
      max_pool_serial_18_out_base_offset_bat <= 0;
      max_pool_serial_18_out_page <= 0;
      max_pool_serial_18_out_page_comp_offset <= 0;
      max_pool_serial_18_out_page_dma_offset <= 0;
      max_pool_serial_18_row_count <= 0;
      max_pool_serial_18_bat_count <= 0;
      max_pool_serial_18_prev_row_count <= 0;
      max_pool_serial_18_prev_bat_count <= 0;
      max_pool_serial_18_skip_read_act <= 0;
      max_pool_serial_18_skip_comp <= 0;
      max_pool_serial_18_skip_write_out <= 0;
      max_pool_serial_18_out_count <= 0;
      axim_flag_1022 <= 0;
      _control_max_pool_serial_18_cond_5_0_1 <= 0;
      axim_flag_1023 <= 0;
      _control_max_pool_serial_18_cond_11_1_1 <= 0;
      axim_flag_1071 <= 0;
      _control_max_pool_serial_18_cond_19_2_1 <= 0;
    end else begin
      _d1_control_max_pool_serial_18 <= control_max_pool_serial_18;
      case(_d1_control_max_pool_serial_18)
        control_max_pool_serial_18_5: begin
          if(_control_max_pool_serial_18_cond_5_0_1) begin
            axim_flag_1022 <= 0;
          end 
        end
        control_max_pool_serial_18_11: begin
          if(_control_max_pool_serial_18_cond_11_1_1) begin
            axim_flag_1023 <= 0;
          end 
        end
        control_max_pool_serial_18_19: begin
          if(_control_max_pool_serial_18_cond_19_2_1) begin
            axim_flag_1071 <= 0;
          end 
        end
      endcase
      case(control_max_pool_serial_18)
        control_max_pool_serial_18_init: begin
          if(main_fsm == 18) begin
            _control_max_pool_serial_18_called <= 1;
          end 
          if(main_fsm == 35) begin
            _control_max_pool_serial_18_called <= 1;
          end 
          if(main_fsm == 52) begin
            _control_max_pool_serial_18_called <= 1;
          end 
          if(main_fsm == 18) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_1;
          end 
          if(main_fsm == 35) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_1;
          end 
          if(main_fsm == 52) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_1;
          end 
        end
        control_max_pool_serial_18_1: begin
          control_max_pool_serial_18 <= control_max_pool_serial_18_2;
        end
        control_max_pool_serial_18_2: begin
          max_pool_serial_18_act_base_offset_row <= 0;
          max_pool_serial_18_act_base_offset_bat <= 0;
          max_pool_serial_18_act_page <= 0;
          max_pool_serial_18_act_page_comp_offset <= 0;
          max_pool_serial_18_act_page_dma_offset <= 0;
          max_pool_serial_18_out_base_offset_row <= 0;
          max_pool_serial_18_out_base_offset_bat <= 0;
          max_pool_serial_18_out_page <= 0;
          max_pool_serial_18_out_page_comp_offset <= 0;
          max_pool_serial_18_out_page_dma_offset <= 0;
          max_pool_serial_18_row_count <= 0;
          max_pool_serial_18_bat_count <= 0;
          max_pool_serial_18_prev_row_count <= 0;
          max_pool_serial_18_prev_bat_count <= 0;
          max_pool_serial_18_skip_read_act <= 0;
          max_pool_serial_18_skip_comp <= 0;
          max_pool_serial_18_skip_write_out <= 1;
          max_pool_serial_18_out_count <= 0;
          control_max_pool_serial_18 <= control_max_pool_serial_18_3;
        end
        control_max_pool_serial_18_3: begin
          control_max_pool_serial_18 <= control_max_pool_serial_18_4;
          if(max_pool_serial_18_dma_pad_mask_0) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_9;
          end 
          if(max_pool_serial_18_skip_read_act) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_16;
          end 
        end
        control_max_pool_serial_18_4: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_5;
          end 
        end
        control_max_pool_serial_18_5: begin
          axim_flag_1022 <= 1;
          _control_max_pool_serial_18_cond_5_0_1 <= 1;
          control_max_pool_serial_18 <= control_max_pool_serial_18_6;
        end
        control_max_pool_serial_18_6: begin
          control_max_pool_serial_18 <= control_max_pool_serial_18_7;
        end
        control_max_pool_serial_18_7: begin
          control_max_pool_serial_18 <= control_max_pool_serial_18_8;
        end
        control_max_pool_serial_18_8: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_9;
          end 
        end
        control_max_pool_serial_18_9: begin
          control_max_pool_serial_18 <= control_max_pool_serial_18_10;
          if(max_pool_serial_18_dma_pad_mask_1) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_15;
          end 
        end
        control_max_pool_serial_18_10: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_11;
          end 
        end
        control_max_pool_serial_18_11: begin
          axim_flag_1023 <= 1;
          _control_max_pool_serial_18_cond_11_1_1 <= 1;
          control_max_pool_serial_18 <= control_max_pool_serial_18_12;
        end
        control_max_pool_serial_18_12: begin
          control_max_pool_serial_18 <= control_max_pool_serial_18_13;
        end
        control_max_pool_serial_18_13: begin
          control_max_pool_serial_18 <= control_max_pool_serial_18_14;
        end
        control_max_pool_serial_18_14: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_15;
          end 
        end
        control_max_pool_serial_18_15: begin
          control_max_pool_serial_18 <= control_max_pool_serial_18_16;
        end
        control_max_pool_serial_18_16: begin
          if(max_pool_serial_18_comp_fsm == 0) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_17;
          end 
        end
        control_max_pool_serial_18_17: begin
          if(max_pool_serial_18_comp_count >= max_pool_serial_18_out_count + cparam_max_pool_serial_18_out_write_size) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_18;
          end 
          if(max_pool_serial_18_skip_write_out) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_23;
          end 
        end
        control_max_pool_serial_18_18: begin
          if(_maxi_write_idle) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_19;
          end 
        end
        control_max_pool_serial_18_19: begin
          axim_flag_1071 <= 1;
          _control_max_pool_serial_18_cond_19_2_1 <= 1;
          control_max_pool_serial_18 <= control_max_pool_serial_18_20;
        end
        control_max_pool_serial_18_20: begin
          control_max_pool_serial_18 <= control_max_pool_serial_18_21;
        end
        control_max_pool_serial_18_21: begin
          control_max_pool_serial_18 <= control_max_pool_serial_18_22;
        end
        control_max_pool_serial_18_22: begin
          max_pool_serial_18_out_count <= max_pool_serial_18_out_count + cparam_max_pool_serial_18_out_write_size;
          control_max_pool_serial_18 <= control_max_pool_serial_18_23;
        end
        control_max_pool_serial_18_23: begin
          max_pool_serial_18_act_base_offset_row <= max_pool_serial_18_act_base_offset_row + cparam_max_pool_serial_18_act_row_step;
          if(max_pool_serial_18_row_count >= cparam_max_pool_serial_18_max_row_count) begin
            max_pool_serial_18_act_base_offset_row <= 0;
            max_pool_serial_18_act_base_offset_bat <= max_pool_serial_18_act_base_offset_bat + cparam_max_pool_serial_18_act_bat_step;
          end 
          if((max_pool_serial_18_row_count >= cparam_max_pool_serial_18_max_row_count) && (max_pool_serial_18_bat_count >= cparam_max_pool_serial_18_max_bat_count)) begin
            max_pool_serial_18_act_base_offset_bat <= 0;
          end 
          max_pool_serial_18_row_count <= max_pool_serial_18_row_count + cparam_max_pool_serial_18_stride_row;
          if(max_pool_serial_18_row_count >= cparam_max_pool_serial_18_max_row_count) begin
            max_pool_serial_18_row_count <= 0;
            max_pool_serial_18_bat_count <= max_pool_serial_18_bat_count + 1;
          end 
          if((max_pool_serial_18_row_count >= cparam_max_pool_serial_18_max_row_count) && (max_pool_serial_18_bat_count >= cparam_max_pool_serial_18_max_bat_count)) begin
            max_pool_serial_18_bat_count <= 0;
          end 
          if(!max_pool_serial_18_act_page) begin
            max_pool_serial_18_act_page_comp_offset <= 1024;
            max_pool_serial_18_act_page_dma_offset <= 1024;
            max_pool_serial_18_act_page <= 1;
          end 
          if(max_pool_serial_18_act_page) begin
            max_pool_serial_18_act_page_comp_offset <= 0;
            max_pool_serial_18_act_page_dma_offset <= 0;
            max_pool_serial_18_act_page <= 0;
          end 
          if(!max_pool_serial_18_skip_write_out) begin
            max_pool_serial_18_out_base_offset_row <= max_pool_serial_18_out_base_offset_row + cparam_max_pool_serial_18_out_row_step;
          end 
          if(!max_pool_serial_18_skip_write_out && (max_pool_serial_18_prev_row_count >= cparam_max_pool_serial_18_max_row_count)) begin
            max_pool_serial_18_out_base_offset_row <= 0;
            max_pool_serial_18_out_base_offset_bat <= max_pool_serial_18_out_base_offset_bat + cparam_max_pool_serial_18_out_bat_step;
          end 
          if(!max_pool_serial_18_skip_write_out && (max_pool_serial_18_prev_row_count >= cparam_max_pool_serial_18_max_row_count) && (max_pool_serial_18_prev_bat_count >= cparam_max_pool_serial_18_max_bat_count)) begin
            max_pool_serial_18_out_base_offset_bat <= 0;
          end 
          if(!max_pool_serial_18_out_page) begin
            max_pool_serial_18_out_page_comp_offset <= 1024;
            max_pool_serial_18_out_page_dma_offset <= 0;
            max_pool_serial_18_out_page <= 1;
          end 
          if(max_pool_serial_18_out_page) begin
            max_pool_serial_18_out_page_comp_offset <= 0;
            max_pool_serial_18_out_page_dma_offset <= 1024;
            max_pool_serial_18_out_page <= 0;
          end 
          max_pool_serial_18_prev_row_count <= max_pool_serial_18_row_count;
          max_pool_serial_18_prev_bat_count <= max_pool_serial_18_bat_count;
          if((max_pool_serial_18_row_count >= cparam_max_pool_serial_18_max_row_count) && (max_pool_serial_18_bat_count >= cparam_max_pool_serial_18_max_bat_count)) begin
            max_pool_serial_18_skip_read_act <= 1;
          end 
          if((max_pool_serial_18_row_count >= cparam_max_pool_serial_18_max_row_count) && (max_pool_serial_18_bat_count >= cparam_max_pool_serial_18_max_bat_count)) begin
            max_pool_serial_18_skip_comp <= 1;
          end 
          if(max_pool_serial_18_skip_write_out && (max_pool_serial_18_prev_row_count == 0) && (max_pool_serial_18_prev_bat_count == 0)) begin
            max_pool_serial_18_skip_write_out <= 0;
          end 
          control_max_pool_serial_18 <= control_max_pool_serial_18_3;
          if(!max_pool_serial_18_skip_write_out && (max_pool_serial_18_prev_row_count >= cparam_max_pool_serial_18_max_row_count) && (max_pool_serial_18_prev_bat_count >= cparam_max_pool_serial_18_max_bat_count)) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_24;
          end 
        end
        control_max_pool_serial_18_24: begin
          if(_maxi_write_idle) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_25;
          end 
        end
        control_max_pool_serial_18_25: begin
          if(main_fsm == 21) begin
            _control_max_pool_serial_18_called <= 0;
          end 
          if(main_fsm == 38) begin
            _control_max_pool_serial_18_called <= 0;
          end 
          if(main_fsm == 55) begin
            _control_max_pool_serial_18_called <= 0;
          end 
          if(main_fsm == 21) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_init;
          end 
          if(main_fsm == 38) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_init;
          end 
          if(main_fsm == 55) begin
            control_max_pool_serial_18 <= control_max_pool_serial_18_init;
          end 
        end
      endcase
    end
  end

  localparam max_pool_serial_18_comp_fsm_1 = 1;
  localparam max_pool_serial_18_comp_fsm_2 = 2;
  localparam max_pool_serial_18_comp_fsm_3 = 3;
  localparam max_pool_serial_18_comp_fsm_4 = 4;
  localparam max_pool_serial_18_comp_fsm_5 = 5;
  localparam max_pool_serial_18_comp_fsm_6 = 6;
  localparam max_pool_serial_18_comp_fsm_7 = 7;

  always @(posedge CLK) begin
    if(RST) begin
      max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_init;
      max_pool_serial_18_stream_act_local <= 0;
      max_pool_serial_18_stream_out_local <= 0;
      max_pool_serial_18_col_count <= 0;
      max_pool_serial_18_act_page_comp_offset_buf <= 0;
      max_pool_serial_18_out_page_comp_offset_buf <= 0;
      max_pool_serial_18_row_count_buf <= 0;
      max_pool_serial_18_stream_pad_masks <= 0;
      max_pool_serial_18_comp_count <= 0;
    end else begin
      if(control_max_pool_serial_18 == 2) begin
        max_pool_serial_18_comp_count <= 0;
      end 
      if(_stream_max_pool_serial_18_end_flag) begin
        max_pool_serial_18_comp_count <= max_pool_serial_18_comp_count + cparam_max_pool_serial_18_inc_out_laddr;
      end 
      case(max_pool_serial_18_comp_fsm)
        max_pool_serial_18_comp_fsm_init: begin
          if((control_max_pool_serial_18 == 16) && !max_pool_serial_18_skip_comp) begin
            max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_1;
          end 
        end
        max_pool_serial_18_comp_fsm_1: begin
          max_pool_serial_18_stream_act_local <= cparam_max_pool_serial_18_local_pad_offset;
          max_pool_serial_18_stream_out_local <= 0;
          max_pool_serial_18_col_count <= 0;
          max_pool_serial_18_act_page_comp_offset_buf <= max_pool_serial_18_act_page_comp_offset;
          max_pool_serial_18_out_page_comp_offset_buf <= max_pool_serial_18_out_page_comp_offset;
          max_pool_serial_18_row_count_buf <= max_pool_serial_18_row_count;
          max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_2;
        end
        max_pool_serial_18_comp_fsm_2: begin
          max_pool_serial_18_stream_pad_masks <= { max_pool_serial_18_stream_pad_mask_1_1, max_pool_serial_18_stream_pad_mask_1_0, max_pool_serial_18_stream_pad_mask_0_1, max_pool_serial_18_stream_pad_mask_0_0 };
          max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_3;
        end
        max_pool_serial_18_comp_fsm_3: begin
          if(!_stream_max_pool_serial_18_source_busy) begin
            max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_4;
          end 
        end
        max_pool_serial_18_comp_fsm_4: begin
          max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_5;
          max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_5;
          max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_5;
          max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_5;
        end
        max_pool_serial_18_comp_fsm_5: begin
          max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_6;
        end
        max_pool_serial_18_comp_fsm_6: begin
          max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_7;
        end
        max_pool_serial_18_comp_fsm_7: begin
          max_pool_serial_18_stream_act_local <= max_pool_serial_18_stream_act_local + cparam_max_pool_serial_18_inc_act_laddr;
          if(max_pool_serial_18_col_count >= cparam_max_pool_serial_18_max_col_count) begin
            max_pool_serial_18_stream_act_local <= cparam_max_pool_serial_18_local_pad_offset;
          end 
          max_pool_serial_18_stream_out_local <= max_pool_serial_18_stream_out_local + cparam_max_pool_serial_18_inc_out_laddr;
          if(max_pool_serial_18_col_count >= cparam_max_pool_serial_18_max_col_count) begin
            max_pool_serial_18_stream_out_local <= 0;
          end 
          max_pool_serial_18_col_count <= max_pool_serial_18_col_count + cparam_max_pool_serial_18_stride_col;
          if(max_pool_serial_18_col_count >= cparam_max_pool_serial_18_max_col_count) begin
            max_pool_serial_18_col_count <= 0;
          end 
          max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_2;
          if(max_pool_serial_18_col_count >= cparam_max_pool_serial_18_max_col_count) begin
            max_pool_serial_18_comp_fsm <= max_pool_serial_18_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_serial_18_source_1_source_pat_fsm_0_1 = 1;
  localparam _stream_max_pool_serial_18_source_1_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_18_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_18_source_1_source_pat_fsm_0_init;
    end else begin
      case(_stream_max_pool_serial_18_source_1_source_pat_fsm_0)
        _stream_max_pool_serial_18_source_1_source_pat_fsm_0_init: begin
          if(_stream_max_pool_serial_18_start && _stream_max_pool_serial_18_source_1_source_mode & 3'b10) begin
            _stream_max_pool_serial_18_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_18_source_1_source_pat_fsm_0_1;
          end 
        end
        _stream_max_pool_serial_18_source_1_source_pat_fsm_0_1: begin
          if((_source_stream_max_pool_serial_18_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_18_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_18_source_1_pat_count_2 == 0) && (_source_stream_max_pool_serial_18_source_1_pat_count_3 == 0)) begin
            _stream_max_pool_serial_18_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_18_source_1_source_pat_fsm_0_2;
          end 
        end
        _stream_max_pool_serial_18_source_1_source_pat_fsm_0_2: begin
          _stream_max_pool_serial_18_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_18_source_1_source_pat_fsm_0_init;
        end
      endcase
    end
  end

  localparam _stream_max_pool_serial_18_sink_3_sink_fsm_1_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_18_sink_3_sink_fsm_1 <= _stream_max_pool_serial_18_sink_3_sink_fsm_1_init;
    end else begin
      case(_stream_max_pool_serial_18_sink_3_sink_fsm_1)
        _stream_max_pool_serial_18_sink_3_sink_fsm_1_init: begin
          if(__stream_max_pool_serial_18_start_10 && _stream_max_pool_serial_18_sink_3_sink_mode & 3'b1) begin
            _stream_max_pool_serial_18_sink_3_sink_fsm_1 <= _stream_max_pool_serial_18_sink_3_sink_fsm_1_1;
          end 
        end
        _stream_max_pool_serial_18_sink_3_sink_fsm_1_1: begin
          if(stream_max_pool_serial_18_sink_4_data && (_stream_max_pool_serial_18_sink_3_sink_count == 1)) begin
            _stream_max_pool_serial_18_sink_3_sink_fsm_1 <= _stream_max_pool_serial_18_sink_3_sink_fsm_1_init;
          end 
          if(_stream_max_pool_serial_18_term_sink) begin
            _stream_max_pool_serial_18_sink_3_sink_fsm_1 <= _stream_max_pool_serial_18_sink_3_sink_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam control_matmul_29_1 = 1;
  localparam control_matmul_29_2 = 2;
  localparam control_matmul_29_3 = 3;
  localparam control_matmul_29_4 = 4;
  localparam control_matmul_29_5 = 5;
  localparam control_matmul_29_6 = 6;
  localparam control_matmul_29_7 = 7;
  localparam control_matmul_29_8 = 8;
  localparam control_matmul_29_9 = 9;
  localparam control_matmul_29_10 = 10;
  localparam control_matmul_29_11 = 11;
  localparam control_matmul_29_12 = 12;
  localparam control_matmul_29_13 = 13;
  localparam control_matmul_29_14 = 14;
  localparam control_matmul_29_15 = 15;
  localparam control_matmul_29_16 = 16;
  localparam control_matmul_29_17 = 17;
  localparam control_matmul_29_18 = 18;
  localparam control_matmul_29_19 = 19;
  localparam control_matmul_29_20 = 20;
  localparam control_matmul_29_21 = 21;
  localparam control_matmul_29_22 = 22;
  localparam control_matmul_29_23 = 23;
  localparam control_matmul_29_24 = 24;
  localparam control_matmul_29_25 = 25;
  localparam control_matmul_29_26 = 26;
  localparam control_matmul_29_27 = 27;
  localparam control_matmul_29_28 = 28;
  localparam control_matmul_29_29 = 29;
  localparam control_matmul_29_30 = 30;
  localparam control_matmul_29_31 = 31;
  localparam control_matmul_29_32 = 32;
  localparam control_matmul_29_33 = 33;
  localparam control_matmul_29_34 = 34;
  localparam control_matmul_29_35 = 35;
  localparam control_matmul_29_36 = 36;
  localparam control_matmul_29_37 = 37;
  localparam control_matmul_29_38 = 38;
  localparam control_matmul_29_39 = 39;

  always @(posedge CLK) begin
    if(RST) begin
      control_matmul_29 <= control_matmul_29_init;
      _d1_control_matmul_29 <= control_matmul_29_init;
      _control_matmul_29_called <= 0;
      matmul_29_filter_base_offset <= 0;
      matmul_29_filter_page_comp_offset <= 0;
      matmul_29_filter_page_dma_offset <= 0;
      matmul_29_act_base_offset_row <= 0;
      matmul_29_act_base_offset_bat <= 0;
      matmul_29_dma_flag_0 <= 0;
      matmul_29_act_page_comp_offset_0 <= 0;
      matmul_29_act_page_dma_offset_0 <= 0;
      matmul_29_out_base_offset_val <= 0;
      matmul_29_out_base_offset_col <= 0;
      matmul_29_out_base_offset_row <= 0;
      matmul_29_out_base_offset_bat <= 0;
      matmul_29_out_base_offset_och <= 0;
      matmul_29_out_page <= 0;
      matmul_29_out_page_comp_offset <= 0;
      matmul_29_out_page_dma_offset <= 0;
      matmul_29_out_laddr_offset <= 0;
      matmul_29_sync_out_count <= 0;
      matmul_29_write_count <= 0;
      matmul_29_next_out_write_size <= 0;
      matmul_29_row_count <= 0;
      matmul_29_bat_count <= 0;
      matmul_29_och_count <= 0;
      matmul_29_row_select <= 0;
      matmul_29_prev_row_count <= 0;
      matmul_29_prev_bat_count <= 0;
      matmul_29_prev_och_count <= 0;
      matmul_29_prev_row_select <= 0;
      matmul_29_out_col_count <= 0;
      matmul_29_out_row_count <= 0;
      matmul_29_out_ram_select <= 0;
      matmul_29_skip_read_filter <= 0;
      matmul_29_skip_read_act <= 0;
      matmul_29_skip_comp <= 0;
      matmul_29_skip_write_out <= 1;
      axim_flag_1121 <= 0;
      _control_matmul_29_cond_3_0_1 <= 0;
      axim_flag_1132 <= 0;
      _control_matmul_29_cond_8_1_1 <= 0;
      axim_flag_1133 <= 0;
      _control_matmul_29_cond_14_2_1 <= 0;
      axim_flag_1152 <= 0;
      _control_matmul_29_cond_22_3_1 <= 0;
      axim_flag_1308 <= 0;
      _control_matmul_29_cond_32_4_1 <= 0;
    end else begin
      _d1_control_matmul_29 <= control_matmul_29;
      case(_d1_control_matmul_29)
        control_matmul_29_3: begin
          if(_control_matmul_29_cond_3_0_1) begin
            axim_flag_1121 <= 0;
          end 
        end
        control_matmul_29_8: begin
          if(_control_matmul_29_cond_8_1_1) begin
            axim_flag_1132 <= 0;
          end 
        end
        control_matmul_29_14: begin
          if(_control_matmul_29_cond_14_2_1) begin
            axim_flag_1133 <= 0;
          end 
        end
        control_matmul_29_22: begin
          if(_control_matmul_29_cond_22_3_1) begin
            axim_flag_1152 <= 0;
          end 
        end
        control_matmul_29_32: begin
          if(_control_matmul_29_cond_32_4_1) begin
            axim_flag_1308 <= 0;
          end 
        end
      endcase
      case(control_matmul_29)
        control_matmul_29_init: begin
          if(main_fsm == 64) begin
            _control_matmul_29_called <= 1;
          end 
          if(main_fsm == 74) begin
            _control_matmul_29_called <= 1;
          end 
          if(main_fsm == 84) begin
            _control_matmul_29_called <= 1;
          end 
          if(main_fsm == 64) begin
            control_matmul_29 <= control_matmul_29_1;
          end 
          if(main_fsm == 74) begin
            control_matmul_29 <= control_matmul_29_1;
          end 
          if(main_fsm == 84) begin
            control_matmul_29 <= control_matmul_29_1;
          end 
        end
        control_matmul_29_1: begin
          control_matmul_29 <= control_matmul_29_2;
        end
        control_matmul_29_2: begin
          matmul_29_filter_base_offset <= 0;
          matmul_29_filter_page_comp_offset <= 0;
          matmul_29_filter_page_dma_offset <= 0;
          matmul_29_act_base_offset_row <= 0;
          matmul_29_act_base_offset_bat <= 0;
          matmul_29_dma_flag_0 <= 1;
          matmul_29_act_page_comp_offset_0 <= 0;
          matmul_29_act_page_dma_offset_0 <= 0;
          matmul_29_out_base_offset_val <= 0;
          matmul_29_out_base_offset_col <= 0;
          matmul_29_out_base_offset_row <= 0;
          matmul_29_out_base_offset_bat <= 0;
          matmul_29_out_base_offset_och <= 0;
          matmul_29_out_page <= 0;
          matmul_29_out_page_comp_offset <= 0;
          matmul_29_out_page_dma_offset <= 0;
          matmul_29_out_laddr_offset <= 0;
          matmul_29_sync_out_count <= 0;
          matmul_29_write_count <= 0;
          matmul_29_next_out_write_size <= (cparam_matmul_29_max_och_count == 0)? cparam_matmul_29_out_write_size_res : cparam_matmul_29_out_write_size;
          matmul_29_row_count <= 0;
          matmul_29_bat_count <= 0;
          matmul_29_och_count <= 0;
          matmul_29_row_select <= 0;
          matmul_29_prev_row_count <= 0;
          matmul_29_prev_bat_count <= 0;
          matmul_29_prev_och_count <= 0;
          matmul_29_prev_row_select <= 0;
          matmul_29_out_col_count <= 0;
          matmul_29_out_row_count <= 0;
          matmul_29_out_ram_select <= 0;
          matmul_29_skip_read_filter <= 0;
          matmul_29_skip_read_act <= 0;
          matmul_29_skip_comp <= 0;
          matmul_29_skip_write_out <= 1;
          if(_maxi_read_idle) begin
            control_matmul_29 <= control_matmul_29_3;
          end 
        end
        control_matmul_29_3: begin
          axim_flag_1121 <= 1;
          _control_matmul_29_cond_3_0_1 <= 1;
          control_matmul_29 <= control_matmul_29_4;
        end
        control_matmul_29_4: begin
          control_matmul_29 <= control_matmul_29_5;
        end
        control_matmul_29_5: begin
          control_matmul_29 <= control_matmul_29_6;
        end
        control_matmul_29_6: begin
          if(_maxi_read_idle) begin
            control_matmul_29 <= control_matmul_29_7;
          end 
        end
        control_matmul_29_7: begin
          if(_maxi_read_idle) begin
            control_matmul_29 <= control_matmul_29_8;
          end 
        end
        control_matmul_29_8: begin
          axim_flag_1132 <= 1;
          _control_matmul_29_cond_8_1_1 <= 1;
          control_matmul_29 <= control_matmul_29_9;
        end
        control_matmul_29_9: begin
          control_matmul_29 <= control_matmul_29_10;
        end
        control_matmul_29_10: begin
          control_matmul_29 <= control_matmul_29_11;
        end
        control_matmul_29_11: begin
          if(_maxi_read_idle) begin
            control_matmul_29 <= control_matmul_29_12;
          end 
        end
        control_matmul_29_12: begin
          if(cparam_matmul_29_data_stationary == 0) begin
            control_matmul_29 <= control_matmul_29_13;
          end 
          if(cparam_matmul_29_data_stationary == 1) begin
            control_matmul_29 <= control_matmul_29_20;
          end 
        end
        control_matmul_29_13: begin
          if(_maxi_read_idle) begin
            control_matmul_29 <= control_matmul_29_14;
          end 
          if(matmul_29_skip_read_filter) begin
            control_matmul_29 <= control_matmul_29_19;
          end 
        end
        control_matmul_29_14: begin
          axim_flag_1133 <= 1;
          _control_matmul_29_cond_14_2_1 <= 1;
          control_matmul_29 <= control_matmul_29_15;
        end
        control_matmul_29_15: begin
          control_matmul_29 <= control_matmul_29_16;
        end
        control_matmul_29_16: begin
          control_matmul_29 <= control_matmul_29_17;
        end
        control_matmul_29_17: begin
          if(_maxi_read_idle) begin
            control_matmul_29 <= control_matmul_29_18;
          end 
        end
        control_matmul_29_18: begin
          control_matmul_29 <= control_matmul_29_19;
        end
        control_matmul_29_19: begin
          if(cparam_matmul_29_data_stationary == 0) begin
            control_matmul_29 <= control_matmul_29_20;
          end 
          if(cparam_matmul_29_data_stationary == 1) begin
            control_matmul_29 <= control_matmul_29_28;
          end 
        end
        control_matmul_29_20: begin
          control_matmul_29 <= control_matmul_29_21;
          if(matmul_29_mux_dma_pad_mask_0 || !matmul_29_mux_dma_flag_0) begin
            control_matmul_29 <= control_matmul_29_26;
          end 
          if(matmul_29_skip_read_act) begin
            control_matmul_29 <= control_matmul_29_27;
          end 
        end
        control_matmul_29_21: begin
          if(_maxi_read_idle) begin
            control_matmul_29 <= control_matmul_29_22;
          end 
        end
        control_matmul_29_22: begin
          axim_flag_1152 <= 1;
          _control_matmul_29_cond_22_3_1 <= 1;
          control_matmul_29 <= control_matmul_29_23;
        end
        control_matmul_29_23: begin
          control_matmul_29 <= control_matmul_29_24;
        end
        control_matmul_29_24: begin
          control_matmul_29 <= control_matmul_29_25;
        end
        control_matmul_29_25: begin
          if(_maxi_read_idle) begin
            control_matmul_29 <= control_matmul_29_26;
          end 
        end
        control_matmul_29_26: begin
          control_matmul_29 <= control_matmul_29_27;
        end
        control_matmul_29_27: begin
          if(cparam_matmul_29_data_stationary == 0) begin
            control_matmul_29 <= control_matmul_29_28;
          end 
          if(cparam_matmul_29_data_stationary == 1) begin
            control_matmul_29 <= control_matmul_29_13;
          end 
        end
        control_matmul_29_28: begin
          if(matmul_29_comp_fsm == 0) begin
            control_matmul_29 <= control_matmul_29_29;
          end 
        end
        control_matmul_29_29: begin
          if(matmul_29_sync_comp_count >= matmul_29_sync_out_count + cparam_matmul_29_inc_sync_out) begin
            control_matmul_29 <= control_matmul_29_30;
          end 
          if(matmul_29_skip_write_out) begin
            control_matmul_29 <= control_matmul_29_37;
          end 
          if((cparam_matmul_29_data_stationary == 1) && (matmul_29_prev_och_count < cparam_matmul_29_max_och_count)) begin
            control_matmul_29 <= control_matmul_29_37;
          end 
        end
        control_matmul_29_30: begin
          if(!matmul_29_dma_out_mask_0) begin
            control_matmul_29 <= control_matmul_29_31;
          end 
          if(matmul_29_dma_out_mask_0) begin
            control_matmul_29 <= control_matmul_29_35;
          end 
        end
        control_matmul_29_31: begin
          if(_maxi_write_idle) begin
            control_matmul_29 <= control_matmul_29_32;
          end 
        end
        control_matmul_29_32: begin
          axim_flag_1308 <= 1;
          _control_matmul_29_cond_32_4_1 <= 1;
          control_matmul_29 <= control_matmul_29_33;
        end
        control_matmul_29_33: begin
          control_matmul_29 <= control_matmul_29_34;
        end
        control_matmul_29_34: begin
          control_matmul_29 <= control_matmul_29_35;
        end
        control_matmul_29_35: begin
          control_matmul_29 <= control_matmul_29_36;
        end
        control_matmul_29_36: begin
          matmul_29_write_count <= matmul_29_write_count + 1;
          if(matmul_29_out_ram_select == 0) begin
            matmul_29_out_laddr_offset <= matmul_29_out_laddr_offset + matmul_29_next_out_write_size;
          end 
          if((cparam_matmul_29_data_stationary == 0) && !cparam_matmul_29_keep_filter) begin
            matmul_29_out_base_offset_col <= matmul_29_out_base_offset_col + cparam_matmul_29_out_col_step;
            matmul_29_out_col_count <= matmul_29_out_col_count + 1;
          end 
          matmul_29_out_ram_select <= matmul_29_out_ram_select + 1;
          if(matmul_29_out_ram_select == 0) begin
            matmul_29_out_ram_select <= 0;
          end 
          matmul_29_sync_out_count <= matmul_29_sync_out_count + cparam_matmul_29_inc_sync_out;
          if((cparam_matmul_29_data_stationary == 0) && !cparam_matmul_29_keep_filter && (matmul_29_write_count >= cparam_matmul_29_out_num_col - 1) || (cparam_matmul_29_data_stationary == 0) && cparam_matmul_29_keep_filter || (cparam_matmul_29_data_stationary == 1)) begin
            matmul_29_sync_out_count <= matmul_29_sync_out_count + (cparam_matmul_29_inc_sync_out + cparam_matmul_29_inc_sync_out_res);
          end 
          if((cparam_matmul_29_data_stationary == 0) && !cparam_matmul_29_keep_filter) begin
            control_matmul_29 <= control_matmul_29_29;
          end 
          if((cparam_matmul_29_data_stationary == 0) && !cparam_matmul_29_keep_filter && (matmul_29_write_count >= cparam_matmul_29_out_num_col - 1) || (cparam_matmul_29_data_stationary == 0) && cparam_matmul_29_keep_filter || (cparam_matmul_29_data_stationary == 1)) begin
            control_matmul_29 <= control_matmul_29_37;
          end 
        end
        control_matmul_29_37: begin
          if(matmul_29_update_filter) begin
            matmul_29_filter_base_offset <= matmul_29_filter_base_offset + cparam_matmul_29_filter_base_step;
          end 
          if((cparam_matmul_29_data_stationary == 1) && (matmul_29_och_count >= cparam_matmul_29_max_och_count)) begin
            matmul_29_filter_base_offset <= 0;
          end 
          if(matmul_29_update_filter) begin
            matmul_29_och_count <= matmul_29_och_count + cparam_matmul_29_och_count_step;
          end 
          if((cparam_matmul_29_data_stationary == 1) && (matmul_29_och_count >= cparam_matmul_29_max_och_count)) begin
            matmul_29_och_count <= 0;
          end 
          if(matmul_29_update_filter) begin
            matmul_29_filter_page_comp_offset <= matmul_29_filter_page_comp_offset + cparam_matmul_29_filter_read_step;
            matmul_29_filter_page_dma_offset <= matmul_29_filter_page_dma_offset + cparam_matmul_29_filter_read_step;
          end 
          if(matmul_29_update_filter && (matmul_29_filter_page_comp_offset + cparam_matmul_29_filter_read_step + cparam_matmul_29_filter_read_step > 8192)) begin
            matmul_29_filter_page_comp_offset <= 0;
            matmul_29_filter_page_dma_offset <= 0;
          end 
          if(matmul_29_update_act) begin
            matmul_29_act_base_offset_row <= matmul_29_act_base_offset_row + cparam_matmul_29_act_row_step;
          end 
          if(matmul_29_update_act && (matmul_29_row_count >= cparam_matmul_29_max_row_count)) begin
            matmul_29_act_base_offset_row <= 0;
            matmul_29_act_base_offset_bat <= matmul_29_act_base_offset_bat + cparam_matmul_29_act_bat_step;
          end 
          if(matmul_29_update_act && (matmul_29_row_count >= cparam_matmul_29_max_row_count) && (matmul_29_bat_count >= cparam_matmul_29_max_bat_count)) begin
            matmul_29_act_base_offset_bat <= 0;
          end 
          if(!matmul_29_update_act) begin
            matmul_29_dma_flag_0 <= 0;
          end 
          if(matmul_29_update_act) begin
            matmul_29_dma_flag_0 <= cparam_matmul_29_dma_flag_conds_0;
          end 
          if(matmul_29_update_act && (matmul_29_row_count >= cparam_matmul_29_max_row_count)) begin
            matmul_29_dma_flag_0 <= 1;
          end 
          if(matmul_29_update_act) begin
            matmul_29_row_count <= matmul_29_row_count + cparam_matmul_29_stride_row_par_row;
          end 
          if(matmul_29_update_act && (matmul_29_row_count >= cparam_matmul_29_max_row_count)) begin
            matmul_29_row_count <= 0;
            matmul_29_bat_count <= matmul_29_bat_count + 1;
          end 
          if(matmul_29_update_act && (matmul_29_row_count >= cparam_matmul_29_max_row_count) && (matmul_29_bat_count >= cparam_matmul_29_max_bat_count)) begin
            matmul_29_bat_count <= 0;
          end 
          if(matmul_29_update_act && (cparam_matmul_29_stride_row_par_row < 1)) begin
            matmul_29_row_select <= matmul_29_row_select + cparam_matmul_29_stride_row_par_row;
            matmul_29_prev_row_select <= matmul_29_row_select;
          end 
          if(matmul_29_update_act && (cparam_matmul_29_stride_row_par_row < 1) && (matmul_29_row_select + cparam_matmul_29_stride_row_par_row >= 1)) begin
            matmul_29_row_select <= matmul_29_row_select - (1 - cparam_matmul_29_stride_row_par_row);
            matmul_29_prev_row_select <= matmul_29_row_select;
          end 
          if(matmul_29_update_act && !(cparam_matmul_29_stride_row_par_row < 1)) begin
            matmul_29_row_select <= 0;
            matmul_29_prev_row_select <= 0;
          end 
          if(matmul_29_update_act && (matmul_29_row_count >= cparam_matmul_29_max_row_count)) begin
            matmul_29_row_select <= 0;
            matmul_29_prev_row_select <= 0;
          end 
          if(matmul_29_update_act && matmul_29_mux_next_dma_flag_0) begin
            matmul_29_act_page_comp_offset_0 <= matmul_29_act_page_comp_offset_0 + cparam_matmul_29_act_read_step;
            matmul_29_act_page_dma_offset_0 <= matmul_29_act_page_dma_offset_0 + cparam_matmul_29_act_read_step;
          end 
          if(matmul_29_update_act && matmul_29_mux_next_dma_flag_0 && (matmul_29_act_page_comp_offset_0 + cparam_matmul_29_act_read_step + cparam_matmul_29_act_read_step > 2048)) begin
            matmul_29_act_page_comp_offset_0 <= 0;
            matmul_29_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_matmul_29_data_stationary == 0) && (matmul_29_row_count >= cparam_matmul_29_max_row_count) && (matmul_29_bat_count >= cparam_matmul_29_max_bat_count) && cparam_matmul_29_keep_input) begin
            matmul_29_act_page_comp_offset_0 <= 0;
            matmul_29_act_page_dma_offset_0 <= 0;
          end 
          matmul_29_next_out_write_size <= (matmul_29_och_count >= cparam_matmul_29_max_och_count)? cparam_matmul_29_out_write_size_res : cparam_matmul_29_out_write_size;
          if(!matmul_29_skip_write_out) begin
            matmul_29_write_count <= 0;
            matmul_29_out_laddr_offset <= 0;
            matmul_29_out_ram_select <= 0;
          end 
          if((cparam_matmul_29_data_stationary == 0) && !matmul_29_skip_write_out) begin
            matmul_29_out_base_offset_col <= 0;
            matmul_29_out_base_offset_row <= matmul_29_out_base_offset_row + cparam_matmul_29_out_row_step;
            matmul_29_out_col_count <= 0;
            matmul_29_out_row_count <= matmul_29_out_row_count + 1;
          end 
          if((cparam_matmul_29_data_stationary == 0) && !matmul_29_skip_write_out && (matmul_29_prev_row_count >= cparam_matmul_29_max_row_count)) begin
            matmul_29_out_base_offset_row <= 0;
            matmul_29_out_base_offset_bat <= matmul_29_out_base_offset_bat + cparam_matmul_29_out_bat_step;
            matmul_29_out_row_count <= 0;
          end 
          if((cparam_matmul_29_data_stationary == 0) && !matmul_29_skip_write_out && (matmul_29_prev_row_count >= cparam_matmul_29_max_row_count) && (matmul_29_prev_bat_count >= cparam_matmul_29_max_bat_count)) begin
            matmul_29_out_base_offset_bat <= 0;
            matmul_29_out_base_offset_och <= matmul_29_out_base_offset_och + cparam_matmul_29_out_och_step;
          end 
          if((cparam_matmul_29_data_stationary == 1) && (matmul_29_prev_och_count >= cparam_matmul_29_max_och_count) && !matmul_29_skip_write_out) begin
            matmul_29_out_base_offset_row <= matmul_29_out_base_offset_row + cparam_matmul_29_out_row_step;
          end 
          if((cparam_matmul_29_data_stationary == 0) && !matmul_29_out_page) begin
            matmul_29_out_page_comp_offset <= 1024;
            matmul_29_out_page_dma_offset <= 0;
            matmul_29_out_page <= 1;
          end 
          if((cparam_matmul_29_data_stationary == 0) && matmul_29_out_page) begin
            matmul_29_out_page_comp_offset <= 0;
            matmul_29_out_page_dma_offset <= 1024;
            matmul_29_out_page <= 0;
          end 
          if((cparam_matmul_29_data_stationary == 1) && (matmul_29_och_count >= cparam_matmul_29_max_och_count) && !matmul_29_out_page) begin
            matmul_29_out_page_comp_offset <= 1024;
            matmul_29_out_page_dma_offset <= 0;
            matmul_29_out_page <= 1;
          end 
          if((cparam_matmul_29_data_stationary == 1) && (matmul_29_och_count >= cparam_matmul_29_max_och_count) && matmul_29_out_page) begin
            matmul_29_out_page_comp_offset <= 0;
            matmul_29_out_page_dma_offset <= 1024;
            matmul_29_out_page <= 0;
          end 
          matmul_29_prev_row_count <= matmul_29_row_count;
          matmul_29_prev_bat_count <= matmul_29_bat_count;
          matmul_29_prev_och_count <= matmul_29_och_count;
          if((matmul_29_row_count >= cparam_matmul_29_max_row_count) && (matmul_29_bat_count >= cparam_matmul_29_max_bat_count) && (matmul_29_och_count >= cparam_matmul_29_max_och_count)) begin
            matmul_29_skip_read_filter <= 1;
          end 
          if((cparam_matmul_29_data_stationary == 1) && cparam_matmul_29_keep_filter) begin
            matmul_29_skip_read_filter <= 1;
          end 
          if((matmul_29_row_count >= cparam_matmul_29_max_row_count) && (matmul_29_bat_count >= cparam_matmul_29_max_bat_count) && (matmul_29_och_count >= cparam_matmul_29_max_och_count)) begin
            matmul_29_skip_read_act <= 1;
          end 
          if((cparam_matmul_29_data_stationary == 0) && (matmul_29_row_count >= cparam_matmul_29_max_row_count) && (matmul_29_bat_count >= cparam_matmul_29_max_bat_count) && cparam_matmul_29_keep_input) begin
            matmul_29_skip_read_act <= 1;
          end 
          if((matmul_29_row_count >= cparam_matmul_29_max_row_count) && (matmul_29_bat_count >= cparam_matmul_29_max_bat_count) && (matmul_29_och_count >= cparam_matmul_29_max_och_count)) begin
            matmul_29_skip_comp <= 1;
          end 
          if(matmul_29_skip_write_out && (matmul_29_prev_row_count == 0) && (matmul_29_prev_bat_count == 0) && (matmul_29_prev_och_count == 0)) begin
            matmul_29_skip_write_out <= 0;
          end 
          if(cparam_matmul_29_data_stationary == 0) begin
            control_matmul_29 <= control_matmul_29_20;
          end 
          if((cparam_matmul_29_data_stationary == 0) && (matmul_29_row_count >= cparam_matmul_29_max_row_count) && (matmul_29_bat_count >= cparam_matmul_29_max_bat_count)) begin
            control_matmul_29 <= control_matmul_29_13;
          end 
          if(cparam_matmul_29_data_stationary == 1) begin
            control_matmul_29 <= control_matmul_29_13;
          end 
          if((cparam_matmul_29_data_stationary == 1) && (matmul_29_och_count >= cparam_matmul_29_max_och_count)) begin
            control_matmul_29 <= control_matmul_29_20;
          end 
          if(!matmul_29_skip_write_out && (matmul_29_prev_och_count >= cparam_matmul_29_max_och_count) && (matmul_29_prev_row_count >= cparam_matmul_29_max_row_count) && (matmul_29_prev_bat_count >= cparam_matmul_29_max_bat_count)) begin
            control_matmul_29 <= control_matmul_29_38;
          end 
        end
        control_matmul_29_38: begin
          if(_maxi_write_idle) begin
            control_matmul_29 <= control_matmul_29_39;
          end 
        end
        control_matmul_29_39: begin
          if(main_fsm == 67) begin
            _control_matmul_29_called <= 0;
          end 
          if(main_fsm == 77) begin
            _control_matmul_29_called <= 0;
          end 
          if(main_fsm == 87) begin
            _control_matmul_29_called <= 0;
          end 
          if(main_fsm == 67) begin
            control_matmul_29 <= control_matmul_29_init;
          end 
          if(main_fsm == 77) begin
            control_matmul_29 <= control_matmul_29_init;
          end 
          if(main_fsm == 87) begin
            control_matmul_29 <= control_matmul_29_init;
          end 
        end
      endcase
    end
  end

  localparam matmul_29_comp_fsm_1 = 1;
  localparam matmul_29_comp_fsm_2 = 2;
  localparam matmul_29_comp_fsm_3 = 3;
  localparam matmul_29_comp_fsm_4 = 4;
  localparam matmul_29_comp_fsm_5 = 5;
  localparam matmul_29_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      matmul_29_comp_fsm <= matmul_29_comp_fsm_init;
      matmul_29_stream_act_local_0 <= 0;
      matmul_29_stream_out_local_col <= 0;
      matmul_29_stream_out_local_val <= 0;
      matmul_29_col_count <= 0;
      matmul_29_col_select <= 0;
      matmul_29_filter_page_comp_offset_buf <= 0;
      matmul_29_act_page_comp_offset_buf_0 <= 0;
      matmul_29_out_page_comp_offset_buf <= 0;
      matmul_29_row_count_buf <= 0;
      matmul_29_row_select_buf <= 0;
      matmul_29_och_count_buf <= 0;
      matmul_29_next_stream_num_ops <= 0;
      matmul_29_stream_pad_masks <= 0;
      matmul_29_sync_comp_count <= 0;
    end else begin
      if(_stream_matmul_29_end_flag) begin
        matmul_29_sync_comp_count <= matmul_29_sync_comp_count + 1;
      end 
      if(control_matmul_29 == 12) begin
        matmul_29_sync_comp_count <= 0;
      end 
      case(matmul_29_comp_fsm)
        matmul_29_comp_fsm_init: begin
          if((control_matmul_29 == 28) && !matmul_29_skip_comp) begin
            matmul_29_comp_fsm <= matmul_29_comp_fsm_1;
          end 
        end
        matmul_29_comp_fsm_1: begin
          matmul_29_stream_act_local_0 <= 0;
          if(cparam_matmul_29_stream_act_local_small_flags_0) begin
            matmul_29_stream_act_local_0 <= cparam_matmul_29_stream_act_local_small_offset;
          end 
          if(cparam_matmul_29_stream_act_local_large_flags_0) begin
            matmul_29_stream_act_local_0 <= cparam_matmul_29_stream_act_local_large_offset;
          end 
          matmul_29_stream_out_local_col <= 0;
          if((cparam_matmul_29_data_stationary == 1) && (matmul_29_och_count == 0)) begin
            matmul_29_stream_out_local_val <= 0;
          end 
          matmul_29_col_count <= 0;
          matmul_29_col_select <= cparam_matmul_29_col_select_initval;
          matmul_29_filter_page_comp_offset_buf <= matmul_29_filter_page_comp_offset;
          matmul_29_act_page_comp_offset_buf_0 <= matmul_29_act_page_comp_offset_0;
          matmul_29_out_page_comp_offset_buf <= matmul_29_out_page_comp_offset;
          matmul_29_row_count_buf <= matmul_29_row_count;
          matmul_29_row_select_buf <= matmul_29_row_select;
          matmul_29_och_count_buf <= matmul_29_och_count;
          matmul_29_next_stream_num_ops <= (matmul_29_och_count >= cparam_matmul_29_max_och_count)? cparam_matmul_29_stream_num_ops_res : cparam_matmul_29_stream_num_ops;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_2;
        end
        matmul_29_comp_fsm_2: begin
          matmul_29_stream_pad_masks <= { matmul_29_stream_pad_mask_0_0 };
          matmul_29_comp_fsm <= matmul_29_comp_fsm_3;
        end
        matmul_29_comp_fsm_3: begin
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
          matmul_29_comp_fsm <= matmul_29_comp_fsm_4;
        end
        matmul_29_comp_fsm_4: begin
          if(!_stream_matmul_29_source_busy) begin
            matmul_29_comp_fsm <= matmul_29_comp_fsm_5;
          end 
        end
        matmul_29_comp_fsm_5: begin
          matmul_29_comp_fsm <= matmul_29_comp_fsm_6;
        end
        matmul_29_comp_fsm_6: begin
          if(!((matmul_29_col_select == 0)? cparam_matmul_29_inc_act_laddr_conds_0 : 0)) begin
            matmul_29_stream_act_local_0 <= matmul_29_stream_act_local_0 + cparam_matmul_29_inc_act_laddr_small;
          end 
          if((matmul_29_col_select == 0)? cparam_matmul_29_inc_act_laddr_conds_0 : 0) begin
            matmul_29_stream_act_local_0 <= matmul_29_stream_act_local_0 + cparam_matmul_29_inc_act_laddr_large;
          end 
          if(matmul_29_col_count >= cparam_matmul_29_max_col_count) begin
            matmul_29_stream_act_local_0 <= 0;
          end 
          if((matmul_29_col_count >= cparam_matmul_29_max_col_count) && cparam_matmul_29_stream_act_local_small_flags_0) begin
            matmul_29_stream_act_local_0 <= cparam_matmul_29_stream_act_local_small_offset;
          end 
          if((matmul_29_col_count >= cparam_matmul_29_max_col_count) && cparam_matmul_29_stream_act_local_large_flags_0) begin
            matmul_29_stream_act_local_0 <= cparam_matmul_29_stream_act_local_large_offset;
          end 
          if(cparam_matmul_29_data_stationary == 0) begin
            matmul_29_stream_out_local_col <= matmul_29_stream_out_local_col + matmul_29_next_stream_num_ops;
          end 
          if((cparam_matmul_29_data_stationary == 0) && (matmul_29_col_count >= cparam_matmul_29_max_col_count)) begin
            matmul_29_stream_out_local_col <= 0;
          end 
          if(cparam_matmul_29_data_stationary == 1) begin
            matmul_29_stream_out_local_col <= matmul_29_stream_out_local_col + cparam_matmul_29_inc_out_laddr_col;
          end 
          if((cparam_matmul_29_data_stationary == 1) && (matmul_29_col_count >= cparam_matmul_29_max_col_count)) begin
            matmul_29_stream_out_local_val <= matmul_29_stream_out_local_val + matmul_29_next_stream_num_ops;
            matmul_29_stream_out_local_col <= 0;
          end 
          matmul_29_col_count <= matmul_29_col_count + cparam_matmul_29_stride_col_par_col;
          if(matmul_29_col_count >= cparam_matmul_29_max_col_count) begin
            matmul_29_col_count <= 0;
          end 
          matmul_29_col_select <= matmul_29_col_select + cparam_matmul_29_stride_col_mod_filter_num;
          if(matmul_29_col_select + cparam_matmul_29_stride_col_mod_filter_num >= 1) begin
            matmul_29_col_select <= matmul_29_col_select - cparam_matmul_29_filter_num_col_minus_stride_col_mod;
          end 
          if(matmul_29_col_count >= cparam_matmul_29_max_col_count) begin
            matmul_29_col_select <= cparam_matmul_29_col_select_initval;
          end 
          matmul_29_comp_fsm <= matmul_29_comp_fsm_2;
          if(matmul_29_col_count >= cparam_matmul_29_max_col_count) begin
            matmul_29_comp_fsm <= matmul_29_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_29_source_6_source_pat_fsm_0_1 = 1;
  localparam _stream_matmul_29_source_6_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_29_source_6_source_pat_fsm_0 <= _stream_matmul_29_source_6_source_pat_fsm_0_init;
    end else begin
      case(_stream_matmul_29_source_6_source_pat_fsm_0)
        _stream_matmul_29_source_6_source_pat_fsm_0_init: begin
          if(_stream_matmul_29_start && _stream_matmul_29_source_6_source_mode & 3'b10) begin
            _stream_matmul_29_source_6_source_pat_fsm_0 <= _stream_matmul_29_source_6_source_pat_fsm_0_1;
          end 
        end
        _stream_matmul_29_source_6_source_pat_fsm_0_1: begin
          if((_source_stream_matmul_29_source_6_pat_count_0 == 0) && (_source_stream_matmul_29_source_6_pat_count_1 == 0) && (_source_stream_matmul_29_source_6_pat_count_2 == 0) && (_source_stream_matmul_29_source_6_pat_count_3 == 0)) begin
            _stream_matmul_29_source_6_source_pat_fsm_0 <= _stream_matmul_29_source_6_source_pat_fsm_0_2;
          end 
        end
        _stream_matmul_29_source_6_source_pat_fsm_0_2: begin
          _stream_matmul_29_source_6_source_pat_fsm_0 <= _stream_matmul_29_source_6_source_pat_fsm_0_init;
        end
      endcase
    end
  end

  localparam _stream_matmul_29_source_8_source_pat_fsm_1_1 = 1;
  localparam _stream_matmul_29_source_8_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_29_source_8_source_pat_fsm_1 <= _stream_matmul_29_source_8_source_pat_fsm_1_init;
    end else begin
      case(_stream_matmul_29_source_8_source_pat_fsm_1)
        _stream_matmul_29_source_8_source_pat_fsm_1_init: begin
          if(_stream_matmul_29_start && _stream_matmul_29_source_8_source_mode & 3'b10) begin
            _stream_matmul_29_source_8_source_pat_fsm_1 <= _stream_matmul_29_source_8_source_pat_fsm_1_1;
          end 
        end
        _stream_matmul_29_source_8_source_pat_fsm_1_1: begin
          if((_source_stream_matmul_29_source_8_pat_count_0 == 0) && (_source_stream_matmul_29_source_8_pat_count_1 == 0) && (_source_stream_matmul_29_source_8_pat_count_2 == 0) && (_source_stream_matmul_29_source_8_pat_count_3 == 0)) begin
            _stream_matmul_29_source_8_source_pat_fsm_1 <= _stream_matmul_29_source_8_source_pat_fsm_1_2;
          end 
        end
        _stream_matmul_29_source_8_source_pat_fsm_1_2: begin
          _stream_matmul_29_source_8_source_pat_fsm_1 <= _stream_matmul_29_source_8_source_pat_fsm_1_init;
        end
      endcase
    end
  end

  localparam _stream_matmul_29_source_19_source_pat_fsm_2_1 = 1;
  localparam _stream_matmul_29_source_19_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_29_source_19_source_pat_fsm_2 <= _stream_matmul_29_source_19_source_pat_fsm_2_init;
    end else begin
      case(_stream_matmul_29_source_19_source_pat_fsm_2)
        _stream_matmul_29_source_19_source_pat_fsm_2_init: begin
          if(_stream_matmul_29_start && _stream_matmul_29_source_19_source_mode & 3'b10) begin
            _stream_matmul_29_source_19_source_pat_fsm_2 <= _stream_matmul_29_source_19_source_pat_fsm_2_1;
          end 
        end
        _stream_matmul_29_source_19_source_pat_fsm_2_1: begin
          if((_source_stream_matmul_29_source_19_pat_count_0 == 0) && (_source_stream_matmul_29_source_19_pat_count_1 == 0) && (_source_stream_matmul_29_source_19_pat_count_2 == 0) && (_source_stream_matmul_29_source_19_pat_count_3 == 0)) begin
            _stream_matmul_29_source_19_source_pat_fsm_2 <= _stream_matmul_29_source_19_source_pat_fsm_2_2;
          end 
        end
        _stream_matmul_29_source_19_source_pat_fsm_2_2: begin
          _stream_matmul_29_source_19_source_pat_fsm_2 <= _stream_matmul_29_source_19_source_pat_fsm_2_init;
        end
      endcase
    end
  end

  localparam _stream_matmul_29_source_20_source_pat_fsm_3_1 = 1;
  localparam _stream_matmul_29_source_20_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_29_source_20_source_pat_fsm_3 <= _stream_matmul_29_source_20_source_pat_fsm_3_init;
    end else begin
      case(_stream_matmul_29_source_20_source_pat_fsm_3)
        _stream_matmul_29_source_20_source_pat_fsm_3_init: begin
          if(_stream_matmul_29_start && _stream_matmul_29_source_20_source_mode & 3'b10) begin
            _stream_matmul_29_source_20_source_pat_fsm_3 <= _stream_matmul_29_source_20_source_pat_fsm_3_1;
          end 
        end
        _stream_matmul_29_source_20_source_pat_fsm_3_1: begin
          if((_source_stream_matmul_29_source_20_pat_count_0 == 0) && (_source_stream_matmul_29_source_20_pat_count_1 == 0) && (_source_stream_matmul_29_source_20_pat_count_2 == 0) && (_source_stream_matmul_29_source_20_pat_count_3 == 0)) begin
            _stream_matmul_29_source_20_source_pat_fsm_3 <= _stream_matmul_29_source_20_source_pat_fsm_3_2;
          end 
        end
        _stream_matmul_29_source_20_source_pat_fsm_3_2: begin
          _stream_matmul_29_source_20_source_pat_fsm_3 <= _stream_matmul_29_source_20_source_pat_fsm_3_init;
        end
      endcase
    end
  end

  localparam _stream_matmul_29_sink_21_sink_fsm_4_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_29_sink_21_sink_fsm_4 <= _stream_matmul_29_sink_21_sink_fsm_4_init;
    end else begin
      case(_stream_matmul_29_sink_21_sink_fsm_4)
        _stream_matmul_29_sink_21_sink_fsm_4_init: begin
          if(__stream_matmul_29_start_42 && _stream_matmul_29_sink_21_sink_mode & 3'b1) begin
            _stream_matmul_29_sink_21_sink_fsm_4 <= _stream_matmul_29_sink_21_sink_fsm_4_1;
          end 
        end
        _stream_matmul_29_sink_21_sink_fsm_4_1: begin
          if(stream_matmul_29_sink_22_data && (_stream_matmul_29_sink_21_sink_count == 1)) begin
            _stream_matmul_29_sink_21_sink_fsm_4 <= _stream_matmul_29_sink_21_sink_fsm_4_init;
          end 
          if(_stream_matmul_29_term_sink) begin
            _stream_matmul_29_sink_21_sink_fsm_4 <= _stream_matmul_29_sink_21_sink_fsm_4_init;
          end 
        end
      endcase
    end
  end


endmodule



module ram_w4_l8192_id0_0
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id0_0_0_addr,
  output [4-1:0] ram_w4_l8192_id0_0_0_rdata,
  input [4-1:0] ram_w4_l8192_id0_0_0_wdata,
  input ram_w4_l8192_id0_0_0_wenable,
  input [10-1:0] ram_w4_l8192_id0_0_1_addr,
  output [4-1:0] ram_w4_l8192_id0_0_1_rdata,
  input [4-1:0] ram_w4_l8192_id0_0_1_wdata,
  input ram_w4_l8192_id0_0_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id0_0_0_daddr;
  reg [10-1:0] ram_w4_l8192_id0_0_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_0_0_wenable) begin
      mem[ram_w4_l8192_id0_0_0_addr] <= ram_w4_l8192_id0_0_0_wdata;
    end 
    ram_w4_l8192_id0_0_0_daddr <= ram_w4_l8192_id0_0_0_addr;
  end

  assign ram_w4_l8192_id0_0_0_rdata = mem[ram_w4_l8192_id0_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_0_1_wenable) begin
      mem[ram_w4_l8192_id0_0_1_addr] <= ram_w4_l8192_id0_0_1_wdata;
    end 
    ram_w4_l8192_id0_0_1_daddr <= ram_w4_l8192_id0_0_1_addr;
  end

  assign ram_w4_l8192_id0_0_1_rdata = mem[ram_w4_l8192_id0_0_1_daddr];

endmodule



module ram_w4_l8192_id0_1
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id0_1_0_addr,
  output [4-1:0] ram_w4_l8192_id0_1_0_rdata,
  input [4-1:0] ram_w4_l8192_id0_1_0_wdata,
  input ram_w4_l8192_id0_1_0_wenable,
  input [10-1:0] ram_w4_l8192_id0_1_1_addr,
  output [4-1:0] ram_w4_l8192_id0_1_1_rdata,
  input [4-1:0] ram_w4_l8192_id0_1_1_wdata,
  input ram_w4_l8192_id0_1_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id0_1_0_daddr;
  reg [10-1:0] ram_w4_l8192_id0_1_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_1_0_wenable) begin
      mem[ram_w4_l8192_id0_1_0_addr] <= ram_w4_l8192_id0_1_0_wdata;
    end 
    ram_w4_l8192_id0_1_0_daddr <= ram_w4_l8192_id0_1_0_addr;
  end

  assign ram_w4_l8192_id0_1_0_rdata = mem[ram_w4_l8192_id0_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_1_1_wenable) begin
      mem[ram_w4_l8192_id0_1_1_addr] <= ram_w4_l8192_id0_1_1_wdata;
    end 
    ram_w4_l8192_id0_1_1_daddr <= ram_w4_l8192_id0_1_1_addr;
  end

  assign ram_w4_l8192_id0_1_1_rdata = mem[ram_w4_l8192_id0_1_1_daddr];

endmodule



module ram_w4_l8192_id0_2
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id0_2_0_addr,
  output [4-1:0] ram_w4_l8192_id0_2_0_rdata,
  input [4-1:0] ram_w4_l8192_id0_2_0_wdata,
  input ram_w4_l8192_id0_2_0_wenable,
  input [10-1:0] ram_w4_l8192_id0_2_1_addr,
  output [4-1:0] ram_w4_l8192_id0_2_1_rdata,
  input [4-1:0] ram_w4_l8192_id0_2_1_wdata,
  input ram_w4_l8192_id0_2_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id0_2_0_daddr;
  reg [10-1:0] ram_w4_l8192_id0_2_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_2_0_wenable) begin
      mem[ram_w4_l8192_id0_2_0_addr] <= ram_w4_l8192_id0_2_0_wdata;
    end 
    ram_w4_l8192_id0_2_0_daddr <= ram_w4_l8192_id0_2_0_addr;
  end

  assign ram_w4_l8192_id0_2_0_rdata = mem[ram_w4_l8192_id0_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_2_1_wenable) begin
      mem[ram_w4_l8192_id0_2_1_addr] <= ram_w4_l8192_id0_2_1_wdata;
    end 
    ram_w4_l8192_id0_2_1_daddr <= ram_w4_l8192_id0_2_1_addr;
  end

  assign ram_w4_l8192_id0_2_1_rdata = mem[ram_w4_l8192_id0_2_1_daddr];

endmodule



module ram_w4_l8192_id0_3
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id0_3_0_addr,
  output [4-1:0] ram_w4_l8192_id0_3_0_rdata,
  input [4-1:0] ram_w4_l8192_id0_3_0_wdata,
  input ram_w4_l8192_id0_3_0_wenable,
  input [10-1:0] ram_w4_l8192_id0_3_1_addr,
  output [4-1:0] ram_w4_l8192_id0_3_1_rdata,
  input [4-1:0] ram_w4_l8192_id0_3_1_wdata,
  input ram_w4_l8192_id0_3_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id0_3_0_daddr;
  reg [10-1:0] ram_w4_l8192_id0_3_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_3_0_wenable) begin
      mem[ram_w4_l8192_id0_3_0_addr] <= ram_w4_l8192_id0_3_0_wdata;
    end 
    ram_w4_l8192_id0_3_0_daddr <= ram_w4_l8192_id0_3_0_addr;
  end

  assign ram_w4_l8192_id0_3_0_rdata = mem[ram_w4_l8192_id0_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_3_1_wenable) begin
      mem[ram_w4_l8192_id0_3_1_addr] <= ram_w4_l8192_id0_3_1_wdata;
    end 
    ram_w4_l8192_id0_3_1_daddr <= ram_w4_l8192_id0_3_1_addr;
  end

  assign ram_w4_l8192_id0_3_1_rdata = mem[ram_w4_l8192_id0_3_1_daddr];

endmodule



module ram_w4_l8192_id0_4
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id0_4_0_addr,
  output [4-1:0] ram_w4_l8192_id0_4_0_rdata,
  input [4-1:0] ram_w4_l8192_id0_4_0_wdata,
  input ram_w4_l8192_id0_4_0_wenable,
  input [10-1:0] ram_w4_l8192_id0_4_1_addr,
  output [4-1:0] ram_w4_l8192_id0_4_1_rdata,
  input [4-1:0] ram_w4_l8192_id0_4_1_wdata,
  input ram_w4_l8192_id0_4_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id0_4_0_daddr;
  reg [10-1:0] ram_w4_l8192_id0_4_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_4_0_wenable) begin
      mem[ram_w4_l8192_id0_4_0_addr] <= ram_w4_l8192_id0_4_0_wdata;
    end 
    ram_w4_l8192_id0_4_0_daddr <= ram_w4_l8192_id0_4_0_addr;
  end

  assign ram_w4_l8192_id0_4_0_rdata = mem[ram_w4_l8192_id0_4_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_4_1_wenable) begin
      mem[ram_w4_l8192_id0_4_1_addr] <= ram_w4_l8192_id0_4_1_wdata;
    end 
    ram_w4_l8192_id0_4_1_daddr <= ram_w4_l8192_id0_4_1_addr;
  end

  assign ram_w4_l8192_id0_4_1_rdata = mem[ram_w4_l8192_id0_4_1_daddr];

endmodule



module ram_w4_l8192_id0_5
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id0_5_0_addr,
  output [4-1:0] ram_w4_l8192_id0_5_0_rdata,
  input [4-1:0] ram_w4_l8192_id0_5_0_wdata,
  input ram_w4_l8192_id0_5_0_wenable,
  input [10-1:0] ram_w4_l8192_id0_5_1_addr,
  output [4-1:0] ram_w4_l8192_id0_5_1_rdata,
  input [4-1:0] ram_w4_l8192_id0_5_1_wdata,
  input ram_w4_l8192_id0_5_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id0_5_0_daddr;
  reg [10-1:0] ram_w4_l8192_id0_5_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_5_0_wenable) begin
      mem[ram_w4_l8192_id0_5_0_addr] <= ram_w4_l8192_id0_5_0_wdata;
    end 
    ram_w4_l8192_id0_5_0_daddr <= ram_w4_l8192_id0_5_0_addr;
  end

  assign ram_w4_l8192_id0_5_0_rdata = mem[ram_w4_l8192_id0_5_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_5_1_wenable) begin
      mem[ram_w4_l8192_id0_5_1_addr] <= ram_w4_l8192_id0_5_1_wdata;
    end 
    ram_w4_l8192_id0_5_1_daddr <= ram_w4_l8192_id0_5_1_addr;
  end

  assign ram_w4_l8192_id0_5_1_rdata = mem[ram_w4_l8192_id0_5_1_daddr];

endmodule



module ram_w4_l8192_id0_6
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id0_6_0_addr,
  output [4-1:0] ram_w4_l8192_id0_6_0_rdata,
  input [4-1:0] ram_w4_l8192_id0_6_0_wdata,
  input ram_w4_l8192_id0_6_0_wenable,
  input [10-1:0] ram_w4_l8192_id0_6_1_addr,
  output [4-1:0] ram_w4_l8192_id0_6_1_rdata,
  input [4-1:0] ram_w4_l8192_id0_6_1_wdata,
  input ram_w4_l8192_id0_6_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id0_6_0_daddr;
  reg [10-1:0] ram_w4_l8192_id0_6_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_6_0_wenable) begin
      mem[ram_w4_l8192_id0_6_0_addr] <= ram_w4_l8192_id0_6_0_wdata;
    end 
    ram_w4_l8192_id0_6_0_daddr <= ram_w4_l8192_id0_6_0_addr;
  end

  assign ram_w4_l8192_id0_6_0_rdata = mem[ram_w4_l8192_id0_6_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_6_1_wenable) begin
      mem[ram_w4_l8192_id0_6_1_addr] <= ram_w4_l8192_id0_6_1_wdata;
    end 
    ram_w4_l8192_id0_6_1_daddr <= ram_w4_l8192_id0_6_1_addr;
  end

  assign ram_w4_l8192_id0_6_1_rdata = mem[ram_w4_l8192_id0_6_1_daddr];

endmodule



module ram_w4_l8192_id0_7
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id0_7_0_addr,
  output [4-1:0] ram_w4_l8192_id0_7_0_rdata,
  input [4-1:0] ram_w4_l8192_id0_7_0_wdata,
  input ram_w4_l8192_id0_7_0_wenable,
  input [10-1:0] ram_w4_l8192_id0_7_1_addr,
  output [4-1:0] ram_w4_l8192_id0_7_1_rdata,
  input [4-1:0] ram_w4_l8192_id0_7_1_wdata,
  input ram_w4_l8192_id0_7_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id0_7_0_daddr;
  reg [10-1:0] ram_w4_l8192_id0_7_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_7_0_wenable) begin
      mem[ram_w4_l8192_id0_7_0_addr] <= ram_w4_l8192_id0_7_0_wdata;
    end 
    ram_w4_l8192_id0_7_0_daddr <= ram_w4_l8192_id0_7_0_addr;
  end

  assign ram_w4_l8192_id0_7_0_rdata = mem[ram_w4_l8192_id0_7_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id0_7_1_wenable) begin
      mem[ram_w4_l8192_id0_7_1_addr] <= ram_w4_l8192_id0_7_1_wdata;
    end 
    ram_w4_l8192_id0_7_1_daddr <= ram_w4_l8192_id0_7_1_addr;
  end

  assign ram_w4_l8192_id0_7_1_rdata = mem[ram_w4_l8192_id0_7_1_daddr];

endmodule



module ram_w4_l8192_id1_0
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id1_0_0_addr,
  output [4-1:0] ram_w4_l8192_id1_0_0_rdata,
  input [4-1:0] ram_w4_l8192_id1_0_0_wdata,
  input ram_w4_l8192_id1_0_0_wenable,
  input [10-1:0] ram_w4_l8192_id1_0_1_addr,
  output [4-1:0] ram_w4_l8192_id1_0_1_rdata,
  input [4-1:0] ram_w4_l8192_id1_0_1_wdata,
  input ram_w4_l8192_id1_0_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id1_0_0_daddr;
  reg [10-1:0] ram_w4_l8192_id1_0_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_0_0_wenable) begin
      mem[ram_w4_l8192_id1_0_0_addr] <= ram_w4_l8192_id1_0_0_wdata;
    end 
    ram_w4_l8192_id1_0_0_daddr <= ram_w4_l8192_id1_0_0_addr;
  end

  assign ram_w4_l8192_id1_0_0_rdata = mem[ram_w4_l8192_id1_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_0_1_wenable) begin
      mem[ram_w4_l8192_id1_0_1_addr] <= ram_w4_l8192_id1_0_1_wdata;
    end 
    ram_w4_l8192_id1_0_1_daddr <= ram_w4_l8192_id1_0_1_addr;
  end

  assign ram_w4_l8192_id1_0_1_rdata = mem[ram_w4_l8192_id1_0_1_daddr];

endmodule



module ram_w4_l8192_id1_1
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id1_1_0_addr,
  output [4-1:0] ram_w4_l8192_id1_1_0_rdata,
  input [4-1:0] ram_w4_l8192_id1_1_0_wdata,
  input ram_w4_l8192_id1_1_0_wenable,
  input [10-1:0] ram_w4_l8192_id1_1_1_addr,
  output [4-1:0] ram_w4_l8192_id1_1_1_rdata,
  input [4-1:0] ram_w4_l8192_id1_1_1_wdata,
  input ram_w4_l8192_id1_1_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id1_1_0_daddr;
  reg [10-1:0] ram_w4_l8192_id1_1_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_1_0_wenable) begin
      mem[ram_w4_l8192_id1_1_0_addr] <= ram_w4_l8192_id1_1_0_wdata;
    end 
    ram_w4_l8192_id1_1_0_daddr <= ram_w4_l8192_id1_1_0_addr;
  end

  assign ram_w4_l8192_id1_1_0_rdata = mem[ram_w4_l8192_id1_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_1_1_wenable) begin
      mem[ram_w4_l8192_id1_1_1_addr] <= ram_w4_l8192_id1_1_1_wdata;
    end 
    ram_w4_l8192_id1_1_1_daddr <= ram_w4_l8192_id1_1_1_addr;
  end

  assign ram_w4_l8192_id1_1_1_rdata = mem[ram_w4_l8192_id1_1_1_daddr];

endmodule



module ram_w4_l8192_id1_2
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id1_2_0_addr,
  output [4-1:0] ram_w4_l8192_id1_2_0_rdata,
  input [4-1:0] ram_w4_l8192_id1_2_0_wdata,
  input ram_w4_l8192_id1_2_0_wenable,
  input [10-1:0] ram_w4_l8192_id1_2_1_addr,
  output [4-1:0] ram_w4_l8192_id1_2_1_rdata,
  input [4-1:0] ram_w4_l8192_id1_2_1_wdata,
  input ram_w4_l8192_id1_2_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id1_2_0_daddr;
  reg [10-1:0] ram_w4_l8192_id1_2_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_2_0_wenable) begin
      mem[ram_w4_l8192_id1_2_0_addr] <= ram_w4_l8192_id1_2_0_wdata;
    end 
    ram_w4_l8192_id1_2_0_daddr <= ram_w4_l8192_id1_2_0_addr;
  end

  assign ram_w4_l8192_id1_2_0_rdata = mem[ram_w4_l8192_id1_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_2_1_wenable) begin
      mem[ram_w4_l8192_id1_2_1_addr] <= ram_w4_l8192_id1_2_1_wdata;
    end 
    ram_w4_l8192_id1_2_1_daddr <= ram_w4_l8192_id1_2_1_addr;
  end

  assign ram_w4_l8192_id1_2_1_rdata = mem[ram_w4_l8192_id1_2_1_daddr];

endmodule



module ram_w4_l8192_id1_3
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id1_3_0_addr,
  output [4-1:0] ram_w4_l8192_id1_3_0_rdata,
  input [4-1:0] ram_w4_l8192_id1_3_0_wdata,
  input ram_w4_l8192_id1_3_0_wenable,
  input [10-1:0] ram_w4_l8192_id1_3_1_addr,
  output [4-1:0] ram_w4_l8192_id1_3_1_rdata,
  input [4-1:0] ram_w4_l8192_id1_3_1_wdata,
  input ram_w4_l8192_id1_3_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id1_3_0_daddr;
  reg [10-1:0] ram_w4_l8192_id1_3_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_3_0_wenable) begin
      mem[ram_w4_l8192_id1_3_0_addr] <= ram_w4_l8192_id1_3_0_wdata;
    end 
    ram_w4_l8192_id1_3_0_daddr <= ram_w4_l8192_id1_3_0_addr;
  end

  assign ram_w4_l8192_id1_3_0_rdata = mem[ram_w4_l8192_id1_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_3_1_wenable) begin
      mem[ram_w4_l8192_id1_3_1_addr] <= ram_w4_l8192_id1_3_1_wdata;
    end 
    ram_w4_l8192_id1_3_1_daddr <= ram_w4_l8192_id1_3_1_addr;
  end

  assign ram_w4_l8192_id1_3_1_rdata = mem[ram_w4_l8192_id1_3_1_daddr];

endmodule



module ram_w4_l8192_id1_4
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id1_4_0_addr,
  output [4-1:0] ram_w4_l8192_id1_4_0_rdata,
  input [4-1:0] ram_w4_l8192_id1_4_0_wdata,
  input ram_w4_l8192_id1_4_0_wenable,
  input [10-1:0] ram_w4_l8192_id1_4_1_addr,
  output [4-1:0] ram_w4_l8192_id1_4_1_rdata,
  input [4-1:0] ram_w4_l8192_id1_4_1_wdata,
  input ram_w4_l8192_id1_4_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id1_4_0_daddr;
  reg [10-1:0] ram_w4_l8192_id1_4_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_4_0_wenable) begin
      mem[ram_w4_l8192_id1_4_0_addr] <= ram_w4_l8192_id1_4_0_wdata;
    end 
    ram_w4_l8192_id1_4_0_daddr <= ram_w4_l8192_id1_4_0_addr;
  end

  assign ram_w4_l8192_id1_4_0_rdata = mem[ram_w4_l8192_id1_4_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_4_1_wenable) begin
      mem[ram_w4_l8192_id1_4_1_addr] <= ram_w4_l8192_id1_4_1_wdata;
    end 
    ram_w4_l8192_id1_4_1_daddr <= ram_w4_l8192_id1_4_1_addr;
  end

  assign ram_w4_l8192_id1_4_1_rdata = mem[ram_w4_l8192_id1_4_1_daddr];

endmodule



module ram_w4_l8192_id1_5
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id1_5_0_addr,
  output [4-1:0] ram_w4_l8192_id1_5_0_rdata,
  input [4-1:0] ram_w4_l8192_id1_5_0_wdata,
  input ram_w4_l8192_id1_5_0_wenable,
  input [10-1:0] ram_w4_l8192_id1_5_1_addr,
  output [4-1:0] ram_w4_l8192_id1_5_1_rdata,
  input [4-1:0] ram_w4_l8192_id1_5_1_wdata,
  input ram_w4_l8192_id1_5_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id1_5_0_daddr;
  reg [10-1:0] ram_w4_l8192_id1_5_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_5_0_wenable) begin
      mem[ram_w4_l8192_id1_5_0_addr] <= ram_w4_l8192_id1_5_0_wdata;
    end 
    ram_w4_l8192_id1_5_0_daddr <= ram_w4_l8192_id1_5_0_addr;
  end

  assign ram_w4_l8192_id1_5_0_rdata = mem[ram_w4_l8192_id1_5_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_5_1_wenable) begin
      mem[ram_w4_l8192_id1_5_1_addr] <= ram_w4_l8192_id1_5_1_wdata;
    end 
    ram_w4_l8192_id1_5_1_daddr <= ram_w4_l8192_id1_5_1_addr;
  end

  assign ram_w4_l8192_id1_5_1_rdata = mem[ram_w4_l8192_id1_5_1_daddr];

endmodule



module ram_w4_l8192_id1_6
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id1_6_0_addr,
  output [4-1:0] ram_w4_l8192_id1_6_0_rdata,
  input [4-1:0] ram_w4_l8192_id1_6_0_wdata,
  input ram_w4_l8192_id1_6_0_wenable,
  input [10-1:0] ram_w4_l8192_id1_6_1_addr,
  output [4-1:0] ram_w4_l8192_id1_6_1_rdata,
  input [4-1:0] ram_w4_l8192_id1_6_1_wdata,
  input ram_w4_l8192_id1_6_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id1_6_0_daddr;
  reg [10-1:0] ram_w4_l8192_id1_6_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_6_0_wenable) begin
      mem[ram_w4_l8192_id1_6_0_addr] <= ram_w4_l8192_id1_6_0_wdata;
    end 
    ram_w4_l8192_id1_6_0_daddr <= ram_w4_l8192_id1_6_0_addr;
  end

  assign ram_w4_l8192_id1_6_0_rdata = mem[ram_w4_l8192_id1_6_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_6_1_wenable) begin
      mem[ram_w4_l8192_id1_6_1_addr] <= ram_w4_l8192_id1_6_1_wdata;
    end 
    ram_w4_l8192_id1_6_1_daddr <= ram_w4_l8192_id1_6_1_addr;
  end

  assign ram_w4_l8192_id1_6_1_rdata = mem[ram_w4_l8192_id1_6_1_daddr];

endmodule



module ram_w4_l8192_id1_7
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id1_7_0_addr,
  output [4-1:0] ram_w4_l8192_id1_7_0_rdata,
  input [4-1:0] ram_w4_l8192_id1_7_0_wdata,
  input ram_w4_l8192_id1_7_0_wenable,
  input [10-1:0] ram_w4_l8192_id1_7_1_addr,
  output [4-1:0] ram_w4_l8192_id1_7_1_rdata,
  input [4-1:0] ram_w4_l8192_id1_7_1_wdata,
  input ram_w4_l8192_id1_7_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id1_7_0_daddr;
  reg [10-1:0] ram_w4_l8192_id1_7_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_7_0_wenable) begin
      mem[ram_w4_l8192_id1_7_0_addr] <= ram_w4_l8192_id1_7_0_wdata;
    end 
    ram_w4_l8192_id1_7_0_daddr <= ram_w4_l8192_id1_7_0_addr;
  end

  assign ram_w4_l8192_id1_7_0_rdata = mem[ram_w4_l8192_id1_7_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id1_7_1_wenable) begin
      mem[ram_w4_l8192_id1_7_1_addr] <= ram_w4_l8192_id1_7_1_wdata;
    end 
    ram_w4_l8192_id1_7_1_daddr <= ram_w4_l8192_id1_7_1_addr;
  end

  assign ram_w4_l8192_id1_7_1_rdata = mem[ram_w4_l8192_id1_7_1_daddr];

endmodule



module ram_w4_l8192_id2_0
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id2_0_0_addr,
  output [4-1:0] ram_w4_l8192_id2_0_0_rdata,
  input [4-1:0] ram_w4_l8192_id2_0_0_wdata,
  input ram_w4_l8192_id2_0_0_wenable,
  input [10-1:0] ram_w4_l8192_id2_0_1_addr,
  output [4-1:0] ram_w4_l8192_id2_0_1_rdata,
  input [4-1:0] ram_w4_l8192_id2_0_1_wdata,
  input ram_w4_l8192_id2_0_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id2_0_0_daddr;
  reg [10-1:0] ram_w4_l8192_id2_0_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_0_0_wenable) begin
      mem[ram_w4_l8192_id2_0_0_addr] <= ram_w4_l8192_id2_0_0_wdata;
    end 
    ram_w4_l8192_id2_0_0_daddr <= ram_w4_l8192_id2_0_0_addr;
  end

  assign ram_w4_l8192_id2_0_0_rdata = mem[ram_w4_l8192_id2_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_0_1_wenable) begin
      mem[ram_w4_l8192_id2_0_1_addr] <= ram_w4_l8192_id2_0_1_wdata;
    end 
    ram_w4_l8192_id2_0_1_daddr <= ram_w4_l8192_id2_0_1_addr;
  end

  assign ram_w4_l8192_id2_0_1_rdata = mem[ram_w4_l8192_id2_0_1_daddr];

endmodule



module ram_w4_l8192_id2_1
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id2_1_0_addr,
  output [4-1:0] ram_w4_l8192_id2_1_0_rdata,
  input [4-1:0] ram_w4_l8192_id2_1_0_wdata,
  input ram_w4_l8192_id2_1_0_wenable,
  input [10-1:0] ram_w4_l8192_id2_1_1_addr,
  output [4-1:0] ram_w4_l8192_id2_1_1_rdata,
  input [4-1:0] ram_w4_l8192_id2_1_1_wdata,
  input ram_w4_l8192_id2_1_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id2_1_0_daddr;
  reg [10-1:0] ram_w4_l8192_id2_1_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_1_0_wenable) begin
      mem[ram_w4_l8192_id2_1_0_addr] <= ram_w4_l8192_id2_1_0_wdata;
    end 
    ram_w4_l8192_id2_1_0_daddr <= ram_w4_l8192_id2_1_0_addr;
  end

  assign ram_w4_l8192_id2_1_0_rdata = mem[ram_w4_l8192_id2_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_1_1_wenable) begin
      mem[ram_w4_l8192_id2_1_1_addr] <= ram_w4_l8192_id2_1_1_wdata;
    end 
    ram_w4_l8192_id2_1_1_daddr <= ram_w4_l8192_id2_1_1_addr;
  end

  assign ram_w4_l8192_id2_1_1_rdata = mem[ram_w4_l8192_id2_1_1_daddr];

endmodule



module ram_w4_l8192_id2_2
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id2_2_0_addr,
  output [4-1:0] ram_w4_l8192_id2_2_0_rdata,
  input [4-1:0] ram_w4_l8192_id2_2_0_wdata,
  input ram_w4_l8192_id2_2_0_wenable,
  input [10-1:0] ram_w4_l8192_id2_2_1_addr,
  output [4-1:0] ram_w4_l8192_id2_2_1_rdata,
  input [4-1:0] ram_w4_l8192_id2_2_1_wdata,
  input ram_w4_l8192_id2_2_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id2_2_0_daddr;
  reg [10-1:0] ram_w4_l8192_id2_2_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_2_0_wenable) begin
      mem[ram_w4_l8192_id2_2_0_addr] <= ram_w4_l8192_id2_2_0_wdata;
    end 
    ram_w4_l8192_id2_2_0_daddr <= ram_w4_l8192_id2_2_0_addr;
  end

  assign ram_w4_l8192_id2_2_0_rdata = mem[ram_w4_l8192_id2_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_2_1_wenable) begin
      mem[ram_w4_l8192_id2_2_1_addr] <= ram_w4_l8192_id2_2_1_wdata;
    end 
    ram_w4_l8192_id2_2_1_daddr <= ram_w4_l8192_id2_2_1_addr;
  end

  assign ram_w4_l8192_id2_2_1_rdata = mem[ram_w4_l8192_id2_2_1_daddr];

endmodule



module ram_w4_l8192_id2_3
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id2_3_0_addr,
  output [4-1:0] ram_w4_l8192_id2_3_0_rdata,
  input [4-1:0] ram_w4_l8192_id2_3_0_wdata,
  input ram_w4_l8192_id2_3_0_wenable,
  input [10-1:0] ram_w4_l8192_id2_3_1_addr,
  output [4-1:0] ram_w4_l8192_id2_3_1_rdata,
  input [4-1:0] ram_w4_l8192_id2_3_1_wdata,
  input ram_w4_l8192_id2_3_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id2_3_0_daddr;
  reg [10-1:0] ram_w4_l8192_id2_3_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_3_0_wenable) begin
      mem[ram_w4_l8192_id2_3_0_addr] <= ram_w4_l8192_id2_3_0_wdata;
    end 
    ram_w4_l8192_id2_3_0_daddr <= ram_w4_l8192_id2_3_0_addr;
  end

  assign ram_w4_l8192_id2_3_0_rdata = mem[ram_w4_l8192_id2_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_3_1_wenable) begin
      mem[ram_w4_l8192_id2_3_1_addr] <= ram_w4_l8192_id2_3_1_wdata;
    end 
    ram_w4_l8192_id2_3_1_daddr <= ram_w4_l8192_id2_3_1_addr;
  end

  assign ram_w4_l8192_id2_3_1_rdata = mem[ram_w4_l8192_id2_3_1_daddr];

endmodule



module ram_w4_l8192_id2_4
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id2_4_0_addr,
  output [4-1:0] ram_w4_l8192_id2_4_0_rdata,
  input [4-1:0] ram_w4_l8192_id2_4_0_wdata,
  input ram_w4_l8192_id2_4_0_wenable,
  input [10-1:0] ram_w4_l8192_id2_4_1_addr,
  output [4-1:0] ram_w4_l8192_id2_4_1_rdata,
  input [4-1:0] ram_w4_l8192_id2_4_1_wdata,
  input ram_w4_l8192_id2_4_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id2_4_0_daddr;
  reg [10-1:0] ram_w4_l8192_id2_4_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_4_0_wenable) begin
      mem[ram_w4_l8192_id2_4_0_addr] <= ram_w4_l8192_id2_4_0_wdata;
    end 
    ram_w4_l8192_id2_4_0_daddr <= ram_w4_l8192_id2_4_0_addr;
  end

  assign ram_w4_l8192_id2_4_0_rdata = mem[ram_w4_l8192_id2_4_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_4_1_wenable) begin
      mem[ram_w4_l8192_id2_4_1_addr] <= ram_w4_l8192_id2_4_1_wdata;
    end 
    ram_w4_l8192_id2_4_1_daddr <= ram_w4_l8192_id2_4_1_addr;
  end

  assign ram_w4_l8192_id2_4_1_rdata = mem[ram_w4_l8192_id2_4_1_daddr];

endmodule



module ram_w4_l8192_id2_5
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id2_5_0_addr,
  output [4-1:0] ram_w4_l8192_id2_5_0_rdata,
  input [4-1:0] ram_w4_l8192_id2_5_0_wdata,
  input ram_w4_l8192_id2_5_0_wenable,
  input [10-1:0] ram_w4_l8192_id2_5_1_addr,
  output [4-1:0] ram_w4_l8192_id2_5_1_rdata,
  input [4-1:0] ram_w4_l8192_id2_5_1_wdata,
  input ram_w4_l8192_id2_5_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id2_5_0_daddr;
  reg [10-1:0] ram_w4_l8192_id2_5_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_5_0_wenable) begin
      mem[ram_w4_l8192_id2_5_0_addr] <= ram_w4_l8192_id2_5_0_wdata;
    end 
    ram_w4_l8192_id2_5_0_daddr <= ram_w4_l8192_id2_5_0_addr;
  end

  assign ram_w4_l8192_id2_5_0_rdata = mem[ram_w4_l8192_id2_5_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_5_1_wenable) begin
      mem[ram_w4_l8192_id2_5_1_addr] <= ram_w4_l8192_id2_5_1_wdata;
    end 
    ram_w4_l8192_id2_5_1_daddr <= ram_w4_l8192_id2_5_1_addr;
  end

  assign ram_w4_l8192_id2_5_1_rdata = mem[ram_w4_l8192_id2_5_1_daddr];

endmodule



module ram_w4_l8192_id2_6
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id2_6_0_addr,
  output [4-1:0] ram_w4_l8192_id2_6_0_rdata,
  input [4-1:0] ram_w4_l8192_id2_6_0_wdata,
  input ram_w4_l8192_id2_6_0_wenable,
  input [10-1:0] ram_w4_l8192_id2_6_1_addr,
  output [4-1:0] ram_w4_l8192_id2_6_1_rdata,
  input [4-1:0] ram_w4_l8192_id2_6_1_wdata,
  input ram_w4_l8192_id2_6_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id2_6_0_daddr;
  reg [10-1:0] ram_w4_l8192_id2_6_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_6_0_wenable) begin
      mem[ram_w4_l8192_id2_6_0_addr] <= ram_w4_l8192_id2_6_0_wdata;
    end 
    ram_w4_l8192_id2_6_0_daddr <= ram_w4_l8192_id2_6_0_addr;
  end

  assign ram_w4_l8192_id2_6_0_rdata = mem[ram_w4_l8192_id2_6_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_6_1_wenable) begin
      mem[ram_w4_l8192_id2_6_1_addr] <= ram_w4_l8192_id2_6_1_wdata;
    end 
    ram_w4_l8192_id2_6_1_daddr <= ram_w4_l8192_id2_6_1_addr;
  end

  assign ram_w4_l8192_id2_6_1_rdata = mem[ram_w4_l8192_id2_6_1_daddr];

endmodule



module ram_w4_l8192_id2_7
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id2_7_0_addr,
  output [4-1:0] ram_w4_l8192_id2_7_0_rdata,
  input [4-1:0] ram_w4_l8192_id2_7_0_wdata,
  input ram_w4_l8192_id2_7_0_wenable,
  input [10-1:0] ram_w4_l8192_id2_7_1_addr,
  output [4-1:0] ram_w4_l8192_id2_7_1_rdata,
  input [4-1:0] ram_w4_l8192_id2_7_1_wdata,
  input ram_w4_l8192_id2_7_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id2_7_0_daddr;
  reg [10-1:0] ram_w4_l8192_id2_7_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_7_0_wenable) begin
      mem[ram_w4_l8192_id2_7_0_addr] <= ram_w4_l8192_id2_7_0_wdata;
    end 
    ram_w4_l8192_id2_7_0_daddr <= ram_w4_l8192_id2_7_0_addr;
  end

  assign ram_w4_l8192_id2_7_0_rdata = mem[ram_w4_l8192_id2_7_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id2_7_1_wenable) begin
      mem[ram_w4_l8192_id2_7_1_addr] <= ram_w4_l8192_id2_7_1_wdata;
    end 
    ram_w4_l8192_id2_7_1_daddr <= ram_w4_l8192_id2_7_1_addr;
  end

  assign ram_w4_l8192_id2_7_1_rdata = mem[ram_w4_l8192_id2_7_1_daddr];

endmodule



module ram_w4_l8192_id3_0
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id3_0_0_addr,
  output [4-1:0] ram_w4_l8192_id3_0_0_rdata,
  input [4-1:0] ram_w4_l8192_id3_0_0_wdata,
  input ram_w4_l8192_id3_0_0_wenable,
  input [10-1:0] ram_w4_l8192_id3_0_1_addr,
  output [4-1:0] ram_w4_l8192_id3_0_1_rdata,
  input [4-1:0] ram_w4_l8192_id3_0_1_wdata,
  input ram_w4_l8192_id3_0_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id3_0_0_daddr;
  reg [10-1:0] ram_w4_l8192_id3_0_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_0_0_wenable) begin
      mem[ram_w4_l8192_id3_0_0_addr] <= ram_w4_l8192_id3_0_0_wdata;
    end 
    ram_w4_l8192_id3_0_0_daddr <= ram_w4_l8192_id3_0_0_addr;
  end

  assign ram_w4_l8192_id3_0_0_rdata = mem[ram_w4_l8192_id3_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_0_1_wenable) begin
      mem[ram_w4_l8192_id3_0_1_addr] <= ram_w4_l8192_id3_0_1_wdata;
    end 
    ram_w4_l8192_id3_0_1_daddr <= ram_w4_l8192_id3_0_1_addr;
  end

  assign ram_w4_l8192_id3_0_1_rdata = mem[ram_w4_l8192_id3_0_1_daddr];

endmodule



module ram_w4_l8192_id3_1
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id3_1_0_addr,
  output [4-1:0] ram_w4_l8192_id3_1_0_rdata,
  input [4-1:0] ram_w4_l8192_id3_1_0_wdata,
  input ram_w4_l8192_id3_1_0_wenable,
  input [10-1:0] ram_w4_l8192_id3_1_1_addr,
  output [4-1:0] ram_w4_l8192_id3_1_1_rdata,
  input [4-1:0] ram_w4_l8192_id3_1_1_wdata,
  input ram_w4_l8192_id3_1_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id3_1_0_daddr;
  reg [10-1:0] ram_w4_l8192_id3_1_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_1_0_wenable) begin
      mem[ram_w4_l8192_id3_1_0_addr] <= ram_w4_l8192_id3_1_0_wdata;
    end 
    ram_w4_l8192_id3_1_0_daddr <= ram_w4_l8192_id3_1_0_addr;
  end

  assign ram_w4_l8192_id3_1_0_rdata = mem[ram_w4_l8192_id3_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_1_1_wenable) begin
      mem[ram_w4_l8192_id3_1_1_addr] <= ram_w4_l8192_id3_1_1_wdata;
    end 
    ram_w4_l8192_id3_1_1_daddr <= ram_w4_l8192_id3_1_1_addr;
  end

  assign ram_w4_l8192_id3_1_1_rdata = mem[ram_w4_l8192_id3_1_1_daddr];

endmodule



module ram_w4_l8192_id3_2
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id3_2_0_addr,
  output [4-1:0] ram_w4_l8192_id3_2_0_rdata,
  input [4-1:0] ram_w4_l8192_id3_2_0_wdata,
  input ram_w4_l8192_id3_2_0_wenable,
  input [10-1:0] ram_w4_l8192_id3_2_1_addr,
  output [4-1:0] ram_w4_l8192_id3_2_1_rdata,
  input [4-1:0] ram_w4_l8192_id3_2_1_wdata,
  input ram_w4_l8192_id3_2_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id3_2_0_daddr;
  reg [10-1:0] ram_w4_l8192_id3_2_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_2_0_wenable) begin
      mem[ram_w4_l8192_id3_2_0_addr] <= ram_w4_l8192_id3_2_0_wdata;
    end 
    ram_w4_l8192_id3_2_0_daddr <= ram_w4_l8192_id3_2_0_addr;
  end

  assign ram_w4_l8192_id3_2_0_rdata = mem[ram_w4_l8192_id3_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_2_1_wenable) begin
      mem[ram_w4_l8192_id3_2_1_addr] <= ram_w4_l8192_id3_2_1_wdata;
    end 
    ram_w4_l8192_id3_2_1_daddr <= ram_w4_l8192_id3_2_1_addr;
  end

  assign ram_w4_l8192_id3_2_1_rdata = mem[ram_w4_l8192_id3_2_1_daddr];

endmodule



module ram_w4_l8192_id3_3
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id3_3_0_addr,
  output [4-1:0] ram_w4_l8192_id3_3_0_rdata,
  input [4-1:0] ram_w4_l8192_id3_3_0_wdata,
  input ram_w4_l8192_id3_3_0_wenable,
  input [10-1:0] ram_w4_l8192_id3_3_1_addr,
  output [4-1:0] ram_w4_l8192_id3_3_1_rdata,
  input [4-1:0] ram_w4_l8192_id3_3_1_wdata,
  input ram_w4_l8192_id3_3_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id3_3_0_daddr;
  reg [10-1:0] ram_w4_l8192_id3_3_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_3_0_wenable) begin
      mem[ram_w4_l8192_id3_3_0_addr] <= ram_w4_l8192_id3_3_0_wdata;
    end 
    ram_w4_l8192_id3_3_0_daddr <= ram_w4_l8192_id3_3_0_addr;
  end

  assign ram_w4_l8192_id3_3_0_rdata = mem[ram_w4_l8192_id3_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_3_1_wenable) begin
      mem[ram_w4_l8192_id3_3_1_addr] <= ram_w4_l8192_id3_3_1_wdata;
    end 
    ram_w4_l8192_id3_3_1_daddr <= ram_w4_l8192_id3_3_1_addr;
  end

  assign ram_w4_l8192_id3_3_1_rdata = mem[ram_w4_l8192_id3_3_1_daddr];

endmodule



module ram_w4_l8192_id3_4
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id3_4_0_addr,
  output [4-1:0] ram_w4_l8192_id3_4_0_rdata,
  input [4-1:0] ram_w4_l8192_id3_4_0_wdata,
  input ram_w4_l8192_id3_4_0_wenable,
  input [10-1:0] ram_w4_l8192_id3_4_1_addr,
  output [4-1:0] ram_w4_l8192_id3_4_1_rdata,
  input [4-1:0] ram_w4_l8192_id3_4_1_wdata,
  input ram_w4_l8192_id3_4_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id3_4_0_daddr;
  reg [10-1:0] ram_w4_l8192_id3_4_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_4_0_wenable) begin
      mem[ram_w4_l8192_id3_4_0_addr] <= ram_w4_l8192_id3_4_0_wdata;
    end 
    ram_w4_l8192_id3_4_0_daddr <= ram_w4_l8192_id3_4_0_addr;
  end

  assign ram_w4_l8192_id3_4_0_rdata = mem[ram_w4_l8192_id3_4_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_4_1_wenable) begin
      mem[ram_w4_l8192_id3_4_1_addr] <= ram_w4_l8192_id3_4_1_wdata;
    end 
    ram_w4_l8192_id3_4_1_daddr <= ram_w4_l8192_id3_4_1_addr;
  end

  assign ram_w4_l8192_id3_4_1_rdata = mem[ram_w4_l8192_id3_4_1_daddr];

endmodule



module ram_w4_l8192_id3_5
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id3_5_0_addr,
  output [4-1:0] ram_w4_l8192_id3_5_0_rdata,
  input [4-1:0] ram_w4_l8192_id3_5_0_wdata,
  input ram_w4_l8192_id3_5_0_wenable,
  input [10-1:0] ram_w4_l8192_id3_5_1_addr,
  output [4-1:0] ram_w4_l8192_id3_5_1_rdata,
  input [4-1:0] ram_w4_l8192_id3_5_1_wdata,
  input ram_w4_l8192_id3_5_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id3_5_0_daddr;
  reg [10-1:0] ram_w4_l8192_id3_5_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_5_0_wenable) begin
      mem[ram_w4_l8192_id3_5_0_addr] <= ram_w4_l8192_id3_5_0_wdata;
    end 
    ram_w4_l8192_id3_5_0_daddr <= ram_w4_l8192_id3_5_0_addr;
  end

  assign ram_w4_l8192_id3_5_0_rdata = mem[ram_w4_l8192_id3_5_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_5_1_wenable) begin
      mem[ram_w4_l8192_id3_5_1_addr] <= ram_w4_l8192_id3_5_1_wdata;
    end 
    ram_w4_l8192_id3_5_1_daddr <= ram_w4_l8192_id3_5_1_addr;
  end

  assign ram_w4_l8192_id3_5_1_rdata = mem[ram_w4_l8192_id3_5_1_daddr];

endmodule



module ram_w4_l8192_id3_6
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id3_6_0_addr,
  output [4-1:0] ram_w4_l8192_id3_6_0_rdata,
  input [4-1:0] ram_w4_l8192_id3_6_0_wdata,
  input ram_w4_l8192_id3_6_0_wenable,
  input [10-1:0] ram_w4_l8192_id3_6_1_addr,
  output [4-1:0] ram_w4_l8192_id3_6_1_rdata,
  input [4-1:0] ram_w4_l8192_id3_6_1_wdata,
  input ram_w4_l8192_id3_6_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id3_6_0_daddr;
  reg [10-1:0] ram_w4_l8192_id3_6_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_6_0_wenable) begin
      mem[ram_w4_l8192_id3_6_0_addr] <= ram_w4_l8192_id3_6_0_wdata;
    end 
    ram_w4_l8192_id3_6_0_daddr <= ram_w4_l8192_id3_6_0_addr;
  end

  assign ram_w4_l8192_id3_6_0_rdata = mem[ram_w4_l8192_id3_6_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_6_1_wenable) begin
      mem[ram_w4_l8192_id3_6_1_addr] <= ram_w4_l8192_id3_6_1_wdata;
    end 
    ram_w4_l8192_id3_6_1_daddr <= ram_w4_l8192_id3_6_1_addr;
  end

  assign ram_w4_l8192_id3_6_1_rdata = mem[ram_w4_l8192_id3_6_1_daddr];

endmodule



module ram_w4_l8192_id3_7
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id3_7_0_addr,
  output [4-1:0] ram_w4_l8192_id3_7_0_rdata,
  input [4-1:0] ram_w4_l8192_id3_7_0_wdata,
  input ram_w4_l8192_id3_7_0_wenable,
  input [10-1:0] ram_w4_l8192_id3_7_1_addr,
  output [4-1:0] ram_w4_l8192_id3_7_1_rdata,
  input [4-1:0] ram_w4_l8192_id3_7_1_wdata,
  input ram_w4_l8192_id3_7_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id3_7_0_daddr;
  reg [10-1:0] ram_w4_l8192_id3_7_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_7_0_wenable) begin
      mem[ram_w4_l8192_id3_7_0_addr] <= ram_w4_l8192_id3_7_0_wdata;
    end 
    ram_w4_l8192_id3_7_0_daddr <= ram_w4_l8192_id3_7_0_addr;
  end

  assign ram_w4_l8192_id3_7_0_rdata = mem[ram_w4_l8192_id3_7_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id3_7_1_wenable) begin
      mem[ram_w4_l8192_id3_7_1_addr] <= ram_w4_l8192_id3_7_1_wdata;
    end 
    ram_w4_l8192_id3_7_1_daddr <= ram_w4_l8192_id3_7_1_addr;
  end

  assign ram_w4_l8192_id3_7_1_rdata = mem[ram_w4_l8192_id3_7_1_daddr];

endmodule



module ram_w4_l8192_id4_0
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id4_0_0_addr,
  output [4-1:0] ram_w4_l8192_id4_0_0_rdata,
  input [4-1:0] ram_w4_l8192_id4_0_0_wdata,
  input ram_w4_l8192_id4_0_0_wenable,
  input [10-1:0] ram_w4_l8192_id4_0_1_addr,
  output [4-1:0] ram_w4_l8192_id4_0_1_rdata,
  input [4-1:0] ram_w4_l8192_id4_0_1_wdata,
  input ram_w4_l8192_id4_0_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id4_0_0_daddr;
  reg [10-1:0] ram_w4_l8192_id4_0_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_0_0_wenable) begin
      mem[ram_w4_l8192_id4_0_0_addr] <= ram_w4_l8192_id4_0_0_wdata;
    end 
    ram_w4_l8192_id4_0_0_daddr <= ram_w4_l8192_id4_0_0_addr;
  end

  assign ram_w4_l8192_id4_0_0_rdata = mem[ram_w4_l8192_id4_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_0_1_wenable) begin
      mem[ram_w4_l8192_id4_0_1_addr] <= ram_w4_l8192_id4_0_1_wdata;
    end 
    ram_w4_l8192_id4_0_1_daddr <= ram_w4_l8192_id4_0_1_addr;
  end

  assign ram_w4_l8192_id4_0_1_rdata = mem[ram_w4_l8192_id4_0_1_daddr];

endmodule



module ram_w4_l8192_id4_1
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id4_1_0_addr,
  output [4-1:0] ram_w4_l8192_id4_1_0_rdata,
  input [4-1:0] ram_w4_l8192_id4_1_0_wdata,
  input ram_w4_l8192_id4_1_0_wenable,
  input [10-1:0] ram_w4_l8192_id4_1_1_addr,
  output [4-1:0] ram_w4_l8192_id4_1_1_rdata,
  input [4-1:0] ram_w4_l8192_id4_1_1_wdata,
  input ram_w4_l8192_id4_1_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id4_1_0_daddr;
  reg [10-1:0] ram_w4_l8192_id4_1_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_1_0_wenable) begin
      mem[ram_w4_l8192_id4_1_0_addr] <= ram_w4_l8192_id4_1_0_wdata;
    end 
    ram_w4_l8192_id4_1_0_daddr <= ram_w4_l8192_id4_1_0_addr;
  end

  assign ram_w4_l8192_id4_1_0_rdata = mem[ram_w4_l8192_id4_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_1_1_wenable) begin
      mem[ram_w4_l8192_id4_1_1_addr] <= ram_w4_l8192_id4_1_1_wdata;
    end 
    ram_w4_l8192_id4_1_1_daddr <= ram_w4_l8192_id4_1_1_addr;
  end

  assign ram_w4_l8192_id4_1_1_rdata = mem[ram_w4_l8192_id4_1_1_daddr];

endmodule



module ram_w4_l8192_id4_2
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id4_2_0_addr,
  output [4-1:0] ram_w4_l8192_id4_2_0_rdata,
  input [4-1:0] ram_w4_l8192_id4_2_0_wdata,
  input ram_w4_l8192_id4_2_0_wenable,
  input [10-1:0] ram_w4_l8192_id4_2_1_addr,
  output [4-1:0] ram_w4_l8192_id4_2_1_rdata,
  input [4-1:0] ram_w4_l8192_id4_2_1_wdata,
  input ram_w4_l8192_id4_2_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id4_2_0_daddr;
  reg [10-1:0] ram_w4_l8192_id4_2_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_2_0_wenable) begin
      mem[ram_w4_l8192_id4_2_0_addr] <= ram_w4_l8192_id4_2_0_wdata;
    end 
    ram_w4_l8192_id4_2_0_daddr <= ram_w4_l8192_id4_2_0_addr;
  end

  assign ram_w4_l8192_id4_2_0_rdata = mem[ram_w4_l8192_id4_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_2_1_wenable) begin
      mem[ram_w4_l8192_id4_2_1_addr] <= ram_w4_l8192_id4_2_1_wdata;
    end 
    ram_w4_l8192_id4_2_1_daddr <= ram_w4_l8192_id4_2_1_addr;
  end

  assign ram_w4_l8192_id4_2_1_rdata = mem[ram_w4_l8192_id4_2_1_daddr];

endmodule



module ram_w4_l8192_id4_3
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id4_3_0_addr,
  output [4-1:0] ram_w4_l8192_id4_3_0_rdata,
  input [4-1:0] ram_w4_l8192_id4_3_0_wdata,
  input ram_w4_l8192_id4_3_0_wenable,
  input [10-1:0] ram_w4_l8192_id4_3_1_addr,
  output [4-1:0] ram_w4_l8192_id4_3_1_rdata,
  input [4-1:0] ram_w4_l8192_id4_3_1_wdata,
  input ram_w4_l8192_id4_3_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id4_3_0_daddr;
  reg [10-1:0] ram_w4_l8192_id4_3_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_3_0_wenable) begin
      mem[ram_w4_l8192_id4_3_0_addr] <= ram_w4_l8192_id4_3_0_wdata;
    end 
    ram_w4_l8192_id4_3_0_daddr <= ram_w4_l8192_id4_3_0_addr;
  end

  assign ram_w4_l8192_id4_3_0_rdata = mem[ram_w4_l8192_id4_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_3_1_wenable) begin
      mem[ram_w4_l8192_id4_3_1_addr] <= ram_w4_l8192_id4_3_1_wdata;
    end 
    ram_w4_l8192_id4_3_1_daddr <= ram_w4_l8192_id4_3_1_addr;
  end

  assign ram_w4_l8192_id4_3_1_rdata = mem[ram_w4_l8192_id4_3_1_daddr];

endmodule



module ram_w4_l8192_id4_4
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id4_4_0_addr,
  output [4-1:0] ram_w4_l8192_id4_4_0_rdata,
  input [4-1:0] ram_w4_l8192_id4_4_0_wdata,
  input ram_w4_l8192_id4_4_0_wenable,
  input [10-1:0] ram_w4_l8192_id4_4_1_addr,
  output [4-1:0] ram_w4_l8192_id4_4_1_rdata,
  input [4-1:0] ram_w4_l8192_id4_4_1_wdata,
  input ram_w4_l8192_id4_4_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id4_4_0_daddr;
  reg [10-1:0] ram_w4_l8192_id4_4_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_4_0_wenable) begin
      mem[ram_w4_l8192_id4_4_0_addr] <= ram_w4_l8192_id4_4_0_wdata;
    end 
    ram_w4_l8192_id4_4_0_daddr <= ram_w4_l8192_id4_4_0_addr;
  end

  assign ram_w4_l8192_id4_4_0_rdata = mem[ram_w4_l8192_id4_4_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_4_1_wenable) begin
      mem[ram_w4_l8192_id4_4_1_addr] <= ram_w4_l8192_id4_4_1_wdata;
    end 
    ram_w4_l8192_id4_4_1_daddr <= ram_w4_l8192_id4_4_1_addr;
  end

  assign ram_w4_l8192_id4_4_1_rdata = mem[ram_w4_l8192_id4_4_1_daddr];

endmodule



module ram_w4_l8192_id4_5
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id4_5_0_addr,
  output [4-1:0] ram_w4_l8192_id4_5_0_rdata,
  input [4-1:0] ram_w4_l8192_id4_5_0_wdata,
  input ram_w4_l8192_id4_5_0_wenable,
  input [10-1:0] ram_w4_l8192_id4_5_1_addr,
  output [4-1:0] ram_w4_l8192_id4_5_1_rdata,
  input [4-1:0] ram_w4_l8192_id4_5_1_wdata,
  input ram_w4_l8192_id4_5_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id4_5_0_daddr;
  reg [10-1:0] ram_w4_l8192_id4_5_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_5_0_wenable) begin
      mem[ram_w4_l8192_id4_5_0_addr] <= ram_w4_l8192_id4_5_0_wdata;
    end 
    ram_w4_l8192_id4_5_0_daddr <= ram_w4_l8192_id4_5_0_addr;
  end

  assign ram_w4_l8192_id4_5_0_rdata = mem[ram_w4_l8192_id4_5_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_5_1_wenable) begin
      mem[ram_w4_l8192_id4_5_1_addr] <= ram_w4_l8192_id4_5_1_wdata;
    end 
    ram_w4_l8192_id4_5_1_daddr <= ram_w4_l8192_id4_5_1_addr;
  end

  assign ram_w4_l8192_id4_5_1_rdata = mem[ram_w4_l8192_id4_5_1_daddr];

endmodule



module ram_w4_l8192_id4_6
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id4_6_0_addr,
  output [4-1:0] ram_w4_l8192_id4_6_0_rdata,
  input [4-1:0] ram_w4_l8192_id4_6_0_wdata,
  input ram_w4_l8192_id4_6_0_wenable,
  input [10-1:0] ram_w4_l8192_id4_6_1_addr,
  output [4-1:0] ram_w4_l8192_id4_6_1_rdata,
  input [4-1:0] ram_w4_l8192_id4_6_1_wdata,
  input ram_w4_l8192_id4_6_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id4_6_0_daddr;
  reg [10-1:0] ram_w4_l8192_id4_6_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_6_0_wenable) begin
      mem[ram_w4_l8192_id4_6_0_addr] <= ram_w4_l8192_id4_6_0_wdata;
    end 
    ram_w4_l8192_id4_6_0_daddr <= ram_w4_l8192_id4_6_0_addr;
  end

  assign ram_w4_l8192_id4_6_0_rdata = mem[ram_w4_l8192_id4_6_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_6_1_wenable) begin
      mem[ram_w4_l8192_id4_6_1_addr] <= ram_w4_l8192_id4_6_1_wdata;
    end 
    ram_w4_l8192_id4_6_1_daddr <= ram_w4_l8192_id4_6_1_addr;
  end

  assign ram_w4_l8192_id4_6_1_rdata = mem[ram_w4_l8192_id4_6_1_daddr];

endmodule



module ram_w4_l8192_id4_7
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id4_7_0_addr,
  output [4-1:0] ram_w4_l8192_id4_7_0_rdata,
  input [4-1:0] ram_w4_l8192_id4_7_0_wdata,
  input ram_w4_l8192_id4_7_0_wenable,
  input [10-1:0] ram_w4_l8192_id4_7_1_addr,
  output [4-1:0] ram_w4_l8192_id4_7_1_rdata,
  input [4-1:0] ram_w4_l8192_id4_7_1_wdata,
  input ram_w4_l8192_id4_7_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id4_7_0_daddr;
  reg [10-1:0] ram_w4_l8192_id4_7_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_7_0_wenable) begin
      mem[ram_w4_l8192_id4_7_0_addr] <= ram_w4_l8192_id4_7_0_wdata;
    end 
    ram_w4_l8192_id4_7_0_daddr <= ram_w4_l8192_id4_7_0_addr;
  end

  assign ram_w4_l8192_id4_7_0_rdata = mem[ram_w4_l8192_id4_7_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id4_7_1_wenable) begin
      mem[ram_w4_l8192_id4_7_1_addr] <= ram_w4_l8192_id4_7_1_wdata;
    end 
    ram_w4_l8192_id4_7_1_daddr <= ram_w4_l8192_id4_7_1_addr;
  end

  assign ram_w4_l8192_id4_7_1_rdata = mem[ram_w4_l8192_id4_7_1_daddr];

endmodule



module ram_w4_l8192_id5_0
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id5_0_0_addr,
  output [4-1:0] ram_w4_l8192_id5_0_0_rdata,
  input [4-1:0] ram_w4_l8192_id5_0_0_wdata,
  input ram_w4_l8192_id5_0_0_wenable,
  input [10-1:0] ram_w4_l8192_id5_0_1_addr,
  output [4-1:0] ram_w4_l8192_id5_0_1_rdata,
  input [4-1:0] ram_w4_l8192_id5_0_1_wdata,
  input ram_w4_l8192_id5_0_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id5_0_0_daddr;
  reg [10-1:0] ram_w4_l8192_id5_0_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_0_0_wenable) begin
      mem[ram_w4_l8192_id5_0_0_addr] <= ram_w4_l8192_id5_0_0_wdata;
    end 
    ram_w4_l8192_id5_0_0_daddr <= ram_w4_l8192_id5_0_0_addr;
  end

  assign ram_w4_l8192_id5_0_0_rdata = mem[ram_w4_l8192_id5_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_0_1_wenable) begin
      mem[ram_w4_l8192_id5_0_1_addr] <= ram_w4_l8192_id5_0_1_wdata;
    end 
    ram_w4_l8192_id5_0_1_daddr <= ram_w4_l8192_id5_0_1_addr;
  end

  assign ram_w4_l8192_id5_0_1_rdata = mem[ram_w4_l8192_id5_0_1_daddr];

endmodule



module ram_w4_l8192_id5_1
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id5_1_0_addr,
  output [4-1:0] ram_w4_l8192_id5_1_0_rdata,
  input [4-1:0] ram_w4_l8192_id5_1_0_wdata,
  input ram_w4_l8192_id5_1_0_wenable,
  input [10-1:0] ram_w4_l8192_id5_1_1_addr,
  output [4-1:0] ram_w4_l8192_id5_1_1_rdata,
  input [4-1:0] ram_w4_l8192_id5_1_1_wdata,
  input ram_w4_l8192_id5_1_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id5_1_0_daddr;
  reg [10-1:0] ram_w4_l8192_id5_1_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_1_0_wenable) begin
      mem[ram_w4_l8192_id5_1_0_addr] <= ram_w4_l8192_id5_1_0_wdata;
    end 
    ram_w4_l8192_id5_1_0_daddr <= ram_w4_l8192_id5_1_0_addr;
  end

  assign ram_w4_l8192_id5_1_0_rdata = mem[ram_w4_l8192_id5_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_1_1_wenable) begin
      mem[ram_w4_l8192_id5_1_1_addr] <= ram_w4_l8192_id5_1_1_wdata;
    end 
    ram_w4_l8192_id5_1_1_daddr <= ram_w4_l8192_id5_1_1_addr;
  end

  assign ram_w4_l8192_id5_1_1_rdata = mem[ram_w4_l8192_id5_1_1_daddr];

endmodule



module ram_w4_l8192_id5_2
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id5_2_0_addr,
  output [4-1:0] ram_w4_l8192_id5_2_0_rdata,
  input [4-1:0] ram_w4_l8192_id5_2_0_wdata,
  input ram_w4_l8192_id5_2_0_wenable,
  input [10-1:0] ram_w4_l8192_id5_2_1_addr,
  output [4-1:0] ram_w4_l8192_id5_2_1_rdata,
  input [4-1:0] ram_w4_l8192_id5_2_1_wdata,
  input ram_w4_l8192_id5_2_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id5_2_0_daddr;
  reg [10-1:0] ram_w4_l8192_id5_2_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_2_0_wenable) begin
      mem[ram_w4_l8192_id5_2_0_addr] <= ram_w4_l8192_id5_2_0_wdata;
    end 
    ram_w4_l8192_id5_2_0_daddr <= ram_w4_l8192_id5_2_0_addr;
  end

  assign ram_w4_l8192_id5_2_0_rdata = mem[ram_w4_l8192_id5_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_2_1_wenable) begin
      mem[ram_w4_l8192_id5_2_1_addr] <= ram_w4_l8192_id5_2_1_wdata;
    end 
    ram_w4_l8192_id5_2_1_daddr <= ram_w4_l8192_id5_2_1_addr;
  end

  assign ram_w4_l8192_id5_2_1_rdata = mem[ram_w4_l8192_id5_2_1_daddr];

endmodule



module ram_w4_l8192_id5_3
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id5_3_0_addr,
  output [4-1:0] ram_w4_l8192_id5_3_0_rdata,
  input [4-1:0] ram_w4_l8192_id5_3_0_wdata,
  input ram_w4_l8192_id5_3_0_wenable,
  input [10-1:0] ram_w4_l8192_id5_3_1_addr,
  output [4-1:0] ram_w4_l8192_id5_3_1_rdata,
  input [4-1:0] ram_w4_l8192_id5_3_1_wdata,
  input ram_w4_l8192_id5_3_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id5_3_0_daddr;
  reg [10-1:0] ram_w4_l8192_id5_3_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_3_0_wenable) begin
      mem[ram_w4_l8192_id5_3_0_addr] <= ram_w4_l8192_id5_3_0_wdata;
    end 
    ram_w4_l8192_id5_3_0_daddr <= ram_w4_l8192_id5_3_0_addr;
  end

  assign ram_w4_l8192_id5_3_0_rdata = mem[ram_w4_l8192_id5_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_3_1_wenable) begin
      mem[ram_w4_l8192_id5_3_1_addr] <= ram_w4_l8192_id5_3_1_wdata;
    end 
    ram_w4_l8192_id5_3_1_daddr <= ram_w4_l8192_id5_3_1_addr;
  end

  assign ram_w4_l8192_id5_3_1_rdata = mem[ram_w4_l8192_id5_3_1_daddr];

endmodule



module ram_w4_l8192_id5_4
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id5_4_0_addr,
  output [4-1:0] ram_w4_l8192_id5_4_0_rdata,
  input [4-1:0] ram_w4_l8192_id5_4_0_wdata,
  input ram_w4_l8192_id5_4_0_wenable,
  input [10-1:0] ram_w4_l8192_id5_4_1_addr,
  output [4-1:0] ram_w4_l8192_id5_4_1_rdata,
  input [4-1:0] ram_w4_l8192_id5_4_1_wdata,
  input ram_w4_l8192_id5_4_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id5_4_0_daddr;
  reg [10-1:0] ram_w4_l8192_id5_4_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_4_0_wenable) begin
      mem[ram_w4_l8192_id5_4_0_addr] <= ram_w4_l8192_id5_4_0_wdata;
    end 
    ram_w4_l8192_id5_4_0_daddr <= ram_w4_l8192_id5_4_0_addr;
  end

  assign ram_w4_l8192_id5_4_0_rdata = mem[ram_w4_l8192_id5_4_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_4_1_wenable) begin
      mem[ram_w4_l8192_id5_4_1_addr] <= ram_w4_l8192_id5_4_1_wdata;
    end 
    ram_w4_l8192_id5_4_1_daddr <= ram_w4_l8192_id5_4_1_addr;
  end

  assign ram_w4_l8192_id5_4_1_rdata = mem[ram_w4_l8192_id5_4_1_daddr];

endmodule



module ram_w4_l8192_id5_5
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id5_5_0_addr,
  output [4-1:0] ram_w4_l8192_id5_5_0_rdata,
  input [4-1:0] ram_w4_l8192_id5_5_0_wdata,
  input ram_w4_l8192_id5_5_0_wenable,
  input [10-1:0] ram_w4_l8192_id5_5_1_addr,
  output [4-1:0] ram_w4_l8192_id5_5_1_rdata,
  input [4-1:0] ram_w4_l8192_id5_5_1_wdata,
  input ram_w4_l8192_id5_5_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id5_5_0_daddr;
  reg [10-1:0] ram_w4_l8192_id5_5_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_5_0_wenable) begin
      mem[ram_w4_l8192_id5_5_0_addr] <= ram_w4_l8192_id5_5_0_wdata;
    end 
    ram_w4_l8192_id5_5_0_daddr <= ram_w4_l8192_id5_5_0_addr;
  end

  assign ram_w4_l8192_id5_5_0_rdata = mem[ram_w4_l8192_id5_5_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_5_1_wenable) begin
      mem[ram_w4_l8192_id5_5_1_addr] <= ram_w4_l8192_id5_5_1_wdata;
    end 
    ram_w4_l8192_id5_5_1_daddr <= ram_w4_l8192_id5_5_1_addr;
  end

  assign ram_w4_l8192_id5_5_1_rdata = mem[ram_w4_l8192_id5_5_1_daddr];

endmodule



module ram_w4_l8192_id5_6
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id5_6_0_addr,
  output [4-1:0] ram_w4_l8192_id5_6_0_rdata,
  input [4-1:0] ram_w4_l8192_id5_6_0_wdata,
  input ram_w4_l8192_id5_6_0_wenable,
  input [10-1:0] ram_w4_l8192_id5_6_1_addr,
  output [4-1:0] ram_w4_l8192_id5_6_1_rdata,
  input [4-1:0] ram_w4_l8192_id5_6_1_wdata,
  input ram_w4_l8192_id5_6_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id5_6_0_daddr;
  reg [10-1:0] ram_w4_l8192_id5_6_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_6_0_wenable) begin
      mem[ram_w4_l8192_id5_6_0_addr] <= ram_w4_l8192_id5_6_0_wdata;
    end 
    ram_w4_l8192_id5_6_0_daddr <= ram_w4_l8192_id5_6_0_addr;
  end

  assign ram_w4_l8192_id5_6_0_rdata = mem[ram_w4_l8192_id5_6_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_6_1_wenable) begin
      mem[ram_w4_l8192_id5_6_1_addr] <= ram_w4_l8192_id5_6_1_wdata;
    end 
    ram_w4_l8192_id5_6_1_daddr <= ram_w4_l8192_id5_6_1_addr;
  end

  assign ram_w4_l8192_id5_6_1_rdata = mem[ram_w4_l8192_id5_6_1_daddr];

endmodule



module ram_w4_l8192_id5_7
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id5_7_0_addr,
  output [4-1:0] ram_w4_l8192_id5_7_0_rdata,
  input [4-1:0] ram_w4_l8192_id5_7_0_wdata,
  input ram_w4_l8192_id5_7_0_wenable,
  input [10-1:0] ram_w4_l8192_id5_7_1_addr,
  output [4-1:0] ram_w4_l8192_id5_7_1_rdata,
  input [4-1:0] ram_w4_l8192_id5_7_1_wdata,
  input ram_w4_l8192_id5_7_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id5_7_0_daddr;
  reg [10-1:0] ram_w4_l8192_id5_7_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_7_0_wenable) begin
      mem[ram_w4_l8192_id5_7_0_addr] <= ram_w4_l8192_id5_7_0_wdata;
    end 
    ram_w4_l8192_id5_7_0_daddr <= ram_w4_l8192_id5_7_0_addr;
  end

  assign ram_w4_l8192_id5_7_0_rdata = mem[ram_w4_l8192_id5_7_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id5_7_1_wenable) begin
      mem[ram_w4_l8192_id5_7_1_addr] <= ram_w4_l8192_id5_7_1_wdata;
    end 
    ram_w4_l8192_id5_7_1_daddr <= ram_w4_l8192_id5_7_1_addr;
  end

  assign ram_w4_l8192_id5_7_1_rdata = mem[ram_w4_l8192_id5_7_1_daddr];

endmodule



module ram_w4_l8192_id6_0
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id6_0_0_addr,
  output [4-1:0] ram_w4_l8192_id6_0_0_rdata,
  input [4-1:0] ram_w4_l8192_id6_0_0_wdata,
  input ram_w4_l8192_id6_0_0_wenable,
  input [10-1:0] ram_w4_l8192_id6_0_1_addr,
  output [4-1:0] ram_w4_l8192_id6_0_1_rdata,
  input [4-1:0] ram_w4_l8192_id6_0_1_wdata,
  input ram_w4_l8192_id6_0_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id6_0_0_daddr;
  reg [10-1:0] ram_w4_l8192_id6_0_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_0_0_wenable) begin
      mem[ram_w4_l8192_id6_0_0_addr] <= ram_w4_l8192_id6_0_0_wdata;
    end 
    ram_w4_l8192_id6_0_0_daddr <= ram_w4_l8192_id6_0_0_addr;
  end

  assign ram_w4_l8192_id6_0_0_rdata = mem[ram_w4_l8192_id6_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_0_1_wenable) begin
      mem[ram_w4_l8192_id6_0_1_addr] <= ram_w4_l8192_id6_0_1_wdata;
    end 
    ram_w4_l8192_id6_0_1_daddr <= ram_w4_l8192_id6_0_1_addr;
  end

  assign ram_w4_l8192_id6_0_1_rdata = mem[ram_w4_l8192_id6_0_1_daddr];

endmodule



module ram_w4_l8192_id6_1
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id6_1_0_addr,
  output [4-1:0] ram_w4_l8192_id6_1_0_rdata,
  input [4-1:0] ram_w4_l8192_id6_1_0_wdata,
  input ram_w4_l8192_id6_1_0_wenable,
  input [10-1:0] ram_w4_l8192_id6_1_1_addr,
  output [4-1:0] ram_w4_l8192_id6_1_1_rdata,
  input [4-1:0] ram_w4_l8192_id6_1_1_wdata,
  input ram_w4_l8192_id6_1_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id6_1_0_daddr;
  reg [10-1:0] ram_w4_l8192_id6_1_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_1_0_wenable) begin
      mem[ram_w4_l8192_id6_1_0_addr] <= ram_w4_l8192_id6_1_0_wdata;
    end 
    ram_w4_l8192_id6_1_0_daddr <= ram_w4_l8192_id6_1_0_addr;
  end

  assign ram_w4_l8192_id6_1_0_rdata = mem[ram_w4_l8192_id6_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_1_1_wenable) begin
      mem[ram_w4_l8192_id6_1_1_addr] <= ram_w4_l8192_id6_1_1_wdata;
    end 
    ram_w4_l8192_id6_1_1_daddr <= ram_w4_l8192_id6_1_1_addr;
  end

  assign ram_w4_l8192_id6_1_1_rdata = mem[ram_w4_l8192_id6_1_1_daddr];

endmodule



module ram_w4_l8192_id6_2
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id6_2_0_addr,
  output [4-1:0] ram_w4_l8192_id6_2_0_rdata,
  input [4-1:0] ram_w4_l8192_id6_2_0_wdata,
  input ram_w4_l8192_id6_2_0_wenable,
  input [10-1:0] ram_w4_l8192_id6_2_1_addr,
  output [4-1:0] ram_w4_l8192_id6_2_1_rdata,
  input [4-1:0] ram_w4_l8192_id6_2_1_wdata,
  input ram_w4_l8192_id6_2_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id6_2_0_daddr;
  reg [10-1:0] ram_w4_l8192_id6_2_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_2_0_wenable) begin
      mem[ram_w4_l8192_id6_2_0_addr] <= ram_w4_l8192_id6_2_0_wdata;
    end 
    ram_w4_l8192_id6_2_0_daddr <= ram_w4_l8192_id6_2_0_addr;
  end

  assign ram_w4_l8192_id6_2_0_rdata = mem[ram_w4_l8192_id6_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_2_1_wenable) begin
      mem[ram_w4_l8192_id6_2_1_addr] <= ram_w4_l8192_id6_2_1_wdata;
    end 
    ram_w4_l8192_id6_2_1_daddr <= ram_w4_l8192_id6_2_1_addr;
  end

  assign ram_w4_l8192_id6_2_1_rdata = mem[ram_w4_l8192_id6_2_1_daddr];

endmodule



module ram_w4_l8192_id6_3
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id6_3_0_addr,
  output [4-1:0] ram_w4_l8192_id6_3_0_rdata,
  input [4-1:0] ram_w4_l8192_id6_3_0_wdata,
  input ram_w4_l8192_id6_3_0_wenable,
  input [10-1:0] ram_w4_l8192_id6_3_1_addr,
  output [4-1:0] ram_w4_l8192_id6_3_1_rdata,
  input [4-1:0] ram_w4_l8192_id6_3_1_wdata,
  input ram_w4_l8192_id6_3_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id6_3_0_daddr;
  reg [10-1:0] ram_w4_l8192_id6_3_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_3_0_wenable) begin
      mem[ram_w4_l8192_id6_3_0_addr] <= ram_w4_l8192_id6_3_0_wdata;
    end 
    ram_w4_l8192_id6_3_0_daddr <= ram_w4_l8192_id6_3_0_addr;
  end

  assign ram_w4_l8192_id6_3_0_rdata = mem[ram_w4_l8192_id6_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_3_1_wenable) begin
      mem[ram_w4_l8192_id6_3_1_addr] <= ram_w4_l8192_id6_3_1_wdata;
    end 
    ram_w4_l8192_id6_3_1_daddr <= ram_w4_l8192_id6_3_1_addr;
  end

  assign ram_w4_l8192_id6_3_1_rdata = mem[ram_w4_l8192_id6_3_1_daddr];

endmodule



module ram_w4_l8192_id6_4
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id6_4_0_addr,
  output [4-1:0] ram_w4_l8192_id6_4_0_rdata,
  input [4-1:0] ram_w4_l8192_id6_4_0_wdata,
  input ram_w4_l8192_id6_4_0_wenable,
  input [10-1:0] ram_w4_l8192_id6_4_1_addr,
  output [4-1:0] ram_w4_l8192_id6_4_1_rdata,
  input [4-1:0] ram_w4_l8192_id6_4_1_wdata,
  input ram_w4_l8192_id6_4_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id6_4_0_daddr;
  reg [10-1:0] ram_w4_l8192_id6_4_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_4_0_wenable) begin
      mem[ram_w4_l8192_id6_4_0_addr] <= ram_w4_l8192_id6_4_0_wdata;
    end 
    ram_w4_l8192_id6_4_0_daddr <= ram_w4_l8192_id6_4_0_addr;
  end

  assign ram_w4_l8192_id6_4_0_rdata = mem[ram_w4_l8192_id6_4_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_4_1_wenable) begin
      mem[ram_w4_l8192_id6_4_1_addr] <= ram_w4_l8192_id6_4_1_wdata;
    end 
    ram_w4_l8192_id6_4_1_daddr <= ram_w4_l8192_id6_4_1_addr;
  end

  assign ram_w4_l8192_id6_4_1_rdata = mem[ram_w4_l8192_id6_4_1_daddr];

endmodule



module ram_w4_l8192_id6_5
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id6_5_0_addr,
  output [4-1:0] ram_w4_l8192_id6_5_0_rdata,
  input [4-1:0] ram_w4_l8192_id6_5_0_wdata,
  input ram_w4_l8192_id6_5_0_wenable,
  input [10-1:0] ram_w4_l8192_id6_5_1_addr,
  output [4-1:0] ram_w4_l8192_id6_5_1_rdata,
  input [4-1:0] ram_w4_l8192_id6_5_1_wdata,
  input ram_w4_l8192_id6_5_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id6_5_0_daddr;
  reg [10-1:0] ram_w4_l8192_id6_5_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_5_0_wenable) begin
      mem[ram_w4_l8192_id6_5_0_addr] <= ram_w4_l8192_id6_5_0_wdata;
    end 
    ram_w4_l8192_id6_5_0_daddr <= ram_w4_l8192_id6_5_0_addr;
  end

  assign ram_w4_l8192_id6_5_0_rdata = mem[ram_w4_l8192_id6_5_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_5_1_wenable) begin
      mem[ram_w4_l8192_id6_5_1_addr] <= ram_w4_l8192_id6_5_1_wdata;
    end 
    ram_w4_l8192_id6_5_1_daddr <= ram_w4_l8192_id6_5_1_addr;
  end

  assign ram_w4_l8192_id6_5_1_rdata = mem[ram_w4_l8192_id6_5_1_daddr];

endmodule



module ram_w4_l8192_id6_6
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id6_6_0_addr,
  output [4-1:0] ram_w4_l8192_id6_6_0_rdata,
  input [4-1:0] ram_w4_l8192_id6_6_0_wdata,
  input ram_w4_l8192_id6_6_0_wenable,
  input [10-1:0] ram_w4_l8192_id6_6_1_addr,
  output [4-1:0] ram_w4_l8192_id6_6_1_rdata,
  input [4-1:0] ram_w4_l8192_id6_6_1_wdata,
  input ram_w4_l8192_id6_6_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id6_6_0_daddr;
  reg [10-1:0] ram_w4_l8192_id6_6_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_6_0_wenable) begin
      mem[ram_w4_l8192_id6_6_0_addr] <= ram_w4_l8192_id6_6_0_wdata;
    end 
    ram_w4_l8192_id6_6_0_daddr <= ram_w4_l8192_id6_6_0_addr;
  end

  assign ram_w4_l8192_id6_6_0_rdata = mem[ram_w4_l8192_id6_6_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_6_1_wenable) begin
      mem[ram_w4_l8192_id6_6_1_addr] <= ram_w4_l8192_id6_6_1_wdata;
    end 
    ram_w4_l8192_id6_6_1_daddr <= ram_w4_l8192_id6_6_1_addr;
  end

  assign ram_w4_l8192_id6_6_1_rdata = mem[ram_w4_l8192_id6_6_1_daddr];

endmodule



module ram_w4_l8192_id6_7
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id6_7_0_addr,
  output [4-1:0] ram_w4_l8192_id6_7_0_rdata,
  input [4-1:0] ram_w4_l8192_id6_7_0_wdata,
  input ram_w4_l8192_id6_7_0_wenable,
  input [10-1:0] ram_w4_l8192_id6_7_1_addr,
  output [4-1:0] ram_w4_l8192_id6_7_1_rdata,
  input [4-1:0] ram_w4_l8192_id6_7_1_wdata,
  input ram_w4_l8192_id6_7_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id6_7_0_daddr;
  reg [10-1:0] ram_w4_l8192_id6_7_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_7_0_wenable) begin
      mem[ram_w4_l8192_id6_7_0_addr] <= ram_w4_l8192_id6_7_0_wdata;
    end 
    ram_w4_l8192_id6_7_0_daddr <= ram_w4_l8192_id6_7_0_addr;
  end

  assign ram_w4_l8192_id6_7_0_rdata = mem[ram_w4_l8192_id6_7_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id6_7_1_wenable) begin
      mem[ram_w4_l8192_id6_7_1_addr] <= ram_w4_l8192_id6_7_1_wdata;
    end 
    ram_w4_l8192_id6_7_1_daddr <= ram_w4_l8192_id6_7_1_addr;
  end

  assign ram_w4_l8192_id6_7_1_rdata = mem[ram_w4_l8192_id6_7_1_daddr];

endmodule



module ram_w4_l8192_id7_0
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id7_0_0_addr,
  output [4-1:0] ram_w4_l8192_id7_0_0_rdata,
  input [4-1:0] ram_w4_l8192_id7_0_0_wdata,
  input ram_w4_l8192_id7_0_0_wenable,
  input [10-1:0] ram_w4_l8192_id7_0_1_addr,
  output [4-1:0] ram_w4_l8192_id7_0_1_rdata,
  input [4-1:0] ram_w4_l8192_id7_0_1_wdata,
  input ram_w4_l8192_id7_0_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id7_0_0_daddr;
  reg [10-1:0] ram_w4_l8192_id7_0_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_0_0_wenable) begin
      mem[ram_w4_l8192_id7_0_0_addr] <= ram_w4_l8192_id7_0_0_wdata;
    end 
    ram_w4_l8192_id7_0_0_daddr <= ram_w4_l8192_id7_0_0_addr;
  end

  assign ram_w4_l8192_id7_0_0_rdata = mem[ram_w4_l8192_id7_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_0_1_wenable) begin
      mem[ram_w4_l8192_id7_0_1_addr] <= ram_w4_l8192_id7_0_1_wdata;
    end 
    ram_w4_l8192_id7_0_1_daddr <= ram_w4_l8192_id7_0_1_addr;
  end

  assign ram_w4_l8192_id7_0_1_rdata = mem[ram_w4_l8192_id7_0_1_daddr];

endmodule



module ram_w4_l8192_id7_1
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id7_1_0_addr,
  output [4-1:0] ram_w4_l8192_id7_1_0_rdata,
  input [4-1:0] ram_w4_l8192_id7_1_0_wdata,
  input ram_w4_l8192_id7_1_0_wenable,
  input [10-1:0] ram_w4_l8192_id7_1_1_addr,
  output [4-1:0] ram_w4_l8192_id7_1_1_rdata,
  input [4-1:0] ram_w4_l8192_id7_1_1_wdata,
  input ram_w4_l8192_id7_1_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id7_1_0_daddr;
  reg [10-1:0] ram_w4_l8192_id7_1_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_1_0_wenable) begin
      mem[ram_w4_l8192_id7_1_0_addr] <= ram_w4_l8192_id7_1_0_wdata;
    end 
    ram_w4_l8192_id7_1_0_daddr <= ram_w4_l8192_id7_1_0_addr;
  end

  assign ram_w4_l8192_id7_1_0_rdata = mem[ram_w4_l8192_id7_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_1_1_wenable) begin
      mem[ram_w4_l8192_id7_1_1_addr] <= ram_w4_l8192_id7_1_1_wdata;
    end 
    ram_w4_l8192_id7_1_1_daddr <= ram_w4_l8192_id7_1_1_addr;
  end

  assign ram_w4_l8192_id7_1_1_rdata = mem[ram_w4_l8192_id7_1_1_daddr];

endmodule



module ram_w4_l8192_id7_2
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id7_2_0_addr,
  output [4-1:0] ram_w4_l8192_id7_2_0_rdata,
  input [4-1:0] ram_w4_l8192_id7_2_0_wdata,
  input ram_w4_l8192_id7_2_0_wenable,
  input [10-1:0] ram_w4_l8192_id7_2_1_addr,
  output [4-1:0] ram_w4_l8192_id7_2_1_rdata,
  input [4-1:0] ram_w4_l8192_id7_2_1_wdata,
  input ram_w4_l8192_id7_2_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id7_2_0_daddr;
  reg [10-1:0] ram_w4_l8192_id7_2_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_2_0_wenable) begin
      mem[ram_w4_l8192_id7_2_0_addr] <= ram_w4_l8192_id7_2_0_wdata;
    end 
    ram_w4_l8192_id7_2_0_daddr <= ram_w4_l8192_id7_2_0_addr;
  end

  assign ram_w4_l8192_id7_2_0_rdata = mem[ram_w4_l8192_id7_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_2_1_wenable) begin
      mem[ram_w4_l8192_id7_2_1_addr] <= ram_w4_l8192_id7_2_1_wdata;
    end 
    ram_w4_l8192_id7_2_1_daddr <= ram_w4_l8192_id7_2_1_addr;
  end

  assign ram_w4_l8192_id7_2_1_rdata = mem[ram_w4_l8192_id7_2_1_daddr];

endmodule



module ram_w4_l8192_id7_3
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id7_3_0_addr,
  output [4-1:0] ram_w4_l8192_id7_3_0_rdata,
  input [4-1:0] ram_w4_l8192_id7_3_0_wdata,
  input ram_w4_l8192_id7_3_0_wenable,
  input [10-1:0] ram_w4_l8192_id7_3_1_addr,
  output [4-1:0] ram_w4_l8192_id7_3_1_rdata,
  input [4-1:0] ram_w4_l8192_id7_3_1_wdata,
  input ram_w4_l8192_id7_3_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id7_3_0_daddr;
  reg [10-1:0] ram_w4_l8192_id7_3_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_3_0_wenable) begin
      mem[ram_w4_l8192_id7_3_0_addr] <= ram_w4_l8192_id7_3_0_wdata;
    end 
    ram_w4_l8192_id7_3_0_daddr <= ram_w4_l8192_id7_3_0_addr;
  end

  assign ram_w4_l8192_id7_3_0_rdata = mem[ram_w4_l8192_id7_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_3_1_wenable) begin
      mem[ram_w4_l8192_id7_3_1_addr] <= ram_w4_l8192_id7_3_1_wdata;
    end 
    ram_w4_l8192_id7_3_1_daddr <= ram_w4_l8192_id7_3_1_addr;
  end

  assign ram_w4_l8192_id7_3_1_rdata = mem[ram_w4_l8192_id7_3_1_daddr];

endmodule



module ram_w4_l8192_id7_4
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id7_4_0_addr,
  output [4-1:0] ram_w4_l8192_id7_4_0_rdata,
  input [4-1:0] ram_w4_l8192_id7_4_0_wdata,
  input ram_w4_l8192_id7_4_0_wenable,
  input [10-1:0] ram_w4_l8192_id7_4_1_addr,
  output [4-1:0] ram_w4_l8192_id7_4_1_rdata,
  input [4-1:0] ram_w4_l8192_id7_4_1_wdata,
  input ram_w4_l8192_id7_4_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id7_4_0_daddr;
  reg [10-1:0] ram_w4_l8192_id7_4_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_4_0_wenable) begin
      mem[ram_w4_l8192_id7_4_0_addr] <= ram_w4_l8192_id7_4_0_wdata;
    end 
    ram_w4_l8192_id7_4_0_daddr <= ram_w4_l8192_id7_4_0_addr;
  end

  assign ram_w4_l8192_id7_4_0_rdata = mem[ram_w4_l8192_id7_4_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_4_1_wenable) begin
      mem[ram_w4_l8192_id7_4_1_addr] <= ram_w4_l8192_id7_4_1_wdata;
    end 
    ram_w4_l8192_id7_4_1_daddr <= ram_w4_l8192_id7_4_1_addr;
  end

  assign ram_w4_l8192_id7_4_1_rdata = mem[ram_w4_l8192_id7_4_1_daddr];

endmodule



module ram_w4_l8192_id7_5
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id7_5_0_addr,
  output [4-1:0] ram_w4_l8192_id7_5_0_rdata,
  input [4-1:0] ram_w4_l8192_id7_5_0_wdata,
  input ram_w4_l8192_id7_5_0_wenable,
  input [10-1:0] ram_w4_l8192_id7_5_1_addr,
  output [4-1:0] ram_w4_l8192_id7_5_1_rdata,
  input [4-1:0] ram_w4_l8192_id7_5_1_wdata,
  input ram_w4_l8192_id7_5_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id7_5_0_daddr;
  reg [10-1:0] ram_w4_l8192_id7_5_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_5_0_wenable) begin
      mem[ram_w4_l8192_id7_5_0_addr] <= ram_w4_l8192_id7_5_0_wdata;
    end 
    ram_w4_l8192_id7_5_0_daddr <= ram_w4_l8192_id7_5_0_addr;
  end

  assign ram_w4_l8192_id7_5_0_rdata = mem[ram_w4_l8192_id7_5_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_5_1_wenable) begin
      mem[ram_w4_l8192_id7_5_1_addr] <= ram_w4_l8192_id7_5_1_wdata;
    end 
    ram_w4_l8192_id7_5_1_daddr <= ram_w4_l8192_id7_5_1_addr;
  end

  assign ram_w4_l8192_id7_5_1_rdata = mem[ram_w4_l8192_id7_5_1_daddr];

endmodule



module ram_w4_l8192_id7_6
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id7_6_0_addr,
  output [4-1:0] ram_w4_l8192_id7_6_0_rdata,
  input [4-1:0] ram_w4_l8192_id7_6_0_wdata,
  input ram_w4_l8192_id7_6_0_wenable,
  input [10-1:0] ram_w4_l8192_id7_6_1_addr,
  output [4-1:0] ram_w4_l8192_id7_6_1_rdata,
  input [4-1:0] ram_w4_l8192_id7_6_1_wdata,
  input ram_w4_l8192_id7_6_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id7_6_0_daddr;
  reg [10-1:0] ram_w4_l8192_id7_6_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_6_0_wenable) begin
      mem[ram_w4_l8192_id7_6_0_addr] <= ram_w4_l8192_id7_6_0_wdata;
    end 
    ram_w4_l8192_id7_6_0_daddr <= ram_w4_l8192_id7_6_0_addr;
  end

  assign ram_w4_l8192_id7_6_0_rdata = mem[ram_w4_l8192_id7_6_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_6_1_wenable) begin
      mem[ram_w4_l8192_id7_6_1_addr] <= ram_w4_l8192_id7_6_1_wdata;
    end 
    ram_w4_l8192_id7_6_1_daddr <= ram_w4_l8192_id7_6_1_addr;
  end

  assign ram_w4_l8192_id7_6_1_rdata = mem[ram_w4_l8192_id7_6_1_daddr];

endmodule



module ram_w4_l8192_id7_7
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id7_7_0_addr,
  output [4-1:0] ram_w4_l8192_id7_7_0_rdata,
  input [4-1:0] ram_w4_l8192_id7_7_0_wdata,
  input ram_w4_l8192_id7_7_0_wenable,
  input [10-1:0] ram_w4_l8192_id7_7_1_addr,
  output [4-1:0] ram_w4_l8192_id7_7_1_rdata,
  input [4-1:0] ram_w4_l8192_id7_7_1_wdata,
  input ram_w4_l8192_id7_7_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id7_7_0_daddr;
  reg [10-1:0] ram_w4_l8192_id7_7_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_7_0_wenable) begin
      mem[ram_w4_l8192_id7_7_0_addr] <= ram_w4_l8192_id7_7_0_wdata;
    end 
    ram_w4_l8192_id7_7_0_daddr <= ram_w4_l8192_id7_7_0_addr;
  end

  assign ram_w4_l8192_id7_7_0_rdata = mem[ram_w4_l8192_id7_7_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id7_7_1_wenable) begin
      mem[ram_w4_l8192_id7_7_1_addr] <= ram_w4_l8192_id7_7_1_wdata;
    end 
    ram_w4_l8192_id7_7_1_daddr <= ram_w4_l8192_id7_7_1_addr;
  end

  assign ram_w4_l8192_id7_7_1_rdata = mem[ram_w4_l8192_id7_7_1_daddr];

endmodule



module ram_w4_l8192_id8_0
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id8_0_0_addr,
  output [4-1:0] ram_w4_l8192_id8_0_0_rdata,
  input [4-1:0] ram_w4_l8192_id8_0_0_wdata,
  input ram_w4_l8192_id8_0_0_wenable,
  input [10-1:0] ram_w4_l8192_id8_0_1_addr,
  output [4-1:0] ram_w4_l8192_id8_0_1_rdata,
  input [4-1:0] ram_w4_l8192_id8_0_1_wdata,
  input ram_w4_l8192_id8_0_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id8_0_0_daddr;
  reg [10-1:0] ram_w4_l8192_id8_0_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_0_0_wenable) begin
      mem[ram_w4_l8192_id8_0_0_addr] <= ram_w4_l8192_id8_0_0_wdata;
    end 
    ram_w4_l8192_id8_0_0_daddr <= ram_w4_l8192_id8_0_0_addr;
  end

  assign ram_w4_l8192_id8_0_0_rdata = mem[ram_w4_l8192_id8_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_0_1_wenable) begin
      mem[ram_w4_l8192_id8_0_1_addr] <= ram_w4_l8192_id8_0_1_wdata;
    end 
    ram_w4_l8192_id8_0_1_daddr <= ram_w4_l8192_id8_0_1_addr;
  end

  assign ram_w4_l8192_id8_0_1_rdata = mem[ram_w4_l8192_id8_0_1_daddr];

endmodule



module ram_w4_l8192_id8_1
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id8_1_0_addr,
  output [4-1:0] ram_w4_l8192_id8_1_0_rdata,
  input [4-1:0] ram_w4_l8192_id8_1_0_wdata,
  input ram_w4_l8192_id8_1_0_wenable,
  input [10-1:0] ram_w4_l8192_id8_1_1_addr,
  output [4-1:0] ram_w4_l8192_id8_1_1_rdata,
  input [4-1:0] ram_w4_l8192_id8_1_1_wdata,
  input ram_w4_l8192_id8_1_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id8_1_0_daddr;
  reg [10-1:0] ram_w4_l8192_id8_1_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_1_0_wenable) begin
      mem[ram_w4_l8192_id8_1_0_addr] <= ram_w4_l8192_id8_1_0_wdata;
    end 
    ram_w4_l8192_id8_1_0_daddr <= ram_w4_l8192_id8_1_0_addr;
  end

  assign ram_w4_l8192_id8_1_0_rdata = mem[ram_w4_l8192_id8_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_1_1_wenable) begin
      mem[ram_w4_l8192_id8_1_1_addr] <= ram_w4_l8192_id8_1_1_wdata;
    end 
    ram_w4_l8192_id8_1_1_daddr <= ram_w4_l8192_id8_1_1_addr;
  end

  assign ram_w4_l8192_id8_1_1_rdata = mem[ram_w4_l8192_id8_1_1_daddr];

endmodule



module ram_w4_l8192_id8_2
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id8_2_0_addr,
  output [4-1:0] ram_w4_l8192_id8_2_0_rdata,
  input [4-1:0] ram_w4_l8192_id8_2_0_wdata,
  input ram_w4_l8192_id8_2_0_wenable,
  input [10-1:0] ram_w4_l8192_id8_2_1_addr,
  output [4-1:0] ram_w4_l8192_id8_2_1_rdata,
  input [4-1:0] ram_w4_l8192_id8_2_1_wdata,
  input ram_w4_l8192_id8_2_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id8_2_0_daddr;
  reg [10-1:0] ram_w4_l8192_id8_2_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_2_0_wenable) begin
      mem[ram_w4_l8192_id8_2_0_addr] <= ram_w4_l8192_id8_2_0_wdata;
    end 
    ram_w4_l8192_id8_2_0_daddr <= ram_w4_l8192_id8_2_0_addr;
  end

  assign ram_w4_l8192_id8_2_0_rdata = mem[ram_w4_l8192_id8_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_2_1_wenable) begin
      mem[ram_w4_l8192_id8_2_1_addr] <= ram_w4_l8192_id8_2_1_wdata;
    end 
    ram_w4_l8192_id8_2_1_daddr <= ram_w4_l8192_id8_2_1_addr;
  end

  assign ram_w4_l8192_id8_2_1_rdata = mem[ram_w4_l8192_id8_2_1_daddr];

endmodule



module ram_w4_l8192_id8_3
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id8_3_0_addr,
  output [4-1:0] ram_w4_l8192_id8_3_0_rdata,
  input [4-1:0] ram_w4_l8192_id8_3_0_wdata,
  input ram_w4_l8192_id8_3_0_wenable,
  input [10-1:0] ram_w4_l8192_id8_3_1_addr,
  output [4-1:0] ram_w4_l8192_id8_3_1_rdata,
  input [4-1:0] ram_w4_l8192_id8_3_1_wdata,
  input ram_w4_l8192_id8_3_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id8_3_0_daddr;
  reg [10-1:0] ram_w4_l8192_id8_3_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_3_0_wenable) begin
      mem[ram_w4_l8192_id8_3_0_addr] <= ram_w4_l8192_id8_3_0_wdata;
    end 
    ram_w4_l8192_id8_3_0_daddr <= ram_w4_l8192_id8_3_0_addr;
  end

  assign ram_w4_l8192_id8_3_0_rdata = mem[ram_w4_l8192_id8_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_3_1_wenable) begin
      mem[ram_w4_l8192_id8_3_1_addr] <= ram_w4_l8192_id8_3_1_wdata;
    end 
    ram_w4_l8192_id8_3_1_daddr <= ram_w4_l8192_id8_3_1_addr;
  end

  assign ram_w4_l8192_id8_3_1_rdata = mem[ram_w4_l8192_id8_3_1_daddr];

endmodule



module ram_w4_l8192_id8_4
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id8_4_0_addr,
  output [4-1:0] ram_w4_l8192_id8_4_0_rdata,
  input [4-1:0] ram_w4_l8192_id8_4_0_wdata,
  input ram_w4_l8192_id8_4_0_wenable,
  input [10-1:0] ram_w4_l8192_id8_4_1_addr,
  output [4-1:0] ram_w4_l8192_id8_4_1_rdata,
  input [4-1:0] ram_w4_l8192_id8_4_1_wdata,
  input ram_w4_l8192_id8_4_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id8_4_0_daddr;
  reg [10-1:0] ram_w4_l8192_id8_4_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_4_0_wenable) begin
      mem[ram_w4_l8192_id8_4_0_addr] <= ram_w4_l8192_id8_4_0_wdata;
    end 
    ram_w4_l8192_id8_4_0_daddr <= ram_w4_l8192_id8_4_0_addr;
  end

  assign ram_w4_l8192_id8_4_0_rdata = mem[ram_w4_l8192_id8_4_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_4_1_wenable) begin
      mem[ram_w4_l8192_id8_4_1_addr] <= ram_w4_l8192_id8_4_1_wdata;
    end 
    ram_w4_l8192_id8_4_1_daddr <= ram_w4_l8192_id8_4_1_addr;
  end

  assign ram_w4_l8192_id8_4_1_rdata = mem[ram_w4_l8192_id8_4_1_daddr];

endmodule



module ram_w4_l8192_id8_5
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id8_5_0_addr,
  output [4-1:0] ram_w4_l8192_id8_5_0_rdata,
  input [4-1:0] ram_w4_l8192_id8_5_0_wdata,
  input ram_w4_l8192_id8_5_0_wenable,
  input [10-1:0] ram_w4_l8192_id8_5_1_addr,
  output [4-1:0] ram_w4_l8192_id8_5_1_rdata,
  input [4-1:0] ram_w4_l8192_id8_5_1_wdata,
  input ram_w4_l8192_id8_5_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id8_5_0_daddr;
  reg [10-1:0] ram_w4_l8192_id8_5_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_5_0_wenable) begin
      mem[ram_w4_l8192_id8_5_0_addr] <= ram_w4_l8192_id8_5_0_wdata;
    end 
    ram_w4_l8192_id8_5_0_daddr <= ram_w4_l8192_id8_5_0_addr;
  end

  assign ram_w4_l8192_id8_5_0_rdata = mem[ram_w4_l8192_id8_5_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_5_1_wenable) begin
      mem[ram_w4_l8192_id8_5_1_addr] <= ram_w4_l8192_id8_5_1_wdata;
    end 
    ram_w4_l8192_id8_5_1_daddr <= ram_w4_l8192_id8_5_1_addr;
  end

  assign ram_w4_l8192_id8_5_1_rdata = mem[ram_w4_l8192_id8_5_1_daddr];

endmodule



module ram_w4_l8192_id8_6
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id8_6_0_addr,
  output [4-1:0] ram_w4_l8192_id8_6_0_rdata,
  input [4-1:0] ram_w4_l8192_id8_6_0_wdata,
  input ram_w4_l8192_id8_6_0_wenable,
  input [10-1:0] ram_w4_l8192_id8_6_1_addr,
  output [4-1:0] ram_w4_l8192_id8_6_1_rdata,
  input [4-1:0] ram_w4_l8192_id8_6_1_wdata,
  input ram_w4_l8192_id8_6_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id8_6_0_daddr;
  reg [10-1:0] ram_w4_l8192_id8_6_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_6_0_wenable) begin
      mem[ram_w4_l8192_id8_6_0_addr] <= ram_w4_l8192_id8_6_0_wdata;
    end 
    ram_w4_l8192_id8_6_0_daddr <= ram_w4_l8192_id8_6_0_addr;
  end

  assign ram_w4_l8192_id8_6_0_rdata = mem[ram_w4_l8192_id8_6_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_6_1_wenable) begin
      mem[ram_w4_l8192_id8_6_1_addr] <= ram_w4_l8192_id8_6_1_wdata;
    end 
    ram_w4_l8192_id8_6_1_daddr <= ram_w4_l8192_id8_6_1_addr;
  end

  assign ram_w4_l8192_id8_6_1_rdata = mem[ram_w4_l8192_id8_6_1_daddr];

endmodule



module ram_w4_l8192_id8_7
(
  input CLK,
  input [10-1:0] ram_w4_l8192_id8_7_0_addr,
  output [4-1:0] ram_w4_l8192_id8_7_0_rdata,
  input [4-1:0] ram_w4_l8192_id8_7_0_wdata,
  input ram_w4_l8192_id8_7_0_wenable,
  input [10-1:0] ram_w4_l8192_id8_7_1_addr,
  output [4-1:0] ram_w4_l8192_id8_7_1_rdata,
  input [4-1:0] ram_w4_l8192_id8_7_1_wdata,
  input ram_w4_l8192_id8_7_1_wenable
);

  reg [10-1:0] ram_w4_l8192_id8_7_0_daddr;
  reg [10-1:0] ram_w4_l8192_id8_7_1_daddr;
  reg [4-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_7_0_wenable) begin
      mem[ram_w4_l8192_id8_7_0_addr] <= ram_w4_l8192_id8_7_0_wdata;
    end 
    ram_w4_l8192_id8_7_0_daddr <= ram_w4_l8192_id8_7_0_addr;
  end

  assign ram_w4_l8192_id8_7_0_rdata = mem[ram_w4_l8192_id8_7_0_daddr];

  always @(posedge CLK) begin
    if(ram_w4_l8192_id8_7_1_wenable) begin
      mem[ram_w4_l8192_id8_7_1_addr] <= ram_w4_l8192_id8_7_1_wdata;
    end 
    ram_w4_l8192_id8_7_1_daddr <= ram_w4_l8192_id8_7_1_addr;
  end

  assign ram_w4_l8192_id8_7_1_rdata = mem[ram_w4_l8192_id8_7_1_daddr];

endmodule



module ram_w8_l2048_id0_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id0_0_0_addr,
  output [8-1:0] ram_w8_l2048_id0_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id0_0_0_wdata,
  input ram_w8_l2048_id0_0_0_wenable,
  input [9-1:0] ram_w8_l2048_id0_0_1_addr,
  output [8-1:0] ram_w8_l2048_id0_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id0_0_1_wdata,
  input ram_w8_l2048_id0_0_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id0_0_0_daddr;
  reg [9-1:0] ram_w8_l2048_id0_0_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_0_0_wenable) begin
      mem[ram_w8_l2048_id0_0_0_addr] <= ram_w8_l2048_id0_0_0_wdata;
    end 
    ram_w8_l2048_id0_0_0_daddr <= ram_w8_l2048_id0_0_0_addr;
  end

  assign ram_w8_l2048_id0_0_0_rdata = mem[ram_w8_l2048_id0_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_0_1_wenable) begin
      mem[ram_w8_l2048_id0_0_1_addr] <= ram_w8_l2048_id0_0_1_wdata;
    end 
    ram_w8_l2048_id0_0_1_daddr <= ram_w8_l2048_id0_0_1_addr;
  end

  assign ram_w8_l2048_id0_0_1_rdata = mem[ram_w8_l2048_id0_0_1_daddr];

endmodule



module ram_w8_l2048_id0_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id0_1_0_addr,
  output [8-1:0] ram_w8_l2048_id0_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id0_1_0_wdata,
  input ram_w8_l2048_id0_1_0_wenable,
  input [9-1:0] ram_w8_l2048_id0_1_1_addr,
  output [8-1:0] ram_w8_l2048_id0_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id0_1_1_wdata,
  input ram_w8_l2048_id0_1_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id0_1_0_daddr;
  reg [9-1:0] ram_w8_l2048_id0_1_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_1_0_wenable) begin
      mem[ram_w8_l2048_id0_1_0_addr] <= ram_w8_l2048_id0_1_0_wdata;
    end 
    ram_w8_l2048_id0_1_0_daddr <= ram_w8_l2048_id0_1_0_addr;
  end

  assign ram_w8_l2048_id0_1_0_rdata = mem[ram_w8_l2048_id0_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_1_1_wenable) begin
      mem[ram_w8_l2048_id0_1_1_addr] <= ram_w8_l2048_id0_1_1_wdata;
    end 
    ram_w8_l2048_id0_1_1_daddr <= ram_w8_l2048_id0_1_1_addr;
  end

  assign ram_w8_l2048_id0_1_1_rdata = mem[ram_w8_l2048_id0_1_1_daddr];

endmodule



module ram_w8_l2048_id0_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id0_2_0_addr,
  output [8-1:0] ram_w8_l2048_id0_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id0_2_0_wdata,
  input ram_w8_l2048_id0_2_0_wenable,
  input [9-1:0] ram_w8_l2048_id0_2_1_addr,
  output [8-1:0] ram_w8_l2048_id0_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id0_2_1_wdata,
  input ram_w8_l2048_id0_2_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id0_2_0_daddr;
  reg [9-1:0] ram_w8_l2048_id0_2_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_2_0_wenable) begin
      mem[ram_w8_l2048_id0_2_0_addr] <= ram_w8_l2048_id0_2_0_wdata;
    end 
    ram_w8_l2048_id0_2_0_daddr <= ram_w8_l2048_id0_2_0_addr;
  end

  assign ram_w8_l2048_id0_2_0_rdata = mem[ram_w8_l2048_id0_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_2_1_wenable) begin
      mem[ram_w8_l2048_id0_2_1_addr] <= ram_w8_l2048_id0_2_1_wdata;
    end 
    ram_w8_l2048_id0_2_1_daddr <= ram_w8_l2048_id0_2_1_addr;
  end

  assign ram_w8_l2048_id0_2_1_rdata = mem[ram_w8_l2048_id0_2_1_daddr];

endmodule



module ram_w8_l2048_id0_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id0_3_0_addr,
  output [8-1:0] ram_w8_l2048_id0_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id0_3_0_wdata,
  input ram_w8_l2048_id0_3_0_wenable,
  input [9-1:0] ram_w8_l2048_id0_3_1_addr,
  output [8-1:0] ram_w8_l2048_id0_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id0_3_1_wdata,
  input ram_w8_l2048_id0_3_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id0_3_0_daddr;
  reg [9-1:0] ram_w8_l2048_id0_3_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_3_0_wenable) begin
      mem[ram_w8_l2048_id0_3_0_addr] <= ram_w8_l2048_id0_3_0_wdata;
    end 
    ram_w8_l2048_id0_3_0_daddr <= ram_w8_l2048_id0_3_0_addr;
  end

  assign ram_w8_l2048_id0_3_0_rdata = mem[ram_w8_l2048_id0_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_3_1_wenable) begin
      mem[ram_w8_l2048_id0_3_1_addr] <= ram_w8_l2048_id0_3_1_wdata;
    end 
    ram_w8_l2048_id0_3_1_daddr <= ram_w8_l2048_id0_3_1_addr;
  end

  assign ram_w8_l2048_id0_3_1_rdata = mem[ram_w8_l2048_id0_3_1_daddr];

endmodule



module ram_w8_l2048_id1_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id1_0_0_addr,
  output [8-1:0] ram_w8_l2048_id1_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id1_0_0_wdata,
  input ram_w8_l2048_id1_0_0_wenable,
  input [9-1:0] ram_w8_l2048_id1_0_1_addr,
  output [8-1:0] ram_w8_l2048_id1_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id1_0_1_wdata,
  input ram_w8_l2048_id1_0_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id1_0_0_daddr;
  reg [9-1:0] ram_w8_l2048_id1_0_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_0_0_wenable) begin
      mem[ram_w8_l2048_id1_0_0_addr] <= ram_w8_l2048_id1_0_0_wdata;
    end 
    ram_w8_l2048_id1_0_0_daddr <= ram_w8_l2048_id1_0_0_addr;
  end

  assign ram_w8_l2048_id1_0_0_rdata = mem[ram_w8_l2048_id1_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_0_1_wenable) begin
      mem[ram_w8_l2048_id1_0_1_addr] <= ram_w8_l2048_id1_0_1_wdata;
    end 
    ram_w8_l2048_id1_0_1_daddr <= ram_w8_l2048_id1_0_1_addr;
  end

  assign ram_w8_l2048_id1_0_1_rdata = mem[ram_w8_l2048_id1_0_1_daddr];

endmodule



module ram_w8_l2048_id1_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id1_1_0_addr,
  output [8-1:0] ram_w8_l2048_id1_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id1_1_0_wdata,
  input ram_w8_l2048_id1_1_0_wenable,
  input [9-1:0] ram_w8_l2048_id1_1_1_addr,
  output [8-1:0] ram_w8_l2048_id1_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id1_1_1_wdata,
  input ram_w8_l2048_id1_1_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id1_1_0_daddr;
  reg [9-1:0] ram_w8_l2048_id1_1_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_1_0_wenable) begin
      mem[ram_w8_l2048_id1_1_0_addr] <= ram_w8_l2048_id1_1_0_wdata;
    end 
    ram_w8_l2048_id1_1_0_daddr <= ram_w8_l2048_id1_1_0_addr;
  end

  assign ram_w8_l2048_id1_1_0_rdata = mem[ram_w8_l2048_id1_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_1_1_wenable) begin
      mem[ram_w8_l2048_id1_1_1_addr] <= ram_w8_l2048_id1_1_1_wdata;
    end 
    ram_w8_l2048_id1_1_1_daddr <= ram_w8_l2048_id1_1_1_addr;
  end

  assign ram_w8_l2048_id1_1_1_rdata = mem[ram_w8_l2048_id1_1_1_daddr];

endmodule



module ram_w8_l2048_id1_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id1_2_0_addr,
  output [8-1:0] ram_w8_l2048_id1_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id1_2_0_wdata,
  input ram_w8_l2048_id1_2_0_wenable,
  input [9-1:0] ram_w8_l2048_id1_2_1_addr,
  output [8-1:0] ram_w8_l2048_id1_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id1_2_1_wdata,
  input ram_w8_l2048_id1_2_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id1_2_0_daddr;
  reg [9-1:0] ram_w8_l2048_id1_2_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_2_0_wenable) begin
      mem[ram_w8_l2048_id1_2_0_addr] <= ram_w8_l2048_id1_2_0_wdata;
    end 
    ram_w8_l2048_id1_2_0_daddr <= ram_w8_l2048_id1_2_0_addr;
  end

  assign ram_w8_l2048_id1_2_0_rdata = mem[ram_w8_l2048_id1_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_2_1_wenable) begin
      mem[ram_w8_l2048_id1_2_1_addr] <= ram_w8_l2048_id1_2_1_wdata;
    end 
    ram_w8_l2048_id1_2_1_daddr <= ram_w8_l2048_id1_2_1_addr;
  end

  assign ram_w8_l2048_id1_2_1_rdata = mem[ram_w8_l2048_id1_2_1_daddr];

endmodule



module ram_w8_l2048_id1_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id1_3_0_addr,
  output [8-1:0] ram_w8_l2048_id1_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id1_3_0_wdata,
  input ram_w8_l2048_id1_3_0_wenable,
  input [9-1:0] ram_w8_l2048_id1_3_1_addr,
  output [8-1:0] ram_w8_l2048_id1_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id1_3_1_wdata,
  input ram_w8_l2048_id1_3_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id1_3_0_daddr;
  reg [9-1:0] ram_w8_l2048_id1_3_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_3_0_wenable) begin
      mem[ram_w8_l2048_id1_3_0_addr] <= ram_w8_l2048_id1_3_0_wdata;
    end 
    ram_w8_l2048_id1_3_0_daddr <= ram_w8_l2048_id1_3_0_addr;
  end

  assign ram_w8_l2048_id1_3_0_rdata = mem[ram_w8_l2048_id1_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_3_1_wenable) begin
      mem[ram_w8_l2048_id1_3_1_addr] <= ram_w8_l2048_id1_3_1_wdata;
    end 
    ram_w8_l2048_id1_3_1_daddr <= ram_w8_l2048_id1_3_1_addr;
  end

  assign ram_w8_l2048_id1_3_1_rdata = mem[ram_w8_l2048_id1_3_1_daddr];

endmodule



module ram_w8_l2048_id2_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id2_0_0_addr,
  output [8-1:0] ram_w8_l2048_id2_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id2_0_0_wdata,
  input ram_w8_l2048_id2_0_0_wenable,
  input [9-1:0] ram_w8_l2048_id2_0_1_addr,
  output [8-1:0] ram_w8_l2048_id2_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id2_0_1_wdata,
  input ram_w8_l2048_id2_0_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id2_0_0_daddr;
  reg [9-1:0] ram_w8_l2048_id2_0_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id2_0_0_wenable) begin
      mem[ram_w8_l2048_id2_0_0_addr] <= ram_w8_l2048_id2_0_0_wdata;
    end 
    ram_w8_l2048_id2_0_0_daddr <= ram_w8_l2048_id2_0_0_addr;
  end

  assign ram_w8_l2048_id2_0_0_rdata = mem[ram_w8_l2048_id2_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id2_0_1_wenable) begin
      mem[ram_w8_l2048_id2_0_1_addr] <= ram_w8_l2048_id2_0_1_wdata;
    end 
    ram_w8_l2048_id2_0_1_daddr <= ram_w8_l2048_id2_0_1_addr;
  end

  assign ram_w8_l2048_id2_0_1_rdata = mem[ram_w8_l2048_id2_0_1_daddr];

endmodule



module ram_w8_l2048_id2_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id2_1_0_addr,
  output [8-1:0] ram_w8_l2048_id2_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id2_1_0_wdata,
  input ram_w8_l2048_id2_1_0_wenable,
  input [9-1:0] ram_w8_l2048_id2_1_1_addr,
  output [8-1:0] ram_w8_l2048_id2_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id2_1_1_wdata,
  input ram_w8_l2048_id2_1_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id2_1_0_daddr;
  reg [9-1:0] ram_w8_l2048_id2_1_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id2_1_0_wenable) begin
      mem[ram_w8_l2048_id2_1_0_addr] <= ram_w8_l2048_id2_1_0_wdata;
    end 
    ram_w8_l2048_id2_1_0_daddr <= ram_w8_l2048_id2_1_0_addr;
  end

  assign ram_w8_l2048_id2_1_0_rdata = mem[ram_w8_l2048_id2_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id2_1_1_wenable) begin
      mem[ram_w8_l2048_id2_1_1_addr] <= ram_w8_l2048_id2_1_1_wdata;
    end 
    ram_w8_l2048_id2_1_1_daddr <= ram_w8_l2048_id2_1_1_addr;
  end

  assign ram_w8_l2048_id2_1_1_rdata = mem[ram_w8_l2048_id2_1_1_daddr];

endmodule



module ram_w8_l2048_id2_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id2_2_0_addr,
  output [8-1:0] ram_w8_l2048_id2_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id2_2_0_wdata,
  input ram_w8_l2048_id2_2_0_wenable,
  input [9-1:0] ram_w8_l2048_id2_2_1_addr,
  output [8-1:0] ram_w8_l2048_id2_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id2_2_1_wdata,
  input ram_w8_l2048_id2_2_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id2_2_0_daddr;
  reg [9-1:0] ram_w8_l2048_id2_2_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id2_2_0_wenable) begin
      mem[ram_w8_l2048_id2_2_0_addr] <= ram_w8_l2048_id2_2_0_wdata;
    end 
    ram_w8_l2048_id2_2_0_daddr <= ram_w8_l2048_id2_2_0_addr;
  end

  assign ram_w8_l2048_id2_2_0_rdata = mem[ram_w8_l2048_id2_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id2_2_1_wenable) begin
      mem[ram_w8_l2048_id2_2_1_addr] <= ram_w8_l2048_id2_2_1_wdata;
    end 
    ram_w8_l2048_id2_2_1_daddr <= ram_w8_l2048_id2_2_1_addr;
  end

  assign ram_w8_l2048_id2_2_1_rdata = mem[ram_w8_l2048_id2_2_1_daddr];

endmodule



module ram_w8_l2048_id2_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id2_3_0_addr,
  output [8-1:0] ram_w8_l2048_id2_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id2_3_0_wdata,
  input ram_w8_l2048_id2_3_0_wenable,
  input [9-1:0] ram_w8_l2048_id2_3_1_addr,
  output [8-1:0] ram_w8_l2048_id2_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id2_3_1_wdata,
  input ram_w8_l2048_id2_3_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id2_3_0_daddr;
  reg [9-1:0] ram_w8_l2048_id2_3_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id2_3_0_wenable) begin
      mem[ram_w8_l2048_id2_3_0_addr] <= ram_w8_l2048_id2_3_0_wdata;
    end 
    ram_w8_l2048_id2_3_0_daddr <= ram_w8_l2048_id2_3_0_addr;
  end

  assign ram_w8_l2048_id2_3_0_rdata = mem[ram_w8_l2048_id2_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id2_3_1_wenable) begin
      mem[ram_w8_l2048_id2_3_1_addr] <= ram_w8_l2048_id2_3_1_wdata;
    end 
    ram_w8_l2048_id2_3_1_daddr <= ram_w8_l2048_id2_3_1_addr;
  end

  assign ram_w8_l2048_id2_3_1_rdata = mem[ram_w8_l2048_id2_3_1_daddr];

endmodule



module ram_w8_l2048_id3_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id3_0_0_addr,
  output [8-1:0] ram_w8_l2048_id3_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id3_0_0_wdata,
  input ram_w8_l2048_id3_0_0_wenable,
  input [9-1:0] ram_w8_l2048_id3_0_1_addr,
  output [8-1:0] ram_w8_l2048_id3_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id3_0_1_wdata,
  input ram_w8_l2048_id3_0_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id3_0_0_daddr;
  reg [9-1:0] ram_w8_l2048_id3_0_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id3_0_0_wenable) begin
      mem[ram_w8_l2048_id3_0_0_addr] <= ram_w8_l2048_id3_0_0_wdata;
    end 
    ram_w8_l2048_id3_0_0_daddr <= ram_w8_l2048_id3_0_0_addr;
  end

  assign ram_w8_l2048_id3_0_0_rdata = mem[ram_w8_l2048_id3_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id3_0_1_wenable) begin
      mem[ram_w8_l2048_id3_0_1_addr] <= ram_w8_l2048_id3_0_1_wdata;
    end 
    ram_w8_l2048_id3_0_1_daddr <= ram_w8_l2048_id3_0_1_addr;
  end

  assign ram_w8_l2048_id3_0_1_rdata = mem[ram_w8_l2048_id3_0_1_daddr];

endmodule



module ram_w8_l2048_id3_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id3_1_0_addr,
  output [8-1:0] ram_w8_l2048_id3_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id3_1_0_wdata,
  input ram_w8_l2048_id3_1_0_wenable,
  input [9-1:0] ram_w8_l2048_id3_1_1_addr,
  output [8-1:0] ram_w8_l2048_id3_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id3_1_1_wdata,
  input ram_w8_l2048_id3_1_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id3_1_0_daddr;
  reg [9-1:0] ram_w8_l2048_id3_1_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id3_1_0_wenable) begin
      mem[ram_w8_l2048_id3_1_0_addr] <= ram_w8_l2048_id3_1_0_wdata;
    end 
    ram_w8_l2048_id3_1_0_daddr <= ram_w8_l2048_id3_1_0_addr;
  end

  assign ram_w8_l2048_id3_1_0_rdata = mem[ram_w8_l2048_id3_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id3_1_1_wenable) begin
      mem[ram_w8_l2048_id3_1_1_addr] <= ram_w8_l2048_id3_1_1_wdata;
    end 
    ram_w8_l2048_id3_1_1_daddr <= ram_w8_l2048_id3_1_1_addr;
  end

  assign ram_w8_l2048_id3_1_1_rdata = mem[ram_w8_l2048_id3_1_1_daddr];

endmodule



module ram_w8_l2048_id3_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id3_2_0_addr,
  output [8-1:0] ram_w8_l2048_id3_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id3_2_0_wdata,
  input ram_w8_l2048_id3_2_0_wenable,
  input [9-1:0] ram_w8_l2048_id3_2_1_addr,
  output [8-1:0] ram_w8_l2048_id3_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id3_2_1_wdata,
  input ram_w8_l2048_id3_2_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id3_2_0_daddr;
  reg [9-1:0] ram_w8_l2048_id3_2_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id3_2_0_wenable) begin
      mem[ram_w8_l2048_id3_2_0_addr] <= ram_w8_l2048_id3_2_0_wdata;
    end 
    ram_w8_l2048_id3_2_0_daddr <= ram_w8_l2048_id3_2_0_addr;
  end

  assign ram_w8_l2048_id3_2_0_rdata = mem[ram_w8_l2048_id3_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id3_2_1_wenable) begin
      mem[ram_w8_l2048_id3_2_1_addr] <= ram_w8_l2048_id3_2_1_wdata;
    end 
    ram_w8_l2048_id3_2_1_daddr <= ram_w8_l2048_id3_2_1_addr;
  end

  assign ram_w8_l2048_id3_2_1_rdata = mem[ram_w8_l2048_id3_2_1_daddr];

endmodule



module ram_w8_l2048_id3_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id3_3_0_addr,
  output [8-1:0] ram_w8_l2048_id3_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id3_3_0_wdata,
  input ram_w8_l2048_id3_3_0_wenable,
  input [9-1:0] ram_w8_l2048_id3_3_1_addr,
  output [8-1:0] ram_w8_l2048_id3_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id3_3_1_wdata,
  input ram_w8_l2048_id3_3_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id3_3_0_daddr;
  reg [9-1:0] ram_w8_l2048_id3_3_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id3_3_0_wenable) begin
      mem[ram_w8_l2048_id3_3_0_addr] <= ram_w8_l2048_id3_3_0_wdata;
    end 
    ram_w8_l2048_id3_3_0_daddr <= ram_w8_l2048_id3_3_0_addr;
  end

  assign ram_w8_l2048_id3_3_0_rdata = mem[ram_w8_l2048_id3_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id3_3_1_wenable) begin
      mem[ram_w8_l2048_id3_3_1_addr] <= ram_w8_l2048_id3_3_1_wdata;
    end 
    ram_w8_l2048_id3_3_1_daddr <= ram_w8_l2048_id3_3_1_addr;
  end

  assign ram_w8_l2048_id3_3_1_rdata = mem[ram_w8_l2048_id3_3_1_daddr];

endmodule



module ram_w8_l2048_id4_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id4_0_0_addr,
  output [8-1:0] ram_w8_l2048_id4_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id4_0_0_wdata,
  input ram_w8_l2048_id4_0_0_wenable,
  input [9-1:0] ram_w8_l2048_id4_0_1_addr,
  output [8-1:0] ram_w8_l2048_id4_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id4_0_1_wdata,
  input ram_w8_l2048_id4_0_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id4_0_0_daddr;
  reg [9-1:0] ram_w8_l2048_id4_0_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id4_0_0_wenable) begin
      mem[ram_w8_l2048_id4_0_0_addr] <= ram_w8_l2048_id4_0_0_wdata;
    end 
    ram_w8_l2048_id4_0_0_daddr <= ram_w8_l2048_id4_0_0_addr;
  end

  assign ram_w8_l2048_id4_0_0_rdata = mem[ram_w8_l2048_id4_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id4_0_1_wenable) begin
      mem[ram_w8_l2048_id4_0_1_addr] <= ram_w8_l2048_id4_0_1_wdata;
    end 
    ram_w8_l2048_id4_0_1_daddr <= ram_w8_l2048_id4_0_1_addr;
  end

  assign ram_w8_l2048_id4_0_1_rdata = mem[ram_w8_l2048_id4_0_1_daddr];

endmodule



module ram_w8_l2048_id4_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id4_1_0_addr,
  output [8-1:0] ram_w8_l2048_id4_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id4_1_0_wdata,
  input ram_w8_l2048_id4_1_0_wenable,
  input [9-1:0] ram_w8_l2048_id4_1_1_addr,
  output [8-1:0] ram_w8_l2048_id4_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id4_1_1_wdata,
  input ram_w8_l2048_id4_1_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id4_1_0_daddr;
  reg [9-1:0] ram_w8_l2048_id4_1_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id4_1_0_wenable) begin
      mem[ram_w8_l2048_id4_1_0_addr] <= ram_w8_l2048_id4_1_0_wdata;
    end 
    ram_w8_l2048_id4_1_0_daddr <= ram_w8_l2048_id4_1_0_addr;
  end

  assign ram_w8_l2048_id4_1_0_rdata = mem[ram_w8_l2048_id4_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id4_1_1_wenable) begin
      mem[ram_w8_l2048_id4_1_1_addr] <= ram_w8_l2048_id4_1_1_wdata;
    end 
    ram_w8_l2048_id4_1_1_daddr <= ram_w8_l2048_id4_1_1_addr;
  end

  assign ram_w8_l2048_id4_1_1_rdata = mem[ram_w8_l2048_id4_1_1_daddr];

endmodule



module ram_w8_l2048_id4_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id4_2_0_addr,
  output [8-1:0] ram_w8_l2048_id4_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id4_2_0_wdata,
  input ram_w8_l2048_id4_2_0_wenable,
  input [9-1:0] ram_w8_l2048_id4_2_1_addr,
  output [8-1:0] ram_w8_l2048_id4_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id4_2_1_wdata,
  input ram_w8_l2048_id4_2_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id4_2_0_daddr;
  reg [9-1:0] ram_w8_l2048_id4_2_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id4_2_0_wenable) begin
      mem[ram_w8_l2048_id4_2_0_addr] <= ram_w8_l2048_id4_2_0_wdata;
    end 
    ram_w8_l2048_id4_2_0_daddr <= ram_w8_l2048_id4_2_0_addr;
  end

  assign ram_w8_l2048_id4_2_0_rdata = mem[ram_w8_l2048_id4_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id4_2_1_wenable) begin
      mem[ram_w8_l2048_id4_2_1_addr] <= ram_w8_l2048_id4_2_1_wdata;
    end 
    ram_w8_l2048_id4_2_1_daddr <= ram_w8_l2048_id4_2_1_addr;
  end

  assign ram_w8_l2048_id4_2_1_rdata = mem[ram_w8_l2048_id4_2_1_daddr];

endmodule



module ram_w8_l2048_id4_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id4_3_0_addr,
  output [8-1:0] ram_w8_l2048_id4_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id4_3_0_wdata,
  input ram_w8_l2048_id4_3_0_wenable,
  input [9-1:0] ram_w8_l2048_id4_3_1_addr,
  output [8-1:0] ram_w8_l2048_id4_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id4_3_1_wdata,
  input ram_w8_l2048_id4_3_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id4_3_0_daddr;
  reg [9-1:0] ram_w8_l2048_id4_3_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id4_3_0_wenable) begin
      mem[ram_w8_l2048_id4_3_0_addr] <= ram_w8_l2048_id4_3_0_wdata;
    end 
    ram_w8_l2048_id4_3_0_daddr <= ram_w8_l2048_id4_3_0_addr;
  end

  assign ram_w8_l2048_id4_3_0_rdata = mem[ram_w8_l2048_id4_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id4_3_1_wenable) begin
      mem[ram_w8_l2048_id4_3_1_addr] <= ram_w8_l2048_id4_3_1_wdata;
    end 
    ram_w8_l2048_id4_3_1_daddr <= ram_w8_l2048_id4_3_1_addr;
  end

  assign ram_w8_l2048_id4_3_1_rdata = mem[ram_w8_l2048_id4_3_1_daddr];

endmodule



module ram_w8_l2048_id5_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id5_0_0_addr,
  output [8-1:0] ram_w8_l2048_id5_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id5_0_0_wdata,
  input ram_w8_l2048_id5_0_0_wenable,
  input [9-1:0] ram_w8_l2048_id5_0_1_addr,
  output [8-1:0] ram_w8_l2048_id5_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id5_0_1_wdata,
  input ram_w8_l2048_id5_0_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id5_0_0_daddr;
  reg [9-1:0] ram_w8_l2048_id5_0_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id5_0_0_wenable) begin
      mem[ram_w8_l2048_id5_0_0_addr] <= ram_w8_l2048_id5_0_0_wdata;
    end 
    ram_w8_l2048_id5_0_0_daddr <= ram_w8_l2048_id5_0_0_addr;
  end

  assign ram_w8_l2048_id5_0_0_rdata = mem[ram_w8_l2048_id5_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id5_0_1_wenable) begin
      mem[ram_w8_l2048_id5_0_1_addr] <= ram_w8_l2048_id5_0_1_wdata;
    end 
    ram_w8_l2048_id5_0_1_daddr <= ram_w8_l2048_id5_0_1_addr;
  end

  assign ram_w8_l2048_id5_0_1_rdata = mem[ram_w8_l2048_id5_0_1_daddr];

endmodule



module ram_w8_l2048_id5_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id5_1_0_addr,
  output [8-1:0] ram_w8_l2048_id5_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id5_1_0_wdata,
  input ram_w8_l2048_id5_1_0_wenable,
  input [9-1:0] ram_w8_l2048_id5_1_1_addr,
  output [8-1:0] ram_w8_l2048_id5_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id5_1_1_wdata,
  input ram_w8_l2048_id5_1_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id5_1_0_daddr;
  reg [9-1:0] ram_w8_l2048_id5_1_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id5_1_0_wenable) begin
      mem[ram_w8_l2048_id5_1_0_addr] <= ram_w8_l2048_id5_1_0_wdata;
    end 
    ram_w8_l2048_id5_1_0_daddr <= ram_w8_l2048_id5_1_0_addr;
  end

  assign ram_w8_l2048_id5_1_0_rdata = mem[ram_w8_l2048_id5_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id5_1_1_wenable) begin
      mem[ram_w8_l2048_id5_1_1_addr] <= ram_w8_l2048_id5_1_1_wdata;
    end 
    ram_w8_l2048_id5_1_1_daddr <= ram_w8_l2048_id5_1_1_addr;
  end

  assign ram_w8_l2048_id5_1_1_rdata = mem[ram_w8_l2048_id5_1_1_daddr];

endmodule



module ram_w8_l2048_id5_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id5_2_0_addr,
  output [8-1:0] ram_w8_l2048_id5_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id5_2_0_wdata,
  input ram_w8_l2048_id5_2_0_wenable,
  input [9-1:0] ram_w8_l2048_id5_2_1_addr,
  output [8-1:0] ram_w8_l2048_id5_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id5_2_1_wdata,
  input ram_w8_l2048_id5_2_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id5_2_0_daddr;
  reg [9-1:0] ram_w8_l2048_id5_2_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id5_2_0_wenable) begin
      mem[ram_w8_l2048_id5_2_0_addr] <= ram_w8_l2048_id5_2_0_wdata;
    end 
    ram_w8_l2048_id5_2_0_daddr <= ram_w8_l2048_id5_2_0_addr;
  end

  assign ram_w8_l2048_id5_2_0_rdata = mem[ram_w8_l2048_id5_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id5_2_1_wenable) begin
      mem[ram_w8_l2048_id5_2_1_addr] <= ram_w8_l2048_id5_2_1_wdata;
    end 
    ram_w8_l2048_id5_2_1_daddr <= ram_w8_l2048_id5_2_1_addr;
  end

  assign ram_w8_l2048_id5_2_1_rdata = mem[ram_w8_l2048_id5_2_1_daddr];

endmodule



module ram_w8_l2048_id5_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id5_3_0_addr,
  output [8-1:0] ram_w8_l2048_id5_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id5_3_0_wdata,
  input ram_w8_l2048_id5_3_0_wenable,
  input [9-1:0] ram_w8_l2048_id5_3_1_addr,
  output [8-1:0] ram_w8_l2048_id5_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id5_3_1_wdata,
  input ram_w8_l2048_id5_3_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id5_3_0_daddr;
  reg [9-1:0] ram_w8_l2048_id5_3_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id5_3_0_wenable) begin
      mem[ram_w8_l2048_id5_3_0_addr] <= ram_w8_l2048_id5_3_0_wdata;
    end 
    ram_w8_l2048_id5_3_0_daddr <= ram_w8_l2048_id5_3_0_addr;
  end

  assign ram_w8_l2048_id5_3_0_rdata = mem[ram_w8_l2048_id5_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id5_3_1_wenable) begin
      mem[ram_w8_l2048_id5_3_1_addr] <= ram_w8_l2048_id5_3_1_wdata;
    end 
    ram_w8_l2048_id5_3_1_daddr <= ram_w8_l2048_id5_3_1_addr;
  end

  assign ram_w8_l2048_id5_3_1_rdata = mem[ram_w8_l2048_id5_3_1_daddr];

endmodule



module ram_w8_l2048_id6_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id6_0_0_addr,
  output [8-1:0] ram_w8_l2048_id6_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id6_0_0_wdata,
  input ram_w8_l2048_id6_0_0_wenable,
  input [9-1:0] ram_w8_l2048_id6_0_1_addr,
  output [8-1:0] ram_w8_l2048_id6_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id6_0_1_wdata,
  input ram_w8_l2048_id6_0_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id6_0_0_daddr;
  reg [9-1:0] ram_w8_l2048_id6_0_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id6_0_0_wenable) begin
      mem[ram_w8_l2048_id6_0_0_addr] <= ram_w8_l2048_id6_0_0_wdata;
    end 
    ram_w8_l2048_id6_0_0_daddr <= ram_w8_l2048_id6_0_0_addr;
  end

  assign ram_w8_l2048_id6_0_0_rdata = mem[ram_w8_l2048_id6_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id6_0_1_wenable) begin
      mem[ram_w8_l2048_id6_0_1_addr] <= ram_w8_l2048_id6_0_1_wdata;
    end 
    ram_w8_l2048_id6_0_1_daddr <= ram_w8_l2048_id6_0_1_addr;
  end

  assign ram_w8_l2048_id6_0_1_rdata = mem[ram_w8_l2048_id6_0_1_daddr];

endmodule



module ram_w8_l2048_id6_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id6_1_0_addr,
  output [8-1:0] ram_w8_l2048_id6_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id6_1_0_wdata,
  input ram_w8_l2048_id6_1_0_wenable,
  input [9-1:0] ram_w8_l2048_id6_1_1_addr,
  output [8-1:0] ram_w8_l2048_id6_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id6_1_1_wdata,
  input ram_w8_l2048_id6_1_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id6_1_0_daddr;
  reg [9-1:0] ram_w8_l2048_id6_1_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id6_1_0_wenable) begin
      mem[ram_w8_l2048_id6_1_0_addr] <= ram_w8_l2048_id6_1_0_wdata;
    end 
    ram_w8_l2048_id6_1_0_daddr <= ram_w8_l2048_id6_1_0_addr;
  end

  assign ram_w8_l2048_id6_1_0_rdata = mem[ram_w8_l2048_id6_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id6_1_1_wenable) begin
      mem[ram_w8_l2048_id6_1_1_addr] <= ram_w8_l2048_id6_1_1_wdata;
    end 
    ram_w8_l2048_id6_1_1_daddr <= ram_w8_l2048_id6_1_1_addr;
  end

  assign ram_w8_l2048_id6_1_1_rdata = mem[ram_w8_l2048_id6_1_1_daddr];

endmodule



module ram_w8_l2048_id6_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id6_2_0_addr,
  output [8-1:0] ram_w8_l2048_id6_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id6_2_0_wdata,
  input ram_w8_l2048_id6_2_0_wenable,
  input [9-1:0] ram_w8_l2048_id6_2_1_addr,
  output [8-1:0] ram_w8_l2048_id6_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id6_2_1_wdata,
  input ram_w8_l2048_id6_2_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id6_2_0_daddr;
  reg [9-1:0] ram_w8_l2048_id6_2_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id6_2_0_wenable) begin
      mem[ram_w8_l2048_id6_2_0_addr] <= ram_w8_l2048_id6_2_0_wdata;
    end 
    ram_w8_l2048_id6_2_0_daddr <= ram_w8_l2048_id6_2_0_addr;
  end

  assign ram_w8_l2048_id6_2_0_rdata = mem[ram_w8_l2048_id6_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id6_2_1_wenable) begin
      mem[ram_w8_l2048_id6_2_1_addr] <= ram_w8_l2048_id6_2_1_wdata;
    end 
    ram_w8_l2048_id6_2_1_daddr <= ram_w8_l2048_id6_2_1_addr;
  end

  assign ram_w8_l2048_id6_2_1_rdata = mem[ram_w8_l2048_id6_2_1_daddr];

endmodule



module ram_w8_l2048_id6_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id6_3_0_addr,
  output [8-1:0] ram_w8_l2048_id6_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id6_3_0_wdata,
  input ram_w8_l2048_id6_3_0_wenable,
  input [9-1:0] ram_w8_l2048_id6_3_1_addr,
  output [8-1:0] ram_w8_l2048_id6_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id6_3_1_wdata,
  input ram_w8_l2048_id6_3_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id6_3_0_daddr;
  reg [9-1:0] ram_w8_l2048_id6_3_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id6_3_0_wenable) begin
      mem[ram_w8_l2048_id6_3_0_addr] <= ram_w8_l2048_id6_3_0_wdata;
    end 
    ram_w8_l2048_id6_3_0_daddr <= ram_w8_l2048_id6_3_0_addr;
  end

  assign ram_w8_l2048_id6_3_0_rdata = mem[ram_w8_l2048_id6_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id6_3_1_wenable) begin
      mem[ram_w8_l2048_id6_3_1_addr] <= ram_w8_l2048_id6_3_1_wdata;
    end 
    ram_w8_l2048_id6_3_1_daddr <= ram_w8_l2048_id6_3_1_addr;
  end

  assign ram_w8_l2048_id6_3_1_rdata = mem[ram_w8_l2048_id6_3_1_daddr];

endmodule



module ram_w8_l2048_id7_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id7_0_0_addr,
  output [8-1:0] ram_w8_l2048_id7_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id7_0_0_wdata,
  input ram_w8_l2048_id7_0_0_wenable,
  input [9-1:0] ram_w8_l2048_id7_0_1_addr,
  output [8-1:0] ram_w8_l2048_id7_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id7_0_1_wdata,
  input ram_w8_l2048_id7_0_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id7_0_0_daddr;
  reg [9-1:0] ram_w8_l2048_id7_0_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id7_0_0_wenable) begin
      mem[ram_w8_l2048_id7_0_0_addr] <= ram_w8_l2048_id7_0_0_wdata;
    end 
    ram_w8_l2048_id7_0_0_daddr <= ram_w8_l2048_id7_0_0_addr;
  end

  assign ram_w8_l2048_id7_0_0_rdata = mem[ram_w8_l2048_id7_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id7_0_1_wenable) begin
      mem[ram_w8_l2048_id7_0_1_addr] <= ram_w8_l2048_id7_0_1_wdata;
    end 
    ram_w8_l2048_id7_0_1_daddr <= ram_w8_l2048_id7_0_1_addr;
  end

  assign ram_w8_l2048_id7_0_1_rdata = mem[ram_w8_l2048_id7_0_1_daddr];

endmodule



module ram_w8_l2048_id7_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id7_1_0_addr,
  output [8-1:0] ram_w8_l2048_id7_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id7_1_0_wdata,
  input ram_w8_l2048_id7_1_0_wenable,
  input [9-1:0] ram_w8_l2048_id7_1_1_addr,
  output [8-1:0] ram_w8_l2048_id7_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id7_1_1_wdata,
  input ram_w8_l2048_id7_1_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id7_1_0_daddr;
  reg [9-1:0] ram_w8_l2048_id7_1_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id7_1_0_wenable) begin
      mem[ram_w8_l2048_id7_1_0_addr] <= ram_w8_l2048_id7_1_0_wdata;
    end 
    ram_w8_l2048_id7_1_0_daddr <= ram_w8_l2048_id7_1_0_addr;
  end

  assign ram_w8_l2048_id7_1_0_rdata = mem[ram_w8_l2048_id7_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id7_1_1_wenable) begin
      mem[ram_w8_l2048_id7_1_1_addr] <= ram_w8_l2048_id7_1_1_wdata;
    end 
    ram_w8_l2048_id7_1_1_daddr <= ram_w8_l2048_id7_1_1_addr;
  end

  assign ram_w8_l2048_id7_1_1_rdata = mem[ram_w8_l2048_id7_1_1_daddr];

endmodule



module ram_w8_l2048_id7_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id7_2_0_addr,
  output [8-1:0] ram_w8_l2048_id7_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id7_2_0_wdata,
  input ram_w8_l2048_id7_2_0_wenable,
  input [9-1:0] ram_w8_l2048_id7_2_1_addr,
  output [8-1:0] ram_w8_l2048_id7_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id7_2_1_wdata,
  input ram_w8_l2048_id7_2_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id7_2_0_daddr;
  reg [9-1:0] ram_w8_l2048_id7_2_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id7_2_0_wenable) begin
      mem[ram_w8_l2048_id7_2_0_addr] <= ram_w8_l2048_id7_2_0_wdata;
    end 
    ram_w8_l2048_id7_2_0_daddr <= ram_w8_l2048_id7_2_0_addr;
  end

  assign ram_w8_l2048_id7_2_0_rdata = mem[ram_w8_l2048_id7_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id7_2_1_wenable) begin
      mem[ram_w8_l2048_id7_2_1_addr] <= ram_w8_l2048_id7_2_1_wdata;
    end 
    ram_w8_l2048_id7_2_1_daddr <= ram_w8_l2048_id7_2_1_addr;
  end

  assign ram_w8_l2048_id7_2_1_rdata = mem[ram_w8_l2048_id7_2_1_daddr];

endmodule



module ram_w8_l2048_id7_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id7_3_0_addr,
  output [8-1:0] ram_w8_l2048_id7_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id7_3_0_wdata,
  input ram_w8_l2048_id7_3_0_wenable,
  input [9-1:0] ram_w8_l2048_id7_3_1_addr,
  output [8-1:0] ram_w8_l2048_id7_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id7_3_1_wdata,
  input ram_w8_l2048_id7_3_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id7_3_0_daddr;
  reg [9-1:0] ram_w8_l2048_id7_3_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id7_3_0_wenable) begin
      mem[ram_w8_l2048_id7_3_0_addr] <= ram_w8_l2048_id7_3_0_wdata;
    end 
    ram_w8_l2048_id7_3_0_daddr <= ram_w8_l2048_id7_3_0_addr;
  end

  assign ram_w8_l2048_id7_3_0_rdata = mem[ram_w8_l2048_id7_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id7_3_1_wenable) begin
      mem[ram_w8_l2048_id7_3_1_addr] <= ram_w8_l2048_id7_3_1_wdata;
    end 
    ram_w8_l2048_id7_3_1_daddr <= ram_w8_l2048_id7_3_1_addr;
  end

  assign ram_w8_l2048_id7_3_1_rdata = mem[ram_w8_l2048_id7_3_1_daddr];

endmodule



module ram_w8_l2048_id8_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id8_0_0_addr,
  output [8-1:0] ram_w8_l2048_id8_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id8_0_0_wdata,
  input ram_w8_l2048_id8_0_0_wenable,
  input [9-1:0] ram_w8_l2048_id8_0_1_addr,
  output [8-1:0] ram_w8_l2048_id8_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id8_0_1_wdata,
  input ram_w8_l2048_id8_0_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id8_0_0_daddr;
  reg [9-1:0] ram_w8_l2048_id8_0_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id8_0_0_wenable) begin
      mem[ram_w8_l2048_id8_0_0_addr] <= ram_w8_l2048_id8_0_0_wdata;
    end 
    ram_w8_l2048_id8_0_0_daddr <= ram_w8_l2048_id8_0_0_addr;
  end

  assign ram_w8_l2048_id8_0_0_rdata = mem[ram_w8_l2048_id8_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id8_0_1_wenable) begin
      mem[ram_w8_l2048_id8_0_1_addr] <= ram_w8_l2048_id8_0_1_wdata;
    end 
    ram_w8_l2048_id8_0_1_daddr <= ram_w8_l2048_id8_0_1_addr;
  end

  assign ram_w8_l2048_id8_0_1_rdata = mem[ram_w8_l2048_id8_0_1_daddr];

endmodule



module ram_w8_l2048_id8_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id8_1_0_addr,
  output [8-1:0] ram_w8_l2048_id8_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id8_1_0_wdata,
  input ram_w8_l2048_id8_1_0_wenable,
  input [9-1:0] ram_w8_l2048_id8_1_1_addr,
  output [8-1:0] ram_w8_l2048_id8_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id8_1_1_wdata,
  input ram_w8_l2048_id8_1_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id8_1_0_daddr;
  reg [9-1:0] ram_w8_l2048_id8_1_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id8_1_0_wenable) begin
      mem[ram_w8_l2048_id8_1_0_addr] <= ram_w8_l2048_id8_1_0_wdata;
    end 
    ram_w8_l2048_id8_1_0_daddr <= ram_w8_l2048_id8_1_0_addr;
  end

  assign ram_w8_l2048_id8_1_0_rdata = mem[ram_w8_l2048_id8_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id8_1_1_wenable) begin
      mem[ram_w8_l2048_id8_1_1_addr] <= ram_w8_l2048_id8_1_1_wdata;
    end 
    ram_w8_l2048_id8_1_1_daddr <= ram_w8_l2048_id8_1_1_addr;
  end

  assign ram_w8_l2048_id8_1_1_rdata = mem[ram_w8_l2048_id8_1_1_daddr];

endmodule



module ram_w8_l2048_id8_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id8_2_0_addr,
  output [8-1:0] ram_w8_l2048_id8_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id8_2_0_wdata,
  input ram_w8_l2048_id8_2_0_wenable,
  input [9-1:0] ram_w8_l2048_id8_2_1_addr,
  output [8-1:0] ram_w8_l2048_id8_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id8_2_1_wdata,
  input ram_w8_l2048_id8_2_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id8_2_0_daddr;
  reg [9-1:0] ram_w8_l2048_id8_2_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id8_2_0_wenable) begin
      mem[ram_w8_l2048_id8_2_0_addr] <= ram_w8_l2048_id8_2_0_wdata;
    end 
    ram_w8_l2048_id8_2_0_daddr <= ram_w8_l2048_id8_2_0_addr;
  end

  assign ram_w8_l2048_id8_2_0_rdata = mem[ram_w8_l2048_id8_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id8_2_1_wenable) begin
      mem[ram_w8_l2048_id8_2_1_addr] <= ram_w8_l2048_id8_2_1_wdata;
    end 
    ram_w8_l2048_id8_2_1_daddr <= ram_w8_l2048_id8_2_1_addr;
  end

  assign ram_w8_l2048_id8_2_1_rdata = mem[ram_w8_l2048_id8_2_1_daddr];

endmodule



module ram_w8_l2048_id8_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id8_3_0_addr,
  output [8-1:0] ram_w8_l2048_id8_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id8_3_0_wdata,
  input ram_w8_l2048_id8_3_0_wenable,
  input [9-1:0] ram_w8_l2048_id8_3_1_addr,
  output [8-1:0] ram_w8_l2048_id8_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id8_3_1_wdata,
  input ram_w8_l2048_id8_3_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id8_3_0_daddr;
  reg [9-1:0] ram_w8_l2048_id8_3_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id8_3_0_wenable) begin
      mem[ram_w8_l2048_id8_3_0_addr] <= ram_w8_l2048_id8_3_0_wdata;
    end 
    ram_w8_l2048_id8_3_0_daddr <= ram_w8_l2048_id8_3_0_addr;
  end

  assign ram_w8_l2048_id8_3_0_rdata = mem[ram_w8_l2048_id8_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id8_3_1_wenable) begin
      mem[ram_w8_l2048_id8_3_1_addr] <= ram_w8_l2048_id8_3_1_wdata;
    end 
    ram_w8_l2048_id8_3_1_daddr <= ram_w8_l2048_id8_3_1_addr;
  end

  assign ram_w8_l2048_id8_3_1_rdata = mem[ram_w8_l2048_id8_3_1_daddr];

endmodule



module ram_w8_l2048_id9_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id9_0_0_addr,
  output [8-1:0] ram_w8_l2048_id9_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id9_0_0_wdata,
  input ram_w8_l2048_id9_0_0_wenable,
  input [9-1:0] ram_w8_l2048_id9_0_1_addr,
  output [8-1:0] ram_w8_l2048_id9_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id9_0_1_wdata,
  input ram_w8_l2048_id9_0_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id9_0_0_daddr;
  reg [9-1:0] ram_w8_l2048_id9_0_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id9_0_0_wenable) begin
      mem[ram_w8_l2048_id9_0_0_addr] <= ram_w8_l2048_id9_0_0_wdata;
    end 
    ram_w8_l2048_id9_0_0_daddr <= ram_w8_l2048_id9_0_0_addr;
  end

  assign ram_w8_l2048_id9_0_0_rdata = mem[ram_w8_l2048_id9_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id9_0_1_wenable) begin
      mem[ram_w8_l2048_id9_0_1_addr] <= ram_w8_l2048_id9_0_1_wdata;
    end 
    ram_w8_l2048_id9_0_1_daddr <= ram_w8_l2048_id9_0_1_addr;
  end

  assign ram_w8_l2048_id9_0_1_rdata = mem[ram_w8_l2048_id9_0_1_daddr];

endmodule



module ram_w8_l2048_id9_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id9_1_0_addr,
  output [8-1:0] ram_w8_l2048_id9_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id9_1_0_wdata,
  input ram_w8_l2048_id9_1_0_wenable,
  input [9-1:0] ram_w8_l2048_id9_1_1_addr,
  output [8-1:0] ram_w8_l2048_id9_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id9_1_1_wdata,
  input ram_w8_l2048_id9_1_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id9_1_0_daddr;
  reg [9-1:0] ram_w8_l2048_id9_1_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id9_1_0_wenable) begin
      mem[ram_w8_l2048_id9_1_0_addr] <= ram_w8_l2048_id9_1_0_wdata;
    end 
    ram_w8_l2048_id9_1_0_daddr <= ram_w8_l2048_id9_1_0_addr;
  end

  assign ram_w8_l2048_id9_1_0_rdata = mem[ram_w8_l2048_id9_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id9_1_1_wenable) begin
      mem[ram_w8_l2048_id9_1_1_addr] <= ram_w8_l2048_id9_1_1_wdata;
    end 
    ram_w8_l2048_id9_1_1_daddr <= ram_w8_l2048_id9_1_1_addr;
  end

  assign ram_w8_l2048_id9_1_1_rdata = mem[ram_w8_l2048_id9_1_1_daddr];

endmodule



module ram_w8_l2048_id9_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id9_2_0_addr,
  output [8-1:0] ram_w8_l2048_id9_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id9_2_0_wdata,
  input ram_w8_l2048_id9_2_0_wenable,
  input [9-1:0] ram_w8_l2048_id9_2_1_addr,
  output [8-1:0] ram_w8_l2048_id9_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id9_2_1_wdata,
  input ram_w8_l2048_id9_2_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id9_2_0_daddr;
  reg [9-1:0] ram_w8_l2048_id9_2_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id9_2_0_wenable) begin
      mem[ram_w8_l2048_id9_2_0_addr] <= ram_w8_l2048_id9_2_0_wdata;
    end 
    ram_w8_l2048_id9_2_0_daddr <= ram_w8_l2048_id9_2_0_addr;
  end

  assign ram_w8_l2048_id9_2_0_rdata = mem[ram_w8_l2048_id9_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id9_2_1_wenable) begin
      mem[ram_w8_l2048_id9_2_1_addr] <= ram_w8_l2048_id9_2_1_wdata;
    end 
    ram_w8_l2048_id9_2_1_daddr <= ram_w8_l2048_id9_2_1_addr;
  end

  assign ram_w8_l2048_id9_2_1_rdata = mem[ram_w8_l2048_id9_2_1_daddr];

endmodule



module ram_w8_l2048_id9_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id9_3_0_addr,
  output [8-1:0] ram_w8_l2048_id9_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id9_3_0_wdata,
  input ram_w8_l2048_id9_3_0_wenable,
  input [9-1:0] ram_w8_l2048_id9_3_1_addr,
  output [8-1:0] ram_w8_l2048_id9_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id9_3_1_wdata,
  input ram_w8_l2048_id9_3_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id9_3_0_daddr;
  reg [9-1:0] ram_w8_l2048_id9_3_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id9_3_0_wenable) begin
      mem[ram_w8_l2048_id9_3_0_addr] <= ram_w8_l2048_id9_3_0_wdata;
    end 
    ram_w8_l2048_id9_3_0_daddr <= ram_w8_l2048_id9_3_0_addr;
  end

  assign ram_w8_l2048_id9_3_0_rdata = mem[ram_w8_l2048_id9_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id9_3_1_wenable) begin
      mem[ram_w8_l2048_id9_3_1_addr] <= ram_w8_l2048_id9_3_1_wdata;
    end 
    ram_w8_l2048_id9_3_1_daddr <= ram_w8_l2048_id9_3_1_addr;
  end

  assign ram_w8_l2048_id9_3_1_rdata = mem[ram_w8_l2048_id9_3_1_daddr];

endmodule



module ram_w8_l2048_id10_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id10_0_0_addr,
  output [8-1:0] ram_w8_l2048_id10_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id10_0_0_wdata,
  input ram_w8_l2048_id10_0_0_wenable,
  input [9-1:0] ram_w8_l2048_id10_0_1_addr,
  output [8-1:0] ram_w8_l2048_id10_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id10_0_1_wdata,
  input ram_w8_l2048_id10_0_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id10_0_0_daddr;
  reg [9-1:0] ram_w8_l2048_id10_0_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id10_0_0_wenable) begin
      mem[ram_w8_l2048_id10_0_0_addr] <= ram_w8_l2048_id10_0_0_wdata;
    end 
    ram_w8_l2048_id10_0_0_daddr <= ram_w8_l2048_id10_0_0_addr;
  end

  assign ram_w8_l2048_id10_0_0_rdata = mem[ram_w8_l2048_id10_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id10_0_1_wenable) begin
      mem[ram_w8_l2048_id10_0_1_addr] <= ram_w8_l2048_id10_0_1_wdata;
    end 
    ram_w8_l2048_id10_0_1_daddr <= ram_w8_l2048_id10_0_1_addr;
  end

  assign ram_w8_l2048_id10_0_1_rdata = mem[ram_w8_l2048_id10_0_1_daddr];

endmodule



module ram_w8_l2048_id10_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id10_1_0_addr,
  output [8-1:0] ram_w8_l2048_id10_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id10_1_0_wdata,
  input ram_w8_l2048_id10_1_0_wenable,
  input [9-1:0] ram_w8_l2048_id10_1_1_addr,
  output [8-1:0] ram_w8_l2048_id10_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id10_1_1_wdata,
  input ram_w8_l2048_id10_1_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id10_1_0_daddr;
  reg [9-1:0] ram_w8_l2048_id10_1_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id10_1_0_wenable) begin
      mem[ram_w8_l2048_id10_1_0_addr] <= ram_w8_l2048_id10_1_0_wdata;
    end 
    ram_w8_l2048_id10_1_0_daddr <= ram_w8_l2048_id10_1_0_addr;
  end

  assign ram_w8_l2048_id10_1_0_rdata = mem[ram_w8_l2048_id10_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id10_1_1_wenable) begin
      mem[ram_w8_l2048_id10_1_1_addr] <= ram_w8_l2048_id10_1_1_wdata;
    end 
    ram_w8_l2048_id10_1_1_daddr <= ram_w8_l2048_id10_1_1_addr;
  end

  assign ram_w8_l2048_id10_1_1_rdata = mem[ram_w8_l2048_id10_1_1_daddr];

endmodule



module ram_w8_l2048_id10_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id10_2_0_addr,
  output [8-1:0] ram_w8_l2048_id10_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id10_2_0_wdata,
  input ram_w8_l2048_id10_2_0_wenable,
  input [9-1:0] ram_w8_l2048_id10_2_1_addr,
  output [8-1:0] ram_w8_l2048_id10_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id10_2_1_wdata,
  input ram_w8_l2048_id10_2_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id10_2_0_daddr;
  reg [9-1:0] ram_w8_l2048_id10_2_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id10_2_0_wenable) begin
      mem[ram_w8_l2048_id10_2_0_addr] <= ram_w8_l2048_id10_2_0_wdata;
    end 
    ram_w8_l2048_id10_2_0_daddr <= ram_w8_l2048_id10_2_0_addr;
  end

  assign ram_w8_l2048_id10_2_0_rdata = mem[ram_w8_l2048_id10_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id10_2_1_wenable) begin
      mem[ram_w8_l2048_id10_2_1_addr] <= ram_w8_l2048_id10_2_1_wdata;
    end 
    ram_w8_l2048_id10_2_1_daddr <= ram_w8_l2048_id10_2_1_addr;
  end

  assign ram_w8_l2048_id10_2_1_rdata = mem[ram_w8_l2048_id10_2_1_daddr];

endmodule



module ram_w8_l2048_id10_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id10_3_0_addr,
  output [8-1:0] ram_w8_l2048_id10_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id10_3_0_wdata,
  input ram_w8_l2048_id10_3_0_wenable,
  input [9-1:0] ram_w8_l2048_id10_3_1_addr,
  output [8-1:0] ram_w8_l2048_id10_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id10_3_1_wdata,
  input ram_w8_l2048_id10_3_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id10_3_0_daddr;
  reg [9-1:0] ram_w8_l2048_id10_3_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id10_3_0_wenable) begin
      mem[ram_w8_l2048_id10_3_0_addr] <= ram_w8_l2048_id10_3_0_wdata;
    end 
    ram_w8_l2048_id10_3_0_daddr <= ram_w8_l2048_id10_3_0_addr;
  end

  assign ram_w8_l2048_id10_3_0_rdata = mem[ram_w8_l2048_id10_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id10_3_1_wenable) begin
      mem[ram_w8_l2048_id10_3_1_addr] <= ram_w8_l2048_id10_3_1_wdata;
    end 
    ram_w8_l2048_id10_3_1_daddr <= ram_w8_l2048_id10_3_1_addr;
  end

  assign ram_w8_l2048_id10_3_1_rdata = mem[ram_w8_l2048_id10_3_1_daddr];

endmodule



module ram_w8_l2048_id11_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id11_0_0_addr,
  output [8-1:0] ram_w8_l2048_id11_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id11_0_0_wdata,
  input ram_w8_l2048_id11_0_0_wenable,
  input [9-1:0] ram_w8_l2048_id11_0_1_addr,
  output [8-1:0] ram_w8_l2048_id11_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id11_0_1_wdata,
  input ram_w8_l2048_id11_0_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id11_0_0_daddr;
  reg [9-1:0] ram_w8_l2048_id11_0_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id11_0_0_wenable) begin
      mem[ram_w8_l2048_id11_0_0_addr] <= ram_w8_l2048_id11_0_0_wdata;
    end 
    ram_w8_l2048_id11_0_0_daddr <= ram_w8_l2048_id11_0_0_addr;
  end

  assign ram_w8_l2048_id11_0_0_rdata = mem[ram_w8_l2048_id11_0_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id11_0_1_wenable) begin
      mem[ram_w8_l2048_id11_0_1_addr] <= ram_w8_l2048_id11_0_1_wdata;
    end 
    ram_w8_l2048_id11_0_1_daddr <= ram_w8_l2048_id11_0_1_addr;
  end

  assign ram_w8_l2048_id11_0_1_rdata = mem[ram_w8_l2048_id11_0_1_daddr];

endmodule



module ram_w8_l2048_id11_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id11_1_0_addr,
  output [8-1:0] ram_w8_l2048_id11_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id11_1_0_wdata,
  input ram_w8_l2048_id11_1_0_wenable,
  input [9-1:0] ram_w8_l2048_id11_1_1_addr,
  output [8-1:0] ram_w8_l2048_id11_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id11_1_1_wdata,
  input ram_w8_l2048_id11_1_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id11_1_0_daddr;
  reg [9-1:0] ram_w8_l2048_id11_1_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id11_1_0_wenable) begin
      mem[ram_w8_l2048_id11_1_0_addr] <= ram_w8_l2048_id11_1_0_wdata;
    end 
    ram_w8_l2048_id11_1_0_daddr <= ram_w8_l2048_id11_1_0_addr;
  end

  assign ram_w8_l2048_id11_1_0_rdata = mem[ram_w8_l2048_id11_1_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id11_1_1_wenable) begin
      mem[ram_w8_l2048_id11_1_1_addr] <= ram_w8_l2048_id11_1_1_wdata;
    end 
    ram_w8_l2048_id11_1_1_daddr <= ram_w8_l2048_id11_1_1_addr;
  end

  assign ram_w8_l2048_id11_1_1_rdata = mem[ram_w8_l2048_id11_1_1_daddr];

endmodule



module ram_w8_l2048_id11_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id11_2_0_addr,
  output [8-1:0] ram_w8_l2048_id11_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id11_2_0_wdata,
  input ram_w8_l2048_id11_2_0_wenable,
  input [9-1:0] ram_w8_l2048_id11_2_1_addr,
  output [8-1:0] ram_w8_l2048_id11_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id11_2_1_wdata,
  input ram_w8_l2048_id11_2_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id11_2_0_daddr;
  reg [9-1:0] ram_w8_l2048_id11_2_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id11_2_0_wenable) begin
      mem[ram_w8_l2048_id11_2_0_addr] <= ram_w8_l2048_id11_2_0_wdata;
    end 
    ram_w8_l2048_id11_2_0_daddr <= ram_w8_l2048_id11_2_0_addr;
  end

  assign ram_w8_l2048_id11_2_0_rdata = mem[ram_w8_l2048_id11_2_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id11_2_1_wenable) begin
      mem[ram_w8_l2048_id11_2_1_addr] <= ram_w8_l2048_id11_2_1_wdata;
    end 
    ram_w8_l2048_id11_2_1_daddr <= ram_w8_l2048_id11_2_1_addr;
  end

  assign ram_w8_l2048_id11_2_1_rdata = mem[ram_w8_l2048_id11_2_1_daddr];

endmodule



module ram_w8_l2048_id11_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id11_3_0_addr,
  output [8-1:0] ram_w8_l2048_id11_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id11_3_0_wdata,
  input ram_w8_l2048_id11_3_0_wenable,
  input [9-1:0] ram_w8_l2048_id11_3_1_addr,
  output [8-1:0] ram_w8_l2048_id11_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id11_3_1_wdata,
  input ram_w8_l2048_id11_3_1_wenable
);

  reg [9-1:0] ram_w8_l2048_id11_3_0_daddr;
  reg [9-1:0] ram_w8_l2048_id11_3_1_daddr;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id11_3_0_wenable) begin
      mem[ram_w8_l2048_id11_3_0_addr] <= ram_w8_l2048_id11_3_0_wdata;
    end 
    ram_w8_l2048_id11_3_0_daddr <= ram_w8_l2048_id11_3_0_addr;
  end

  assign ram_w8_l2048_id11_3_0_rdata = mem[ram_w8_l2048_id11_3_0_daddr];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id11_3_1_wenable) begin
      mem[ram_w8_l2048_id11_3_1_addr] <= ram_w8_l2048_id11_3_1_wdata;
    end 
    ram_w8_l2048_id11_3_1_daddr <= ram_w8_l2048_id11_3_1_addr;
  end

  assign ram_w8_l2048_id11_3_1_rdata = mem[ram_w8_l2048_id11_3_1_daddr];

endmodule



module madd_0
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);


  madd_core_0
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_0
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [4-1:0] _b;
  reg signed [12-1:0] _c;
  wire signed [12-1:0] _mul;
  wire signed [12-1:0] _madd;
  reg signed [12-1:0] _pipe_madd0;
  reg signed [12-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_1
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);


  madd_core_1
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_1
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [4-1:0] _b;
  reg signed [12-1:0] _c;
  wire signed [12-1:0] _mul;
  wire signed [12-1:0] _madd;
  reg signed [12-1:0] _pipe_madd0;
  reg signed [12-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_2
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);


  madd_core_2
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_2
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [4-1:0] _b;
  reg signed [12-1:0] _c;
  wire signed [12-1:0] _mul;
  wire signed [12-1:0] _madd;
  reg signed [12-1:0] _pipe_madd0;
  reg signed [12-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_3
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);


  madd_core_3
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_3
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [4-1:0] _b;
  reg signed [12-1:0] _c;
  wire signed [12-1:0] _mul;
  wire signed [12-1:0] _madd;
  reg signed [12-1:0] _pipe_madd0;
  reg signed [12-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_4
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);


  madd_core_4
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_4
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [4-1:0] _b;
  reg signed [12-1:0] _c;
  wire signed [12-1:0] _mul;
  wire signed [12-1:0] _madd;
  reg signed [12-1:0] _pipe_madd0;
  reg signed [12-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_5
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);


  madd_core_5
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_5
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [4-1:0] _b;
  reg signed [12-1:0] _c;
  wire signed [12-1:0] _mul;
  wire signed [12-1:0] _madd;
  reg signed [12-1:0] _pipe_madd0;
  reg signed [12-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_6
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);


  madd_core_6
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_6
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [4-1:0] _b;
  reg signed [12-1:0] _c;
  wire signed [12-1:0] _mul;
  wire signed [12-1:0] _madd;
  reg signed [12-1:0] _pipe_madd0;
  reg signed [12-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_7
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);


  madd_core_7
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_7
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [4-1:0] _b;
  reg signed [12-1:0] _c;
  wire signed [12-1:0] _mul;
  wire signed [12-1:0] _madd;
  reg signed [12-1:0] _pipe_madd0;
  reg signed [12-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_8
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);


  madd_core_8
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_8
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [4-1:0] b,
  input [12-1:0] c,
  output [12-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [4-1:0] _b;
  reg signed [12-1:0] _c;
  wire signed [12-1:0] _mul;
  wire signed [12-1:0] _madd;
  reg signed [12-1:0] _pipe_madd0;
  reg signed [12-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module multiplier_0
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [8-1:0] b,
  output [40-1:0] c
);


  multiplier_core_0
  mult
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c)
  );


endmodule



module multiplier_core_0
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [8-1:0] b,
  output [40-1:0] c
);

  reg signed [32-1:0] _a;
  reg signed [8-1:0] _b;
  wire signed [40-1:0] _mul;
  reg signed [40-1:0] _pipe_mul0;
  reg signed [40-1:0] _pipe_mul1;
  assign _mul = _a * _b;
  assign c = _pipe_mul1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _pipe_mul0 <= _mul;
      _pipe_mul1 <= _pipe_mul0;
    end 
  end


endmodule

