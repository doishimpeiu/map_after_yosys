module nngenmod(CLK, RESETN, maxi_awaddr, maxi_awlen, maxi_awsize, maxi_awburst, maxi_awlock, maxi_awcache, maxi_awprot, maxi_awqos, maxi_awuser, maxi_awvalid, maxi_awready, maxi_wdata, maxi_wstrb, maxi_wlast, maxi_wvalid, maxi_wready, maxi_bresp, maxi_bvalid, maxi_bready, maxi_araddr, maxi_arlen, maxi_arsize, maxi_arburst, maxi_arlock, maxi_arcache, maxi_arprot, maxi_arqos, maxi_aruser, maxi_arvalid, maxi_arready, maxi_rdata, maxi_rresp, maxi_rlast, maxi_rvalid, maxi_rready, saxi_awaddr, saxi_awcache, saxi_awprot, saxi_awvalid, saxi_awready, saxi_wdata, saxi_wstrb, saxi_wvalid, saxi_wready, saxi_bresp, saxi_bvalid, saxi_bready, saxi_araddr, saxi_arcache, saxi_arprot, saxi_arvalid, saxi_arready, saxi_rdata, saxi_rresp, saxi_rvalid, saxi_rready);
  input CLK;
  input RESETN;
  input maxi_arready;
  input maxi_awready;
  input [1:0] maxi_bresp;
  input maxi_bvalid;
  input [31:0] maxi_rdata;
  input maxi_rlast;
  input [1:0] maxi_rresp;
  input maxi_rvalid;
  input maxi_wready;
  input [5:0] saxi_araddr;
  input [3:0] saxi_arcache;
  input [2:0] saxi_arprot;
  input saxi_arvalid;
  input [5:0] saxi_awaddr;
  input [3:0] saxi_awcache;
  input [2:0] saxi_awprot;
  input saxi_awvalid;
  input saxi_bready;
  input saxi_rready;
  input [31:0] saxi_wdata;
  input [3:0] saxi_wstrb;
  input saxi_wvalid;
  output [31:0] maxi_araddr;
  output [1:0] maxi_arburst;
  output [3:0] maxi_arcache;
  output [7:0] maxi_arlen;
  output maxi_arlock;
  output [2:0] maxi_arprot;
  output [3:0] maxi_arqos;
  output [2:0] maxi_arsize;
  output [1:0] maxi_aruser;
  output maxi_arvalid;
  output [31:0] maxi_awaddr;
  output [1:0] maxi_awburst;
  output [3:0] maxi_awcache;
  output [7:0] maxi_awlen;
  output maxi_awlock;
  output [2:0] maxi_awprot;
  output [3:0] maxi_awqos;
  output [2:0] maxi_awsize;
  output [1:0] maxi_awuser;
  output maxi_awvalid;
  output maxi_bready;
  output maxi_rready;
  output [31:0] maxi_wdata;
  output maxi_wlast;
  output [3:0] maxi_wstrb;
  output maxi_wvalid;
  output saxi_arready;
  output saxi_awready;
  output [1:0] saxi_bresp;
  output saxi_bvalid;
  output [31:0] saxi_rdata;
  output [1:0] saxi_rresp;
  output saxi_rvalid;
  output saxi_wready;
  wire _00000_;
  wire [3:0] _00001_;
  wire [3:0] _00002_;
  wire [3:0] _00003_;
  wire [3:0] _00004_;
  wire [3:0] _00005_;
  wire [3:0] _00006_;
  wire [3:0] _00007_;
  wire [7:0] _00008_;
  wire [7:0] _00009_;
  wire [7:0] _00010_;
  wire [7:0] _00011_;
  wire [7:0] _00012_;
  wire [7:0] _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire [7:0] _00017_;
  wire [7:0] _00018_;
  wire [7:0] _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire [7:0] _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire [7:0] _00033_;
  wire [7:0] _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire [3:0] _00042_;
  wire [3:0] _00043_;
  wire [3:0] _00044_;
  wire [3:0] _00045_;
  wire [3:0] _00046_;
  wire [3:0] _00047_;
  wire [3:0] _00048_;
  wire [3:0] _00049_;
  wire [7:0] _00050_;
  wire [7:0] _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire [3:0] _00059_;
  wire [3:0] _00060_;
  wire [3:0] _00061_;
  wire [3:0] _00062_;
  wire [3:0] _00063_;
  wire [3:0] _00064_;
  wire [3:0] _00065_;
  wire [3:0] _00066_;
  wire [7:0] _00067_;
  wire [7:0] _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire [3:0] _00076_;
  wire [3:0] _00077_;
  wire [3:0] _00078_;
  wire [3:0] _00079_;
  wire [3:0] _00080_;
  wire [3:0] _00081_;
  wire [3:0] _00082_;
  wire [3:0] _00083_;
  wire [7:0] _00084_;
  wire [7:0] _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire [3:0] _00093_;
  wire [3:0] _00094_;
  wire [3:0] _00095_;
  wire [3:0] _00096_;
  wire [3:0] _00097_;
  wire [3:0] _00098_;
  wire [3:0] _00099_;
  wire [3:0] _00100_;
  wire [7:0] _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire [3:0] _00109_;
  wire [3:0] _00110_;
  wire [3:0] _00111_;
  wire [3:0] _00112_;
  wire [3:0] _00113_;
  wire [3:0] _00114_;
  wire [3:0] _00115_;
  wire [3:0] _00116_;
  wire [7:0] _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire [3:0] _00125_;
  wire [3:0] _00126_;
  wire [3:0] _00127_;
  wire [3:0] _00128_;
  wire [3:0] _00129_;
  wire [3:0] _00130_;
  wire [3:0] _00131_;
  wire [3:0] _00132_;
  wire [7:0] _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire [3:0] _00141_;
  wire [3:0] _00142_;
  wire [3:0] _00143_;
  wire [3:0] _00144_;
  wire [3:0] _00145_;
  wire [3:0] _00146_;
  wire [3:0] _00147_;
  wire [3:0] _00148_;
  wire _00149_;
  wire [7:0] _00150_;
  wire [7:0] _00151_;
  wire [7:0] _00152_;
  wire [7:0] _00153_;
  wire [7:0] _00154_;
  wire [7:0] _00155_;
  wire [7:0] _00156_;
  wire [7:0] _00157_;
  wire [7:0] _00158_;
  wire [7:0] _00159_;
  wire [7:0] _00160_;
  wire [7:0] _00161_;
  wire [7:0] _00162_;
  wire [7:0] _00163_;
  wire [7:0] _00164_;
  wire [7:0] _00165_;
  wire [7:0] _00166_;
  wire [7:0] _00167_;
  wire [7:0] _00168_;
  wire [7:0] _00169_;
  wire [5:0] _00170_;
  wire [5:0] _00171_;
  wire [5:0] _00172_;
  wire [5:0] _00173_;
  wire [5:0] _00174_;
  wire [5:0] _00175_;
  wire [5:0] _00176_;
  wire [5:0] _00177_;
  wire [5:0] _00178_;
  wire [5:0] _00179_;
  wire [5:0] _00180_;
  wire [5:0] _00181_;
  wire [5:0] _00182_;
  wire [5:0] _00183_;
  wire [5:0] _00184_;
  wire [5:0] _00185_;
  wire [5:0] _00186_;
  wire [5:0] _00187_;
  wire [5:0] _00188_;
  wire [5:0] _00189_;
  wire [5:0] _00190_;
  wire [5:0] _00191_;
  wire [7:0] _00192_;
  wire [7:0] _00193_;
  wire [7:0] _00194_;
  wire [7:0] _00195_;
  wire [7:0] _00196_;
  wire [7:0] _00197_;
  wire [7:0] _00198_;
  wire [7:0] _00199_;
  wire [7:0] _00200_;
  wire [7:0] _00201_;
  wire [7:0] _00202_;
  wire [7:0] _00203_;
  wire [7:0] _00204_;
  wire [7:0] _00205_;
  wire [7:0] _00206_;
  wire [7:0] _00207_;
  wire [7:0] _00208_;
  wire [7:0] _00209_;
  wire [7:0] _00210_;
  wire [7:0] _00211_;
  wire [7:0] _00212_;
  wire [7:0] _00213_;
  wire [7:0] _00214_;
  wire [7:0] _00215_;
  wire [7:0] _00216_;
  wire [7:0] _00217_;
  wire [7:0] _00218_;
  wire [7:0] _00219_;
  wire [3:0] _00220_;
  wire [7:0] _00221_;
  wire [7:0] _00222_;
  wire [7:0] _00223_;
  wire [7:0] _00224_;
  wire [7:0] _00225_;
  wire [7:0] _00226_;
  wire [7:0] _00227_;
  wire [7:0] _00228_;
  wire [7:0] _00229_;
  wire [7:0] _00230_;
  wire [7:0] _00231_;
  wire [7:0] _00232_;
  wire [7:0] _00233_;
  wire [7:0] _00234_;
  wire [7:0] _00235_;
  wire [7:0] _00236_;
  wire [7:0] _00237_;
  wire [7:0] _00238_;
  wire [7:0] _00239_;
  wire [7:0] _00240_;
  wire [7:0] _00241_;
  wire [7:0] _00242_;
  wire [7:0] _00243_;
  wire [7:0] _00244_;
  wire [7:0] _00245_;
  wire [7:0] _00246_;
  wire [7:0] _00247_;
  wire [7:0] _00248_;
  wire [7:0] _00249_;
  wire [7:0] _00250_;
  wire [7:0] _00251_;
  wire [7:0] _00252_;
  wire [7:0] _00253_;
  wire [7:0] _00254_;
  wire [7:0] _00255_;
  wire [7:0] _00256_;
  wire [7:0] _00257_;
  wire [7:0] _00258_;
  wire [7:0] _00259_;
  wire [7:0] _00260_;
  wire [7:0] _00261_;
  wire [7:0] _00262_;
  wire [7:0] _00263_;
  wire [7:0] _00264_;
  wire [7:0] _00265_;
  wire [7:0] _00266_;
  wire [7:0] _00267_;
  wire [7:0] _00268_;
  wire [7:0] _00269_;
  wire [7:0] _00270_;
  wire [7:0] _00271_;
  wire [7:0] _00272_;
  wire [7:0] _00273_;
  wire [7:0] _00274_;
  wire [7:0] _00275_;
  wire [7:0] _00276_;
  wire [7:0] _00277_;
  wire [7:0] _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire [3:0] _00292_;
  wire [7:0] _00293_;
  wire [7:0] _00294_;
  wire [2:0] _00295_;
  wire [2:0] _00296_;
  wire [2:0] _00297_;
  wire [7:0] _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire [3:0] _00304_;
  wire [3:0] _00305_;
  wire [3:0] _00306_;
  wire [3:0] _00307_;
  wire [7:0] _00308_;
  wire [7:0] _00309_;
  wire _00310_;
  wire [7:0] _00311_;
  wire [7:0] _00312_;
  wire [7:0] _00313_;
  wire [7:0] _00314_;
  wire [7:0] _00315_;
  wire [7:0] _00316_;
  wire [7:0] _00317_;
  wire [7:0] _00318_;
  wire [7:0] _00319_;
  wire [7:0] _00320_;
  wire [7:0] _00321_;
  wire [7:0] _00322_;
  wire [7:0] _00323_;
  wire [7:0] _00324_;
  wire [10:0] _00325_;
  wire [10:0] _00326_;
  wire [10:0] _00327_;
  wire [10:0] _00328_;
  wire [10:0] _00329_;
  wire [10:0] _00330_;
  wire [10:0] _00331_;
  wire [10:0] _00332_;
  wire [10:0] _00333_;
  wire [10:0] _00334_;
  wire [10:0] _00335_;
  wire [10:0] _00336_;
  wire [10:0] _00337_;
  wire [10:0] _00338_;
  wire [10:0] _00339_;
  wire [10:0] _00340_;
  wire [7:0] _00341_;
  wire [7:0] _00342_;
  wire [7:0] _00343_;
  wire [7:0] _00344_;
  wire [7:0] _00345_;
  wire [7:0] _00346_;
  wire [7:0] _00347_;
  wire [7:0] _00348_;
  wire [7:0] _00349_;
  wire [7:0] _00350_;
  wire [7:0] _00351_;
  wire [7:0] _00352_;
  wire [7:0] _00353_;
  wire [7:0] _00354_;
  wire [7:0] _00355_;
  wire [7:0] _00356_;
  wire [7:0] _00357_;
  wire [7:0] _00358_;
  wire [7:0] _00359_;
  wire [7:0] _00360_;
  wire [7:0] _00361_;
  wire [7:0] _00362_;
  wire [3:0] _00363_;
  wire [7:0] _00364_;
  wire [7:0] _00365_;
  wire [7:0] _00366_;
  wire [7:0] _00367_;
  wire [7:0] _00368_;
  wire [7:0] _00369_;
  wire [7:0] _00370_;
  wire [7:0] _00371_;
  wire [7:0] _00372_;
  wire [7:0] _00373_;
  wire [7:0] _00374_;
  wire [7:0] _00375_;
  wire [7:0] _00376_;
  wire [7:0] _00377_;
  wire [7:0] _00378_;
  wire [7:0] _00379_;
  wire [7:0] _00380_;
  wire [7:0] _00381_;
  wire [7:0] _00382_;
  wire [7:0] _00383_;
  wire [7:0] _00384_;
  wire [7:0] _00385_;
  wire [7:0] _00386_;
  wire [7:0] _00387_;
  wire [7:0] _00388_;
  wire [7:0] _00389_;
  wire [7:0] _00390_;
  wire [7:0] _00391_;
  wire [7:0] _00392_;
  wire [7:0] _00393_;
  wire [7:0] _00394_;
  wire [7:0] _00395_;
  wire [7:0] _00396_;
  wire [7:0] _00397_;
  wire [7:0] _00398_;
  wire [7:0] _00399_;
  wire [7:0] _00400_;
  wire [7:0] _00401_;
  wire [7:0] _00402_;
  wire [7:0] _00403_;
  wire [7:0] _00404_;
  wire [7:0] _00405_;
  wire [7:0] _00406_;
  wire [7:0] _00407_;
  wire [7:0] _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire [7:0] _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire [7:0] _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire [7:0] _00485_;
  wire [7:0] _00486_;
  wire [7:0] _00487_;
  wire [3:0] _00488_;
  wire [3:0] _00489_;
  wire [3:0] _00490_;
  wire [3:0] _00491_;
  wire [3:0] _00492_;
  wire [3:0] _00493_;
  wire [3:0] _00494_;
  wire [3:0] _00495_;
  wire [3:0] _00496_;
  wire [3:0] _00497_;
  wire _00498_;
  wire [7:0] _00499_;
  wire [7:0] _00500_;
  wire [7:0] _00501_;
  wire [3:0] _00502_;
  wire [3:0] _00503_;
  wire [3:0] _00504_;
  wire [3:0] _00505_;
  wire [3:0] _00506_;
  wire [3:0] _00507_;
  wire [3:0] _00508_;
  wire [3:0] _00509_;
  wire [3:0] _00510_;
  wire [3:0] _00511_;
  wire _00512_;
  wire [7:0] _00513_;
  wire [7:0] _00514_;
  wire [7:0] _00515_;
  wire [3:0] _00516_;
  wire [3:0] _00517_;
  wire [3:0] _00518_;
  wire [3:0] _00519_;
  wire [3:0] _00520_;
  wire [3:0] _00521_;
  wire [3:0] _00522_;
  wire [3:0] _00523_;
  wire [3:0] _00524_;
  wire [3:0] _00525_;
  wire _00526_;
  wire [7:0] _00527_;
  wire [7:0] _00528_;
  wire [7:0] _00529_;
  wire [3:0] _00530_;
  wire [3:0] _00531_;
  wire [3:0] _00532_;
  wire [3:0] _00533_;
  wire [3:0] _00534_;
  wire [3:0] _00535_;
  wire [3:0] _00536_;
  wire [3:0] _00537_;
  wire [3:0] _00538_;
  wire [3:0] _00539_;
  wire _00540_;
  wire [7:0] _00541_;
  wire [7:0] _00542_;
  wire [7:0] _00543_;
  wire [3:0] _00544_;
  wire [3:0] _00545_;
  wire [3:0] _00546_;
  wire [3:0] _00547_;
  wire [3:0] _00548_;
  wire [3:0] _00549_;
  wire [3:0] _00550_;
  wire [3:0] _00551_;
  wire [3:0] _00552_;
  wire [3:0] _00553_;
  wire _00554_;
  wire [7:0] _00555_;
  wire [7:0] _00556_;
  wire [7:0] _00557_;
  wire [3:0] _00558_;
  wire [3:0] _00559_;
  wire [3:0] _00560_;
  wire [3:0] _00561_;
  wire [3:0] _00562_;
  wire [3:0] _00563_;
  wire [3:0] _00564_;
  wire [3:0] _00565_;
  wire [3:0] _00566_;
  wire [3:0] _00567_;
  wire _00568_;
  wire [7:0] _00569_;
  wire [7:0] _00570_;
  wire [7:0] _00571_;
  wire [3:0] _00572_;
  wire [3:0] _00573_;
  wire [3:0] _00574_;
  wire [3:0] _00575_;
  wire [3:0] _00576_;
  wire [3:0] _00577_;
  wire [3:0] _00578_;
  wire [3:0] _00579_;
  wire [3:0] _00580_;
  wire [3:0] _00581_;
  wire _00582_;
  wire [7:0] _00583_;
  wire [7:0] _00584_;
  wire [7:0] _00585_;
  wire [3:0] _00586_;
  wire [3:0] _00587_;
  wire [3:0] _00588_;
  wire [3:0] _00589_;
  wire [3:0] _00590_;
  wire [3:0] _00591_;
  wire [3:0] _00592_;
  wire [3:0] _00593_;
  wire [3:0] _00594_;
  wire [3:0] _00595_;
  wire _00596_;
  wire [7:0] _00597_;
  wire [7:0] _00598_;
  wire [7:0] _00599_;
  wire [3:0] _00600_;
  wire [3:0] _00601_;
  wire [3:0] _00602_;
  wire [3:0] _00603_;
  wire [3:0] _00604_;
  wire [3:0] _00605_;
  wire [3:0] _00606_;
  wire [3:0] _00607_;
  wire [3:0] _00608_;
  wire [3:0] _00609_;
  wire _00610_;
  wire [31:0] _00611_;
  wire [31:0] _00612_;
  wire [5:0] _00613_;
  wire [5:0] _00614_;
  wire [5:0] _00615_;
  wire [5:0] _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire [5:0] _00621_;
  wire [5:0] _00622_;
  wire [5:0] _00623_;
  wire [5:0] _00624_;
  wire [39:0] _00625_;
  wire _00626_;
  wire [7:0] _00627_;
  wire [7:0] _00628_;
  wire [7:0] _00629_;
  wire [7:0] _00630_;
  wire [7:0] _00631_;
  wire [7:0] _00632_;
  wire [7:0] _00633_;
  wire [7:0] _00634_;
  wire [7:0] _00635_;
  wire [7:0] _00636_;
  wire [7:0] _00637_;
  wire [7:0] _00638_;
  wire [7:0] _00639_;
  wire [7:0] _00640_;
  wire [7:0] _00641_;
  wire [7:0] _00642_;
  wire [7:0] _00643_;
  wire [7:0] _00644_;
  wire [7:0] _00645_;
  wire [7:0] _00646_;
  wire [7:0] _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire [3:0] _00656_;
  wire [3:0] _00657_;
  wire [3:0] _00658_;
  wire [3:0] _00659_;
  wire [3:0] _00660_;
  wire [3:0] _00661_;
  wire [3:0] _00662_;
  wire [3:0] _00663_;
  wire [7:0] _00664_;
  wire [7:0] _00665_;
  wire [7:0] _00666_;
  wire [7:0] _00667_;
  wire [7:0] _00668_;
  wire [7:0] _00669_;
  wire [7:0] _00670_;
  wire [7:0] _00671_;
  wire [7:0] _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire [3:0] _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire [11:0] _00692_;
  wire [11:0] _00693_;
  wire [11:0] _00694_;
  wire [11:0] _00695_;
  wire [11:0] _00696_;
  wire [11:0] _00697_;
  wire [11:0] _00698_;
  wire [11:0] _00699_;
  wire [11:0] _00700_;
  wire [31:0] _00701_;
  wire [31:0] _00702_;
  wire [31:0] _00703_;
  wire [31:0] _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire [31:0] _00801_;
  wire [31:0] _00802_;
  wire [31:0] _00803_;
  wire [31:0] _00804_;
  wire [31:0] _00805_;
  wire [31:0] _00806_;
  wire [31:0] _00807_;
  wire [31:0] _00808_;
  wire [31:0] _00809_;
  wire [31:0] _00810_;
  wire [31:0] _00811_;
  wire [31:0] _00812_;
  wire [31:0] _00813_;
  wire [31:0] _00814_;
  wire [31:0] _00815_;
  wire [31:0] _00816_;
  wire [31:0] _00817_;
  wire [31:0] _00818_;
  wire [31:0] _00819_;
  wire [31:0] _00820_;
  wire [31:0] _00821_;
  wire [31:0] _00822_;
  wire [31:0] _00823_;
  wire [31:0] _00824_;
  wire [31:0] _00825_;
  wire [31:0] _00826_;
  wire [31:0] _00827_;
  wire [31:0] _00828_;
  wire [31:0] _00829_;
  wire [31:0] _00830_;
  wire [31:0] _00831_;
  wire [31:0] _00832_;
  wire [31:0] _00833_;
  wire [31:0] _00834_;
  wire [31:0] _00835_;
  wire [31:0] _00836_;
  wire [31:0] _00837_;
  wire [31:0] _00838_;
  wire [31:0] _00839_;
  wire [31:0] _00840_;
  wire [31:0] _00841_;
  wire [31:0] _00842_;
  wire [31:0] _00843_;
  wire [31:0] _00844_;
  wire [31:0] _00845_;
  wire [32:0] _00846_;
  wire [32:0] _00847_;
  wire [32:0] _00848_;
  wire [32:0] _00849_;
  wire [32:0] _00850_;
  wire [32:0] _00851_;
  wire [32:0] _00852_;
  wire [32:0] _00853_;
  wire [32:0] _00854_;
  wire [32:0] _00855_;
  wire [32:0] _00856_;
  wire [32:0] _00857_;
  wire [32:0] _00858_;
  wire [32:0] _00859_;
  wire [32:0] _00860_;
  wire [32:0] _00861_;
  wire [32:0] _00862_;
  wire [32:0] _00863_;
  wire [32:0] _00864_;
  wire [32:0] _00865_;
  wire [32:0] _00866_;
  wire [32:0] _00867_;
  wire [32:0] _00868_;
  wire [32:0] _00869_;
  wire [32:0] _00870_;
  wire [32:0] _00871_;
  wire [32:0] _00872_;
  wire [32:0] _00873_;
  wire [32:0] _00874_;
  wire [32:0] _00875_;
  wire [32:0] _00876_;
  wire [32:0] _00877_;
  wire [32:0] _00878_;
  wire [32:0] _00879_;
  wire [32:0] _00880_;
  wire [32:0] _00881_;
  wire [32:0] _00882_;
  wire [32:0] _00883_;
  wire [32:0] _00884_;
  wire [32:0] _00885_;
  wire [32:0] _00886_;
  wire [32:0] _00887_;
  wire [32:0] _00888_;
  wire [32:0] _00889_;
  wire [32:0] _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire [31:0] _00937_;
  wire [31:0] _00938_;
  wire [31:0] _00939_;
  wire [31:0] _00940_;
  wire [31:0] _00941_;
  wire [31:0] _00942_;
  wire [31:0] _00943_;
  wire [31:0] _00944_;
  wire [31:0] _00945_;
  wire [31:0] _00946_;
  wire [31:0] _00947_;
  wire [31:0] _00948_;
  wire [31:0] _00949_;
  wire [31:0] _00950_;
  wire [31:0] _00951_;
  wire [31:0] _00952_;
  wire [31:0] _00953_;
  wire [31:0] _00954_;
  wire [31:0] _00955_;
  wire [31:0] _00956_;
  wire [31:0] _00957_;
  wire [31:0] _00958_;
  wire [31:0] _00959_;
  wire [31:0] _00960_;
  wire [31:0] _00961_;
  wire [31:0] _00962_;
  wire [31:0] _00963_;
  wire [31:0] _00964_;
  wire [31:0] _00965_;
  wire [31:0] _00966_;
  wire [31:0] _00967_;
  wire [31:0] _00968_;
  wire [31:0] _00969_;
  wire [31:0] _00970_;
  wire [31:0] _00971_;
  wire [31:0] _00972_;
  wire [31:0] _00973_;
  wire [31:0] _00974_;
  wire [31:0] _00975_;
  wire [31:0] _00976_;
  wire [31:0] _00977_;
  wire [32:0] _00978_;
  wire [32:0] _00979_;
  wire [32:0] _00980_;
  wire [32:0] _00981_;
  wire [32:0] _00982_;
  wire [32:0] _00983_;
  wire [32:0] _00984_;
  wire [32:0] _00985_;
  wire [32:0] _00986_;
  wire [32:0] _00987_;
  wire [32:0] _00988_;
  wire [32:0] _00989_;
  wire [32:0] _00990_;
  wire [32:0] _00991_;
  wire [32:0] _00992_;
  wire [32:0] _00993_;
  wire [32:0] _00994_;
  wire [32:0] _00995_;
  wire [32:0] _00996_;
  wire [32:0] _00997_;
  wire [32:0] _00998_;
  wire [32:0] _00999_;
  wire [32:0] _01000_;
  wire [32:0] _01001_;
  wire [32:0] _01002_;
  wire [32:0] _01003_;
  wire [32:0] _01004_;
  wire [32:0] _01005_;
  wire [32:0] _01006_;
  wire [32:0] _01007_;
  wire [32:0] _01008_;
  wire [32:0] _01009_;
  wire [32:0] _01010_;
  wire [32:0] _01011_;
  wire [32:0] _01012_;
  wire [32:0] _01013_;
  wire [32:0] _01014_;
  wire [32:0] _01015_;
  wire [32:0] _01016_;
  wire [32:0] _01017_;
  wire [32:0] _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire [31:0] _01061_;
  wire [31:0] _01062_;
  wire [31:0] _01063_;
  wire [31:0] _01064_;
  wire [31:0] _01065_;
  wire [31:0] _01066_;
  wire [31:0] _01067_;
  wire [31:0] _01068_;
  wire [31:0] _01069_;
  wire [32:0] _01070_;
  wire [32:0] _01071_;
  wire [32:0] _01072_;
  wire [32:0] _01073_;
  wire [32:0] _01074_;
  wire [32:0] _01075_;
  wire [32:0] _01076_;
  wire [32:0] _01077_;
  wire [32:0] _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire [11:0] _01089_;
  wire [11:0] _01090_;
  wire [11:0] _01091_;
  wire [11:0] _01092_;
  wire [11:0] _01093_;
  wire [11:0] _01094_;
  wire [11:0] _01095_;
  wire [11:0] _01096_;
  wire [11:0] _01097_;
  wire [31:0] _01098_;
  wire [31:0] _01099_;
  wire _01100_;
  wire [7:0] _01101_;
  wire [7:0] _01102_;
  wire _01103_;
  wire [31:0] _01104_;
  wire _01105_;
  wire [7:0] _01106_;
  wire _01107_;
  wire [7:0] _01108_;
  wire [1:0] _01109_;
  wire [1:0] _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire [7:0] _01132_;
  wire _01133_;
  wire [7:0] _01134_;
  wire _01135_;
  wire [7:0] _01136_;
  wire _01137_;
  wire [7:0] _01138_;
  wire [1:0] _01139_;
  wire [1:0] _01140_;
  wire _01141_;
  wire [1:0] _01142_;
  wire [1:0] _01143_;
  wire _01144_;
  wire [1:0] _01145_;
  wire [1:0] _01146_;
  wire _01147_;
  wire [2:0] _01148_;
  wire [2:0] _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire [7:0] _01222_;
  wire _01223_;
  wire [7:0] _01224_;
  wire _01225_;
  wire [7:0] _01226_;
  wire _01227_;
  wire [7:0] _01228_;
  wire [1:0] _01229_;
  wire [1:0] _01230_;
  wire _01231_;
  wire [1:0] _01232_;
  wire [1:0] _01233_;
  wire _01234_;
  wire [1:0] _01235_;
  wire [1:0] _01236_;
  wire _01237_;
  wire [1:0] _01238_;
  wire [1:0] _01239_;
  wire _01240_;
  wire [1:0] _01241_;
  wire [1:0] _01242_;
  wire _01243_;
  wire [1:0] _01244_;
  wire [1:0] _01245_;
  wire _01246_;
  wire [1:0] _01247_;
  wire [1:0] _01248_;
  wire _01249_;
  wire [1:0] _01250_;
  wire [1:0] _01251_;
  wire _01252_;
  wire [1:0] _01253_;
  wire [1:0] _01254_;
  wire _01255_;
  wire [1:0] _01256_;
  wire [1:0] _01257_;
  wire _01258_;
  wire [1:0] _01259_;
  wire [1:0] _01260_;
  wire _01261_;
  wire [2:0] _01262_;
  wire [2:0] _01263_;
  wire _01264_;
  wire [2:0] _01265_;
  wire [2:0] _01266_;
  wire _01267_;
  wire [2:0] _01268_;
  wire [2:0] _01269_;
  wire _01270_;
  wire [2:0] _01271_;
  wire [2:0] _01272_;
  wire _01273_;
  wire [2:0] _01274_;
  wire [2:0] _01275_;
  wire _01276_;
  wire [2:0] _01277_;
  wire [2:0] _01278_;
  wire _01279_;
  wire [2:0] _01280_;
  wire [2:0] _01281_;
  wire _01282_;
  wire [2:0] _01283_;
  wire [2:0] _01284_;
  wire _01285_;
  wire [2:0] _01286_;
  wire [2:0] _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire [7:0] _01370_;
  wire _01371_;
  wire [7:0] _01372_;
  wire [31:0] _01373_;
  wire [7:0] _01374_;
  wire [3:0] _01375_;
  wire [3:0] _01376_;
  wire [7:0] _01377_;
  wire [3:0] _01378_;
  wire [3:0] _01379_;
  wire [7:0] _01380_;
  wire [3:0] _01381_;
  wire [3:0] _01382_;
  wire [7:0] _01383_;
  wire [3:0] _01384_;
  wire [3:0] _01385_;
  wire [7:0] _01386_;
  wire [3:0] _01387_;
  wire [3:0] _01388_;
  wire [7:0] _01389_;
  wire [3:0] _01390_;
  wire [3:0] _01391_;
  wire [5:0] _01392_;
  wire [7:0] _01393_;
  wire [7:0] _01394_;
  wire [5:0] _01395_;
  wire [1:0] _01396_;
  wire [1:0] _01397_;
  wire [8:0] _01398_;
  wire [31:0] _01399_;
  wire [7:0] _01400_;
  wire [7:0] _01401_;
  wire [7:0] _01402_;
  wire [31:0] _01403_;
  wire [7:0] _01404_;
  wire [7:0] _01405_;
  wire [31:0] _01406_;
  wire _01407_;
  wire _01408_;
  wire [3:0] _01409_;
  wire [7:0] _01410_;
  wire [7:0] _01411_;
  wire [31:0] _01412_;
  wire [7:0] _01413_;
  wire [7:0] _01414_;
  wire [7:0] _01415_;
  wire [7:0] _01416_;
  wire [7:0] _01417_;
  wire [7:0] _01418_;
  wire [7:0] _01419_;
  wire [31:0] _01420_;
  wire [31:0] _01421_;
  wire [31:0] _01422_;
  wire [31:0] _01423_;
  wire [31:0] _01424_;
  wire [31:0] _01425_;
  wire [31:0] _01426_;
  wire [31:0] _01427_;
  wire [7:0] _01428_;
  wire [5:0] _01429_;
  wire [3:0] _01430_;
  wire [3:0] _01431_;
  wire [3:0] _01432_;
  wire [3:0] _01433_;
  wire [3:0] _01434_;
  wire [3:0] _01435_;
  wire [3:0] _01436_;
  wire [3:0] _01437_;
  wire [3:0] _01438_;
  wire [7:0] _01439_;
  wire [3:0] _01440_;
  wire [3:0] _01441_;
  wire [7:0] _01442_;
  wire [3:0] _01443_;
  wire [3:0] _01444_;
  wire [2:0] _01445_;
  wire [7:0] _01446_;
  wire [3:0] _01447_;
  wire [10:0] _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire [7:0] _01452_;
  wire [7:0] _01453_;
  wire [7:0] _01454_;
  wire [7:0] _01455_;
  wire [7:0] _01456_;
  wire _01457_;
  wire _01458_;
  wire [3:0] _01459_;
  wire [1:0] _01460_;
  wire [7:0] _01461_;
  wire [3:0] _01462_;
  wire [7:0] _01463_;
  wire [3:0] _01464_;
  wire [3:0] _01465_;
  wire _01466_;
  wire [11:0] _01467_;
  wire [11:0] _01468_;
  wire [11:0] _01469_;
  wire [31:0] _01470_;
  wire [11:0] _01471_;
  wire [11:0] _01472_;
  wire [11:0] _01473_;
  wire [11:0] _01474_;
  wire [7:0] _01475_;
  wire [7:0] _01476_;
  wire [7:0] _01477_;
  wire [7:0] _01478_;
  wire [7:0] _01479_;
  wire [7:0] _01480_;
  wire [7:0] _01481_;
  wire [7:0] _01482_;
  wire [7:0] _01483_;
  wire [7:0] _01484_;
  wire [7:0] _01485_;
  wire [7:0] _01486_;
  wire [7:0] _01487_;
  wire [7:0] _01488_;
  wire [7:0] _01489_;
  wire [7:0] _01490_;
  wire [7:0] _01491_;
  wire [7:0] _01492_;
  wire [7:0] _01493_;
  wire [7:0] _01494_;
  wire [7:0] _01495_;
  wire [7:0] _01496_;
  wire [7:0] _01497_;
  wire [7:0] _01498_;
  wire [7:0] _01499_;
  wire [7:0] _01500_;
  wire [7:0] _01501_;
  wire [7:0] _01502_;
  wire [7:0] _01503_;
  wire [7:0] _01504_;
  wire [7:0] _01505_;
  wire [7:0] _01506_;
  wire [7:0] _01507_;
  wire [7:0] _01508_;
  wire [7:0] _01509_;
  wire [7:0] _01510_;
  wire [7:0] _01511_;
  wire [7:0] _01512_;
  wire [7:0] _01513_;
  wire [7:0] _01514_;
  wire [7:0] _01515_;
  wire [7:0] _01516_;
  wire [7:0] _01517_;
  wire [7:0] _01518_;
  wire [7:0] _01519_;
  wire [7:0] _01520_;
  wire [7:0] _01521_;
  wire [7:0] _01522_;
  wire [7:0] _01523_;
  wire [7:0] _01524_;
  wire [7:0] _01525_;
  wire [7:0] _01526_;
  wire [7:0] _01527_;
  wire [7:0] _01528_;
  wire [7:0] _01529_;
  wire [7:0] _01530_;
  wire [7:0] _01531_;
  wire [7:0] _01532_;
  wire [7:0] _01533_;
  wire [39:0] _01534_;
  wire [39:0] _01535_;
  wire [7:0] _01536_;
  wire [7:0] _01537_;
  wire [7:0] _01538_;
  wire [7:0] _01539_;
  wire [7:0] _01540_;
  wire [7:0] _01541_;
  wire [7:0] _01542_;
  wire [7:0] _01543_;
  wire [7:0] _01544_;
  wire [7:0] _01545_;
  wire [11:0] _01546_;
  wire [7:0] _01547_;
  wire [8:0] _01548_;
  wire [7:0] _01549_;
  wire [7:0] _01550_;
  wire [7:0] _01551_;
  wire [7:0] _01552_;
  wire [7:0] _01553_;
  wire [11:0] _01554_;
  wire [7:0] _01555_;
  wire [7:0] _01556_;
  wire [7:0] _01557_;
  wire [7:0] _01558_;
  wire [7:0] _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire [31:0] _01579_;
  wire [31:0] _01580_;
  wire [31:0] _01581_;
  wire [31:0] _01582_;
  wire [31:0] _01583_;
  wire [31:0] _01584_;
  wire [31:0] _01585_;
  wire [31:0] _01586_;
  wire [31:0] _01587_;
  wire [31:0] _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire [7:0] _01592_;
  wire [7:0] _01593_;
  wire [7:0] _01594_;
  wire [7:0] _01595_;
  wire [3:0] _01596_;
  wire [3:0] _01597_;
  wire [7:0] _01598_;
  wire [3:0] _01599_;
  wire [3:0] _01600_;
  wire [3:0] _01601_;
  wire [3:0] _01602_;
  wire [3:0] _01603_;
  wire [3:0] _01604_;
  wire [7:0] _01605_;
  wire [7:0] _01606_;
  wire [7:0] _01607_;
  wire [7:0] _01608_;
  wire [7:0] _01609_;
  wire [7:0] _01610_;
  wire [7:0] _01611_;
  wire [7:0] _01612_;
  wire [3:0] _01613_;
  wire [3:0] _01614_;
  wire [3:0] _01615_;
  wire [3:0] _01616_;
  wire [7:0] _01617_;
  wire [3:0] _01618_;
  wire [3:0] _01619_;
  wire [3:0] _01620_;
  wire [3:0] _01621_;
  wire [7:0] _01622_;
  wire [7:0] _01623_;
  wire [7:0] _01624_;
  wire [7:0] _01625_;
  wire [7:0] _01626_;
  wire [7:0] _01627_;
  wire [7:0] _01628_;
  wire [7:0] _01629_;
  wire [7:0] _01630_;
  wire [7:0] _01631_;
  wire [7:0] _01632_;
  wire [7:0] _01633_;
  wire [7:0] _01634_;
  wire [7:0] _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire [31:0] _01705_;
  wire [31:0] _01706_;
  wire [31:0] _01707_;
  wire [31:0] _01708_;
  wire [7:0] _01709_;
  wire [32:0] _01710_;
  wire _01711_;
  wire [31:0] _01712_;
  wire [31:0] _01713_;
  wire [31:0] _01714_;
  wire [7:0] _01715_;
  wire [32:0] _01716_;
  wire _01717_;
  wire [31:0] _01718_;
  wire [31:0] _01719_;
  wire [31:0] _01720_;
  wire [7:0] _01721_;
  wire [32:0] _01722_;
  wire _01723_;
  wire [31:0] _01724_;
  wire [31:0] _01725_;
  wire [31:0] _01726_;
  wire [7:0] _01727_;
  wire [32:0] _01728_;
  wire _01729_;
  wire [31:0] _01730_;
  wire [31:0] _01731_;
  wire [31:0] _01732_;
  wire [7:0] _01733_;
  wire [32:0] _01734_;
  wire _01735_;
  wire [31:0] _01736_;
  wire [31:0] _01737_;
  wire [31:0] _01738_;
  wire [7:0] _01739_;
  wire [32:0] _01740_;
  wire _01741_;
  wire [31:0] _01742_;
  wire [31:0] _01743_;
  wire [31:0] _01744_;
  wire [7:0] _01745_;
  wire [32:0] _01746_;
  wire _01747_;
  wire [31:0] _01748_;
  wire [31:0] _01749_;
  wire [31:0] _01750_;
  wire [7:0] _01751_;
  wire [32:0] _01752_;
  wire _01753_;
  wire [31:0] _01754_;
  wire [31:0] _01755_;
  wire [31:0] _01756_;
  wire [7:0] _01757_;
  wire [32:0] _01758_;
  wire _01759_;
  wire [31:0] _01760_;
  wire [31:0] _01761_;
  wire [31:0] _01762_;
  wire [7:0] _01763_;
  wire [32:0] _01764_;
  wire _01765_;
  wire [31:0] _01766_;
  wire [31:0] _01767_;
  wire [31:0] _01768_;
  wire [7:0] _01769_;
  wire [32:0] _01770_;
  wire _01771_;
  wire [31:0] _01772_;
  wire [31:0] _01773_;
  wire [31:0] _01774_;
  wire [7:0] _01775_;
  wire [32:0] _01776_;
  wire _01777_;
  wire [31:0] _01778_;
  wire [32:0] _01779_;
  wire [31:0] _01780_;
  wire [31:0] _01781_;
  wire _01782_;
  wire [31:0] _01783_;
  wire [31:0] _01784_;
  wire [7:0] _01785_;
  wire [32:0] _01786_;
  wire [32:0] _01787_;
  wire _01788_;
  wire [31:0] _01789_;
  wire [32:0] _01790_;
  wire [31:0] _01791_;
  wire [31:0] _01792_;
  wire _01793_;
  wire [31:0] _01794_;
  wire [31:0] _01795_;
  wire [7:0] _01796_;
  wire [32:0] _01797_;
  wire [32:0] _01798_;
  wire _01799_;
  wire [3:0] _01800_;
  wire [3:0] _01801_;
  wire [3:0] _01802_;
  wire [3:0] _01803_;
  wire [3:0] _01804_;
  wire [3:0] _01805_;
  wire [3:0] _01806_;
  wire [5:0] _01807_;
  wire [3:0] _01808_;
  wire [3:0] _01809_;
  wire [31:0] _01810_;
  wire [7:0] _01811_;
  wire [7:0] _01812_;
  wire [31:0] _01813_;
  wire [7:0] _01814_;
  wire [7:0] _01815_;
  wire [7:0] _01816_;
  wire [31:0] _01817_;
  wire [7:0] _01818_;
  wire _01819_;
  wire [32:0] _01820_;
  wire [8:0] _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire [32:0] _01837_;
  wire [31:0] _01838_;
  wire [8:0] _01839_;
  wire [7:0] _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire [31:0] _01855_;
  wire [31:0] _01856_;
  wire [31:0] _01857_;
  wire [31:0] _01858_;
  wire [31:0] _01859_;
  wire [31:0] _01860_;
  wire [31:0] _01861_;
  wire [31:0] _01862_;
  wire [31:0] _01863_;
  wire [31:0] _01864_;
  wire [31:0] _01865_;
  wire [31:0] _01866_;
  wire [31:0] _01867_;
  wire [31:0] _01868_;
  wire [31:0] _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire [17:0] _01874_;
  wire [17:0] _01875_;
  wire [17:0] _01876_;
  wire [17:0] _01877_;
  wire [17:0] _01878_;
  wire [17:0] _01879_;
  wire [17:0] _01880_;
  wire [17:0] _01881_;
  wire [65:0] _01882_;
  wire [17:0] _01883_;
  wire [32:0] _01884_;
  wire [32:0] _01885_;
  wire [32:0] _01886_;
  wire [32:0] _01887_;
  wire [31:0] _01888_;
  wire [31:0] _01889_;
  wire [31:0] _01890_;
  wire [31:0] _01891_;
  wire [32:0] _01892_;
  wire [32:0] _01893_;
  wire [32:0] _01894_;
  wire [32:0] _01895_;
  wire [32:0] _01896_;
  wire [32:0] _01897_;
  wire [32:0] _01898_;
  wire [32:0] _01899_;
  wire [31:0] _01900_;
  wire [31:0] _01901_;
  wire [31:0] _01902_;
  wire [31:0] _01903_;
  wire [31:0] _01904_;
  wire [31:0] _01905_;
  wire [31:0] _01906_;
  wire [31:0] _01907_;
  wire [32:0] _01908_;
  wire [32:0] _01909_;
  wire [32:0] _01910_;
  wire [32:0] _01911_;
  wire [31:0] _01912_;
  wire [31:0] _01913_;
  wire [31:0] _01914_;
  wire [31:0] _01915_;
  wire [32:0] _01916_;
  wire [32:0] _01917_;
  wire [32:0] _01918_;
  wire [32:0] _01919_;
  wire [32:0] _01920_;
  wire [32:0] _01921_;
  wire [32:0] _01922_;
  wire [32:0] _01923_;
  wire [31:0] _01924_;
  wire [31:0] _01925_;
  wire [31:0] _01926_;
  wire [31:0] _01927_;
  wire [31:0] _01928_;
  wire [31:0] _01929_;
  wire [31:0] _01930_;
  wire [31:0] _01931_;
  wire [32:0] _01932_;
  wire [32:0] _01933_;
  wire [32:0] _01934_;
  wire [32:0] _01935_;
  wire [31:0] _01936_;
  wire [31:0] _01937_;
  wire [31:0] _01938_;
  wire [31:0] _01939_;
  wire [32:0] _01940_;
  wire [32:0] _01941_;
  wire [32:0] _01942_;
  wire [32:0] _01943_;
  wire [32:0] _01944_;
  wire [32:0] _01945_;
  wire [32:0] _01946_;
  wire [32:0] _01947_;
  wire [31:0] _01948_;
  wire [31:0] _01949_;
  wire [31:0] _01950_;
  wire [31:0] _01951_;
  wire [31:0] _01952_;
  wire [31:0] _01953_;
  wire [31:0] _01954_;
  wire [31:0] _01955_;
  wire [32:0] _01956_;
  wire [32:0] _01957_;
  wire [32:0] _01958_;
  wire [32:0] _01959_;
  wire [31:0] _01960_;
  wire [31:0] _01961_;
  wire [31:0] _01962_;
  wire [31:0] _01963_;
  wire [32:0] _01964_;
  wire [32:0] _01965_;
  wire [32:0] _01966_;
  wire [32:0] _01967_;
  wire [32:0] _01968_;
  wire [32:0] _01969_;
  wire [32:0] _01970_;
  wire [32:0] _01971_;
  wire [31:0] _01972_;
  wire [31:0] _01973_;
  wire [31:0] _01974_;
  wire [31:0] _01975_;
  wire [31:0] _01976_;
  wire [31:0] _01977_;
  wire [31:0] _01978_;
  wire [31:0] _01979_;
  wire [32:0] _01980_;
  wire [32:0] _01981_;
  wire [32:0] _01982_;
  wire [32:0] _01983_;
  wire [31:0] _01984_;
  wire [31:0] _01985_;
  wire [31:0] _01986_;
  wire [31:0] _01987_;
  wire [32:0] _01988_;
  wire [32:0] _01989_;
  wire [32:0] _01990_;
  wire [32:0] _01991_;
  wire [32:0] _01992_;
  wire [32:0] _01993_;
  wire [32:0] _01994_;
  wire [32:0] _01995_;
  wire [31:0] _01996_;
  wire [31:0] _01997_;
  wire [31:0] _01998_;
  wire [31:0] _01999_;
  wire [31:0] _02000_;
  wire [31:0] _02001_;
  wire [31:0] _02002_;
  wire [31:0] _02003_;
  wire [32:0] _02004_;
  wire [32:0] _02005_;
  wire [32:0] _02006_;
  wire [32:0] _02007_;
  wire [31:0] _02008_;
  wire [31:0] _02009_;
  wire [31:0] _02010_;
  wire [31:0] _02011_;
  wire [32:0] _02012_;
  wire [32:0] _02013_;
  wire [32:0] _02014_;
  wire [32:0] _02015_;
  wire [32:0] _02016_;
  wire [32:0] _02017_;
  wire [32:0] _02018_;
  wire [32:0] _02019_;
  wire [31:0] _02020_;
  wire [31:0] _02021_;
  wire [31:0] _02022_;
  wire [31:0] _02023_;
  wire [31:0] _02024_;
  wire [31:0] _02025_;
  wire [31:0] _02026_;
  wire [31:0] _02027_;
  wire [32:0] _02028_;
  wire [32:0] _02029_;
  wire [32:0] _02030_;
  wire [32:0] _02031_;
  wire [31:0] _02032_;
  wire [31:0] _02033_;
  wire [31:0] _02034_;
  wire [31:0] _02035_;
  wire [32:0] _02036_;
  wire [32:0] _02037_;
  wire [32:0] _02038_;
  wire [32:0] _02039_;
  wire [32:0] _02040_;
  wire [32:0] _02041_;
  wire [32:0] _02042_;
  wire [32:0] _02043_;
  wire [31:0] _02044_;
  wire [31:0] _02045_;
  wire [31:0] _02046_;
  wire [31:0] _02047_;
  wire [31:0] _02048_;
  wire [31:0] _02049_;
  wire [31:0] _02050_;
  wire [31:0] _02051_;
  wire [32:0] _02052_;
  wire [32:0] _02053_;
  wire [32:0] _02054_;
  wire [32:0] _02055_;
  wire [31:0] _02056_;
  wire [31:0] _02057_;
  wire [31:0] _02058_;
  wire [31:0] _02059_;
  wire [32:0] _02060_;
  wire [32:0] _02061_;
  wire [32:0] _02062_;
  wire [32:0] _02063_;
  wire [32:0] _02064_;
  wire [32:0] _02065_;
  wire [32:0] _02066_;
  wire [32:0] _02067_;
  wire [31:0] _02068_;
  wire [31:0] _02069_;
  wire [31:0] _02070_;
  wire [31:0] _02071_;
  wire [31:0] _02072_;
  wire [31:0] _02073_;
  wire [31:0] _02074_;
  wire [31:0] _02075_;
  wire [32:0] _02076_;
  wire [32:0] _02077_;
  wire [32:0] _02078_;
  wire [32:0] _02079_;
  wire [31:0] _02080_;
  wire [31:0] _02081_;
  wire [31:0] _02082_;
  wire [31:0] _02083_;
  wire [32:0] _02084_;
  wire [32:0] _02085_;
  wire [32:0] _02086_;
  wire [32:0] _02087_;
  wire [32:0] _02088_;
  wire [32:0] _02089_;
  wire [32:0] _02090_;
  wire [32:0] _02091_;
  wire [31:0] _02092_;
  wire [31:0] _02093_;
  wire [31:0] _02094_;
  wire [31:0] _02095_;
  wire [31:0] _02096_;
  wire [31:0] _02097_;
  wire [31:0] _02098_;
  wire [31:0] _02099_;
  wire [32:0] _02100_;
  wire [32:0] _02101_;
  wire [32:0] _02102_;
  wire [32:0] _02103_;
  wire [31:0] _02104_;
  wire [31:0] _02105_;
  wire [31:0] _02106_;
  wire [31:0] _02107_;
  wire [32:0] _02108_;
  wire [32:0] _02109_;
  wire [32:0] _02110_;
  wire [32:0] _02111_;
  wire [32:0] _02112_;
  wire [32:0] _02113_;
  wire [32:0] _02114_;
  wire [32:0] _02115_;
  wire [31:0] _02116_;
  wire [31:0] _02117_;
  wire [31:0] _02118_;
  wire [31:0] _02119_;
  wire [31:0] _02120_;
  wire [31:0] _02121_;
  wire [31:0] _02122_;
  wire [31:0] _02123_;
  wire [32:0] _02124_;
  wire [32:0] _02125_;
  wire [32:0] _02126_;
  wire [32:0] _02127_;
  wire [31:0] _02128_;
  wire [31:0] _02129_;
  wire [31:0] _02130_;
  wire [31:0] _02131_;
  wire [32:0] _02132_;
  wire [32:0] _02133_;
  wire [32:0] _02134_;
  wire [32:0] _02135_;
  wire [32:0] _02136_;
  wire [32:0] _02137_;
  wire [32:0] _02138_;
  wire [32:0] _02139_;
  wire [31:0] _02140_;
  wire [31:0] _02141_;
  wire [31:0] _02142_;
  wire [31:0] _02143_;
  wire [31:0] _02144_;
  wire [31:0] _02145_;
  wire [31:0] _02146_;
  wire [31:0] _02147_;
  wire [32:0] _02148_;
  wire [32:0] _02149_;
  wire [32:0] _02150_;
  wire [32:0] _02151_;
  wire [31:0] _02152_;
  wire [31:0] _02153_;
  wire [31:0] _02154_;
  wire [31:0] _02155_;
  wire [32:0] _02156_;
  wire [32:0] _02157_;
  wire [32:0] _02158_;
  wire [32:0] _02159_;
  wire [32:0] _02160_;
  wire [32:0] _02161_;
  wire [32:0] _02162_;
  wire [32:0] _02163_;
  wire [31:0] _02164_;
  wire [31:0] _02165_;
  wire [31:0] _02166_;
  wire [31:0] _02167_;
  wire [31:0] _02168_;
  wire [31:0] _02169_;
  wire [31:0] _02170_;
  wire [31:0] _02171_;
  wire [32:0] _02172_;
  wire [32:0] _02173_;
  wire [32:0] _02174_;
  wire [32:0] _02175_;
  wire [31:0] _02176_;
  wire [31:0] _02177_;
  wire [31:0] _02178_;
  wire [31:0] _02179_;
  wire [32:0] _02180_;
  wire [32:0] _02181_;
  wire [32:0] _02182_;
  wire [32:0] _02183_;
  wire [32:0] _02184_;
  wire [32:0] _02185_;
  wire [32:0] _02186_;
  wire [32:0] _02187_;
  wire [31:0] _02188_;
  wire [31:0] _02189_;
  wire [31:0] _02190_;
  wire [31:0] _02191_;
  wire [31:0] _02192_;
  wire [31:0] _02193_;
  wire [31:0] _02194_;
  wire [31:0] _02195_;
  wire [32:0] _02196_;
  wire [32:0] _02197_;
  wire [32:0] _02198_;
  wire [32:0] _02199_;
  wire [31:0] _02200_;
  wire [31:0] _02201_;
  wire [31:0] _02202_;
  wire [31:0] _02203_;
  wire [32:0] _02204_;
  wire [32:0] _02205_;
  wire [32:0] _02206_;
  wire [32:0] _02207_;
  wire [32:0] _02208_;
  wire [32:0] _02209_;
  wire [32:0] _02210_;
  wire [32:0] _02211_;
  wire [31:0] _02212_;
  wire [31:0] _02213_;
  wire [31:0] _02214_;
  wire [31:0] _02215_;
  wire [31:0] _02216_;
  wire [31:0] _02217_;
  wire [31:0] _02218_;
  wire [31:0] _02219_;
  wire [32:0] _02220_;
  wire [32:0] _02221_;
  wire [32:0] _02222_;
  wire [32:0] _02223_;
  wire [31:0] _02224_;
  wire [31:0] _02225_;
  wire [31:0] _02226_;
  wire [31:0] _02227_;
  wire [32:0] _02228_;
  wire [32:0] _02229_;
  wire [32:0] _02230_;
  wire [32:0] _02231_;
  wire [32:0] _02232_;
  wire [32:0] _02233_;
  wire [32:0] _02234_;
  wire [32:0] _02235_;
  wire [31:0] _02236_;
  wire [31:0] _02237_;
  wire [31:0] _02238_;
  wire [31:0] _02239_;
  wire [31:0] _02240_;
  wire [31:0] _02241_;
  wire [31:0] _02242_;
  wire [31:0] _02243_;
  wire [32:0] _02244_;
  wire [32:0] _02245_;
  wire [32:0] _02246_;
  wire [32:0] _02247_;
  wire [31:0] _02248_;
  wire [31:0] _02249_;
  wire [31:0] _02250_;
  wire [31:0] _02251_;
  wire [32:0] _02252_;
  wire [32:0] _02253_;
  wire [32:0] _02254_;
  wire [32:0] _02255_;
  wire [32:0] _02256_;
  wire [32:0] _02257_;
  wire [32:0] _02258_;
  wire [32:0] _02259_;
  wire [31:0] _02260_;
  wire [31:0] _02261_;
  wire [31:0] _02262_;
  wire [31:0] _02263_;
  wire [31:0] _02264_;
  wire [31:0] _02265_;
  wire [31:0] _02266_;
  wire [31:0] _02267_;
  wire [32:0] _02268_;
  wire [32:0] _02269_;
  wire [32:0] _02270_;
  wire [32:0] _02271_;
  wire [31:0] _02272_;
  wire [31:0] _02273_;
  wire [31:0] _02274_;
  wire [31:0] _02275_;
  wire [32:0] _02276_;
  wire [32:0] _02277_;
  wire [32:0] _02278_;
  wire [32:0] _02279_;
  wire [32:0] _02280_;
  wire [32:0] _02281_;
  wire [32:0] _02282_;
  wire [32:0] _02283_;
  wire [31:0] _02284_;
  wire [31:0] _02285_;
  wire [31:0] _02286_;
  wire [31:0] _02287_;
  wire [31:0] _02288_;
  wire [31:0] _02289_;
  wire [31:0] _02290_;
  wire [31:0] _02291_;
  wire [32:0] _02292_;
  wire [32:0] _02293_;
  wire [32:0] _02294_;
  wire [32:0] _02295_;
  wire [31:0] _02296_;
  wire [31:0] _02297_;
  wire [31:0] _02298_;
  wire [31:0] _02299_;
  wire [32:0] _02300_;
  wire [32:0] _02301_;
  wire [32:0] _02302_;
  wire [32:0] _02303_;
  wire [32:0] _02304_;
  wire [32:0] _02305_;
  wire [32:0] _02306_;
  wire [32:0] _02307_;
  wire [31:0] _02308_;
  wire [31:0] _02309_;
  wire [31:0] _02310_;
  wire [31:0] _02311_;
  wire [31:0] _02312_;
  wire [31:0] _02313_;
  wire [31:0] _02314_;
  wire [31:0] _02315_;
  wire [32:0] _02316_;
  wire [32:0] _02317_;
  wire [32:0] _02318_;
  wire [32:0] _02319_;
  wire [31:0] _02320_;
  wire [31:0] _02321_;
  wire [31:0] _02322_;
  wire [31:0] _02323_;
  wire [32:0] _02324_;
  wire [32:0] _02325_;
  wire [32:0] _02326_;
  wire [32:0] _02327_;
  wire [32:0] _02328_;
  wire [32:0] _02329_;
  wire [32:0] _02330_;
  wire [32:0] _02331_;
  wire [31:0] _02332_;
  wire [31:0] _02333_;
  wire [31:0] _02334_;
  wire [31:0] _02335_;
  wire [31:0] _02336_;
  wire [31:0] _02337_;
  wire [31:0] _02338_;
  wire [31:0] _02339_;
  wire [32:0] _02340_;
  wire [32:0] _02341_;
  wire [32:0] _02342_;
  wire [32:0] _02343_;
  wire [31:0] _02344_;
  wire [31:0] _02345_;
  wire [31:0] _02346_;
  wire [31:0] _02347_;
  wire [32:0] _02348_;
  wire [32:0] _02349_;
  wire [32:0] _02350_;
  wire [32:0] _02351_;
  wire [32:0] _02352_;
  wire [32:0] _02353_;
  wire [32:0] _02354_;
  wire [32:0] _02355_;
  wire [31:0] _02356_;
  wire [31:0] _02357_;
  wire [31:0] _02358_;
  wire [31:0] _02359_;
  wire [31:0] _02360_;
  wire [31:0] _02361_;
  wire [31:0] _02362_;
  wire [31:0] _02363_;
  wire [32:0] _02364_;
  wire [32:0] _02365_;
  wire [32:0] _02366_;
  wire [32:0] _02367_;
  wire [31:0] _02368_;
  wire [31:0] _02369_;
  wire [31:0] _02370_;
  wire [31:0] _02371_;
  wire [32:0] _02372_;
  wire [32:0] _02373_;
  wire [32:0] _02374_;
  wire [32:0] _02375_;
  wire [32:0] _02376_;
  wire [32:0] _02377_;
  wire [32:0] _02378_;
  wire [32:0] _02379_;
  wire [31:0] _02380_;
  wire [31:0] _02381_;
  wire [31:0] _02382_;
  wire [31:0] _02383_;
  wire [31:0] _02384_;
  wire [31:0] _02385_;
  wire [31:0] _02386_;
  wire [31:0] _02387_;
  wire [32:0] _02388_;
  wire [32:0] _02389_;
  wire [32:0] _02390_;
  wire [32:0] _02391_;
  wire [31:0] _02392_;
  wire [31:0] _02393_;
  wire [31:0] _02394_;
  wire [31:0] _02395_;
  wire [32:0] _02396_;
  wire [32:0] _02397_;
  wire [32:0] _02398_;
  wire [32:0] _02399_;
  wire [32:0] _02400_;
  wire [32:0] _02401_;
  wire [32:0] _02402_;
  wire [32:0] _02403_;
  wire [31:0] _02404_;
  wire [31:0] _02405_;
  wire [31:0] _02406_;
  wire [31:0] _02407_;
  wire [31:0] _02408_;
  wire [31:0] _02409_;
  wire [31:0] _02410_;
  wire [31:0] _02411_;
  wire [32:0] _02412_;
  wire [32:0] _02413_;
  wire [32:0] _02414_;
  wire [32:0] _02415_;
  wire [31:0] _02416_;
  wire [31:0] _02417_;
  wire [31:0] _02418_;
  wire [31:0] _02419_;
  wire [32:0] _02420_;
  wire [32:0] _02421_;
  wire [32:0] _02422_;
  wire [32:0] _02423_;
  wire [32:0] _02424_;
  wire [32:0] _02425_;
  wire [32:0] _02426_;
  wire [32:0] _02427_;
  wire [31:0] _02428_;
  wire [31:0] _02429_;
  wire [31:0] _02430_;
  wire [31:0] _02431_;
  wire [31:0] _02432_;
  wire [31:0] _02433_;
  wire [31:0] _02434_;
  wire [31:0] _02435_;
  wire [32:0] _02436_;
  wire [32:0] _02437_;
  wire [32:0] _02438_;
  wire [32:0] _02439_;
  wire [31:0] _02440_;
  wire [31:0] _02441_;
  wire [31:0] _02442_;
  wire [31:0] _02443_;
  wire [32:0] _02444_;
  wire [32:0] _02445_;
  wire [32:0] _02446_;
  wire [32:0] _02447_;
  wire [32:0] _02448_;
  wire [32:0] _02449_;
  wire [32:0] _02450_;
  wire [32:0] _02451_;
  wire [31:0] _02452_;
  wire [31:0] _02453_;
  wire [31:0] _02454_;
  wire [31:0] _02455_;
  wire [31:0] _02456_;
  wire [31:0] _02457_;
  wire [31:0] _02458_;
  wire [31:0] _02459_;
  wire [32:0] _02460_;
  wire [32:0] _02461_;
  wire [32:0] _02462_;
  wire [32:0] _02463_;
  wire [31:0] _02464_;
  wire [31:0] _02465_;
  wire [31:0] _02466_;
  wire [31:0] _02467_;
  wire [32:0] _02468_;
  wire [32:0] _02469_;
  wire [32:0] _02470_;
  wire [32:0] _02471_;
  wire [32:0] _02472_;
  wire [32:0] _02473_;
  wire [32:0] _02474_;
  wire [32:0] _02475_;
  wire [31:0] _02476_;
  wire [31:0] _02477_;
  wire [31:0] _02478_;
  wire [31:0] _02479_;
  wire [31:0] _02480_;
  wire [31:0] _02481_;
  wire [31:0] _02482_;
  wire [31:0] _02483_;
  wire [11:0] _02484_;
  wire [11:0] _02485_;
  wire [11:0] _02486_;
  wire [11:0] _02487_;
  wire [11:0] _02488_;
  wire [11:0] _02489_;
  wire [11:0] _02490_;
  wire [31:0] _02491_;
  wire [39:0] _02492_;
  wire [11:0] _02493_;
  wire [11:0] _02494_;
  wire [5:0] _02495_;
  wire _02496_;
  wire _02497_;
  wire [3:0] _02498_;
  wire [1:0] _02499_;
  wire [1:0] _02500_;
  wire [8:0] _02501_;
  wire _02502_;
  wire [31:0] _02503_;
  wire [32:0] _02504_;
  wire [31:0] _02505_;
  wire [2:0] _02506_;
  wire [31:0] _02507_;
  wire [7:0] _02508_;
  wire [32:0] _02509_;
  wire [31:0] _02510_;
  wire [31:0] _02511_;
  wire [31:0] _02512_;
  wire [7:0] _02513_;
  wire _02514_;
  wire _02515_;
  wire [7:0] _02516_;
  wire _02517_;
  wire [7:0] _02518_;
  wire _02519_;
  wire [7:0] _02520_;
  wire _02521_;
  wire [2:0] _02522_;
  wire [31:0] _02523_;
  wire [31:0] _02524_;
  wire [31:0] _02525_;
  wire [31:0] _02526_;
  wire _02527_;
  wire _02528_;
  wire [7:0] _02529_;
  wire _02530_;
  wire [2:0] _02531_;
  wire [31:0] _02532_;
  wire [31:0] _02533_;
  wire [31:0] _02534_;
  wire [31:0] _02535_;
  wire _02536_;
  wire _02537_;
  wire [7:0] _02538_;
  wire _02539_;
  wire [2:0] _02540_;
  wire [31:0] _02541_;
  wire [31:0] _02542_;
  wire [31:0] _02543_;
  wire [31:0] _02544_;
  wire _02545_;
  wire _02546_;
  wire [7:0] _02547_;
  wire _02548_;
  wire [2:0] _02549_;
  wire [31:0] _02550_;
  wire [31:0] _02551_;
  wire [31:0] _02552_;
  wire [31:0] _02553_;
  wire _02554_;
  wire _02555_;
  wire [7:0] _02556_;
  wire _02557_;
  wire [2:0] _02558_;
  wire [31:0] _02559_;
  wire [31:0] _02560_;
  wire [31:0] _02561_;
  wire [31:0] _02562_;
  wire _02563_;
  wire _02564_;
  wire [7:0] _02565_;
  wire _02566_;
  wire [2:0] _02567_;
  wire [31:0] _02568_;
  wire [31:0] _02569_;
  wire [31:0] _02570_;
  wire [31:0] _02571_;
  wire _02572_;
  wire _02573_;
  wire [7:0] _02574_;
  wire _02575_;
  wire [2:0] _02576_;
  wire [31:0] _02577_;
  wire [31:0] _02578_;
  wire [31:0] _02579_;
  wire [31:0] _02580_;
  wire _02581_;
  wire _02582_;
  wire [7:0] _02583_;
  wire _02584_;
  wire [2:0] _02585_;
  wire [31:0] _02586_;
  wire [31:0] _02587_;
  wire [31:0] _02588_;
  wire [31:0] _02589_;
  wire _02590_;
  wire _02591_;
  wire [7:0] _02592_;
  wire _02593_;
  wire [2:0] _02594_;
  wire [31:0] _02595_;
  wire [31:0] _02596_;
  wire [31:0] _02597_;
  wire [31:0] _02598_;
  wire _02599_;
  wire _02600_;
  wire [7:0] _02601_;
  wire _02602_;
  wire [2:0] _02603_;
  wire [31:0] _02604_;
  wire [31:0] _02605_;
  wire [31:0] _02606_;
  wire [31:0] _02607_;
  wire _02608_;
  wire _02609_;
  wire [7:0] _02610_;
  wire _02611_;
  wire [2:0] _02612_;
  wire [31:0] _02613_;
  wire [31:0] _02614_;
  wire [31:0] _02615_;
  wire [31:0] _02616_;
  wire _02617_;
  wire _02618_;
  wire [7:0] _02619_;
  wire _02620_;
  wire [2:0] _02621_;
  wire [31:0] _02622_;
  wire [31:0] _02623_;
  wire [31:0] _02624_;
  wire [31:0] _02625_;
  wire _02626_;
  wire _02627_;
  wire [7:0] _02628_;
  wire _02629_;
  wire [2:0] _02630_;
  wire [31:0] _02631_;
  wire [31:0] _02632_;
  wire [31:0] _02633_;
  wire [31:0] _02634_;
  wire _02635_;
  wire _02636_;
  wire [7:0] _02637_;
  wire _02638_;
  wire [2:0] _02639_;
  wire [31:0] _02640_;
  wire [31:0] _02641_;
  wire [31:0] _02642_;
  wire [31:0] _02643_;
  wire _02644_;
  wire _02645_;
  wire [7:0] _02646_;
  wire _02647_;
  wire [2:0] _02648_;
  wire [31:0] _02649_;
  wire [31:0] _02650_;
  wire [31:0] _02651_;
  wire [31:0] _02652_;
  wire _02653_;
  wire _02654_;
  wire [7:0] _02655_;
  wire _02656_;
  wire [2:0] _02657_;
  wire [31:0] _02658_;
  wire [31:0] _02659_;
  wire [31:0] _02660_;
  wire [31:0] _02661_;
  wire _02662_;
  wire _02663_;
  wire [7:0] _02664_;
  wire _02665_;
  wire [2:0] _02666_;
  wire [31:0] _02667_;
  wire [31:0] _02668_;
  wire [31:0] _02669_;
  wire [31:0] _02670_;
  wire _02671_;
  wire _02672_;
  wire [7:0] _02673_;
  wire _02674_;
  wire [2:0] _02675_;
  wire [31:0] _02676_;
  wire [31:0] _02677_;
  wire [31:0] _02678_;
  wire [31:0] _02679_;
  wire _02680_;
  wire _02681_;
  wire [7:0] _02682_;
  wire _02683_;
  wire [2:0] _02684_;
  wire [31:0] _02685_;
  wire [31:0] _02686_;
  wire [31:0] _02687_;
  wire [31:0] _02688_;
  wire _02689_;
  wire _02690_;
  wire [7:0] _02691_;
  wire _02692_;
  wire [2:0] _02693_;
  wire [31:0] _02694_;
  wire [31:0] _02695_;
  wire [31:0] _02696_;
  wire [31:0] _02697_;
  wire _02698_;
  wire _02699_;
  wire [7:0] _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire [10:0] _02704_;
  wire _02705_;
  wire _02706_;
  wire [3:0] _02707_;
  wire [1:0] _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire [31:0] _02713_;
  wire [32:0] _02714_;
  wire [31:0] _02715_;
  wire [2:0] _02716_;
  wire [31:0] _02717_;
  wire [7:0] _02718_;
  wire [32:0] _02719_;
  wire [31:0] _02720_;
  wire [31:0] _02721_;
  wire [31:0] _02722_;
  wire [7:0] _02723_;
  wire _02724_;
  wire _02725_;
  wire [7:0] _02726_;
  wire _02727_;
  wire [7:0] _02728_;
  wire _02729_;
  wire [7:0] _02730_;
  wire _02731_;
  wire [2:0] _02732_;
  wire [31:0] _02733_;
  wire [31:0] _02734_;
  wire [31:0] _02735_;
  wire [31:0] _02736_;
  wire _02737_;
  wire _02738_;
  wire [7:0] _02739_;
  wire _02740_;
  wire [2:0] _02741_;
  wire [31:0] _02742_;
  wire [31:0] _02743_;
  wire [31:0] _02744_;
  wire [31:0] _02745_;
  wire _02746_;
  wire _02747_;
  wire [7:0] _02748_;
  wire _02749_;
  wire [2:0] _02750_;
  wire [31:0] _02751_;
  wire [31:0] _02752_;
  wire [31:0] _02753_;
  wire [31:0] _02754_;
  wire _02755_;
  wire _02756_;
  wire [7:0] _02757_;
  wire _02758_;
  wire [2:0] _02759_;
  wire [31:0] _02760_;
  wire [31:0] _02761_;
  wire [31:0] _02762_;
  wire [31:0] _02763_;
  wire _02764_;
  wire _02765_;
  wire [7:0] _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire [2:0] _02770_;
  wire [3:0] _02771_;
  wire _02772_;
  wire [31:0] _02773_;
  wire _02774_;
  wire [32:0] _02775_;
  wire [31:0] _02776_;
  wire [2:0] _02777_;
  wire [31:0] _02778_;
  wire [7:0] _02779_;
  wire [32:0] _02780_;
  wire [31:0] _02781_;
  wire [31:0] _02782_;
  wire [31:0] _02783_;
  wire [7:0] _02784_;
  wire _02785_;
  wire _02786_;
  wire [2:0] _02787_;
  wire [31:0] _02788_;
  wire [31:0] _02789_;
  wire [31:0] _02790_;
  wire [31:0] _02791_;
  wire _02792_;
  wire _02793_;
  wire [7:0] _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire [39:0] _02852_;
  wire [5:0] _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire [33:0] _02858_;
  wire _02859_;
  wire [10:0] _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire [33:0] _02865_;
  wire [8:0] _02866_;
  wire [33:0] _02867_;
  wire _02868_;
  wire _02869_;
  wire [9:0] _02870_;
  wire [9:0] _02871_;
  wire [9:0] _02872_;
  wire [9:0] _02873_;
  wire _02874_;
  wire _02875_;
  wire [9:0] _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire [33:0] _02880_;
  wire _02881_;
  wire [9:0] _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire [33:0] _02887_;
  wire _02888_;
  wire [9:0] _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire [33:0] _02894_;
  wire _02895_;
  wire [9:0] _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire [33:0] _02901_;
  wire [9:0] _02902_;
  wire _02903_;
  wire [33:0] _02904_;
  wire _02905_;
  wire [33:0] _02906_;
  wire _02907_;
  wire [33:0] _02908_;
  wire _02909_;
  wire [33:0] _02910_;
  wire _02911_;
  wire [33:0] _02912_;
  wire _02913_;
  wire [33:0] _02914_;
  wire _02915_;
  wire [33:0] _02916_;
  wire _02917_;
  wire [33:0] _02918_;
  wire _02919_;
  wire [33:0] _02920_;
  wire _02921_;
  wire [33:0] _02922_;
  wire _02923_;
  wire [33:0] _02924_;
  wire _02925_;
  wire [33:0] _02926_;
  wire _02927_;
  wire [33:0] _02928_;
  wire _02929_;
  wire [33:0] _02930_;
  wire _02931_;
  wire [33:0] _02932_;
  wire _02933_;
  wire [33:0] _02934_;
  wire _02935_;
  wire [33:0] _02936_;
  wire _02937_;
  wire [3:0] _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire [10:0] _02943_;
  wire [33:0] _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire [33:0] _02948_;
  wire _02949_;
  wire _02950_;
  wire [33:0] _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire [33:0] _02958_;
  wire _02959_;
  wire [9:0] _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire [33:0] _02965_;
  wire _02966_;
  wire [9:0] _02967_;
  wire [9:0] _02968_;
  wire [9:0] _02969_;
  wire [9:0] _02970_;
  wire [9:0] _02971_;
  wire _02972_;
  wire [9:0] _02973_;
  wire [9:0] _02974_;
  wire [9:0] _02975_;
  wire [33:0] _02976_;
  wire _02977_;
  wire [3:0] _02978_;
  wire [10:0] _02979_;
  wire [33:0] _02980_;
  wire _02981_;
  wire [9:0] _02982_;
  wire [9:0] _02983_;
  wire [9:0] _02984_;
  wire [9:0] _02985_;
  wire [9:0] _02986_;
  wire [33:0] _02987_;
  wire [9:0] _02988_;
  wire [9:0] _02989_;
  wire [9:0] _02990_;
  wire [9:0] _02991_;
  wire _02992_;
  wire [33:0] _02993_;
  wire [3:0] _02994_;
  wire [10:0] _02995_;
  wire [33:0] _02996_;
  wire _02997_;
  wire [9:0] _02998_;
  wire [9:0] _02999_;
  wire [9:0] _03000_;
  wire [9:0] _03001_;
  wire _03002_;
  wire _03003_;
  wire [9:0] _03004_;
  wire [9:0] _03005_;
  wire [9:0] _03006_;
  wire [9:0] _03007_;
  wire [9:0] _03008_;
  wire [8:0] _03009_;
  wire [3:0] _03010_;
  wire [10:0] _03011_;
  wire [33:0] _03012_;
  wire _03013_;
  wire [9:0] _03014_;
  wire [9:0] _03015_;
  wire [9:0] _03016_;
  wire [9:0] _03017_;
  wire [9:0] _03018_;
  wire [9:0] _03019_;
  wire [9:0] _03020_;
  wire [9:0] _03021_;
  wire [9:0] _03022_;
  wire [3:0] _03023_;
  wire [10:0] _03024_;
  wire [33:0] _03025_;
  wire _03026_;
  wire [9:0] _03027_;
  wire [9:0] _03028_;
  wire [33:0] _03029_;
  wire [9:0] _03030_;
  wire [9:0] _03031_;
  wire [9:0] _03032_;
  wire [9:0] _03033_;
  wire [9:0] _03034_;
  wire [9:0] _03035_;
  wire [9:0] _03036_;
  wire _03037_;
  wire [33:0] _03038_;
  wire [3:0] _03039_;
  wire _03040_;
  wire [9:0] _03041_;
  wire [33:0] _03042_;
  wire _03043_;
  wire [8:0] _03044_;
  wire [8:0] _03045_;
  wire [8:0] _03046_;
  wire [33:0] _03047_;
  wire _03048_;
  wire [1:0] _03049_;
  wire [9:0] _03050_;
  wire [33:0] _03051_;
  wire _03052_;
  wire [8:0] _03053_;
  wire [8:0] _03054_;
  wire [8:0] _03055_;
  wire _03056_;
  wire [1:0] _03057_;
  wire [9:0] _03058_;
  wire [33:0] _03059_;
  wire _03060_;
  wire [33:0] _03061_;
  wire [8:0] _03062_;
  wire [8:0] _03063_;
  wire [8:0] _03064_;
  wire [1:0] _03065_;
  wire _03066_;
  wire [9:0] _03067_;
  wire [33:0] _03068_;
  wire _03069_;
  wire [8:0] _03070_;
  wire [8:0] _03071_;
  wire [8:0] _03072_;
  wire [1:0] _03073_;
  wire [9:0] _03074_;
  wire [33:0] _03075_;
  wire _03076_;
  wire [8:0] _03077_;
  wire [8:0] _03078_;
  wire [8:0] _03079_;
  wire [1:0] _03080_;
  wire [9:0] _03081_;
  wire [33:0] _03082_;
  wire _03083_;
  wire [8:0] _03084_;
  wire [8:0] _03085_;
  wire [8:0] _03086_;
  wire [1:0] _03087_;
  wire [9:0] _03088_;
  wire [33:0] _03089_;
  wire _03090_;
  wire [8:0] _03091_;
  wire [8:0] _03092_;
  wire [8:0] _03093_;
  wire [1:0] _03094_;
  wire [9:0] _03095_;
  wire [33:0] _03096_;
  wire _03097_;
  wire [10:0] _03098_;
  wire [8:0] _03099_;
  wire [8:0] _03100_;
  wire [8:0] _03101_;
  wire [1:0] _03102_;
  wire [33:0] _03103_;
  wire _03104_;
  wire [9:0] _03105_;
  wire [33:0] _03106_;
  wire _03107_;
  wire [8:0] _03108_;
  wire [8:0] _03109_;
  wire _03110_;
  wire [8:0] _03111_;
  wire [1:0] _03112_;
  wire [9:0] _03113_;
  wire [33:0] _03114_;
  wire [9:0] _03115_;
  wire _03116_;
  wire [8:0] _03117_;
  wire [8:0] _03118_;
  wire [8:0] _03119_;
  wire [9:0] _03120_;
  wire [1:0] _03121_;
  wire [9:0] _03122_;
  wire [33:0] _03123_;
  wire _03124_;
  wire [8:0] _03125_;
  wire [8:0] _03126_;
  wire [8:0] _03127_;
  wire [9:0] _03128_;
  wire [1:0] _03129_;
  wire [9:0] _03130_;
  wire [33:0] _03131_;
  wire _03132_;
  wire [8:0] _03133_;
  wire [8:0] _03134_;
  wire [8:0] _03135_;
  wire [9:0] _03136_;
  wire [1:0] _03137_;
  wire [9:0] _03138_;
  wire [9:0] _03139_;
  wire [9:0] _03140_;
  wire [9:0] _03141_;
  wire [9:0] _03142_;
  wire _03143_;
  wire [3:0] _03144_;
  wire [3:0] _03145_;
  wire [10:0] _03146_;
  wire [33:0] _03147_;
  wire _03148_;
  wire [9:0] _03149_;
  wire [9:0] _03150_;
  wire [9:0] _03151_;
  wire [9:0] _03152_;
  wire [9:0] _03153_;
  wire [9:0] _03154_;
  wire [9:0] _03155_;
  wire [9:0] _03156_;
  wire [9:0] _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire [33:0] _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire [33:0] _03169_;
  wire _03170_;
  wire [3:0] _03171_;
  wire [31:0] _03172_;
  wire [31:0] _03173_;
  wire [31:0] _03174_;
  wire [31:0] _03175_;
  wire [31:0] _03176_;
  wire [31:0] _03177_;
  wire [31:0] _03178_;
  wire [31:0] _03179_;
  wire [31:0] _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire [31:0] _03207_;
  wire [31:0] _03208_;
  wire [31:0] _03209_;
  wire [31:0] _03210_;
  wire [31:0] _03211_;
  wire [31:0] _03212_;
  wire [31:0] _03213_;
  wire [31:0] _03214_;
  wire [31:0] _03215_;
  wire [31:0] _03216_;
  wire [31:0] _03217_;
  wire [31:0] _03218_;
  wire [31:0] _03219_;
  wire [31:0] _03220_;
  wire [31:0] _03221_;
  wire [31:0] _03222_;
  wire [31:0] _03223_;
  wire [31:0] _03224_;
  wire [31:0] _03225_;
  wire [31:0] _03226_;
  wire [1:0] _03227_;
  wire [31:0] _03228_;
  wire [1:0] _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire [31:0] _03233_;
  wire [31:0] _03234_;
  wire [31:0] _03235_;
  wire [31:0] _03236_;
  wire [31:0] _03237_;
  wire [31:0] _03238_;
  wire [31:0] _03239_;
  wire [31:0] _03240_;
  wire [31:0] _03241_;
  wire [31:0] _03242_;
  wire [31:0] _03243_;
  wire [31:0] _03244_;
  wire [31:0] _03245_;
  wire [31:0] _03246_;
  wire [31:0] _03247_;
  wire _03248_;
  wire [31:0] _03249_;
  wire [31:0] _03250_;
  wire [31:0] _03251_;
  wire [31:0] _03252_;
  wire [31:0] _03253_;
  wire [31:0] _03254_;
  wire [31:0] _03255_;
  wire [31:0] _03256_;
  wire [1:0] _03257_;
  wire [31:0] _03258_;
  wire [31:0] _03259_;
  wire [1:0] _03260_;
  wire [1:0] _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire [31:0] _03266_;
  wire [31:0] _03267_;
  wire [31:0] _03268_;
  wire [31:0] _03269_;
  wire [31:0] _03270_;
  wire [31:0] _03271_;
  wire [31:0] _03272_;
  wire [31:0] _03273_;
  wire [31:0] _03274_;
  wire [31:0] _03275_;
  wire [8:0] _03276_;
  wire [31:0] _03277_;
  wire [31:0] _03278_;
  wire [31:0] _03279_;
  wire [31:0] _03280_;
  wire [31:0] _03281_;
  wire [31:0] _03282_;
  wire [31:0] _03283_;
  wire [31:0] _03284_;
  wire [31:0] _03285_;
  wire [31:0] _03286_;
  wire [31:0] _03287_;
  wire [31:0] _03288_;
  wire [31:0] _03289_;
  wire [31:0] _03290_;
  wire _03291_;
  wire [31:0] _03292_;
  wire [1:0] _03293_;
  wire _03294_;
  wire [31:0] _03295_;
  wire [31:0] _03296_;
  wire [31:0] _03297_;
  wire [31:0] _03298_;
  wire [31:0] _03299_;
  wire [31:0] _03300_;
  wire [31:0] _03301_;
  wire [31:0] _03302_;
  wire [31:0] _03303_;
  wire [31:0] _03304_;
  wire [31:0] _03305_;
  wire [31:0] _03306_;
  wire [31:0] _03307_;
  wire [31:0] _03308_;
  wire [31:0] _03309_;
  wire _03310_;
  wire [31:0] _03311_;
  wire [31:0] _03312_;
  wire [31:0] _03313_;
  wire [31:0] _03314_;
  wire [31:0] _03315_;
  wire [31:0] _03316_;
  wire [31:0] _03317_;
  wire [31:0] _03318_;
  wire _03319_;
  wire [31:0] _03320_;
  wire [31:0] _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire [31:0] _03328_;
  wire [31:0] _03329_;
  wire _03330_;
  wire [31:0] _03331_;
  wire [31:0] _03332_;
  wire [31:0] _03333_;
  wire [31:0] _03334_;
  wire _03335_;
  wire [31:0] _03336_;
  wire [31:0] _03337_;
  wire [31:0] _03338_;
  wire [31:0] _03339_;
  wire [31:0] _03340_;
  wire [31:0] _03341_;
  wire [31:0] _03342_;
  wire [31:0] _03343_;
  wire [1:0] _03344_;
  wire [31:0] _03345_;
  wire [31:0] _03346_;
  wire [31:0] _03347_;
  wire [31:0] _03348_;
  wire _03349_;
  wire [31:0] _03350_;
  wire [31:0] _03351_;
  wire [31:0] _03352_;
  wire [31:0] _03353_;
  wire [31:0] _03354_;
  wire [31:0] _03355_;
  wire [31:0] _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire [31:0] _03360_;
  wire [31:0] _03361_;
  wire [3:0] _03362_;
  wire [31:0] _03363_;
  wire [7:0] _03364_;
  wire _03365_;
  wire [31:0] _03366_;
  wire [7:0] _03367_;
  wire _03368_;
  wire [31:0] _03369_;
  wire _03370_;
  wire [3:0] _03371_;
  wire _03372_;
  wire [9:0] _03373_;
  wire [9:0] _03374_;
  wire [3:0] _03375_;
  wire _03376_;
  wire [9:0] _03377_;
  wire [9:0] _03378_;
  wire [3:0] _03379_;
  wire _03380_;
  wire [9:0] _03381_;
  wire [9:0] _03382_;
  wire [3:0] _03383_;
  wire _03384_;
  wire [9:0] _03385_;
  wire [9:0] _03386_;
  wire [3:0] _03387_;
  wire _03388_;
  wire [9:0] _03389_;
  wire [9:0] _03390_;
  wire [3:0] _03391_;
  wire _03392_;
  wire [9:0] _03393_;
  wire [9:0] _03394_;
  wire [3:0] _03395_;
  wire _03396_;
  wire [9:0] _03397_;
  wire [9:0] _03398_;
  wire [3:0] _03399_;
  wire _03400_;
  wire [9:0] _03401_;
  wire [9:0] _03402_;
  wire [3:0] _03403_;
  wire _03404_;
  wire [9:0] _03405_;
  wire [9:0] _03406_;
  wire [3:0] _03407_;
  wire _03408_;
  wire [9:0] _03409_;
  wire [9:0] _03410_;
  wire [3:0] _03411_;
  wire _03412_;
  wire [9:0] _03413_;
  wire [9:0] _03414_;
  wire [3:0] _03415_;
  wire _03416_;
  wire [9:0] _03417_;
  wire [9:0] _03418_;
  wire [3:0] _03419_;
  wire _03420_;
  wire [9:0] _03421_;
  wire [9:0] _03422_;
  wire [3:0] _03423_;
  wire _03424_;
  wire [9:0] _03425_;
  wire [9:0] _03426_;
  wire [3:0] _03427_;
  wire _03428_;
  wire [9:0] _03429_;
  wire [9:0] _03430_;
  wire [3:0] _03431_;
  wire _03432_;
  wire [9:0] _03433_;
  wire [9:0] _03434_;
  wire [3:0] _03435_;
  wire _03436_;
  wire [9:0] _03437_;
  wire [9:0] _03438_;
  wire [3:0] _03439_;
  wire _03440_;
  wire [9:0] _03441_;
  wire [9:0] _03442_;
  wire [3:0] _03443_;
  wire _03444_;
  wire [9:0] _03445_;
  wire [9:0] _03446_;
  wire [3:0] _03447_;
  wire _03448_;
  wire [9:0] _03449_;
  wire [9:0] _03450_;
  wire [3:0] _03451_;
  wire _03452_;
  wire [9:0] _03453_;
  wire [9:0] _03454_;
  wire [3:0] _03455_;
  wire _03456_;
  wire [9:0] _03457_;
  wire [9:0] _03458_;
  wire [3:0] _03459_;
  wire _03460_;
  wire [9:0] _03461_;
  wire [9:0] _03462_;
  wire [3:0] _03463_;
  wire _03464_;
  wire [9:0] _03465_;
  wire [9:0] _03466_;
  wire [3:0] _03467_;
  wire _03468_;
  wire [9:0] _03469_;
  wire [9:0] _03470_;
  wire [3:0] _03471_;
  wire _03472_;
  wire [9:0] _03473_;
  wire [9:0] _03474_;
  wire [3:0] _03475_;
  wire _03476_;
  wire [9:0] _03477_;
  wire [9:0] _03478_;
  wire [3:0] _03479_;
  wire _03480_;
  wire [9:0] _03481_;
  wire [9:0] _03482_;
  wire [3:0] _03483_;
  wire _03484_;
  wire [9:0] _03485_;
  wire [9:0] _03486_;
  wire [3:0] _03487_;
  wire _03488_;
  wire [9:0] _03489_;
  wire [9:0] _03490_;
  wire [3:0] _03491_;
  wire _03492_;
  wire [9:0] _03493_;
  wire [9:0] _03494_;
  wire [3:0] _03495_;
  wire _03496_;
  wire [9:0] _03497_;
  wire [9:0] _03498_;
  wire [3:0] _03499_;
  wire _03500_;
  wire [9:0] _03501_;
  wire [9:0] _03502_;
  wire [3:0] _03503_;
  wire _03504_;
  wire [9:0] _03505_;
  wire [9:0] _03506_;
  wire [3:0] _03507_;
  wire _03508_;
  wire [9:0] _03509_;
  wire [9:0] _03510_;
  wire [3:0] _03511_;
  wire _03512_;
  wire [9:0] _03513_;
  wire [9:0] _03514_;
  wire [3:0] _03515_;
  wire _03516_;
  wire [9:0] _03517_;
  wire [9:0] _03518_;
  wire [3:0] _03519_;
  wire _03520_;
  wire [9:0] _03521_;
  wire [9:0] _03522_;
  wire [3:0] _03523_;
  wire _03524_;
  wire [9:0] _03525_;
  wire [9:0] _03526_;
  wire [3:0] _03527_;
  wire _03528_;
  wire [9:0] _03529_;
  wire [9:0] _03530_;
  wire [3:0] _03531_;
  wire _03532_;
  wire [9:0] _03533_;
  wire [9:0] _03534_;
  wire [3:0] _03535_;
  wire _03536_;
  wire [9:0] _03537_;
  wire [9:0] _03538_;
  wire [3:0] _03539_;
  wire _03540_;
  wire [9:0] _03541_;
  wire [9:0] _03542_;
  wire [3:0] _03543_;
  wire _03544_;
  wire [9:0] _03545_;
  wire [9:0] _03546_;
  wire [3:0] _03547_;
  wire _03548_;
  wire [9:0] _03549_;
  wire [9:0] _03550_;
  wire [3:0] _03551_;
  wire _03552_;
  wire [9:0] _03553_;
  wire [9:0] _03554_;
  wire [3:0] _03555_;
  wire _03556_;
  wire [9:0] _03557_;
  wire [9:0] _03558_;
  wire [3:0] _03559_;
  wire _03560_;
  wire [9:0] _03561_;
  wire [9:0] _03562_;
  wire [3:0] _03563_;
  wire _03564_;
  wire [9:0] _03565_;
  wire [9:0] _03566_;
  wire [3:0] _03567_;
  wire _03568_;
  wire [9:0] _03569_;
  wire [9:0] _03570_;
  wire [3:0] _03571_;
  wire _03572_;
  wire [9:0] _03573_;
  wire [9:0] _03574_;
  wire [3:0] _03575_;
  wire _03576_;
  wire [9:0] _03577_;
  wire [9:0] _03578_;
  wire [3:0] _03579_;
  wire _03580_;
  wire [9:0] _03581_;
  wire [9:0] _03582_;
  wire [3:0] _03583_;
  wire _03584_;
  wire [9:0] _03585_;
  wire [9:0] _03586_;
  wire [3:0] _03587_;
  wire _03588_;
  wire [9:0] _03589_;
  wire [9:0] _03590_;
  wire [3:0] _03591_;
  wire _03592_;
  wire [9:0] _03593_;
  wire [9:0] _03594_;
  wire [3:0] _03595_;
  wire _03596_;
  wire [9:0] _03597_;
  wire [9:0] _03598_;
  wire [3:0] _03599_;
  wire _03600_;
  wire [9:0] _03601_;
  wire [9:0] _03602_;
  wire [3:0] _03603_;
  wire _03604_;
  wire [9:0] _03605_;
  wire [9:0] _03606_;
  wire [3:0] _03607_;
  wire _03608_;
  wire [9:0] _03609_;
  wire [9:0] _03610_;
  wire [3:0] _03611_;
  wire _03612_;
  wire [9:0] _03613_;
  wire [9:0] _03614_;
  wire [3:0] _03615_;
  wire _03616_;
  wire [9:0] _03617_;
  wire [9:0] _03618_;
  wire [3:0] _03619_;
  wire _03620_;
  wire [9:0] _03621_;
  wire [9:0] _03622_;
  wire [3:0] _03623_;
  wire _03624_;
  wire [9:0] _03625_;
  wire [9:0] _03626_;
  wire [3:0] _03627_;
  wire _03628_;
  wire [9:0] _03629_;
  wire [9:0] _03630_;
  wire [3:0] _03631_;
  wire _03632_;
  wire [9:0] _03633_;
  wire [9:0] _03634_;
  wire [3:0] _03635_;
  wire _03636_;
  wire [9:0] _03637_;
  wire [9:0] _03638_;
  wire [3:0] _03639_;
  wire _03640_;
  wire [9:0] _03641_;
  wire [9:0] _03642_;
  wire [3:0] _03643_;
  wire _03644_;
  wire [9:0] _03645_;
  wire [9:0] _03646_;
  wire [3:0] _03647_;
  wire _03648_;
  wire [9:0] _03649_;
  wire [9:0] _03650_;
  wire [3:0] _03651_;
  wire _03652_;
  wire [9:0] _03653_;
  wire [9:0] _03654_;
  wire [3:0] _03655_;
  wire _03656_;
  wire [9:0] _03657_;
  wire [9:0] _03658_;
  wire [3:0] _03659_;
  wire _03660_;
  wire [8:0] _03661_;
  wire [7:0] _03662_;
  wire _03663_;
  wire [8:0] _03664_;
  wire [7:0] _03665_;
  wire _03666_;
  wire [8:0] _03667_;
  wire [7:0] _03668_;
  wire _03669_;
  wire [8:0] _03670_;
  wire [7:0] _03671_;
  wire _03672_;
  wire [8:0] _03673_;
  wire [7:0] _03674_;
  wire _03675_;
  wire [8:0] _03676_;
  wire [7:0] _03677_;
  wire _03678_;
  wire [8:0] _03679_;
  wire [7:0] _03680_;
  wire _03681_;
  wire [8:0] _03682_;
  wire [7:0] _03683_;
  wire _03684_;
  wire [8:0] _03685_;
  wire [8:0] _03686_;
  wire [7:0] _03687_;
  wire _03688_;
  wire [8:0] _03689_;
  wire [8:0] _03690_;
  wire [7:0] _03691_;
  wire _03692_;
  wire [8:0] _03693_;
  wire [8:0] _03694_;
  wire [7:0] _03695_;
  wire _03696_;
  wire [8:0] _03697_;
  wire [8:0] _03698_;
  wire [7:0] _03699_;
  wire _03700_;
  wire [8:0] _03701_;
  wire [7:0] _03702_;
  wire _03703_;
  wire [8:0] _03704_;
  wire [8:0] _03705_;
  wire [7:0] _03706_;
  wire _03707_;
  wire [8:0] _03708_;
  wire [8:0] _03709_;
  wire [7:0] _03710_;
  wire _03711_;
  wire [8:0] _03712_;
  wire [8:0] _03713_;
  wire [7:0] _03714_;
  wire _03715_;
  wire [8:0] _03716_;
  wire [8:0] _03717_;
  wire [7:0] _03718_;
  wire _03719_;
  wire [8:0] _03720_;
  wire [7:0] _03721_;
  wire _03722_;
  wire [8:0] _03723_;
  wire [7:0] _03724_;
  wire _03725_;
  wire [8:0] _03726_;
  wire [7:0] _03727_;
  wire _03728_;
  wire [8:0] _03729_;
  wire [7:0] _03730_;
  wire _03731_;
  wire [8:0] _03732_;
  wire [7:0] _03733_;
  wire _03734_;
  wire [8:0] _03735_;
  wire [7:0] _03736_;
  wire _03737_;
  wire [8:0] _03738_;
  wire [7:0] _03739_;
  wire _03740_;
  wire [8:0] _03741_;
  wire [8:0] _03742_;
  wire [7:0] _03743_;
  wire _03744_;
  wire [8:0] _03745_;
  wire [8:0] _03746_;
  wire [7:0] _03747_;
  wire _03748_;
  wire [8:0] _03749_;
  wire [8:0] _03750_;
  wire [7:0] _03751_;
  wire _03752_;
  wire [8:0] _03753_;
  wire [8:0] _03754_;
  wire [7:0] _03755_;
  wire _03756_;
  wire [8:0] _03757_;
  wire [8:0] _03758_;
  wire [7:0] _03759_;
  wire _03760_;
  wire [8:0] _03761_;
  wire [8:0] _03762_;
  wire [7:0] _03763_;
  wire _03764_;
  wire [8:0] _03765_;
  wire [8:0] _03766_;
  wire [7:0] _03767_;
  wire _03768_;
  wire [8:0] _03769_;
  wire [8:0] _03770_;
  wire [7:0] _03771_;
  wire _03772_;
  wire [8:0] _03773_;
  wire [8:0] _03774_;
  wire [7:0] _03775_;
  wire _03776_;
  wire [8:0] _03777_;
  wire [8:0] _03778_;
  wire [7:0] _03779_;
  wire _03780_;
  wire [8:0] _03781_;
  wire [8:0] _03782_;
  wire [7:0] _03783_;
  wire _03784_;
  wire [8:0] _03785_;
  wire [8:0] _03786_;
  wire [7:0] _03787_;
  wire _03788_;
  wire [8:0] _03789_;
  wire [8:0] _03790_;
  wire [7:0] _03791_;
  wire _03792_;
  wire [8:0] _03793_;
  wire [8:0] _03794_;
  wire [7:0] _03795_;
  wire _03796_;
  wire [8:0] _03797_;
  wire [8:0] _03798_;
  wire [7:0] _03799_;
  wire _03800_;
  wire [8:0] _03801_;
  wire [8:0] _03802_;
  wire [7:0] _03803_;
  wire _03804_;
  wire [8:0] _03805_;
  wire [8:0] _03806_;
  wire [7:0] _03807_;
  wire _03808_;
  wire [8:0] _03809_;
  wire [8:0] _03810_;
  wire [7:0] _03811_;
  wire _03812_;
  wire [8:0] _03813_;
  wire [8:0] _03814_;
  wire [7:0] _03815_;
  wire _03816_;
  wire [8:0] _03817_;
  wire [8:0] _03818_;
  wire [7:0] _03819_;
  wire _03820_;
  wire [8:0] _03821_;
  wire [8:0] _03822_;
  wire [7:0] _03823_;
  wire _03824_;
  wire [8:0] _03825_;
  wire [8:0] _03826_;
  wire [7:0] _03827_;
  wire _03828_;
  wire [8:0] _03829_;
  wire [8:0] _03830_;
  wire [7:0] _03831_;
  wire _03832_;
  wire [8:0] _03833_;
  wire [8:0] _03834_;
  wire [7:0] _03835_;
  wire _03836_;
  wire [8:0] _03837_;
  wire [8:0] _03838_;
  wire [7:0] _03839_;
  wire _03840_;
  wire [8:0] _03841_;
  wire [8:0] _03842_;
  wire [7:0] _03843_;
  wire _03844_;
  wire [8:0] _03845_;
  wire [8:0] _03846_;
  wire [7:0] _03847_;
  wire _03848_;
  wire [8:0] _03849_;
  wire [8:0] _03850_;
  wire [7:0] _03851_;
  wire _03852_;
  wire [8:0] _03853_;
  wire [8:0] _03854_;
  wire [7:0] _03855_;
  wire _03856_;
  wire [8:0] _03857_;
  wire [8:0] _03858_;
  wire [7:0] _03859_;
  wire _03860_;
  wire [8:0] _03861_;
  wire [8:0] _03862_;
  wire [7:0] _03863_;
  wire _03864_;
  wire [8:0] _03865_;
  wire [8:0] _03866_;
  wire [7:0] _03867_;
  wire _03868_;
  wire [8:0] _03869_;
  wire [9:0] _03870_;
  wire [8:0] _03871_;
  wire [8:0] _03872_;
  wire _03873_;
  wire [31:0] _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire [31:0] _24196_;
  wire [31:0] _24197_;
  wire [31:0] _24198_;
  wire [31:0] _24199_;
  wire [31:0] _24200_;
  wire [31:0] _24201_;
  wire [31:0] _24202_;
  wire [31:0] _24203_;
  wire [31:0] _24204_;
  wire [31:0] _24205_;
  wire [31:0] _24206_;
  wire [31:0] _24207_;
  wire [31:0] _24208_;
  wire [31:0] _24209_;
  wire [31:0] _24210_;
  wire [31:0] _24211_;
  wire [31:0] _24212_;
  wire [31:0] _24213_;
  wire [31:0] _24214_;
  wire [32:0] _24215_;
  wire [31:0] _24216_;
  wire [32:0] _24217_;
  wire [32:0] _24218_;
  wire [31:0] _24219_;
  wire [31:0] _24220_;
  wire [32:0] _24221_;
  wire [31:0] _24222_;
  wire [31:0] _24223_;
  wire [31:0] _24224_;
  wire [31:0] _24225_;
  wire [31:0] _24226_;
  wire [32:0] _24227_;
  wire [31:0] _24228_;
  wire [32:0] _24229_;
  wire [32:0] _24230_;
  wire [31:0] _24231_;
  wire [31:0] _24232_;
  wire [32:0] _24233_;
  wire [31:0] _24234_;
  wire [31:0] _24235_;
  wire [31:0] _24236_;
  wire [31:0] _24237_;
  wire [31:0] _24238_;
  wire [31:0] _24239_;
  wire [31:0] _24240_;
  wire [31:0] _24241_;
  wire [31:0] _24242_;
  wire [31:0] _24243_;
  wire [31:0] _24244_;
  wire [31:0] _24245_;
  wire [31:0] _24246_;
  wire [31:0] _24247_;
  wire [31:0] _24248_;
  wire [31:0] _24249_;
  wire [31:0] _24250_;
  wire [31:0] _24251_;
  wire [31:0] _24252_;
  wire [31:0] _24253_;
  wire [31:0] _24254_;
  wire [31:0] _24255_;
  wire [31:0] _24256_;
  wire [31:0] _24257_;
  wire [31:0] _24258_;
  wire [31:0] _24259_;
  wire [31:0] _24260_;
  wire [31:0] _24261_;
  wire [31:0] _24262_;
  wire [31:0] _24263_;
  wire [31:0] _24264_;
  wire [31:0] _24265_;
  wire [31:0] _24266_;
  wire [31:0] _24267_;
  wire [31:0] _24268_;
  wire [31:0] _24269_;
  wire [31:0] _24270_;
  wire [31:0] _24271_;
  wire [31:0] _24272_;
  wire [31:0] _24273_;
  wire [31:0] _24274_;
  wire [31:0] _24275_;
  wire [31:0] _24276_;
  wire [31:0] _24277_;
  wire [31:0] _24278_;
  wire [31:0] _24279_;
  wire [31:0] _24280_;
  wire [31:0] _24281_;
  wire [31:0] _24282_;
  wire [31:0] _24283_;
  wire [31:0] _24284_;
  wire [31:0] _24285_;
  wire [31:0] _24286_;
  wire [31:0] _24287_;
  wire [31:0] _24288_;
  wire [31:0] _24289_;
  wire [31:0] _24290_;
  wire [32:0] _24291_;
  wire [32:0] _24292_;
  wire [31:0] _24293_;
  wire [31:0] _24294_;
  wire [31:0] _24295_;
  wire [31:0] _24296_;
  wire [31:0] _24297_;
  wire [31:0] _24298_;
  wire [31:0] _24299_;
  wire [31:0] _24300_;
  wire [31:0] _24301_;
  wire [31:0] _24302_;
  wire [31:0] _24303_;
  wire [7:0] _24304_;
  wire [7:0] _24305_;
  wire [7:0] _24306_;
  wire [31:0] _24307_;
  wire [31:0] _24308_;
  wire [31:0] _24309_;
  wire [31:0] _24310_;
  wire [31:0] _24311_;
  wire [31:0] _24312_;
  wire [31:0] _24313_;
  wire [31:0] _24314_;
  wire [31:0] _24315_;
  wire [31:0] _24316_;
  wire [31:0] _24317_;
  wire [31:0] _24318_;
  wire [31:0] _24319_;
  wire [31:0] _24320_;
  wire [31:0] _24321_;
  wire [31:0] _24322_;
  wire [31:0] _24323_;
  wire [31:0] _24324_;
  wire [31:0] _24325_;
  wire [31:0] _24326_;
  wire [31:0] _24327_;
  wire [31:0] _24328_;
  wire [31:0] _24329_;
  wire [31:0] _24330_;
  wire [31:0] _24331_;
  wire [31:0] _24332_;
  wire [31:0] _24333_;
  wire [31:0] _24334_;
  wire [31:0] _24335_;
  wire [31:0] _24336_;
  wire [31:0] _24337_;
  wire [31:0] _24338_;
  wire [31:0] _24339_;
  wire [31:0] _24340_;
  wire [31:0] _24341_;
  wire [31:0] _24342_;
  wire [31:0] _24343_;
  wire [31:0] _24344_;
  wire [31:0] _24345_;
  wire [31:0] _24346_;
  wire [31:0] _24347_;
  wire [31:0] _24348_;
  wire [31:0] _24349_;
  wire [31:0] _24350_;
  wire [31:0] _24351_;
  wire [31:0] _24352_;
  wire [31:0] _24353_;
  wire [31:0] _24354_;
  wire [31:0] _24355_;
  wire [31:0] _24356_;
  wire [31:0] _24357_;
  wire [31:0] _24358_;
  wire [31:0] _24359_;
  wire [31:0] _24360_;
  wire [31:0] _24361_;
  wire [31:0] _24362_;
  wire [31:0] _24363_;
  wire [31:0] _24364_;
  wire [31:0] _24365_;
  wire [31:0] _24366_;
  wire [31:0] _24367_;
  wire [31:0] _24368_;
  wire [31:0] _24369_;
  wire [31:0] _24370_;
  wire [31:0] _24371_;
  wire [31:0] _24372_;
  wire [31:0] _24373_;
  wire [31:0] _24374_;
  wire [31:0] _24375_;
  wire [31:0] _24376_;
  wire [31:0] _24377_;
  wire [31:0] _24378_;
  wire [31:0] _24379_;
  wire [31:0] _24380_;
  wire [31:0] _24381_;
  wire [31:0] _24382_;
  wire [31:0] _24383_;
  wire [31:0] _24384_;
  wire [31:0] _24385_;
  wire [31:0] _24386_;
  wire [31:0] _24387_;
  wire [31:0] _24388_;
  wire [31:0] _24389_;
  wire [31:0] _24390_;
  wire [31:0] _24391_;
  wire [31:0] _24392_;
  wire [31:0] _24393_;
  wire [31:0] _24394_;
  wire [31:0] _24395_;
  wire [31:0] _24396_;
  wire [31:0] _24397_;
  wire [31:0] _24398_;
  wire [31:0] _24399_;
  wire [31:0] _24400_;
  wire [31:0] _24401_;
  wire [31:0] _24402_;
  wire [31:0] _24403_;
  wire [31:0] _24404_;
  wire [31:0] _24405_;
  wire [31:0] _24406_;
  wire [7:0] _24407_;
  wire [7:0] _24408_;
  wire [7:0] _24409_;
  wire [31:0] _24410_;
  wire [31:0] _24411_;
  wire [31:0] _24412_;
  wire [31:0] _24413_;
  wire [31:0] _24414_;
  wire [31:0] _24415_;
  wire [31:0] _24416_;
  wire [31:0] _24417_;
  wire [31:0] _24418_;
  wire [31:0] _24419_;
  wire [31:0] _24420_;
  wire [31:0] _24421_;
  wire [31:0] _24422_;
  wire [31:0] _24423_;
  wire [31:0] _24424_;
  wire [31:0] _24425_;
  wire [31:0] _24426_;
  wire [31:0] _24427_;
  wire [31:0] _24428_;
  wire [31:0] _24429_;
  wire [31:0] _24430_;
  wire [31:0] _24431_;
  wire [31:0] _24432_;
  wire [31:0] _24433_;
  wire [31:0] _24434_;
  wire [31:0] _24435_;
  wire [31:0] _24436_;
  wire [31:0] _24437_;
  wire [1:0] _24438_;
  wire [31:0] _24439_;
  wire [31:0] _24440_;
  wire [31:0] _24441_;
  wire [31:0] _24442_;
  wire [31:0] _24443_;
  wire [31:0] _24444_;
  wire [31:0] _24445_;
  wire [31:0] _24446_;
  wire [31:0] _24447_;
  wire [31:0] _24448_;
  wire [32:0] _24449_;
  wire [31:0] _24450_;
  wire [31:0] _24451_;
  wire [31:0] _24452_;
  wire [31:0] _24453_;
  wire [31:0] _24454_;
  wire [31:0] _24455_;
  wire [31:0] _24456_;
  wire [31:0] _24457_;
  wire [31:0] _24458_;
  wire [31:0] _24459_;
  wire [31:0] _24460_;
  wire [31:0] _24461_;
  wire [1:0] _24462_;
  wire [31:0] _24463_;
  wire [32:0] _24464_;
  wire [31:0] _24465_;
  wire [31:0] _24466_;
  wire [31:0] _24467_;
  wire [31:0] _24468_;
  wire [31:0] _24469_;
  wire [31:0] _24470_;
  wire [31:0] _24471_;
  wire [31:0] _24472_;
  wire [31:0] _24473_;
  wire [31:0] _24474_;
  wire [31:0] _24475_;
  wire [31:0] _24476_;
  wire [31:0] _24477_;
  wire [31:0] _24478_;
  wire [31:0] _24479_;
  wire [31:0] _24480_;
  wire [31:0] _24481_;
  wire [31:0] _24482_;
  wire [31:0] _24483_;
  wire [31:0] _24484_;
  wire [31:0] _24485_;
  wire [31:0] _24486_;
  wire [31:0] _24487_;
  wire [31:0] _24488_;
  wire [31:0] _24489_;
  wire [31:0] _24490_;
  wire [31:0] _24491_;
  wire [31:0] _24492_;
  wire [31:0] _24493_;
  wire [31:0] _24494_;
  wire [31:0] _24495_;
  wire [31:0] _24496_;
  wire [31:0] _24497_;
  wire [31:0] _24498_;
  wire [31:0] _24499_;
  wire [31:0] _24500_;
  wire [31:0] _24501_;
  wire [31:0] _24502_;
  wire [31:0] _24503_;
  wire [31:0] _24504_;
  wire [31:0] _24505_;
  wire [31:0] _24506_;
  wire [31:0] _24507_;
  wire [31:0] _24508_;
  wire [31:0] _24509_;
  wire [31:0] _24510_;
  wire [31:0] _24511_;
  wire [31:0] _24512_;
  wire [31:0] _24513_;
  wire [31:0] _24514_;
  wire [31:0] _24515_;
  wire [31:0] _24516_;
  wire [31:0] _24517_;
  wire [31:0] _24518_;
  wire [31:0] _24519_;
  wire [31:0] _24520_;
  wire [31:0] _24521_;
  wire [31:0] _24522_;
  wire [31:0] _24523_;
  wire [31:0] _24524_;
  wire [31:0] _24525_;
  wire [31:0] _24526_;
  wire [31:0] _24527_;
  wire [31:0] _24528_;
  wire [31:0] _24529_;
  wire [31:0] _24530_;
  wire [31:0] _24531_;
  wire [31:0] _24532_;
  wire [31:0] _24533_;
  wire [31:0] _24534_;
  wire [31:0] _24535_;
  wire [31:0] _24536_;
  wire [31:0] _24537_;
  wire [31:0] _24538_;
  wire [31:0] _24539_;
  wire [31:0] _24540_;
  wire [31:0] _24541_;
  wire [31:0] _24542_;
  wire [31:0] _24543_;
  wire [31:0] _24544_;
  wire [31:0] _24545_;
  wire [31:0] _24546_;
  wire [31:0] _24547_;
  wire [31:0] _24548_;
  wire [31:0] _24549_;
  wire [31:0] _24550_;
  wire [31:0] _24551_;
  wire [31:0] _24552_;
  wire [31:0] _24553_;
  wire [31:0] _24554_;
  wire [31:0] _24555_;
  wire [31:0] _24556_;
  wire [31:0] _24557_;
  wire [31:0] _24558_;
  wire [31:0] _24559_;
  wire [31:0] _24560_;
  wire [31:0] _24561_;
  wire [31:0] _24562_;
  wire [31:0] _24563_;
  wire [31:0] _24564_;
  wire [31:0] _24565_;
  wire [31:0] _24566_;
  wire [31:0] _24567_;
  wire [31:0] _24568_;
  wire [31:0] _24569_;
  wire [31:0] _24570_;
  wire [31:0] _24571_;
  wire [31:0] _24572_;
  wire [31:0] _24573_;
  wire [31:0] _24574_;
  wire [31:0] _24575_;
  wire [31:0] _24576_;
  wire [31:0] _24577_;
  wire [31:0] _24578_;
  wire [31:0] _24579_;
  wire [31:0] _24580_;
  wire [31:0] _24581_;
  wire [31:0] _24582_;
  wire [31:0] _24583_;
  wire [31:0] _24584_;
  wire [31:0] _24585_;
  wire [31:0] _24586_;
  wire [31:0] _24587_;
  wire [31:0] _24588_;
  wire [31:0] _24589_;
  wire [31:0] _24590_;
  wire [31:0] _24591_;
  wire [31:0] _24592_;
  wire [31:0] _24593_;
  wire [31:0] _24594_;
  wire [31:0] _24595_;
  wire [31:0] _24596_;
  wire [31:0] _24597_;
  wire [31:0] _24598_;
  wire [31:0] _24599_;
  wire [31:0] _24600_;
  wire [31:0] _24601_;
  wire [31:0] _24602_;
  wire [31:0] _24603_;
  wire [31:0] _24604_;
  wire [31:0] _24605_;
  wire [31:0] _24606_;
  wire [31:0] _24607_;
  wire [31:0] _24608_;
  wire [31:0] _24609_;
  wire [31:0] _24610_;
  wire [31:0] _24611_;
  wire [31:0] _24612_;
  wire [31:0] _24613_;
  wire [31:0] _24614_;
  wire [31:0] _24615_;
  wire [31:0] _24616_;
  wire [31:0] _24617_;
  wire [31:0] _24618_;
  wire [31:0] _24619_;
  wire [31:0] _24620_;
  wire [31:0] _24621_;
  wire [31:0] _24622_;
  wire [31:0] _24623_;
  wire [31:0] _24624_;
  wire [31:0] _24625_;
  wire [31:0] _24626_;
  wire [31:0] _24627_;
  wire [31:0] _24628_;
  wire [31:0] _24629_;
  wire [31:0] _24630_;
  wire [31:0] _24631_;
  wire [31:0] _24632_;
  wire [31:0] _24633_;
  wire [31:0] _24634_;
  wire [31:0] _24635_;
  wire [31:0] _24636_;
  wire [31:0] _24637_;
  wire [31:0] _24638_;
  wire [31:0] _24639_;
  wire [31:0] _24640_;
  wire [31:0] _24641_;
  wire [31:0] _24642_;
  wire [31:0] _24643_;
  wire [31:0] _24644_;
  wire [31:0] _24645_;
  wire [31:0] _24646_;
  wire [31:0] _24647_;
  wire [31:0] _24648_;
  wire [31:0] _24649_;
  wire [31:0] _24650_;
  wire [31:0] _24651_;
  wire [31:0] _24652_;
  wire [31:0] _24653_;
  wire [31:0] _24654_;
  wire [31:0] _24655_;
  wire [31:0] _24656_;
  wire [31:0] _24657_;
  wire [31:0] _24658_;
  wire [31:0] _24659_;
  wire [31:0] _24660_;
  wire _24661_;
  wire [31:0] _24662_;
  wire _24663_;
  wire [31:0] _24664_;
  wire [31:0] _24665_;
  wire [31:0] _24666_;
  wire [31:0] _24667_;
  wire [31:0] _24668_;
  wire [31:0] _24669_;
  wire [31:0] _24670_;
  wire _24671_;
  wire [31:0] _24672_;
  wire [31:0] _24673_;
  wire [31:0] _24674_;
  wire [31:0] _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire [31:0] _24700_;
  wire [31:0] _24701_;
  wire [31:0] _24702_;
  wire _24703_;
  wire [31:0] _24704_;
  wire [31:0] _24705_;
  wire [31:0] _24706_;
  wire [31:0] _24707_;
  wire _24708_;
  wire [31:0] _24709_;
  wire [31:0] _24710_;
  wire [31:0] _24711_;
  wire [31:0] _24712_;
  wire [31:0] _24713_;
  wire _24714_;
  wire [31:0] _24715_;
  wire [31:0] _24716_;
  wire [31:0] _24717_;
  wire [31:0] _24718_;
  wire [31:0] _24719_;
  wire _24720_;
  wire [31:0] _24721_;
  wire [31:0] _24722_;
  wire [31:0] _24723_;
  wire [31:0] _24724_;
  wire [31:0] _24725_;
  wire [31:0] _24726_;
  wire [31:0] _24727_;
  wire [31:0] _24728_;
  wire [31:0] _24729_;
  wire [31:0] _24730_;
  wire [31:0] _24731_;
  wire [31:0] _24732_;
  wire [31:0] _24733_;
  wire [31:0] _24734_;
  wire [31:0] _24735_;
  wire [31:0] _24736_;
  wire [31:0] _24737_;
  wire [31:0] _24738_;
  wire [31:0] _24739_;
  wire [3:0] _24740_;
  wire [31:0] _24741_;
  wire [31:0] _24742_;
  wire [31:0] _24743_;
  wire [31:0] _24744_;
  wire [31:0] _24745_;
  wire [31:0] _24746_;
  wire [31:0] _24747_;
  wire [31:0] _24748_;
  wire [31:0] _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire [31:0] _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire [31:0] _24766_;
  wire [31:0] _24767_;
  wire _24768_;
  wire [31:0] _24769_;
  wire [31:0] _24770_;
  wire _24771_;
  wire [31:0] _24772_;
  wire [31:0] _24773_;
  wire [31:0] _24774_;
  wire [31:0] _24775_;
  wire [31:0] _24776_;
  wire [31:0] _24777_;
  wire [31:0] _24778_;
  wire [31:0] _24779_;
  wire [31:0] _24780_;
  wire [31:0] _24781_;
  wire [31:0] _24782_;
  wire [31:0] _24783_;
  wire [31:0] _24784_;
  wire [31:0] _24785_;
  wire [31:0] _24786_;
  wire [31:0] _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire [32:0] _24792_;
  wire [32:0] _24793_;
  wire [32:0] _24794_;
  wire [32:0] _24795_;
  wire [32:0] _24796_;
  wire [32:0] _24797_;
  wire [32:0] _24798_;
  wire [31:0] _24799_;
  wire [31:0] _24800_;
  wire [31:0] _24801_;
  wire [31:0] _24802_;
  wire [31:0] _24803_;
  wire [31:0] _24804_;
  wire [31:0] _24805_;
  wire [31:0] _24806_;
  wire [31:0] _24807_;
  wire [31:0] _24808_;
  wire [31:0] _24809_;
  wire [31:0] _24810_;
  wire [31:0] _24811_;
  wire [31:0] _24812_;
  wire [31:0] _24813_;
  wire [31:0] _24814_;
  wire [31:0] _24815_;
  wire [31:0] _24816_;
  wire [31:0] _24817_;
  wire [31:0] _24818_;
  wire [31:0] _24819_;
  wire [31:0] _24820_;
  wire [31:0] _24821_;
  wire [31:0] _24822_;
  wire [31:0] _24823_;
  wire [31:0] _24824_;
  wire [31:0] _24825_;
  wire [8:0] _24826_;
  wire [31:0] _24827_;
  wire [1:0] _24828_;
  wire [31:0] _24829_;
  wire [31:0] _24830_;
  wire [31:0] _24831_;
  wire [31:0] _24832_;
  wire [31:0] _24833_;
  wire [31:0] _24834_;
  wire [31:0] _24835_;
  wire [31:0] _24836_;
  wire [31:0] _24837_;
  wire [31:0] _24838_;
  wire [31:0] _24839_;
  wire [31:0] _24840_;
  wire [31:0] _24841_;
  wire [31:0] _24842_;
  wire [31:0] _24843_;
  wire [31:0] _24844_;
  wire [31:0] _24845_;
  wire [31:0] _24846_;
  wire [31:0] _24847_;
  wire [31:0] _24848_;
  wire [31:0] _24849_;
  wire [31:0] _24850_;
  wire [31:0] _24851_;
  wire [31:0] _24852_;
  wire [31:0] _24853_;
  wire [31:0] _24854_;
  wire [1:0] _24855_;
  wire [1:0] _24856_;
  wire [31:0] _24857_;
  wire [31:0] _24858_;
  wire [31:0] _24859_;
  wire [31:0] _24860_;
  wire [8:0] _24861_;
  wire [8:0] _24862_;
  wire [8:0] _24863_;
  wire [9:0] _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire [31:0] _24870_;
  wire [31:0] _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire [31:0] _24877_;
  wire [31:0] _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire [31:0] _24884_;
  wire [31:0] _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire [31:0] _24891_;
  wire [31:0] _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire [31:0] _24898_;
  wire [31:0] _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire [31:0] _24905_;
  wire [31:0] _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire [31:0] _24912_;
  wire [31:0] _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire [31:0] _24919_;
  wire [31:0] _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire [31:0] _24930_;
  wire [31:0] _24931_;
  wire [32:0] _24932_;
  wire [32:0] _24933_;
  wire [32:0] _24934_;
  wire [32:0] _24935_;
  wire [32:0] _24936_;
  wire [32:0] _24937_;
  wire [32:0] _24938_;
  wire [31:0] _24939_;
  wire [31:0] _24940_;
  wire [31:0] _24941_;
  wire [31:0] _24942_;
  wire [31:0] _24943_;
  wire [31:0] _24944_;
  wire [31:0] _24945_;
  wire [31:0] _24946_;
  wire [31:0] _24947_;
  wire [31:0] _24948_;
  wire [31:0] _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire [31:0] _24998_;
  wire [31:0] _24999_;
  wire [31:0] _25000_;
  wire _25001_;
  wire [31:0] _25002_;
  wire [31:0] _25003_;
  wire [31:0] _25004_;
  wire [31:0] _25005_;
  wire [31:0] _25006_;
  wire [31:0] _25007_;
  wire [31:0] _25008_;
  wire [31:0] _25009_;
  wire [31:0] _25010_;
  wire [31:0] _25011_;
  wire [31:0] _25012_;
  wire [31:0] _25013_;
  wire [31:0] _25014_;
  wire [31:0] _25015_;
  wire [31:0] _25016_;
  wire [31:0] _25017_;
  wire [31:0] _25018_;
  wire [31:0] _25019_;
  wire [31:0] _25020_;
  wire [31:0] _25021_;
  wire [31:0] _25022_;
  wire [31:0] _25023_;
  wire [1:0] _25024_;
  wire [31:0] _25025_;
  wire [31:0] _25026_;
  wire [31:0] _25027_;
  wire [31:0] _25028_;
  wire [31:0] _25029_;
  wire [31:0] _25030_;
  wire [1:0] _25031_;
  wire [1:0] _25032_;
  wire [31:0] _25033_;
  wire [31:0] _25034_;
  wire [31:0] _25035_;
  wire [31:0] _25036_;
  wire [31:0] _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire [31:0] _25041_;
  wire [31:0] _25042_;
  wire [31:0] _25043_;
  wire [31:0] _25044_;
  wire [31:0] _25045_;
  wire [31:0] _25046_;
  wire [31:0] _25047_;
  wire [31:0] _25048_;
  wire [31:0] _25049_;
  wire [31:0] _25050_;
  wire [31:0] _25051_;
  wire [31:0] _25052_;
  wire [31:0] _25053_;
  wire [31:0] _25054_;
  wire [31:0] _25055_;
  wire [31:0] _25056_;
  wire [31:0] _25057_;
  wire [31:0] _25058_;
  wire [31:0] _25059_;
  wire [31:0] _25060_;
  wire [31:0] _25061_;
  wire [31:0] _25062_;
  wire [31:0] _25063_;
  wire [31:0] _25064_;
  wire [31:0] _25065_;
  wire [31:0] _25066_;
  wire [31:0] _25067_;
  wire [31:0] _25068_;
  wire [31:0] _25069_;
  wire [31:0] _25070_;
  wire [31:0] _25071_;
  wire [1:0] _25072_;
  wire [1:0] _25073_;
  wire [1:0] _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire [31:0] _25080_;
  wire _25081_;
  wire [3:0] _25082_;
  wire [31:0] _25083_;
  wire [31:0] _25084_;
  wire [31:0] _25085_;
  wire [31:0] _25086_;
  wire [32:0] _25087_;
  wire [32:0] _25088_;
  wire [32:0] _25089_;
  wire [32:0] _25090_;
  wire [32:0] _25091_;
  wire [32:0] _25092_;
  wire [32:0] _25093_;
  wire [32:0] _25094_;
  wire [32:0] _25095_;
  wire [32:0] _25096_;
  wire [32:0] _25097_;
  wire [32:0] _25098_;
  wire [32:0] _25099_;
  wire [32:0] _25100_;
  wire [32:0] _25101_;
  wire [32:0] _25102_;
  wire [31:0] _25103_;
  wire [31:0] _25104_;
  wire [31:0] _25105_;
  wire [31:0] _25106_;
  wire [32:0] _25107_;
  wire [32:0] _25108_;
  wire [32:0] _25109_;
  wire [32:0] _25110_;
  wire [31:0] _25111_;
  wire [31:0] _25112_;
  wire [31:0] _25113_;
  wire [31:0] _25114_;
  wire [31:0] _25115_;
  wire [31:0] _25116_;
  wire [31:0] _25117_;
  wire [31:0] _25118_;
  wire [31:0] _25119_;
  wire [31:0] _25120_;
  wire [31:0] _25121_;
  wire [31:0] _25122_;
  wire [7:0] _25123_;
  wire [31:0] _25124_;
  wire [31:0] _25125_;
  wire [31:0] _25126_;
  wire [31:0] _25127_;
  wire [32:0] _25128_;
  wire [32:0] _25129_;
  wire [32:0] _25130_;
  wire [32:0] _25131_;
  wire [32:0] _25132_;
  wire [32:0] _25133_;
  wire [32:0] _25134_;
  wire [32:0] _25135_;
  wire [32:0] _25136_;
  wire [32:0] _25137_;
  wire [32:0] _25138_;
  wire [32:0] _25139_;
  wire [32:0] _25140_;
  wire [32:0] _25141_;
  wire [32:0] _25142_;
  wire [32:0] _25143_;
  wire [31:0] _25144_;
  wire [31:0] _25145_;
  wire [31:0] _25146_;
  wire [31:0] _25147_;
  wire [32:0] _25148_;
  wire [32:0] _25149_;
  wire [32:0] _25150_;
  wire [32:0] _25151_;
  wire [31:0] _25152_;
  wire [31:0] _25153_;
  wire [31:0] _25154_;
  wire [31:0] _25155_;
  wire [31:0] _25156_;
  wire [31:0] _25157_;
  wire [31:0] _25158_;
  wire [31:0] _25159_;
  wire [31:0] _25160_;
  wire [31:0] _25161_;
  wire [31:0] _25162_;
  wire [31:0] _25163_;
  wire [1:0] _25164_;
  wire [3:0] _25165_;
  wire _25166_;
  wire _25167_;
  wire [7:0] _25168_;
  wire [7:0] _25169_;
  wire [7:0] _25170_;
  wire [7:0] _25171_;
  wire [31:0] _25172_;
  wire [31:0] _25173_;
  wire [31:0] _25174_;
  wire [31:0] _25175_;
  wire [32:0] _25176_;
  wire [32:0] _25177_;
  wire [32:0] _25178_;
  wire [32:0] _25179_;
  wire [32:0] _25180_;
  wire [32:0] _25181_;
  wire [32:0] _25182_;
  wire [32:0] _25183_;
  wire [32:0] _25184_;
  wire [32:0] _25185_;
  wire [32:0] _25186_;
  wire [32:0] _25187_;
  wire [32:0] _25188_;
  wire [32:0] _25189_;
  wire [32:0] _25190_;
  wire [32:0] _25191_;
  wire [31:0] _25192_;
  wire [31:0] _25193_;
  wire [31:0] _25194_;
  wire [31:0] _25195_;
  wire [32:0] _25196_;
  wire [32:0] _25197_;
  wire [32:0] _25198_;
  wire [32:0] _25199_;
  wire [31:0] _25200_;
  wire [31:0] _25201_;
  wire [31:0] _25202_;
  wire [31:0] _25203_;
  wire [31:0] _25204_;
  wire [31:0] _25205_;
  wire [31:0] _25206_;
  wire [31:0] _25207_;
  wire [31:0] _25208_;
  wire [31:0] _25209_;
  wire [31:0] _25210_;
  wire [31:0] _25211_;
  wire [7:0] _25212_;
  wire [31:0] _25213_;
  wire [31:0] _25214_;
  wire [31:0] _25215_;
  wire [31:0] _25216_;
  wire [32:0] _25217_;
  wire [32:0] _25218_;
  wire [32:0] _25219_;
  wire [32:0] _25220_;
  wire [32:0] _25221_;
  wire [32:0] _25222_;
  wire [32:0] _25223_;
  wire [32:0] _25224_;
  wire [32:0] _25225_;
  wire [32:0] _25226_;
  wire [32:0] _25227_;
  wire [32:0] _25228_;
  wire [32:0] _25229_;
  wire [32:0] _25230_;
  wire [32:0] _25231_;
  wire [32:0] _25232_;
  wire [31:0] _25233_;
  wire [31:0] _25234_;
  wire [31:0] _25235_;
  wire [31:0] _25236_;
  wire [32:0] _25237_;
  wire [32:0] _25238_;
  wire [32:0] _25239_;
  wire [32:0] _25240_;
  wire [31:0] _25241_;
  wire [31:0] _25242_;
  wire [31:0] _25243_;
  wire [31:0] _25244_;
  wire [31:0] _25245_;
  wire [31:0] _25246_;
  wire [31:0] _25247_;
  wire [31:0] _25248_;
  wire [31:0] _25249_;
  wire [31:0] _25250_;
  wire [31:0] _25251_;
  wire [31:0] _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire [10:0] _25256_;
  wire [7:0] _25257_;
  wire _25258_;
  wire [31:0] _25259_;
  wire [31:0] _25260_;
  wire [7:0] _25261_;
  wire [31:0] _25262_;
  wire [32:0] _25263_;
  wire [32:0] _25264_;
  wire [31:0] _25265_;
  wire [32:0] _25266_;
  wire [31:0] _25267_;
  wire [2:0] _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire [31:0] _25272_;
  wire [7:0] _25273_;
  wire [31:0] _25274_;
  wire [31:0] _25275_;
  wire [2:0] _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire [31:0] _25282_;
  wire [7:0] _25283_;
  wire [31:0] _25284_;
  wire [31:0] _25285_;
  wire [2:0] _25286_;
  wire _25287_;
  wire _25288_;
  wire [1:0] _25289_;
  wire [3:0] _25290_;
  wire _25291_;
  wire _25292_;
  wire [7:0] _25293_;
  wire _25294_;
  wire [7:0] _25295_;
  wire _25296_;
  wire [7:0] _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire [31:0] _25302_;
  wire [7:0] _25303_;
  wire [31:0] _25304_;
  wire [31:0] _25305_;
  wire [2:0] _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire [31:0] _25312_;
  wire [7:0] _25313_;
  wire [31:0] _25314_;
  wire [31:0] _25315_;
  wire [2:0] _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire [10:0] _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire [31:0] _25330_;
  wire _25331_;
  wire _25332_;
  wire [7:0] _25333_;
  wire [31:0] _25334_;
  wire [31:0] _25335_;
  wire [31:0] _25336_;
  wire [31:0] _25337_;
  wire [32:0] _25338_;
  wire [32:0] _25339_;
  wire [32:0] _25340_;
  wire [32:0] _25341_;
  wire [32:0] _25342_;
  wire [32:0] _25343_;
  wire [32:0] _25344_;
  wire [32:0] _25345_;
  wire [32:0] _25346_;
  wire [32:0] _25347_;
  wire [32:0] _25348_;
  wire [32:0] _25349_;
  wire [32:0] _25350_;
  wire [32:0] _25351_;
  wire [32:0] _25352_;
  wire [32:0] _25353_;
  wire [31:0] _25354_;
  wire [31:0] _25355_;
  wire [31:0] _25356_;
  wire [31:0] _25357_;
  wire [32:0] _25358_;
  wire [32:0] _25359_;
  wire [32:0] _25360_;
  wire [32:0] _25361_;
  wire [31:0] _25362_;
  wire [31:0] _25363_;
  wire [31:0] _25364_;
  wire [31:0] _25365_;
  wire [31:0] _25366_;
  wire [31:0] _25367_;
  wire [31:0] _25368_;
  wire [31:0] _25369_;
  wire [31:0] _25370_;
  wire [31:0] _25371_;
  wire [31:0] _25372_;
  wire [31:0] _25373_;
  wire [3:0] _25374_;
  wire [2:0] _25375_;
  wire [31:0] _25376_;
  wire [31:0] _25377_;
  wire [7:0] _25378_;
  wire _25379_;
  wire [31:0] _25380_;
  wire [31:0] _25381_;
  wire [7:0] _25382_;
  wire [31:0] _25383_;
  wire [32:0] _25384_;
  wire [32:0] _25385_;
  wire [31:0] _25386_;
  wire [32:0] _25387_;
  wire [31:0] _25388_;
  wire [2:0] _25389_;
  wire [3:0] _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire [31:0] _25394_;
  wire [7:0] _25395_;
  wire [31:0] _25396_;
  wire [31:0] _25397_;
  wire [2:0] _25398_;
  wire _25399_;
  wire _25400_;
  wire [2:0] _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire [31:0] _25407_;
  wire _25408_;
  wire [3:0] _25409_;
  wire [31:0] _25410_;
  wire [31:0] _25411_;
  wire [31:0] _25412_;
  wire [31:0] _25413_;
  wire [32:0] _25414_;
  wire [32:0] _25415_;
  wire [32:0] _25416_;
  wire [32:0] _25417_;
  wire [32:0] _25418_;
  wire [32:0] _25419_;
  wire [32:0] _25420_;
  wire [32:0] _25421_;
  wire [32:0] _25422_;
  wire [32:0] _25423_;
  wire [32:0] _25424_;
  wire [32:0] _25425_;
  wire [32:0] _25426_;
  wire [32:0] _25427_;
  wire [32:0] _25428_;
  wire [32:0] _25429_;
  wire [31:0] _25430_;
  wire [31:0] _25431_;
  wire [31:0] _25432_;
  wire [31:0] _25433_;
  wire [32:0] _25434_;
  wire [32:0] _25435_;
  wire [32:0] _25436_;
  wire [32:0] _25437_;
  wire [31:0] _25438_;
  wire [31:0] _25439_;
  wire [31:0] _25440_;
  wire [31:0] _25441_;
  wire [31:0] _25442_;
  wire [31:0] _25443_;
  wire [31:0] _25444_;
  wire [31:0] _25445_;
  wire [31:0] _25446_;
  wire [31:0] _25447_;
  wire [31:0] _25448_;
  wire [31:0] _25449_;
  wire [3:0] _25450_;
  wire [31:0] _25451_;
  wire [31:0] _25452_;
  wire [31:0] _25453_;
  wire [31:0] _25454_;
  wire [32:0] _25455_;
  wire [32:0] _25456_;
  wire [32:0] _25457_;
  wire [32:0] _25458_;
  wire [32:0] _25459_;
  wire [32:0] _25460_;
  wire [32:0] _25461_;
  wire [32:0] _25462_;
  wire [32:0] _25463_;
  wire [32:0] _25464_;
  wire [32:0] _25465_;
  wire [32:0] _25466_;
  wire [32:0] _25467_;
  wire [32:0] _25468_;
  wire [32:0] _25469_;
  wire [32:0] _25470_;
  wire [31:0] _25471_;
  wire [31:0] _25472_;
  wire [31:0] _25473_;
  wire [31:0] _25474_;
  wire [32:0] _25475_;
  wire [32:0] _25476_;
  wire [32:0] _25477_;
  wire [32:0] _25478_;
  wire [31:0] _25479_;
  wire [31:0] _25480_;
  wire [31:0] _25481_;
  wire [31:0] _25482_;
  wire [31:0] _25483_;
  wire [31:0] _25484_;
  wire [31:0] _25485_;
  wire [31:0] _25486_;
  wire [31:0] _25487_;
  wire [31:0] _25488_;
  wire [31:0] _25489_;
  wire [31:0] _25490_;
  wire [3:0] _25491_;
  wire [31:0] _25492_;
  wire [31:0] _25493_;
  wire [31:0] _25494_;
  wire [31:0] _25495_;
  wire [32:0] _25496_;
  wire [32:0] _25497_;
  wire [32:0] _25498_;
  wire [32:0] _25499_;
  wire [32:0] _25500_;
  wire [32:0] _25501_;
  wire [32:0] _25502_;
  wire [32:0] _25503_;
  wire [32:0] _25504_;
  wire [32:0] _25505_;
  wire [32:0] _25506_;
  wire [32:0] _25507_;
  wire [32:0] _25508_;
  wire [32:0] _25509_;
  wire [32:0] _25510_;
  wire [32:0] _25511_;
  wire [31:0] _25512_;
  wire [31:0] _25513_;
  wire [31:0] _25514_;
  wire [31:0] _25515_;
  wire [32:0] _25516_;
  wire [32:0] _25517_;
  wire [32:0] _25518_;
  wire [32:0] _25519_;
  wire [31:0] _25520_;
  wire [31:0] _25521_;
  wire [31:0] _25522_;
  wire [31:0] _25523_;
  wire [31:0] _25524_;
  wire [31:0] _25525_;
  wire [31:0] _25526_;
  wire [31:0] _25527_;
  wire [31:0] _25528_;
  wire [31:0] _25529_;
  wire [31:0] _25530_;
  wire [31:0] _25531_;
  wire [3:0] _25532_;
  wire [31:0] _25533_;
  wire [31:0] _25534_;
  wire [31:0] _25535_;
  wire [31:0] _25536_;
  wire [32:0] _25537_;
  wire [32:0] _25538_;
  wire [32:0] _25539_;
  wire [32:0] _25540_;
  wire [32:0] _25541_;
  wire [32:0] _25542_;
  wire [32:0] _25543_;
  wire [32:0] _25544_;
  wire [32:0] _25545_;
  wire [32:0] _25546_;
  wire [32:0] _25547_;
  wire [32:0] _25548_;
  wire [32:0] _25549_;
  wire [32:0] _25550_;
  wire [32:0] _25551_;
  wire [32:0] _25552_;
  wire [31:0] _25553_;
  wire [31:0] _25554_;
  wire [31:0] _25555_;
  wire [31:0] _25556_;
  wire [32:0] _25557_;
  wire [32:0] _25558_;
  wire [32:0] _25559_;
  wire [32:0] _25560_;
  wire [31:0] _25561_;
  wire [31:0] _25562_;
  wire [31:0] _25563_;
  wire [31:0] _25564_;
  wire [31:0] _25565_;
  wire [31:0] _25566_;
  wire [31:0] _25567_;
  wire [31:0] _25568_;
  wire [31:0] _25569_;
  wire [31:0] _25570_;
  wire [31:0] _25571_;
  wire [31:0] _25572_;
  wire [3:0] _25573_;
  wire [31:0] _25574_;
  wire [31:0] _25575_;
  wire [31:0] _25576_;
  wire [31:0] _25577_;
  wire [32:0] _25578_;
  wire [32:0] _25579_;
  wire [32:0] _25580_;
  wire [32:0] _25581_;
  wire [32:0] _25582_;
  wire [32:0] _25583_;
  wire [32:0] _25584_;
  wire [32:0] _25585_;
  wire [32:0] _25586_;
  wire [32:0] _25587_;
  wire [32:0] _25588_;
  wire [32:0] _25589_;
  wire [32:0] _25590_;
  wire [32:0] _25591_;
  wire [32:0] _25592_;
  wire [32:0] _25593_;
  wire [31:0] _25594_;
  wire [31:0] _25595_;
  wire [31:0] _25596_;
  wire [31:0] _25597_;
  wire [32:0] _25598_;
  wire [32:0] _25599_;
  wire [32:0] _25600_;
  wire [32:0] _25601_;
  wire [31:0] _25602_;
  wire [31:0] _25603_;
  wire [31:0] _25604_;
  wire [31:0] _25605_;
  wire [31:0] _25606_;
  wire [31:0] _25607_;
  wire [31:0] _25608_;
  wire [31:0] _25609_;
  wire [31:0] _25610_;
  wire [31:0] _25611_;
  wire [31:0] _25612_;
  wire [31:0] _25613_;
  wire [3:0] _25614_;
  wire [31:0] _25615_;
  wire [31:0] _25616_;
  wire [31:0] _25617_;
  wire [31:0] _25618_;
  wire [32:0] _25619_;
  wire [32:0] _25620_;
  wire [32:0] _25621_;
  wire [32:0] _25622_;
  wire [32:0] _25623_;
  wire [32:0] _25624_;
  wire [32:0] _25625_;
  wire [32:0] _25626_;
  wire [32:0] _25627_;
  wire [32:0] _25628_;
  wire [32:0] _25629_;
  wire [32:0] _25630_;
  wire [32:0] _25631_;
  wire [32:0] _25632_;
  wire [32:0] _25633_;
  wire [32:0] _25634_;
  wire [31:0] _25635_;
  wire [31:0] _25636_;
  wire [31:0] _25637_;
  wire [31:0] _25638_;
  wire [32:0] _25639_;
  wire [32:0] _25640_;
  wire [32:0] _25641_;
  wire [32:0] _25642_;
  wire [31:0] _25643_;
  wire [31:0] _25644_;
  wire [31:0] _25645_;
  wire [31:0] _25646_;
  wire [31:0] _25647_;
  wire [31:0] _25648_;
  wire [31:0] _25649_;
  wire [31:0] _25650_;
  wire [31:0] _25651_;
  wire [31:0] _25652_;
  wire [31:0] _25653_;
  wire [31:0] _25654_;
  wire [3:0] _25655_;
  wire [31:0] _25656_;
  wire [31:0] _25657_;
  wire [31:0] _25658_;
  wire [31:0] _25659_;
  wire [32:0] _25660_;
  wire [32:0] _25661_;
  wire [32:0] _25662_;
  wire [32:0] _25663_;
  wire [32:0] _25664_;
  wire [32:0] _25665_;
  wire [32:0] _25666_;
  wire [32:0] _25667_;
  wire [32:0] _25668_;
  wire [32:0] _25669_;
  wire [32:0] _25670_;
  wire [32:0] _25671_;
  wire [32:0] _25672_;
  wire [32:0] _25673_;
  wire [32:0] _25674_;
  wire [32:0] _25675_;
  wire [31:0] _25676_;
  wire [31:0] _25677_;
  wire [31:0] _25678_;
  wire [31:0] _25679_;
  wire [32:0] _25680_;
  wire [32:0] _25681_;
  wire [32:0] _25682_;
  wire [32:0] _25683_;
  wire [31:0] _25684_;
  wire [31:0] _25685_;
  wire [31:0] _25686_;
  wire [31:0] _25687_;
  wire [31:0] _25688_;
  wire [31:0] _25689_;
  wire [31:0] _25690_;
  wire [31:0] _25691_;
  wire [31:0] _25692_;
  wire [31:0] _25693_;
  wire [31:0] _25694_;
  wire [31:0] _25695_;
  wire [3:0] _25696_;
  wire [31:0] _25697_;
  wire [31:0] _25698_;
  wire [31:0] _25699_;
  wire [31:0] _25700_;
  wire [32:0] _25701_;
  wire [32:0] _25702_;
  wire [32:0] _25703_;
  wire [32:0] _25704_;
  wire [32:0] _25705_;
  wire [32:0] _25706_;
  wire [32:0] _25707_;
  wire [32:0] _25708_;
  wire [32:0] _25709_;
  wire [32:0] _25710_;
  wire [32:0] _25711_;
  wire [32:0] _25712_;
  wire [32:0] _25713_;
  wire [32:0] _25714_;
  wire [32:0] _25715_;
  wire [32:0] _25716_;
  wire [31:0] _25717_;
  wire [31:0] _25718_;
  wire [31:0] _25719_;
  wire [31:0] _25720_;
  wire [32:0] _25721_;
  wire [32:0] _25722_;
  wire [32:0] _25723_;
  wire [32:0] _25724_;
  wire [31:0] _25725_;
  wire [31:0] _25726_;
  wire [31:0] _25727_;
  wire [31:0] _25728_;
  wire [31:0] _25729_;
  wire [31:0] _25730_;
  wire [31:0] _25731_;
  wire [31:0] _25732_;
  wire [31:0] _25733_;
  wire [31:0] _25734_;
  wire [31:0] _25735_;
  wire [31:0] _25736_;
  wire [3:0] _25737_;
  wire [31:0] _25738_;
  wire [31:0] _25739_;
  wire [31:0] _25740_;
  wire [31:0] _25741_;
  wire [32:0] _25742_;
  wire [32:0] _25743_;
  wire [32:0] _25744_;
  wire [32:0] _25745_;
  wire [32:0] _25746_;
  wire [32:0] _25747_;
  wire [32:0] _25748_;
  wire [32:0] _25749_;
  wire [32:0] _25750_;
  wire [32:0] _25751_;
  wire [32:0] _25752_;
  wire [32:0] _25753_;
  wire [32:0] _25754_;
  wire [32:0] _25755_;
  wire [32:0] _25756_;
  wire [32:0] _25757_;
  wire [31:0] _25758_;
  wire [31:0] _25759_;
  wire [31:0] _25760_;
  wire [31:0] _25761_;
  wire [32:0] _25762_;
  wire [32:0] _25763_;
  wire [32:0] _25764_;
  wire [32:0] _25765_;
  wire [31:0] _25766_;
  wire [31:0] _25767_;
  wire [31:0] _25768_;
  wire [31:0] _25769_;
  wire [31:0] _25770_;
  wire [31:0] _25771_;
  wire [31:0] _25772_;
  wire [31:0] _25773_;
  wire [31:0] _25774_;
  wire [31:0] _25775_;
  wire [31:0] _25776_;
  wire [31:0] _25777_;
  wire [7:0] _25778_;
  wire [31:0] _25779_;
  wire [31:0] _25780_;
  wire [31:0] _25781_;
  wire [31:0] _25782_;
  wire [32:0] _25783_;
  wire [32:0] _25784_;
  wire [32:0] _25785_;
  wire [32:0] _25786_;
  wire [32:0] _25787_;
  wire [32:0] _25788_;
  wire [32:0] _25789_;
  wire [32:0] _25790_;
  wire [32:0] _25791_;
  wire [32:0] _25792_;
  wire [32:0] _25793_;
  wire [32:0] _25794_;
  wire [32:0] _25795_;
  wire [32:0] _25796_;
  wire [32:0] _25797_;
  wire [32:0] _25798_;
  wire [31:0] _25799_;
  wire [31:0] _25800_;
  wire [31:0] _25801_;
  wire [31:0] _25802_;
  wire [32:0] _25803_;
  wire [32:0] _25804_;
  wire [32:0] _25805_;
  wire [32:0] _25806_;
  wire [31:0] _25807_;
  wire [31:0] _25808_;
  wire [31:0] _25809_;
  wire [31:0] _25810_;
  wire [31:0] _25811_;
  wire [31:0] _25812_;
  wire [31:0] _25813_;
  wire [31:0] _25814_;
  wire [31:0] _25815_;
  wire [31:0] _25816_;
  wire [31:0] _25817_;
  wire [31:0] _25818_;
  wire [7:0] _25819_;
  wire [31:0] _25820_;
  wire [31:0] _25821_;
  wire [31:0] _25822_;
  wire [31:0] _25823_;
  wire [32:0] _25824_;
  wire [32:0] _25825_;
  wire [32:0] _25826_;
  wire [32:0] _25827_;
  wire [32:0] _25828_;
  wire [32:0] _25829_;
  wire [32:0] _25830_;
  wire [32:0] _25831_;
  wire [32:0] _25832_;
  wire [32:0] _25833_;
  wire [32:0] _25834_;
  wire [32:0] _25835_;
  wire [32:0] _25836_;
  wire [32:0] _25837_;
  wire [32:0] _25838_;
  wire [32:0] _25839_;
  wire [31:0] _25840_;
  wire [31:0] _25841_;
  wire [31:0] _25842_;
  wire [31:0] _25843_;
  wire [32:0] _25844_;
  wire [32:0] _25845_;
  wire [32:0] _25846_;
  wire [32:0] _25847_;
  wire [31:0] _25848_;
  wire [31:0] _25849_;
  wire [31:0] _25850_;
  wire [31:0] _25851_;
  wire [31:0] _25852_;
  wire [31:0] _25853_;
  wire [31:0] _25854_;
  wire [31:0] _25855_;
  wire [31:0] _25856_;
  wire [31:0] _25857_;
  wire [31:0] _25858_;
  wire [31:0] _25859_;
  wire [7:0] _25860_;
  wire [31:0] _25861_;
  wire [31:0] _25862_;
  wire [31:0] _25863_;
  wire [31:0] _25864_;
  wire [32:0] _25865_;
  wire [32:0] _25866_;
  wire [32:0] _25867_;
  wire [32:0] _25868_;
  wire [32:0] _25869_;
  wire [32:0] _25870_;
  wire [32:0] _25871_;
  wire [32:0] _25872_;
  wire [32:0] _25873_;
  wire [32:0] _25874_;
  wire [32:0] _25875_;
  wire [32:0] _25876_;
  wire [32:0] _25877_;
  wire [32:0] _25878_;
  wire [32:0] _25879_;
  wire [32:0] _25880_;
  wire [31:0] _25881_;
  wire [31:0] _25882_;
  wire [31:0] _25883_;
  wire [31:0] _25884_;
  wire [32:0] _25885_;
  wire [32:0] _25886_;
  wire [32:0] _25887_;
  wire [32:0] _25888_;
  wire [31:0] _25889_;
  wire [31:0] _25890_;
  wire [31:0] _25891_;
  wire [31:0] _25892_;
  wire [31:0] _25893_;
  wire [31:0] _25894_;
  wire [31:0] _25895_;
  wire [31:0] _25896_;
  wire [31:0] _25897_;
  wire [31:0] _25898_;
  wire [31:0] _25899_;
  wire [31:0] _25900_;
  wire [7:0] _25901_;
  wire [31:0] _25902_;
  wire [31:0] _25903_;
  wire [31:0] _25904_;
  wire [31:0] _25905_;
  wire [32:0] _25906_;
  wire [32:0] _25907_;
  wire [32:0] _25908_;
  wire [32:0] _25909_;
  wire [32:0] _25910_;
  wire [32:0] _25911_;
  wire [32:0] _25912_;
  wire [32:0] _25913_;
  wire [32:0] _25914_;
  wire [32:0] _25915_;
  wire [32:0] _25916_;
  wire [32:0] _25917_;
  wire [32:0] _25918_;
  wire [32:0] _25919_;
  wire [32:0] _25920_;
  wire [32:0] _25921_;
  wire [31:0] _25922_;
  wire [31:0] _25923_;
  wire [31:0] _25924_;
  wire [31:0] _25925_;
  wire [32:0] _25926_;
  wire [32:0] _25927_;
  wire [32:0] _25928_;
  wire [32:0] _25929_;
  wire [31:0] _25930_;
  wire [31:0] _25931_;
  wire [31:0] _25932_;
  wire [31:0] _25933_;
  wire [31:0] _25934_;
  wire [31:0] _25935_;
  wire [31:0] _25936_;
  wire [31:0] _25937_;
  wire [31:0] _25938_;
  wire [31:0] _25939_;
  wire [31:0] _25940_;
  wire [31:0] _25941_;
  wire [7:0] _25942_;
  wire [31:0] _25943_;
  wire [31:0] _25944_;
  wire [31:0] _25945_;
  wire [31:0] _25946_;
  wire [32:0] _25947_;
  wire [32:0] _25948_;
  wire [32:0] _25949_;
  wire [32:0] _25950_;
  wire [32:0] _25951_;
  wire [32:0] _25952_;
  wire [32:0] _25953_;
  wire [32:0] _25954_;
  wire [32:0] _25955_;
  wire [32:0] _25956_;
  wire [32:0] _25957_;
  wire [32:0] _25958_;
  wire [32:0] _25959_;
  wire [32:0] _25960_;
  wire [32:0] _25961_;
  wire [32:0] _25962_;
  wire [31:0] _25963_;
  wire [31:0] _25964_;
  wire [31:0] _25965_;
  wire [31:0] _25966_;
  wire [32:0] _25967_;
  wire [32:0] _25968_;
  wire [32:0] _25969_;
  wire [32:0] _25970_;
  wire [31:0] _25971_;
  wire [31:0] _25972_;
  wire [31:0] _25973_;
  wire [31:0] _25974_;
  wire [31:0] _25975_;
  wire [31:0] _25976_;
  wire [31:0] _25977_;
  wire [31:0] _25978_;
  wire [31:0] _25979_;
  wire [31:0] _25980_;
  wire [31:0] _25981_;
  wire [31:0] _25982_;
  wire [7:0] _25983_;
  wire [31:0] _25984_;
  wire [31:0] _25985_;
  wire [31:0] _25986_;
  wire [31:0] _25987_;
  wire [32:0] _25988_;
  wire [32:0] _25989_;
  wire [32:0] _25990_;
  wire [32:0] _25991_;
  wire [32:0] _25992_;
  wire [32:0] _25993_;
  wire [32:0] _25994_;
  wire [32:0] _25995_;
  wire [32:0] _25996_;
  wire [32:0] _25997_;
  wire [32:0] _25998_;
  wire [32:0] _25999_;
  wire [32:0] _26000_;
  wire [32:0] _26001_;
  wire [32:0] _26002_;
  wire [32:0] _26003_;
  wire [31:0] _26004_;
  wire [31:0] _26005_;
  wire [31:0] _26006_;
  wire [31:0] _26007_;
  wire [32:0] _26008_;
  wire [32:0] _26009_;
  wire [32:0] _26010_;
  wire [32:0] _26011_;
  wire [31:0] _26012_;
  wire [31:0] _26013_;
  wire [31:0] _26014_;
  wire [31:0] _26015_;
  wire [31:0] _26016_;
  wire [31:0] _26017_;
  wire [31:0] _26018_;
  wire [31:0] _26019_;
  wire [31:0] _26020_;
  wire [31:0] _26021_;
  wire [31:0] _26022_;
  wire [31:0] _26023_;
  wire [7:0] _26024_;
  wire [31:0] _26025_;
  wire [31:0] _26026_;
  wire [31:0] _26027_;
  wire [31:0] _26028_;
  wire [32:0] _26029_;
  wire [32:0] _26030_;
  wire [32:0] _26031_;
  wire [32:0] _26032_;
  wire [32:0] _26033_;
  wire [32:0] _26034_;
  wire [32:0] _26035_;
  wire [32:0] _26036_;
  wire [32:0] _26037_;
  wire [32:0] _26038_;
  wire [32:0] _26039_;
  wire [32:0] _26040_;
  wire [32:0] _26041_;
  wire [32:0] _26042_;
  wire [32:0] _26043_;
  wire [32:0] _26044_;
  wire [31:0] _26045_;
  wire [31:0] _26046_;
  wire [31:0] _26047_;
  wire [31:0] _26048_;
  wire [32:0] _26049_;
  wire [32:0] _26050_;
  wire [32:0] _26051_;
  wire [32:0] _26052_;
  wire [31:0] _26053_;
  wire [31:0] _26054_;
  wire [31:0] _26055_;
  wire [31:0] _26056_;
  wire [31:0] _26057_;
  wire [31:0] _26058_;
  wire [31:0] _26059_;
  wire [31:0] _26060_;
  wire [31:0] _26061_;
  wire [31:0] _26062_;
  wire [31:0] _26063_;
  wire [31:0] _26064_;
  wire [7:0] _26065_;
  wire [31:0] _26066_;
  wire [31:0] _26067_;
  wire [31:0] _26068_;
  wire [31:0] _26069_;
  wire [32:0] _26070_;
  wire [32:0] _26071_;
  wire [32:0] _26072_;
  wire [32:0] _26073_;
  wire [32:0] _26074_;
  wire [32:0] _26075_;
  wire [32:0] _26076_;
  wire [32:0] _26077_;
  wire [32:0] _26078_;
  wire [32:0] _26079_;
  wire [32:0] _26080_;
  wire [32:0] _26081_;
  wire [32:0] _26082_;
  wire [32:0] _26083_;
  wire [32:0] _26084_;
  wire [32:0] _26085_;
  wire [31:0] _26086_;
  wire [31:0] _26087_;
  wire [31:0] _26088_;
  wire [31:0] _26089_;
  wire [32:0] _26090_;
  wire [32:0] _26091_;
  wire [32:0] _26092_;
  wire [32:0] _26093_;
  wire [31:0] _26094_;
  wire [31:0] _26095_;
  wire [31:0] _26096_;
  wire [31:0] _26097_;
  wire [31:0] _26098_;
  wire [31:0] _26099_;
  wire [31:0] _26100_;
  wire [31:0] _26101_;
  wire [31:0] _26102_;
  wire [31:0] _26103_;
  wire [31:0] _26104_;
  wire [31:0] _26105_;
  wire [7:0] _26106_;
  wire [31:0] _26107_;
  wire [31:0] _26108_;
  wire [31:0] _26109_;
  wire [31:0] _26110_;
  wire [32:0] _26111_;
  wire [32:0] _26112_;
  wire [32:0] _26113_;
  wire [32:0] _26114_;
  wire [32:0] _26115_;
  wire [32:0] _26116_;
  wire [32:0] _26117_;
  wire [32:0] _26118_;
  wire [32:0] _26119_;
  wire [32:0] _26120_;
  wire [32:0] _26121_;
  wire [32:0] _26122_;
  wire [32:0] _26123_;
  wire [32:0] _26124_;
  wire [32:0] _26125_;
  wire [32:0] _26126_;
  wire [31:0] _26127_;
  wire [31:0] _26128_;
  wire [31:0] _26129_;
  wire [31:0] _26130_;
  wire [32:0] _26131_;
  wire [32:0] _26132_;
  wire [32:0] _26133_;
  wire [32:0] _26134_;
  wire [31:0] _26135_;
  wire [31:0] _26136_;
  wire [31:0] _26137_;
  wire [31:0] _26138_;
  wire [31:0] _26139_;
  wire [31:0] _26140_;
  wire [31:0] _26141_;
  wire [31:0] _26142_;
  wire [31:0] _26143_;
  wire [31:0] _26144_;
  wire [31:0] _26145_;
  wire [31:0] _26146_;
  wire [3:0] _26147_;
  wire _26148_;
  wire _26149_;
  wire [7:0] _26150_;
  wire [7:0] _26151_;
  wire [7:0] _26152_;
  wire [7:0] _26153_;
  wire [31:0] _26154_;
  wire [31:0] _26155_;
  wire [31:0] _26156_;
  wire [31:0] _26157_;
  wire [32:0] _26158_;
  wire [32:0] _26159_;
  wire [32:0] _26160_;
  wire [32:0] _26161_;
  wire [32:0] _26162_;
  wire [32:0] _26163_;
  wire [32:0] _26164_;
  wire [32:0] _26165_;
  wire [32:0] _26166_;
  wire [32:0] _26167_;
  wire [32:0] _26168_;
  wire [32:0] _26169_;
  wire [32:0] _26170_;
  wire [32:0] _26171_;
  wire [32:0] _26172_;
  wire [32:0] _26173_;
  wire [31:0] _26174_;
  wire [31:0] _26175_;
  wire [31:0] _26176_;
  wire [31:0] _26177_;
  wire [32:0] _26178_;
  wire [32:0] _26179_;
  wire [32:0] _26180_;
  wire [32:0] _26181_;
  wire [31:0] _26182_;
  wire [31:0] _26183_;
  wire [31:0] _26184_;
  wire [31:0] _26185_;
  wire [31:0] _26186_;
  wire [31:0] _26187_;
  wire [31:0] _26188_;
  wire [31:0] _26189_;
  wire [31:0] _26190_;
  wire [31:0] _26191_;
  wire [31:0] _26192_;
  wire [31:0] _26193_;
  wire [7:0] _26194_;
  wire [31:0] _26195_;
  wire [31:0] _26196_;
  wire [31:0] _26197_;
  wire [31:0] _26198_;
  wire [32:0] _26199_;
  wire [32:0] _26200_;
  wire [32:0] _26201_;
  wire [32:0] _26202_;
  wire [32:0] _26203_;
  wire [32:0] _26204_;
  wire [32:0] _26205_;
  wire [32:0] _26206_;
  wire [32:0] _26207_;
  wire [32:0] _26208_;
  wire [32:0] _26209_;
  wire [32:0] _26210_;
  wire [32:0] _26211_;
  wire [32:0] _26212_;
  wire [32:0] _26213_;
  wire [32:0] _26214_;
  wire [31:0] _26215_;
  wire [31:0] _26216_;
  wire [31:0] _26217_;
  wire [31:0] _26218_;
  wire [32:0] _26219_;
  wire [32:0] _26220_;
  wire [32:0] _26221_;
  wire [32:0] _26222_;
  wire [31:0] _26223_;
  wire [31:0] _26224_;
  wire [31:0] _26225_;
  wire [31:0] _26226_;
  wire [31:0] _26227_;
  wire [31:0] _26228_;
  wire [31:0] _26229_;
  wire [31:0] _26230_;
  wire [31:0] _26231_;
  wire [31:0] _26232_;
  wire [31:0] _26233_;
  wire [31:0] _26234_;
  wire [8:0] _26235_;
  wire [1:0] _26236_;
  wire [1:0] _26237_;
  wire [5:0] _26238_;
  wire [7:0] _26239_;
  wire _26240_;
  wire [31:0] _26241_;
  wire [31:0] _26242_;
  wire [7:0] _26243_;
  wire [31:0] _26244_;
  wire [32:0] _26245_;
  wire [32:0] _26246_;
  wire [31:0] _26247_;
  wire [32:0] _26248_;
  wire [31:0] _26249_;
  wire [2:0] _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire [31:0] _26254_;
  wire [7:0] _26255_;
  wire [31:0] _26256_;
  wire [31:0] _26257_;
  wire [2:0] _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire [31:0] _26264_;
  wire [7:0] _26265_;
  wire [31:0] _26266_;
  wire [31:0] _26267_;
  wire [2:0] _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire [31:0] _26274_;
  wire [7:0] _26275_;
  wire [31:0] _26276_;
  wire [31:0] _26277_;
  wire [2:0] _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire [31:0] _26284_;
  wire [7:0] _26285_;
  wire [31:0] _26286_;
  wire [31:0] _26287_;
  wire [2:0] _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire [31:0] _26294_;
  wire [7:0] _26295_;
  wire [31:0] _26296_;
  wire [31:0] _26297_;
  wire [2:0] _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire [31:0] _26304_;
  wire [7:0] _26305_;
  wire [31:0] _26306_;
  wire [31:0] _26307_;
  wire [2:0] _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire [31:0] _26314_;
  wire [7:0] _26315_;
  wire [31:0] _26316_;
  wire [31:0] _26317_;
  wire [2:0] _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire [31:0] _26324_;
  wire [7:0] _26325_;
  wire [31:0] _26326_;
  wire [31:0] _26327_;
  wire [2:0] _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire [31:0] _26334_;
  wire [7:0] _26335_;
  wire [31:0] _26336_;
  wire [31:0] _26337_;
  wire [2:0] _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire [31:0] _26344_;
  wire [7:0] _26345_;
  wire [31:0] _26346_;
  wire [31:0] _26347_;
  wire [2:0] _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire [31:0] _26354_;
  wire [7:0] _26355_;
  wire [31:0] _26356_;
  wire [31:0] _26357_;
  wire [2:0] _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire [31:0] _26364_;
  wire [7:0] _26365_;
  wire [31:0] _26366_;
  wire [31:0] _26367_;
  wire [2:0] _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire [31:0] _26374_;
  wire [7:0] _26375_;
  wire [31:0] _26376_;
  wire [31:0] _26377_;
  wire [2:0] _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire [31:0] _26384_;
  wire [7:0] _26385_;
  wire [31:0] _26386_;
  wire [31:0] _26387_;
  wire [2:0] _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire [31:0] _26394_;
  wire [7:0] _26395_;
  wire [31:0] _26396_;
  wire [31:0] _26397_;
  wire [2:0] _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire [31:0] _26404_;
  wire [7:0] _26405_;
  wire [31:0] _26406_;
  wire [31:0] _26407_;
  wire [2:0] _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire [31:0] _26414_;
  wire [7:0] _26415_;
  wire [31:0] _26416_;
  wire [31:0] _26417_;
  wire [2:0] _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire [31:0] _26424_;
  wire [7:0] _26425_;
  wire [31:0] _26426_;
  wire [31:0] _26427_;
  wire [2:0] _26428_;
  wire _26429_;
  wire _26430_;
  wire [3:0] _26431_;
  wire _26432_;
  wire _26433_;
  wire [7:0] _26434_;
  wire _26435_;
  wire [7:0] _26436_;
  wire _26437_;
  wire [7:0] _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire [31:0] _26443_;
  wire [7:0] _26444_;
  wire [31:0] _26445_;
  wire [31:0] _26446_;
  wire [2:0] _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire [31:0] _26453_;
  wire [7:0] _26454_;
  wire [31:0] _26455_;
  wire [31:0] _26456_;
  wire [2:0] _26457_;
  wire _26458_;
  wire _26459_;
  wire [8:0] _26460_;
  wire [1:0] _26461_;
  wire [1:0] _26462_;
  wire [5:0] _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire [7:0] _26470_;
  wire [7:0] _26471_;
  wire [8:0] _26472_;
  wire [8:0] _26473_;
  wire [7:0] _26474_;
  wire [7:0] _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire [3:0] _26482_;
  wire [3:0] _26483_;
  wire [7:0] _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire [3:0] _26491_;
  wire [3:0] _26492_;
  wire [7:0] _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire [3:0] _26500_;
  wire [3:0] _26501_;
  wire [7:0] _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire [3:0] _26509_;
  wire [3:0] _26510_;
  wire [7:0] _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire [3:0] _26518_;
  wire [3:0] _26519_;
  wire [7:0] _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire [3:0] _26527_;
  wire [3:0] _26528_;
  wire [7:0] _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire [3:0] _26536_;
  wire [3:0] _26537_;
  wire [7:0] _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire [3:0] _26545_;
  wire [3:0] _26546_;
  wire [7:0] _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire [3:0] _26560_;
  wire [3:0] _26561_;
  wire [3:0] _26562_;
  wire [3:0] _26563_;
  wire [7:0] _26564_;
  wire [7:0] _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire [5:0] _26578_;
  wire [5:0] _26579_;
  wire [7:0] _26580_;
  wire [7:0] _26581_;
  wire [31:0] _26582_;
  wire [31:0] _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire [31:0] _26602_;
  wire [31:0] _26603_;
  wire [31:0] _26604_;
  wire [31:0] _26605_;
  wire [31:0] _26606_;
  wire [31:0] _26607_;
  wire [31:0] _26608_;
  wire [31:0] _26609_;
  wire [31:0] _26610_;
  wire _26611_;
  wire _26612_;
  wire [31:0] _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire [31:0] _26630_;
  wire [31:0] _26631_;
  wire [5:0] _26632_;
  wire [5:0] _26633_;
  wire [31:0] _26634_;
  wire [31:0] _26635_;
  wire [32:0] _26636_;
  wire [32:0] _26637_;
  wire [31:0] _26638_;
  wire [31:0] _26639_;
  wire [33:0] _26640_;
  wire [33:0] _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire [8:0] _26655_;
  wire [8:0] _26656_;
  wire _26657_;
  wire _26658_;
  wire [7:0] _26659_;
  wire [8:0] _26660_;
  wire [33:0] _26661_;
  wire [33:0] _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire [8:0] _26676_;
  wire [8:0] _26677_;
  wire _26678_;
  wire _26679_;
  wire [7:0] _26680_;
  wire [8:0] _26681_;
  wire [33:0] _26682_;
  wire [33:0] _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire [8:0] _26697_;
  wire [8:0] _26698_;
  wire _26699_;
  wire _26700_;
  wire [7:0] _26701_;
  wire [8:0] _26702_;
  wire _26703_;
  wire _26704_;
  wire [31:0] _26705_;
  wire [33:0] _26706_;
  wire [33:0] _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire [8:0] _26721_;
  wire [8:0] _26722_;
  wire _26723_;
  wire _26724_;
  wire [7:0] _26725_;
  wire [8:0] _26726_;
  wire _26727_;
  wire _26728_;
  wire [7:0] _26729_;
  wire [8:0] _26730_;
  wire [8:0] _26731_;
  wire _26732_;
  wire _26733_;
  wire [7:0] _26734_;
  wire [8:0] _26735_;
  wire [8:0] _26736_;
  wire _26737_;
  wire _26738_;
  wire [7:0] _26739_;
  wire [8:0] _26740_;
  wire [8:0] _26741_;
  wire _26742_;
  wire _26743_;
  wire [7:0] _26744_;
  wire [8:0] _26745_;
  wire [8:0] _26746_;
  wire _26747_;
  wire _26748_;
  wire [7:0] _26749_;
  wire [8:0] _26750_;
  wire [8:0] _26751_;
  wire _26752_;
  wire _26753_;
  wire [7:0] _26754_;
  wire [8:0] _26755_;
  wire [8:0] _26756_;
  wire _26757_;
  wire _26758_;
  wire [7:0] _26759_;
  wire [8:0] _26760_;
  wire [8:0] _26761_;
  wire _26762_;
  wire _26763_;
  wire [7:0] _26764_;
  wire [8:0] _26765_;
  wire [8:0] _26766_;
  wire [1:0] _26767_;
  wire [1:0] _26768_;
  wire [1:0] _26769_;
  wire [8:0] _26770_;
  wire [8:0] _26771_;
  wire [8:0] _26772_;
  wire [8:0] _26773_;
  wire [8:0] _26774_;
  wire [8:0] _26775_;
  wire _26776_;
  wire _26777_;
  wire [33:0] _26778_;
  wire [33:0] _26779_;
  wire [9:0] _26780_;
  wire [9:0] _26781_;
  wire [9:0] _26782_;
  wire _26783_;
  wire _26784_;
  wire [7:0] _26785_;
  wire [8:0] _26786_;
  wire [8:0] _26787_;
  wire [1:0] _26788_;
  wire [1:0] _26789_;
  wire [1:0] _26790_;
  wire [8:0] _26791_;
  wire [8:0] _26792_;
  wire [8:0] _26793_;
  wire [8:0] _26794_;
  wire [8:0] _26795_;
  wire [8:0] _26796_;
  wire _26797_;
  wire _26798_;
  wire [33:0] _26799_;
  wire [33:0] _26800_;
  wire [9:0] _26801_;
  wire [9:0] _26802_;
  wire [9:0] _26803_;
  wire _26804_;
  wire _26805_;
  wire [7:0] _26806_;
  wire [8:0] _26807_;
  wire [8:0] _26808_;
  wire [1:0] _26809_;
  wire [1:0] _26810_;
  wire [1:0] _26811_;
  wire [8:0] _26812_;
  wire [8:0] _26813_;
  wire [8:0] _26814_;
  wire [8:0] _26815_;
  wire [8:0] _26816_;
  wire [8:0] _26817_;
  wire _26818_;
  wire _26819_;
  wire [33:0] _26820_;
  wire [33:0] _26821_;
  wire [9:0] _26822_;
  wire [9:0] _26823_;
  wire [9:0] _26824_;
  wire _26825_;
  wire _26826_;
  wire [7:0] _26827_;
  wire [8:0] _26828_;
  wire [8:0] _26829_;
  wire [1:0] _26830_;
  wire [1:0] _26831_;
  wire [1:0] _26832_;
  wire [8:0] _26833_;
  wire [8:0] _26834_;
  wire [8:0] _26835_;
  wire [8:0] _26836_;
  wire [8:0] _26837_;
  wire [8:0] _26838_;
  wire _26839_;
  wire _26840_;
  wire [33:0] _26841_;
  wire [33:0] _26842_;
  wire [9:0] _26843_;
  wire [9:0] _26844_;
  wire [9:0] _26845_;
  wire _26846_;
  wire _26847_;
  wire [7:0] _26848_;
  wire [8:0] _26849_;
  wire [8:0] _26850_;
  wire _26851_;
  wire _26852_;
  wire [7:0] _26853_;
  wire [8:0] _26854_;
  wire [8:0] _26855_;
  wire _26856_;
  wire _26857_;
  wire [7:0] _26858_;
  wire [8:0] _26859_;
  wire [8:0] _26860_;
  wire _26861_;
  wire _26862_;
  wire [7:0] _26863_;
  wire [8:0] _26864_;
  wire [8:0] _26865_;
  wire _26866_;
  wire _26867_;
  wire [7:0] _26868_;
  wire [8:0] _26869_;
  wire [8:0] _26870_;
  wire _26871_;
  wire _26872_;
  wire [7:0] _26873_;
  wire [8:0] _26874_;
  wire [8:0] _26875_;
  wire _26876_;
  wire _26877_;
  wire [7:0] _26878_;
  wire [8:0] _26879_;
  wire [8:0] _26880_;
  wire _26881_;
  wire _26882_;
  wire [7:0] _26883_;
  wire [8:0] _26884_;
  wire [8:0] _26885_;
  wire _26886_;
  wire _26887_;
  wire [7:0] _26888_;
  wire [8:0] _26889_;
  wire [8:0] _26890_;
  wire [1:0] _26891_;
  wire [1:0] _26892_;
  wire [1:0] _26893_;
  wire [8:0] _26894_;
  wire [8:0] _26895_;
  wire [8:0] _26896_;
  wire [8:0] _26897_;
  wire [8:0] _26898_;
  wire [8:0] _26899_;
  wire _26900_;
  wire _26901_;
  wire [33:0] _26902_;
  wire [33:0] _26903_;
  wire [9:0] _26904_;
  wire [9:0] _26905_;
  wire [9:0] _26906_;
  wire _26907_;
  wire _26908_;
  wire [7:0] _26909_;
  wire [8:0] _26910_;
  wire [8:0] _26911_;
  wire [1:0] _26912_;
  wire [1:0] _26913_;
  wire [1:0] _26914_;
  wire [8:0] _26915_;
  wire [8:0] _26916_;
  wire [8:0] _26917_;
  wire [8:0] _26918_;
  wire [8:0] _26919_;
  wire [8:0] _26920_;
  wire _26921_;
  wire _26922_;
  wire [33:0] _26923_;
  wire [33:0] _26924_;
  wire [9:0] _26925_;
  wire [9:0] _26926_;
  wire [9:0] _26927_;
  wire _26928_;
  wire _26929_;
  wire [7:0] _26930_;
  wire [8:0] _26931_;
  wire [8:0] _26932_;
  wire [1:0] _26933_;
  wire [1:0] _26934_;
  wire [1:0] _26935_;
  wire [8:0] _26936_;
  wire [8:0] _26937_;
  wire [8:0] _26938_;
  wire [8:0] _26939_;
  wire [8:0] _26940_;
  wire [8:0] _26941_;
  wire _26942_;
  wire _26943_;
  wire [33:0] _26944_;
  wire [33:0] _26945_;
  wire [9:0] _26946_;
  wire [9:0] _26947_;
  wire [9:0] _26948_;
  wire _26949_;
  wire _26950_;
  wire [7:0] _26951_;
  wire [8:0] _26952_;
  wire [8:0] _26953_;
  wire [1:0] _26954_;
  wire [1:0] _26955_;
  wire [1:0] _26956_;
  wire [8:0] _26957_;
  wire [8:0] _26958_;
  wire [8:0] _26959_;
  wire [8:0] _26960_;
  wire [8:0] _26961_;
  wire [8:0] _26962_;
  wire _26963_;
  wire _26964_;
  wire [33:0] _26965_;
  wire [33:0] _26966_;
  wire [9:0] _26967_;
  wire [9:0] _26968_;
  wire [9:0] _26969_;
  wire _26970_;
  wire _26971_;
  wire [7:0] _26972_;
  wire [8:0] _26973_;
  wire [8:0] _26974_;
  wire _26975_;
  wire _26976_;
  wire [7:0] _26977_;
  wire [8:0] _26978_;
  wire [8:0] _26979_;
  wire _26980_;
  wire _26981_;
  wire [7:0] _26982_;
  wire [8:0] _26983_;
  wire [8:0] _26984_;
  wire _26985_;
  wire _26986_;
  wire [7:0] _26987_;
  wire [8:0] _26988_;
  wire [8:0] _26989_;
  wire _26990_;
  wire _26991_;
  wire [7:0] _26992_;
  wire [8:0] _26993_;
  wire [8:0] _26994_;
  wire _26995_;
  wire _26996_;
  wire [33:0] _26997_;
  wire [33:0] _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire [7:0] _27002_;
  wire [7:0] _27003_;
  wire [8:0] _27004_;
  wire [8:0] _27005_;
  wire [8:0] _27006_;
  wire [8:0] _27007_;
  wire [8:0] _27008_;
  wire _27009_;
  wire _27010_;
  wire [33:0] _27011_;
  wire [33:0] _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire [7:0] _27016_;
  wire [7:0] _27017_;
  wire [8:0] _27018_;
  wire [8:0] _27019_;
  wire [8:0] _27020_;
  wire [8:0] _27021_;
  wire [8:0] _27022_;
  wire _27023_;
  wire _27024_;
  wire [33:0] _27025_;
  wire [33:0] _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire [7:0] _27030_;
  wire [7:0] _27031_;
  wire [8:0] _27032_;
  wire [8:0] _27033_;
  wire [8:0] _27034_;
  wire [8:0] _27035_;
  wire [8:0] _27036_;
  wire _27037_;
  wire _27038_;
  wire [33:0] _27039_;
  wire [33:0] _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire [7:0] _27044_;
  wire [7:0] _27045_;
  wire [8:0] _27046_;
  wire [8:0] _27047_;
  wire [8:0] _27048_;
  wire [8:0] _27049_;
  wire [8:0] _27050_;
  wire _27051_;
  wire _27052_;
  wire [33:0] _27053_;
  wire [33:0] _27054_;
  wire [1:0] _27055_;
  wire [1:0] _27056_;
  wire [1:0] _27057_;
  wire [8:0] _27058_;
  wire [8:0] _27059_;
  wire [8:0] _27060_;
  wire [8:0] _27061_;
  wire [8:0] _27062_;
  wire [8:0] _27063_;
  wire _27064_;
  wire _27065_;
  wire [33:0] _27066_;
  wire [33:0] _27067_;
  wire [9:0] _27068_;
  wire [9:0] _27069_;
  wire [9:0] _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire [7:0] _27074_;
  wire [7:0] _27075_;
  wire [8:0] _27076_;
  wire [8:0] _27077_;
  wire [8:0] _27078_;
  wire [8:0] _27079_;
  wire [8:0] _27080_;
  wire _27081_;
  wire _27082_;
  wire [33:0] _27083_;
  wire [33:0] _27084_;
  wire [1:0] _27085_;
  wire [1:0] _27086_;
  wire [1:0] _27087_;
  wire [8:0] _27088_;
  wire [8:0] _27089_;
  wire [8:0] _27090_;
  wire [8:0] _27091_;
  wire [8:0] _27092_;
  wire [8:0] _27093_;
  wire _27094_;
  wire _27095_;
  wire [33:0] _27096_;
  wire [33:0] _27097_;
  wire [9:0] _27098_;
  wire [9:0] _27099_;
  wire [9:0] _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire [7:0] _27104_;
  wire [7:0] _27105_;
  wire [8:0] _27106_;
  wire [8:0] _27107_;
  wire [8:0] _27108_;
  wire [8:0] _27109_;
  wire [8:0] _27110_;
  wire _27111_;
  wire _27112_;
  wire [33:0] _27113_;
  wire [33:0] _27114_;
  wire [1:0] _27115_;
  wire [1:0] _27116_;
  wire [1:0] _27117_;
  wire [8:0] _27118_;
  wire [8:0] _27119_;
  wire [8:0] _27120_;
  wire [8:0] _27121_;
  wire [8:0] _27122_;
  wire [8:0] _27123_;
  wire _27124_;
  wire _27125_;
  wire [33:0] _27126_;
  wire [33:0] _27127_;
  wire [9:0] _27128_;
  wire [9:0] _27129_;
  wire [9:0] _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire [7:0] _27134_;
  wire [7:0] _27135_;
  wire [8:0] _27136_;
  wire [8:0] _27137_;
  wire [8:0] _27138_;
  wire [8:0] _27139_;
  wire [8:0] _27140_;
  wire _27141_;
  wire _27142_;
  wire [33:0] _27143_;
  wire [33:0] _27144_;
  wire [1:0] _27145_;
  wire [1:0] _27146_;
  wire [1:0] _27147_;
  wire [8:0] _27148_;
  wire [8:0] _27149_;
  wire [8:0] _27150_;
  wire [8:0] _27151_;
  wire [8:0] _27152_;
  wire [8:0] _27153_;
  wire _27154_;
  wire _27155_;
  wire [33:0] _27156_;
  wire [33:0] _27157_;
  wire [9:0] _27158_;
  wire [9:0] _27159_;
  wire [9:0] _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire [7:0] _27164_;
  wire [7:0] _27165_;
  wire [8:0] _27166_;
  wire [8:0] _27167_;
  wire [8:0] _27168_;
  wire [8:0] _27169_;
  wire [8:0] _27170_;
  wire [33:0] _27171_;
  wire [33:0] _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire [33:0] _27188_;
  wire [33:0] _27189_;
  wire _27190_;
  wire _27191_;
  wire [7:0] _27192_;
  wire [8:0] _27193_;
  wire [8:0] _27194_;
  wire [8:0] _27195_;
  wire [8:0] _27196_;
  wire _27197_;
  wire _27198_;
  wire [7:0] _27199_;
  wire [8:0] _27200_;
  wire [8:0] _27201_;
  wire [8:0] _27202_;
  wire [33:0] _27203_;
  wire [33:0] _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire [33:0] _27220_;
  wire [33:0] _27221_;
  wire _27222_;
  wire _27223_;
  wire [7:0] _27224_;
  wire [8:0] _27225_;
  wire [8:0] _27226_;
  wire [8:0] _27227_;
  wire [8:0] _27228_;
  wire _27229_;
  wire _27230_;
  wire [7:0] _27231_;
  wire [8:0] _27232_;
  wire [8:0] _27233_;
  wire [8:0] _27234_;
  wire [33:0] _27235_;
  wire [33:0] _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire [33:0] _27252_;
  wire [33:0] _27253_;
  wire _27254_;
  wire _27255_;
  wire [7:0] _27256_;
  wire [8:0] _27257_;
  wire [8:0] _27258_;
  wire [8:0] _27259_;
  wire [8:0] _27260_;
  wire _27261_;
  wire _27262_;
  wire [7:0] _27263_;
  wire [8:0] _27264_;
  wire [8:0] _27265_;
  wire [8:0] _27266_;
  wire _27267_;
  wire _27268_;
  wire [31:0] _27269_;
  wire [33:0] _27270_;
  wire [33:0] _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire [33:0] _27287_;
  wire [33:0] _27288_;
  wire _27289_;
  wire _27290_;
  wire [7:0] _27291_;
  wire [8:0] _27292_;
  wire [8:0] _27293_;
  wire [8:0] _27294_;
  wire [8:0] _27295_;
  wire _27296_;
  wire _27297_;
  wire [7:0] _27298_;
  wire [8:0] _27299_;
  wire [8:0] _27300_;
  wire [8:0] _27301_;
  wire [33:0] _27302_;
  wire [33:0] _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire [33:0] _27319_;
  wire [33:0] _27320_;
  wire _27321_;
  wire _27322_;
  wire [7:0] _27323_;
  wire [8:0] _27324_;
  wire [8:0] _27325_;
  wire [8:0] _27326_;
  wire [8:0] _27327_;
  wire _27328_;
  wire _27329_;
  wire [7:0] _27330_;
  wire [8:0] _27331_;
  wire [8:0] _27332_;
  wire [8:0] _27333_;
  wire [33:0] _27334_;
  wire [33:0] _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire [33:0] _27351_;
  wire [33:0] _27352_;
  wire _27353_;
  wire _27354_;
  wire [7:0] _27355_;
  wire [8:0] _27356_;
  wire [8:0] _27357_;
  wire [8:0] _27358_;
  wire [8:0] _27359_;
  wire _27360_;
  wire _27361_;
  wire [7:0] _27362_;
  wire [8:0] _27363_;
  wire [8:0] _27364_;
  wire [8:0] _27365_;
  wire [33:0] _27366_;
  wire [33:0] _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire [33:0] _27383_;
  wire [33:0] _27384_;
  wire _27385_;
  wire _27386_;
  wire [7:0] _27387_;
  wire [8:0] _27388_;
  wire [8:0] _27389_;
  wire [8:0] _27390_;
  wire [8:0] _27391_;
  wire _27392_;
  wire _27393_;
  wire [7:0] _27394_;
  wire [8:0] _27395_;
  wire [8:0] _27396_;
  wire [8:0] _27397_;
  wire _27398_;
  wire _27399_;
  wire [31:0] _27400_;
  wire [33:0] _27401_;
  wire [33:0] _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire [33:0] _27418_;
  wire [33:0] _27419_;
  wire _27420_;
  wire _27421_;
  wire [7:0] _27422_;
  wire [8:0] _27423_;
  wire [8:0] _27424_;
  wire [8:0] _27425_;
  wire [8:0] _27426_;
  wire _27427_;
  wire _27428_;
  wire [7:0] _27429_;
  wire [8:0] _27430_;
  wire [8:0] _27431_;
  wire [8:0] _27432_;
  wire _27433_;
  wire _27434_;
  wire [3:0] _27435_;
  wire [9:0] _27436_;
  wire [9:0] _27437_;
  wire _27438_;
  wire _27439_;
  wire [3:0] _27440_;
  wire [9:0] _27441_;
  wire [9:0] _27442_;
  wire _27443_;
  wire _27444_;
  wire [3:0] _27445_;
  wire [9:0] _27446_;
  wire [9:0] _27447_;
  wire _27448_;
  wire _27449_;
  wire [3:0] _27450_;
  wire [9:0] _27451_;
  wire [9:0] _27452_;
  wire _27453_;
  wire _27454_;
  wire [3:0] _27455_;
  wire [9:0] _27456_;
  wire [9:0] _27457_;
  wire _27458_;
  wire _27459_;
  wire [3:0] _27460_;
  wire [9:0] _27461_;
  wire [9:0] _27462_;
  wire _27463_;
  wire _27464_;
  wire [3:0] _27465_;
  wire [9:0] _27466_;
  wire [9:0] _27467_;
  wire _27468_;
  wire _27469_;
  wire [3:0] _27470_;
  wire [9:0] _27471_;
  wire [9:0] _27472_;
  wire _27473_;
  wire _27474_;
  wire [3:0] _27475_;
  wire [9:0] _27476_;
  wire [9:0] _27477_;
  wire _27478_;
  wire _27479_;
  wire [3:0] _27480_;
  wire [9:0] _27481_;
  wire [9:0] _27482_;
  wire _27483_;
  wire _27484_;
  wire [3:0] _27485_;
  wire [9:0] _27486_;
  wire [9:0] _27487_;
  wire _27488_;
  wire _27489_;
  wire [3:0] _27490_;
  wire [9:0] _27491_;
  wire [9:0] _27492_;
  wire _27493_;
  wire _27494_;
  wire [3:0] _27495_;
  wire [9:0] _27496_;
  wire [9:0] _27497_;
  wire _27498_;
  wire _27499_;
  wire [3:0] _27500_;
  wire [9:0] _27501_;
  wire [9:0] _27502_;
  wire _27503_;
  wire _27504_;
  wire [3:0] _27505_;
  wire [9:0] _27506_;
  wire [9:0] _27507_;
  wire _27508_;
  wire _27509_;
  wire [3:0] _27510_;
  wire [9:0] _27511_;
  wire [9:0] _27512_;
  wire _27513_;
  wire _27514_;
  wire [3:0] _27515_;
  wire [9:0] _27516_;
  wire [9:0] _27517_;
  wire _27518_;
  wire _27519_;
  wire [3:0] _27520_;
  wire [9:0] _27521_;
  wire [9:0] _27522_;
  wire _27523_;
  wire _27524_;
  wire [3:0] _27525_;
  wire [9:0] _27526_;
  wire [9:0] _27527_;
  wire _27528_;
  wire _27529_;
  wire [3:0] _27530_;
  wire [9:0] _27531_;
  wire [9:0] _27532_;
  wire _27533_;
  wire _27534_;
  wire [3:0] _27535_;
  wire [9:0] _27536_;
  wire [9:0] _27537_;
  wire _27538_;
  wire _27539_;
  wire [3:0] _27540_;
  wire [9:0] _27541_;
  wire [9:0] _27542_;
  wire _27543_;
  wire _27544_;
  wire [3:0] _27545_;
  wire [9:0] _27546_;
  wire [9:0] _27547_;
  wire _27548_;
  wire _27549_;
  wire [3:0] _27550_;
  wire [9:0] _27551_;
  wire [9:0] _27552_;
  wire _27553_;
  wire _27554_;
  wire [3:0] _27555_;
  wire [9:0] _27556_;
  wire [9:0] _27557_;
  wire _27558_;
  wire _27559_;
  wire [3:0] _27560_;
  wire [9:0] _27561_;
  wire [9:0] _27562_;
  wire _27563_;
  wire _27564_;
  wire [3:0] _27565_;
  wire [9:0] _27566_;
  wire [9:0] _27567_;
  wire _27568_;
  wire _27569_;
  wire [3:0] _27570_;
  wire [9:0] _27571_;
  wire [9:0] _27572_;
  wire _27573_;
  wire _27574_;
  wire [3:0] _27575_;
  wire [9:0] _27576_;
  wire [9:0] _27577_;
  wire _27578_;
  wire _27579_;
  wire [3:0] _27580_;
  wire [9:0] _27581_;
  wire [9:0] _27582_;
  wire _27583_;
  wire _27584_;
  wire [3:0] _27585_;
  wire [9:0] _27586_;
  wire [9:0] _27587_;
  wire _27588_;
  wire _27589_;
  wire [3:0] _27590_;
  wire [9:0] _27591_;
  wire [9:0] _27592_;
  wire _27593_;
  wire _27594_;
  wire [3:0] _27595_;
  wire [9:0] _27596_;
  wire [9:0] _27597_;
  wire _27598_;
  wire _27599_;
  wire [3:0] _27600_;
  wire [9:0] _27601_;
  wire [9:0] _27602_;
  wire _27603_;
  wire _27604_;
  wire [3:0] _27605_;
  wire [9:0] _27606_;
  wire [9:0] _27607_;
  wire _27608_;
  wire _27609_;
  wire [3:0] _27610_;
  wire [9:0] _27611_;
  wire [9:0] _27612_;
  wire _27613_;
  wire _27614_;
  wire [3:0] _27615_;
  wire [9:0] _27616_;
  wire [9:0] _27617_;
  wire _27618_;
  wire _27619_;
  wire [3:0] _27620_;
  wire [9:0] _27621_;
  wire [9:0] _27622_;
  wire _27623_;
  wire _27624_;
  wire [3:0] _27625_;
  wire [9:0] _27626_;
  wire [9:0] _27627_;
  wire _27628_;
  wire _27629_;
  wire [3:0] _27630_;
  wire [9:0] _27631_;
  wire [9:0] _27632_;
  wire _27633_;
  wire _27634_;
  wire [3:0] _27635_;
  wire [9:0] _27636_;
  wire [9:0] _27637_;
  wire _27638_;
  wire _27639_;
  wire [3:0] _27640_;
  wire [9:0] _27641_;
  wire [9:0] _27642_;
  wire _27643_;
  wire _27644_;
  wire [3:0] _27645_;
  wire [9:0] _27646_;
  wire [9:0] _27647_;
  wire _27648_;
  wire _27649_;
  wire [3:0] _27650_;
  wire [9:0] _27651_;
  wire [9:0] _27652_;
  wire _27653_;
  wire _27654_;
  wire [3:0] _27655_;
  wire [9:0] _27656_;
  wire [9:0] _27657_;
  wire _27658_;
  wire _27659_;
  wire [3:0] _27660_;
  wire [9:0] _27661_;
  wire [9:0] _27662_;
  wire _27663_;
  wire _27664_;
  wire [3:0] _27665_;
  wire [9:0] _27666_;
  wire [9:0] _27667_;
  wire _27668_;
  wire _27669_;
  wire [3:0] _27670_;
  wire [9:0] _27671_;
  wire [9:0] _27672_;
  wire _27673_;
  wire _27674_;
  wire [3:0] _27675_;
  wire [9:0] _27676_;
  wire [9:0] _27677_;
  wire _27678_;
  wire _27679_;
  wire [3:0] _27680_;
  wire [9:0] _27681_;
  wire [9:0] _27682_;
  wire _27683_;
  wire _27684_;
  wire [3:0] _27685_;
  wire [9:0] _27686_;
  wire [9:0] _27687_;
  wire _27688_;
  wire _27689_;
  wire [3:0] _27690_;
  wire [9:0] _27691_;
  wire [9:0] _27692_;
  wire _27693_;
  wire _27694_;
  wire [3:0] _27695_;
  wire [9:0] _27696_;
  wire [9:0] _27697_;
  wire _27698_;
  wire _27699_;
  wire [3:0] _27700_;
  wire [9:0] _27701_;
  wire [9:0] _27702_;
  wire _27703_;
  wire _27704_;
  wire [3:0] _27705_;
  wire [9:0] _27706_;
  wire [9:0] _27707_;
  wire _27708_;
  wire _27709_;
  wire [3:0] _27710_;
  wire [9:0] _27711_;
  wire [9:0] _27712_;
  wire _27713_;
  wire _27714_;
  wire [3:0] _27715_;
  wire [9:0] _27716_;
  wire [9:0] _27717_;
  wire _27718_;
  wire _27719_;
  wire [3:0] _27720_;
  wire [9:0] _27721_;
  wire [9:0] _27722_;
  wire _27723_;
  wire _27724_;
  wire [3:0] _27725_;
  wire [9:0] _27726_;
  wire [9:0] _27727_;
  wire _27728_;
  wire _27729_;
  wire [3:0] _27730_;
  wire [9:0] _27731_;
  wire [9:0] _27732_;
  wire _27733_;
  wire _27734_;
  wire [3:0] _27735_;
  wire [9:0] _27736_;
  wire [9:0] _27737_;
  wire _27738_;
  wire _27739_;
  wire [3:0] _27740_;
  wire [9:0] _27741_;
  wire [9:0] _27742_;
  wire _27743_;
  wire _27744_;
  wire [3:0] _27745_;
  wire [9:0] _27746_;
  wire [9:0] _27747_;
  wire _27748_;
  wire _27749_;
  wire [3:0] _27750_;
  wire [9:0] _27751_;
  wire [9:0] _27752_;
  wire _27753_;
  wire _27754_;
  wire [33:0] _27755_;
  wire [33:0] _27756_;
  wire [3:0] _27757_;
  wire [3:0] _27758_;
  wire [3:0] _27759_;
  wire [9:0] _27760_;
  wire [9:0] _27761_;
  wire [9:0] _27762_;
  wire [9:0] _27763_;
  wire [9:0] _27764_;
  wire [9:0] _27765_;
  wire [9:0] _27766_;
  wire [9:0] _27767_;
  wire [9:0] _27768_;
  wire [9:0] _27769_;
  wire [9:0] _27770_;
  wire [9:0] _27771_;
  wire [9:0] _27772_;
  wire [9:0] _27773_;
  wire [9:0] _27774_;
  wire [9:0] _27775_;
  wire [9:0] _27776_;
  wire [9:0] _27777_;
  wire _27778_;
  wire _27779_;
  wire [33:0] _27780_;
  wire [33:0] _27781_;
  wire [10:0] _27782_;
  wire [10:0] _27783_;
  wire [10:0] _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire [3:0] _27788_;
  wire [3:0] _27789_;
  wire [9:0] _27790_;
  wire [9:0] _27791_;
  wire [9:0] _27792_;
  wire [9:0] _27793_;
  wire [9:0] _27794_;
  wire _27795_;
  wire _27796_;
  wire [33:0] _27797_;
  wire [33:0] _27798_;
  wire [3:0] _27799_;
  wire [3:0] _27800_;
  wire [3:0] _27801_;
  wire [9:0] _27802_;
  wire [9:0] _27803_;
  wire [9:0] _27804_;
  wire [9:0] _27805_;
  wire [9:0] _27806_;
  wire [9:0] _27807_;
  wire [9:0] _27808_;
  wire [9:0] _27809_;
  wire [9:0] _27810_;
  wire [9:0] _27811_;
  wire [9:0] _27812_;
  wire [9:0] _27813_;
  wire [9:0] _27814_;
  wire [9:0] _27815_;
  wire [9:0] _27816_;
  wire [9:0] _27817_;
  wire [9:0] _27818_;
  wire [9:0] _27819_;
  wire _27820_;
  wire _27821_;
  wire [33:0] _27822_;
  wire [33:0] _27823_;
  wire [10:0] _27824_;
  wire [10:0] _27825_;
  wire [10:0] _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire [3:0] _27830_;
  wire [3:0] _27831_;
  wire [9:0] _27832_;
  wire [9:0] _27833_;
  wire [9:0] _27834_;
  wire [9:0] _27835_;
  wire [9:0] _27836_;
  wire _27837_;
  wire _27838_;
  wire [33:0] _27839_;
  wire [33:0] _27840_;
  wire [3:0] _27841_;
  wire [3:0] _27842_;
  wire [3:0] _27843_;
  wire [9:0] _27844_;
  wire [9:0] _27845_;
  wire [9:0] _27846_;
  wire [9:0] _27847_;
  wire [9:0] _27848_;
  wire [9:0] _27849_;
  wire [9:0] _27850_;
  wire [9:0] _27851_;
  wire [9:0] _27852_;
  wire [9:0] _27853_;
  wire [9:0] _27854_;
  wire [9:0] _27855_;
  wire [9:0] _27856_;
  wire [9:0] _27857_;
  wire [9:0] _27858_;
  wire [9:0] _27859_;
  wire [9:0] _27860_;
  wire [9:0] _27861_;
  wire _27862_;
  wire _27863_;
  wire [33:0] _27864_;
  wire [33:0] _27865_;
  wire [10:0] _27866_;
  wire [10:0] _27867_;
  wire [10:0] _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire [3:0] _27872_;
  wire [3:0] _27873_;
  wire [9:0] _27874_;
  wire [9:0] _27875_;
  wire [9:0] _27876_;
  wire [9:0] _27877_;
  wire [9:0] _27878_;
  wire _27879_;
  wire _27880_;
  wire [33:0] _27881_;
  wire [33:0] _27882_;
  wire [3:0] _27883_;
  wire [3:0] _27884_;
  wire [3:0] _27885_;
  wire [9:0] _27886_;
  wire [9:0] _27887_;
  wire [9:0] _27888_;
  wire [9:0] _27889_;
  wire [9:0] _27890_;
  wire [9:0] _27891_;
  wire [9:0] _27892_;
  wire [9:0] _27893_;
  wire [9:0] _27894_;
  wire [9:0] _27895_;
  wire [9:0] _27896_;
  wire [9:0] _27897_;
  wire [9:0] _27898_;
  wire [9:0] _27899_;
  wire [9:0] _27900_;
  wire [9:0] _27901_;
  wire [9:0] _27902_;
  wire [9:0] _27903_;
  wire _27904_;
  wire _27905_;
  wire [33:0] _27906_;
  wire [33:0] _27907_;
  wire [10:0] _27908_;
  wire [10:0] _27909_;
  wire [10:0] _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire [3:0] _27914_;
  wire [3:0] _27915_;
  wire [9:0] _27916_;
  wire [9:0] _27917_;
  wire [9:0] _27918_;
  wire [9:0] _27919_;
  wire [9:0] _27920_;
  wire _27921_;
  wire _27922_;
  wire [33:0] _27923_;
  wire [33:0] _27924_;
  wire [3:0] _27925_;
  wire [3:0] _27926_;
  wire [3:0] _27927_;
  wire [9:0] _27928_;
  wire [9:0] _27929_;
  wire [9:0] _27930_;
  wire [9:0] _27931_;
  wire [9:0] _27932_;
  wire [9:0] _27933_;
  wire [9:0] _27934_;
  wire [9:0] _27935_;
  wire [9:0] _27936_;
  wire [9:0] _27937_;
  wire [9:0] _27938_;
  wire [9:0] _27939_;
  wire [9:0] _27940_;
  wire [9:0] _27941_;
  wire [9:0] _27942_;
  wire [9:0] _27943_;
  wire [9:0] _27944_;
  wire [9:0] _27945_;
  wire _27946_;
  wire _27947_;
  wire [33:0] _27948_;
  wire [33:0] _27949_;
  wire [10:0] _27950_;
  wire [10:0] _27951_;
  wire [10:0] _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire [3:0] _27956_;
  wire [3:0] _27957_;
  wire [9:0] _27958_;
  wire [9:0] _27959_;
  wire [9:0] _27960_;
  wire [9:0] _27961_;
  wire [9:0] _27962_;
  wire _27963_;
  wire _27964_;
  wire [33:0] _27965_;
  wire [33:0] _27966_;
  wire [3:0] _27967_;
  wire [3:0] _27968_;
  wire [3:0] _27969_;
  wire [9:0] _27970_;
  wire [9:0] _27971_;
  wire [9:0] _27972_;
  wire [9:0] _27973_;
  wire [9:0] _27974_;
  wire [9:0] _27975_;
  wire [9:0] _27976_;
  wire [9:0] _27977_;
  wire [9:0] _27978_;
  wire [9:0] _27979_;
  wire [9:0] _27980_;
  wire [9:0] _27981_;
  wire [9:0] _27982_;
  wire [9:0] _27983_;
  wire [9:0] _27984_;
  wire [9:0] _27985_;
  wire [9:0] _27986_;
  wire [9:0] _27987_;
  wire _27988_;
  wire _27989_;
  wire [33:0] _27990_;
  wire [33:0] _27991_;
  wire [10:0] _27992_;
  wire [10:0] _27993_;
  wire [10:0] _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire [3:0] _27998_;
  wire [3:0] _27999_;
  wire [9:0] _28000_;
  wire [9:0] _28001_;
  wire [9:0] _28002_;
  wire [9:0] _28003_;
  wire [9:0] _28004_;
  wire _28005_;
  wire _28006_;
  wire [33:0] _28007_;
  wire [33:0] _28008_;
  wire [3:0] _28009_;
  wire [3:0] _28010_;
  wire [3:0] _28011_;
  wire [9:0] _28012_;
  wire [9:0] _28013_;
  wire [9:0] _28014_;
  wire [9:0] _28015_;
  wire [9:0] _28016_;
  wire [9:0] _28017_;
  wire [9:0] _28018_;
  wire [9:0] _28019_;
  wire [9:0] _28020_;
  wire [9:0] _28021_;
  wire [9:0] _28022_;
  wire [9:0] _28023_;
  wire [9:0] _28024_;
  wire [9:0] _28025_;
  wire [9:0] _28026_;
  wire [9:0] _28027_;
  wire [9:0] _28028_;
  wire [9:0] _28029_;
  wire _28030_;
  wire _28031_;
  wire [33:0] _28032_;
  wire [33:0] _28033_;
  wire [10:0] _28034_;
  wire [10:0] _28035_;
  wire [10:0] _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire [3:0] _28040_;
  wire [3:0] _28041_;
  wire [9:0] _28042_;
  wire [9:0] _28043_;
  wire [9:0] _28044_;
  wire [9:0] _28045_;
  wire [9:0] _28046_;
  wire _28047_;
  wire _28048_;
  wire [33:0] _28049_;
  wire [33:0] _28050_;
  wire [3:0] _28051_;
  wire [3:0] _28052_;
  wire [3:0] _28053_;
  wire [9:0] _28054_;
  wire [9:0] _28055_;
  wire [9:0] _28056_;
  wire [9:0] _28057_;
  wire [9:0] _28058_;
  wire [9:0] _28059_;
  wire [9:0] _28060_;
  wire [9:0] _28061_;
  wire [9:0] _28062_;
  wire [9:0] _28063_;
  wire [9:0] _28064_;
  wire [9:0] _28065_;
  wire [9:0] _28066_;
  wire [9:0] _28067_;
  wire [9:0] _28068_;
  wire [9:0] _28069_;
  wire [9:0] _28070_;
  wire [9:0] _28071_;
  wire _28072_;
  wire _28073_;
  wire [33:0] _28074_;
  wire [33:0] _28075_;
  wire [10:0] _28076_;
  wire [10:0] _28077_;
  wire [10:0] _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire [3:0] _28082_;
  wire [3:0] _28083_;
  wire [9:0] _28084_;
  wire [9:0] _28085_;
  wire [9:0] _28086_;
  wire [9:0] _28087_;
  wire [9:0] _28088_;
  wire [3:0] _28089_;
  wire [3:0] _28090_;
  wire [31:0] _28091_;
  wire [31:0] _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire [5:0] _28096_;
  wire [5:0] _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire [31:0] _28115_;
  wire [31:0] _28116_;
  wire [31:0] _28117_;
  wire [31:0] _28118_;
  wire [31:0] _28119_;
  wire [31:0] _28120_;
  wire [31:0] _28121_;
  wire [31:0] _28122_;
  wire [31:0] _28123_;
  wire [31:0] _28124_;
  wire [31:0] _28125_;
  wire [31:0] _28126_;
  wire [31:0] _28127_;
  wire [31:0] _28128_;
  wire [31:0] _28129_;
  wire [31:0] _28130_;
  wire [31:0] _28131_;
  wire [31:0] _28132_;
  wire [31:0] _28133_;
  wire [31:0] _28134_;
  wire [31:0] _28135_;
  wire [31:0] _28136_;
  wire [31:0] _28137_;
  wire [31:0] _28138_;
  wire [31:0] _28139_;
  wire [31:0] _28140_;
  wire [31:0] _28141_;
  wire [31:0] _28142_;
  wire [31:0] _28143_;
  wire [31:0] _28144_;
  wire [31:0] _28145_;
  wire [31:0] _28146_;
  wire [31:0] _28147_;
  wire [31:0] _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire [31:0] _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire [7:0] _28157_;
  wire _28158_;
  wire _28159_;
  wire [7:0] _28160_;
  wire _28161_;
  wire _28162_;
  wire [7:0] _28163_;
  wire _28164_;
  wire _28165_;
  wire [7:0] _28166_;
  wire _28167_;
  wire _28168_;
  wire [3:0] _28169_;
  wire _28170_;
  wire _28171_;
  wire [3:0] _28172_;
  wire _28173_;
  wire _28174_;
  wire [3:0] _28175_;
  wire _28176_;
  wire _28177_;
  wire [3:0] _28178_;
  wire _28179_;
  wire _28180_;
  wire [3:0] _28181_;
  wire _28182_;
  wire _28183_;
  wire [3:0] _28184_;
  wire _28185_;
  wire _28186_;
  wire [3:0] _28187_;
  wire _28188_;
  wire _28189_;
  wire [3:0] _28190_;
  wire _28191_;
  wire _28192_;
  wire [7:0] _28193_;
  wire _28194_;
  wire _28195_;
  wire [7:0] _28196_;
  wire _28197_;
  wire _28198_;
  wire [7:0] _28199_;
  wire _28200_;
  wire _28201_;
  wire [7:0] _28202_;
  wire _28203_;
  wire _28204_;
  wire [7:0] _28205_;
  wire _28206_;
  wire _28207_;
  wire [7:0] _28208_;
  wire _28209_;
  wire _28210_;
  wire [7:0] _28211_;
  wire _28212_;
  wire _28213_;
  wire [7:0] _28214_;
  wire _28215_;
  wire _28216_;
  wire [7:0] _28217_;
  wire _28218_;
  wire _28219_;
  wire [7:0] _28220_;
  wire _28221_;
  wire _28222_;
  wire [7:0] _28223_;
  wire _28224_;
  wire _28225_;
  wire [7:0] _28226_;
  wire _28227_;
  wire _28228_;
  wire [7:0] _28229_;
  wire _28230_;
  wire _28231_;
  wire [7:0] _28232_;
  wire _28233_;
  wire _28234_;
  wire [7:0] _28235_;
  wire _28236_;
  wire _28237_;
  wire [7:0] _28238_;
  wire _28239_;
  wire _28240_;
  wire [3:0] _28241_;
  wire _28242_;
  wire _28243_;
  wire [3:0] _28244_;
  wire _28245_;
  wire _28246_;
  wire [3:0] _28247_;
  wire _28248_;
  wire _28249_;
  wire [3:0] _28250_;
  wire _28251_;
  wire _28252_;
  wire [3:0] _28253_;
  wire _28254_;
  wire _28255_;
  wire [3:0] _28256_;
  wire _28257_;
  wire _28258_;
  wire [3:0] _28259_;
  wire _28260_;
  wire _28261_;
  wire [3:0] _28262_;
  wire _28263_;
  wire _28264_;
  wire [7:0] _28265_;
  wire _28266_;
  wire _28267_;
  wire [7:0] _28268_;
  wire _28269_;
  wire _28270_;
  wire [7:0] _28271_;
  wire _28272_;
  wire _28273_;
  wire [7:0] _28274_;
  wire _28275_;
  wire _28276_;
  wire [7:0] _28277_;
  wire _28278_;
  wire _28279_;
  wire [7:0] _28280_;
  wire _28281_;
  wire _28282_;
  wire [7:0] _28283_;
  wire _28284_;
  wire _28285_;
  wire [7:0] _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire [31:0] _28290_;
  wire [32:0] _28291_;
  wire [31:0] _28292_;
  wire [31:0] _28293_;
  wire [7:0] _28294_;
  wire _28295_;
  wire [31:0] _28296_;
  wire [32:0] _28297_;
  wire [31:0] _28298_;
  wire [31:0] _28299_;
  wire [7:0] _28300_;
  wire _28301_;
  wire [31:0] _28302_;
  wire [32:0] _28303_;
  wire [31:0] _28304_;
  wire [31:0] _28305_;
  wire [7:0] _28306_;
  wire _28307_;
  wire [31:0] _28308_;
  wire [32:0] _28309_;
  wire [31:0] _28310_;
  wire [31:0] _28311_;
  wire [7:0] _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire [31:0] _28317_;
  wire [32:0] _28318_;
  wire [31:0] _28319_;
  wire [31:0] _28320_;
  wire [7:0] _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire [8:0] _28326_;
  wire [8:0] _28327_;
  wire [8:0] _28328_;
  wire [8:0] _28329_;
  wire [31:0] _28330_;
  wire [32:0] _28331_;
  wire [31:0] _28332_;
  wire [31:0] _28333_;
  wire [7:0] _28334_;
  wire _28335_;
  wire [31:0] _28336_;
  wire [32:0] _28337_;
  wire [31:0] _28338_;
  wire [31:0] _28339_;
  wire [7:0] _28340_;
  wire _28341_;
  wire [31:0] _28342_;
  wire [32:0] _28343_;
  wire [31:0] _28344_;
  wire [31:0] _28345_;
  wire [7:0] _28346_;
  wire _28347_;
  wire [31:0] _28348_;
  wire [32:0] _28349_;
  wire [31:0] _28350_;
  wire [31:0] _28351_;
  wire [7:0] _28352_;
  wire _28353_;
  wire [31:0] _28354_;
  wire [32:0] _28355_;
  wire [31:0] _28356_;
  wire [31:0] _28357_;
  wire [7:0] _28358_;
  wire _28359_;
  wire [31:0] _28360_;
  wire [31:0] _28361_;
  wire [32:0] _28362_;
  wire [32:0] _28363_;
  wire [31:0] _28364_;
  wire [31:0] _28365_;
  wire [31:0] _28366_;
  wire [31:0] _28367_;
  wire [7:0] _28368_;
  wire [7:0] _28369_;
  wire _28370_;
  wire _28371_;
  wire [8:0] _28372_;
  wire [8:0] _28373_;
  wire [31:0] _28374_;
  wire [31:0] _28375_;
  wire [31:0] _28376_;
  wire [32:0] _28377_;
  wire [32:0] _28378_;
  wire [32:0] _28379_;
  wire [31:0] _28380_;
  wire [31:0] _28381_;
  wire [31:0] _28382_;
  wire [31:0] _28383_;
  wire [31:0] _28384_;
  wire [31:0] _28385_;
  wire [7:0] _28386_;
  wire [7:0] _28387_;
  wire [7:0] _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire [31:0] _28396_;
  wire [31:0] _28397_;
  wire [31:0] _28398_;
  wire [32:0] _28399_;
  wire [32:0] _28400_;
  wire [32:0] _28401_;
  wire [31:0] _28402_;
  wire [31:0] _28403_;
  wire [31:0] _28404_;
  wire [31:0] _28405_;
  wire [31:0] _28406_;
  wire [31:0] _28407_;
  wire [7:0] _28408_;
  wire [7:0] _28409_;
  wire [7:0] _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire [31:0] _28424_;
  wire [31:0] _28425_;
  wire [31:0] _28426_;
  wire [31:0] _28427_;
  wire [31:0] _28428_;
  wire [31:0] _28429_;
  wire [31:0] _28430_;
  wire [31:0] _28431_;
  wire [31:0] _28432_;
  wire [32:0] _28433_;
  wire [32:0] _28434_;
  wire [32:0] _28435_;
  wire [32:0] _28436_;
  wire [32:0] _28437_;
  wire [32:0] _28438_;
  wire [32:0] _28439_;
  wire [32:0] _28440_;
  wire [32:0] _28441_;
  wire [31:0] _28442_;
  wire [31:0] _28443_;
  wire [31:0] _28444_;
  wire [31:0] _28445_;
  wire [31:0] _28446_;
  wire [31:0] _28447_;
  wire [31:0] _28448_;
  wire [31:0] _28449_;
  wire [31:0] _28450_;
  wire [31:0] _28451_;
  wire [31:0] _28452_;
  wire [31:0] _28453_;
  wire [31:0] _28454_;
  wire [31:0] _28455_;
  wire [31:0] _28456_;
  wire [31:0] _28457_;
  wire [31:0] _28458_;
  wire [31:0] _28459_;
  wire [7:0] _28460_;
  wire [7:0] _28461_;
  wire [7:0] _28462_;
  wire [7:0] _28463_;
  wire [7:0] _28464_;
  wire [7:0] _28465_;
  wire [7:0] _28466_;
  wire [7:0] _28467_;
  wire [7:0] _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire [7:0] _28481_;
  wire [31:0] _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire [3:0] _28496_;
  wire [3:0] _28497_;
  wire [3:0] _28498_;
  wire [31:0] _28499_;
  wire [31:0] _28500_;
  wire [31:0] _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire [7:0] _28506_;
  wire [31:0] _28507_;
  wire [1:0] _28508_;
  wire [65:0] _28509_;
  wire [17:0] _28510_;
  wire [17:0] _28511_;
  wire [17:0] _28512_;
  wire [17:0] _28513_;
  wire [17:0] _28514_;
  wire [17:0] _28515_;
  wire [17:0] _28516_;
  wire [17:0] _28517_;
  wire [17:0] _28518_;
  wire [32:0] _28519_;
  wire [32:0] _28520_;
  wire [31:0] _28521_;
  wire [39:0] _28522_;
  wire [11:0] _28523_;
  wire [11:0] _28524_;
  wire [11:0] _28525_;
  wire [11:0] _28526_;
  wire [11:0] _28527_;
  wire [11:0] _28528_;
  wire [11:0] _28529_;
  wire [11:0] _28530_;
  wire [11:0] _28531_;
  wire [32:0] _28532_;
  wire [31:0] _28533_;
  wire [32:0] _28534_;
  wire [31:0] _28535_;
  wire [31:0] _28536_;
  wire [31:0] _28537_;
  wire [31:0] _28538_;
  wire [33:0] _28539_;
  wire [33:0] _28540_;
  wire [31:0] _28541_;
  wire [33:0] _28542_;
  wire [33:0] _28543_;
  wire [31:0] _28544_;
  wire [33:0] _28545_;
  wire [33:0] _28546_;
  wire [31:0] _28547_;
  wire [33:0] _28548_;
  wire [33:0] _28549_;
  wire [31:0] _28550_;
  wire [33:0] _28551_;
  wire [33:0] _28552_;
  wire [31:0] _28553_;
  wire [33:0] _28554_;
  wire [33:0] _28555_;
  wire [31:0] _28556_;
  wire [33:0] _28557_;
  wire [33:0] _28558_;
  wire [31:0] _28559_;
  wire [33:0] _28560_;
  wire [33:0] _28561_;
  wire [33:0] _28562_;
  wire [33:0] _28563_;
  wire [33:0] _28564_;
  wire [33:0] _28565_;
  wire [33:0] _28566_;
  wire [33:0] _28567_;
  wire [33:0] _28568_;
  wire [33:0] _28569_;
  wire [33:0] _28570_;
  wire [33:0] _28571_;
  wire [33:0] _28572_;
  wire [33:0] _28573_;
  wire [33:0] _28574_;
  wire [33:0] _28575_;
  wire [33:0] _28576_;
  wire [33:0] _28577_;
  wire [33:0] _28578_;
  wire [31:0] _28579_;
  wire [31:0] _28580_;
  wire [33:0] _28581_;
  wire [33:0] _28582_;
  wire [31:0] _28583_;
  wire [33:0] _28584_;
  wire [33:0] _28585_;
  wire [31:0] _28586_;
  wire [33:0] _28587_;
  wire [33:0] _28588_;
  wire [31:0] _28589_;
  wire [33:0] _28590_;
  wire [33:0] _28591_;
  wire [33:0] _28592_;
  wire [33:0] _28593_;
  wire [33:0] _28594_;
  wire [33:0] _28595_;
  wire [31:0] _28596_;
  wire [31:0] _28597_;
  wire [33:0] _28598_;
  wire [31:0] _28599_;
  wire [33:0] _28600_;
  wire [31:0] _28601_;
  wire [33:0] _28602_;
  wire [31:0] _28603_;
  wire [33:0] _28604_;
  wire [31:0] _28605_;
  wire [31:0] _28606_;
  wire [33:0] _28607_;
  wire [31:0] _28608_;
  wire [33:0] _28609_;
  wire [31:0] _28610_;
  wire [33:0] _28611_;
  wire [31:0] _28612_;
  wire [33:0] _28613_;
  wire [33:0] _28614_;
  wire [33:0] _28615_;
  wire [33:0] _28616_;
  wire [33:0] _28617_;
  wire [5:0] _28618_;
  wire [3:0] _28619_;
  wire [3:0] _28620_;
  wire [3:0] _28621_;
  wire [3:0] _28622_;
  wire [3:0] _28623_;
  wire [3:0] _28624_;
  wire [3:0] _28625_;
  wire [3:0] _28626_;
  wire [3:0] _28627_;
  wire [32:0] _28628_;
  wire [32:0] _28629_;
  wire [32:0] _28630_;
  wire [32:0] _28631_;
  wire [32:0] _28632_;
  wire [32:0] _28633_;
  wire [32:0] _28634_;
  wire [32:0] _28635_;
  wire [32:0] _28636_;
  wire [32:0] _28637_;
  wire [32:0] _28638_;
  wire [32:0] _28639_;
  wire [32:0] _28640_;
  wire [32:0] _28641_;
  wire [32:0] _28642_;
  wire [32:0] _28643_;
  wire [32:0] _28644_;
  wire [32:0] _28645_;
  wire [32:0] _28646_;
  wire [32:0] _28647_;
  wire [32:0] _28648_;
  wire [32:0] _28649_;
  wire [32:0] _28650_;
  wire [32:0] _28651_;
  wire [32:0] _28652_;
  wire [32:0] _28653_;
  wire [32:0] _28654_;
  wire [32:0] _28655_;
  wire [32:0] _28656_;
  wire [32:0] _28657_;
  wire [32:0] _28658_;
  wire [32:0] _28659_;
  wire [32:0] _28660_;
  wire [32:0] _28661_;
  wire [32:0] _28662_;
  wire [32:0] _28663_;
  wire [32:0] _28664_;
  wire [32:0] _28665_;
  wire [32:0] _28666_;
  wire [32:0] _28667_;
  wire [32:0] _28668_;
  wire [32:0] _28669_;
  wire [32:0] _28670_;
  wire [32:0] _28671_;
  wire [32:0] _28672_;
  wire [32:0] _28673_;
  wire [32:0] _28674_;
  wire [32:0] _28675_;
  wire [32:0] _28676_;
  wire [32:0] _28677_;
  wire [32:0] _28678_;
  wire [32:0] _28679_;
  wire [32:0] _28680_;
  wire [32:0] _28681_;
  wire [32:0] _28682_;
  wire [32:0] _28683_;
  wire [32:0] _28684_;
  wire [32:0] _28685_;
  wire [32:0] _28686_;
  wire [32:0] _28687_;
  wire [32:0] _28688_;
  wire [32:0] _28689_;
  wire [32:0] _28690_;
  wire [32:0] _28691_;
  wire [32:0] _28692_;
  wire [32:0] _28693_;
  wire [32:0] _28694_;
  wire [32:0] _28695_;
  wire [32:0] _28696_;
  wire [32:0] _28697_;
  wire [32:0] _28698_;
  wire [32:0] _28699_;
  wire [32:0] _28700_;
  wire [32:0] _28701_;
  wire [32:0] _28702_;
  wire [32:0] _28703_;
  wire [32:0] _28704_;
  wire [32:0] _28705_;
  wire [32:0] _28706_;
  wire [32:0] _28707_;
  wire [32:0] _28708_;
  wire [32:0] _28709_;
  wire [32:0] _28710_;
  wire [32:0] _28711_;
  wire [32:0] _28712_;
  wire [32:0] _28713_;
  wire [32:0] _28714_;
  wire [32:0] _28715_;
  wire [32:0] _28716_;
  wire [32:0] _28717_;
  wire [32:0] _28718_;
  wire [32:0] _28719_;
  wire [32:0] _28720_;
  wire [32:0] _28721_;
  wire [32:0] _28722_;
  wire [32:0] _28723_;
  wire [32:0] _28724_;
  wire [32:0] _28725_;
  wire [32:0] _28726_;
  wire [32:0] _28727_;
  wire [32:0] _28728_;
  wire [32:0] _28729_;
  wire [32:0] _28730_;
  wire [32:0] _28731_;
  wire [32:0] _28732_;
  wire [32:0] _28733_;
  wire [32:0] _28734_;
  wire [32:0] _28735_;
  wire [32:0] _28736_;
  wire [32:0] _28737_;
  wire [32:0] _28738_;
  wire [32:0] _28739_;
  wire [32:0] _28740_;
  wire [32:0] _28741_;
  wire [32:0] _28742_;
  wire [32:0] _28743_;
  wire [32:0] _28744_;
  wire [32:0] _28745_;
  wire [32:0] _28746_;
  wire [32:0] _28747_;
  wire [32:0] _28748_;
  wire [32:0] _28749_;
  wire [32:0] _28750_;
  wire [32:0] _28751_;
  wire [32:0] _28752_;
  wire [32:0] _28753_;
  wire [32:0] _28754_;
  wire [32:0] _28755_;
  wire [32:0] _28756_;
  wire [32:0] _28757_;
  wire [32:0] _28758_;
  wire [32:0] _28759_;
  wire [32:0] _28760_;
  wire [32:0] _28761_;
  wire [32:0] _28762_;
  wire [32:0] _28763_;
  wire [32:0] _28764_;
  wire [32:0] _28765_;
  wire [32:0] _28766_;
  wire [32:0] _28767_;
  wire [32:0] _28768_;
  wire [32:0] _28769_;
  wire [32:0] _28770_;
  wire [32:0] _28771_;
  wire [32:0] _28772_;
  wire [32:0] _28773_;
  wire [32:0] _28774_;
  wire [32:0] _28775_;
  wire [32:0] _28776_;
  wire [32:0] _28777_;
  wire [32:0] _28778_;
  wire [32:0] _28779_;
  wire [32:0] _28780_;
  wire [32:0] _28781_;
  wire [32:0] _28782_;
  wire [32:0] _28783_;
  wire [32:0] _28784_;
  wire [32:0] _28785_;
  wire [32:0] _28786_;
  wire [32:0] _28787_;
  wire [32:0] _28788_;
  wire [32:0] _28789_;
  wire [32:0] _28790_;
  wire [32:0] _28791_;
  wire [32:0] _28792_;
  wire [32:0] _28793_;
  wire [32:0] _28794_;
  wire [32:0] _28795_;
  wire [32:0] _28796_;
  wire [32:0] _28797_;
  wire [32:0] _28798_;
  wire [32:0] _28799_;
  wire [32:0] _28800_;
  wire [32:0] _28801_;
  wire [32:0] _28802_;
  wire [32:0] _28803_;
  wire [32:0] _28804_;
  wire [32:0] _28805_;
  wire [32:0] _28806_;
  wire [32:0] _28807_;
  wire [32:0] _28808_;
  wire [32:0] _28809_;
  wire [32:0] _28810_;
  wire [32:0] _28811_;
  wire [32:0] _28812_;
  wire [32:0] _28813_;
  wire [32:0] _28814_;
  wire [32:0] _28815_;
  wire [32:0] _28816_;
  wire [32:0] _28817_;
  wire [32:0] _28818_;
  wire [32:0] _28819_;
  wire [32:0] _28820_;
  wire [32:0] _28821_;
  wire [32:0] _28822_;
  wire [32:0] _28823_;
  wire [32:0] _28824_;
  wire [32:0] _28825_;
  wire [32:0] _28826_;
  wire [32:0] _28827_;
  wire [32:0] _28828_;
  wire [32:0] _28829_;
  wire [32:0] _28830_;
  wire [32:0] _28831_;
  wire [32:0] _28832_;
  wire [32:0] _28833_;
  wire [32:0] _28834_;
  wire [32:0] _28835_;
  wire [32:0] _28836_;
  wire [32:0] _28837_;
  wire [32:0] _28838_;
  wire [32:0] _28839_;
  wire [32:0] _28840_;
  wire [32:0] _28841_;
  wire [32:0] _28842_;
  wire [32:0] _28843_;
  wire [32:0] _28844_;
  wire [32:0] _28845_;
  wire [32:0] _28846_;
  wire [32:0] _28847_;
  wire [32:0] _28848_;
  wire [32:0] _28849_;
  wire [32:0] _28850_;
  wire [32:0] _28851_;
  wire [32:0] _28852_;
  wire [32:0] _28853_;
  wire [32:0] _28854_;
  wire [32:0] _28855_;
  wire [32:0] _28856_;
  wire [32:0] _28857_;
  wire [32:0] _28858_;
  wire [32:0] _28859_;
  wire [32:0] _28860_;
  wire [32:0] _28861_;
  wire [32:0] _28862_;
  wire [32:0] _28863_;
  wire [32:0] _28864_;
  wire [32:0] _28865_;
  wire [32:0] _28866_;
  wire [32:0] _28867_;
  wire [31:0] _28868_;
  wire [32:0] _28869_;
  wire [31:0] _28870_;
  wire [32:0] _28871_;
  wire [32:0] _28872_;
  wire [32:0] _28873_;
  wire [32:0] _28874_;
  wire [32:0] _28875_;
  wire [32:0] _28876_;
  wire [32:0] _28877_;
  wire [32:0] _28878_;
  wire [32:0] _28879_;
  wire [32:0] _28880_;
  wire [32:0] _28881_;
  wire [32:0] _28882_;
  wire [31:0] _28883_;
  wire [32:0] _28884_;
  wire [32:0] _28885_;
  wire [32:0] _28886_;
  wire [32:0] _28887_;
  wire [32:0] _28888_;
  wire [32:0] _28889_;
  wire [32:0] _28890_;
  wire [32:0] _28891_;
  wire [32:0] _28892_;
  wire [32:0] _28893_;
  wire [32:0] _28894_;
  wire [32:0] _28895_;
  wire [32:0] _28896_;
  wire [32:0] _28897_;
  wire [32:0] _28898_;
  wire [32:0] _28899_;
  wire [32:0] _28900_;
  wire [32:0] _28901_;
  wire [32:0] _28902_;
  wire [32:0] _28903_;
  wire [32:0] _28904_;
  wire [32:0] _28905_;
  wire [32:0] _28906_;
  wire [32:0] _28907_;
  wire [32:0] _28908_;
  wire [32:0] _28909_;
  wire [32:0] _28910_;
  wire [32:0] _28911_;
  wire [32:0] _28912_;
  wire [32:0] _28913_;
  wire [32:0] _28914_;
  wire [32:0] _28915_;
  wire [32:0] _28916_;
  wire [32:0] _28917_;
  wire [32:0] _28918_;
  wire [32:0] _28919_;
  wire [32:0] _28920_;
  wire [32:0] _28921_;
  wire [32:0] _28922_;
  wire [32:0] _28923_;
  wire [32:0] _28924_;
  wire [32:0] _28925_;
  wire [32:0] _28926_;
  wire [32:0] _28927_;
  wire [32:0] _28928_;
  wire [32:0] _28929_;
  wire [32:0] _28930_;
  wire [32:0] _28931_;
  wire [32:0] _28932_;
  wire [31:0] _28933_;
  wire [32:0] _28934_;
  wire [31:0] _28935_;
  wire [32:0] _28936_;
  wire [32:0] _28937_;
  wire [32:0] _28938_;
  wire [1:0] _28939_;
  wire [32:0] _28940_;
  wire [32:0] _28941_;
  wire [32:0] _28942_;
  wire [65:0] _28943_;
  wire [65:0] _28944_;
  wire [65:0] _28945_;
  wire [65:0] _28946_;
  wire [65:0] _28947_;
  wire [65:0] _28948_;
  wire [65:0] _28949_;
  wire [17:0] _28950_;
  wire [17:0] _28951_;
  wire [17:0] _28952_;
  wire [17:0] _28953_;
  wire [17:0] _28954_;
  wire [17:0] _28955_;
  wire [17:0] _28956_;
  wire [17:0] _28957_;
  wire [17:0] _28958_;
  wire [17:0] _28959_;
  wire [17:0] _28960_;
  wire [17:0] _28961_;
  wire [17:0] _28962_;
  wire [17:0] _28963_;
  wire [17:0] _28964_;
  wire [17:0] _28965_;
  wire [17:0] _28966_;
  wire [17:0] _28967_;
  wire [17:0] _28968_;
  wire [17:0] _28969_;
  wire [17:0] _28970_;
  wire [17:0] _28971_;
  wire [17:0] _28972_;
  wire [17:0] _28973_;
  wire [17:0] _28974_;
  wire [17:0] _28975_;
  wire [17:0] _28976_;
  wire [31:0] _28977_;
  wire [31:0] _28978_;
  wire [31:0] _28979_;
  wire [31:0] _28980_;
  wire [31:0] _28981_;
  wire [31:0] _28982_;
  wire [39:0] _28983_;
  wire [39:0] _28984_;
  wire [39:0] _28985_;
  wire [39:0] _28986_;
  wire [39:0] _28987_;
  wire [39:0] _28988_;
  wire [11:0] _28989_;
  wire [11:0] _28990_;
  wire [11:0] _28991_;
  wire [11:0] _28992_;
  wire [11:0] _28993_;
  wire [11:0] _28994_;
  wire [11:0] _28995_;
  wire [11:0] _28996_;
  wire [11:0] _28997_;
  wire [11:0] _28998_;
  wire [11:0] _28999_;
  wire [11:0] _29000_;
  wire [11:0] _29001_;
  wire [11:0] _29002_;
  wire [11:0] _29003_;
  wire [11:0] _29004_;
  wire [11:0] _29005_;
  wire [11:0] _29006_;
  wire [11:0] _29007_;
  wire [11:0] _29008_;
  wire [11:0] _29009_;
  wire [11:0] _29010_;
  wire [11:0] _29011_;
  wire [11:0] _29012_;
  wire [11:0] _29013_;
  wire [11:0] _29014_;
  wire [11:0] _29015_;
  wire [11:0] _29016_;
  wire [11:0] _29017_;
  wire [11:0] _29018_;
  wire [11:0] _29019_;
  wire [11:0] _29020_;
  wire [11:0] _29021_;
  wire [11:0] _29022_;
  wire [11:0] _29023_;
  wire [11:0] _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire [31:0] _29057_;
  wire [31:0] _29058_;
  wire [31:0] _29059_;
  wire [31:0] _29060_;
  wire [31:0] _29061_;
  wire [31:0] _29062_;
  wire [31:0] _29063_;
  wire [31:0] _29064_;
  wire [31:0] _29065_;
  wire [31:0] _29066_;
  wire [31:0] _29067_;
  wire [31:0] _29068_;
  wire [31:0] _29069_;
  wire [31:0] _29070_;
  wire [31:0] _29071_;
  wire [31:0] _29072_;
  wire [31:0] _29073_;
  wire [31:0] _29074_;
  wire [31:0] _29075_;
  wire [31:0] _29076_;
  wire [31:0] _29077_;
  wire [31:0] _29078_;
  wire [31:0] _29079_;
  wire [31:0] _29080_;
  wire [31:0] _29081_;
  wire [31:0] _29082_;
  wire [31:0] _29083_;
  wire [31:0] _29084_;
  wire [31:0] _29085_;
  wire [31:0] _29086_;
  wire [31:0] _29087_;
  wire [31:0] _29088_;
  wire [31:0] _29089_;
  wire [31:0] _29090_;
  wire [31:0] _29091_;
  wire [31:0] _29092_;
  wire [31:0] _29093_;
  wire [31:0] _29094_;
  wire [31:0] _29095_;
  wire [31:0] _29096_;
  wire [31:0] _29097_;
  wire [31:0] _29098_;
  wire [31:0] _29099_;
  wire [31:0] _29100_;
  wire [31:0] _29101_;
  wire [31:0] _29102_;
  wire [31:0] _29103_;
  wire [31:0] _29104_;
  wire [31:0] _29105_;
  wire [31:0] _29106_;
  wire [31:0] _29107_;
  wire [31:0] _29108_;
  wire [31:0] _29109_;
  wire [31:0] _29110_;
  wire [31:0] _29111_;
  wire [31:0] _29112_;
  wire [31:0] _29113_;
  wire [31:0] _29114_;
  wire [31:0] _29115_;
  wire [31:0] _29116_;
  wire [31:0] _29117_;
  wire [31:0] _29118_;
  wire [31:0] _29119_;
  wire [31:0] _29120_;
  wire [31:0] _29121_;
  wire [31:0] _29122_;
  wire [31:0] _29123_;
  wire [31:0] _29124_;
  wire [31:0] _29125_;
  wire [31:0] _29126_;
  wire [31:0] _29127_;
  wire [31:0] _29128_;
  wire [31:0] _29129_;
  wire [31:0] _29130_;
  wire [31:0] _29131_;
  wire [31:0] _29132_;
  wire [31:0] _29133_;
  wire [31:0] _29134_;
  wire [31:0] _29135_;
  wire [31:0] _29136_;
  wire [31:0] _29137_;
  wire [31:0] _29138_;
  wire [31:0] _29139_;
  wire [31:0] _29140_;
  wire [31:0] _29141_;
  wire [31:0] _29142_;
  wire [31:0] _29143_;
  wire [31:0] _29144_;
  wire [31:0] _29145_;
  wire [31:0] _29146_;
  wire [31:0] _29147_;
  wire [32:0] _29148_;
  wire [32:0] _29149_;
  wire [65:0] _29150_;
  wire [39:0] _29151_;
  wire [39:0] _29152_;
  wire [39:0] _29153_;
  wire [17:0] _29154_;
  wire [17:0] _29155_;
  wire [17:0] _29156_;
  wire [17:0] _29157_;
  wire [17:0] _29158_;
  wire [17:0] _29159_;
  wire [17:0] _29160_;
  wire [17:0] _29161_;
  wire [17:0] _29162_;
  wire [7:0] _29163_;
  wire [31:0] _29164_;
  wire [8:0] _29165_;
  wire [31:0] _29166_;
  wire [7:0] _29167_;
  wire [7:0] _29168_;
  wire [7:0] _29169_;
  wire [7:0] _29170_;
  wire [7:0] _29171_;
  wire [7:0] _29172_;
  wire [7:0] _29173_;
  wire [7:0] _29174_;
  wire [7:0] _29175_;
  wire [7:0] _29176_;
  wire [7:0] _29177_;
  wire [7:0] _29178_;
  wire [7:0] _29179_;
  wire [7:0] _29180_;
  wire [7:0] _29181_;
  wire [7:0] _29182_;
  wire [7:0] _29183_;
  wire [7:0] _29184_;
  wire [7:0] _29185_;
  wire [7:0] _29186_;
  wire [7:0] _29187_;
  wire [7:0] _29188_;
  wire [7:0] _29189_;
  wire [7:0] _29190_;
  wire [7:0] _29191_;
  wire [7:0] _29192_;
  wire [7:0] _29193_;
  wire [7:0] _29194_;
  wire [7:0] _29195_;
  wire [7:0] _29196_;
  wire [7:0] _29197_;
  wire [7:0] _29198_;
  wire [7:0] _29199_;
  wire [7:0] _29200_;
  wire [7:0] _29201_;
  wire [7:0] _29202_;
  wire [7:0] _29203_;
  wire [7:0] _29204_;
  wire [7:0] _29205_;
  wire [7:0] _29206_;
  wire [7:0] _29207_;
  wire [7:0] _29208_;
  wire [7:0] _29209_;
  wire [7:0] _29210_;
  wire [7:0] _29211_;
  wire [7:0] _29212_;
  wire [7:0] _29213_;
  wire [7:0] _29214_;
  wire [7:0] _29215_;
  wire [7:0] _29216_;
  wire [7:0] _29217_;
  wire [7:0] _29218_;
  wire [7:0] _29219_;
  wire [7:0] _29220_;
  wire [7:0] _29221_;
  wire [7:0] _29222_;
  wire [7:0] _29223_;
  wire [7:0] _29224_;
  wire [7:0] _29225_;
  wire [7:0] _29226_;
  wire [7:0] _29227_;
  wire [7:0] _29228_;
  wire [7:0] _29229_;
  wire [7:0] _29230_;
  wire [31:0] _29231_;
  wire [31:0] _29232_;
  wire [31:0] _29233_;
  wire [31:0] _29234_;
  wire [31:0] _29235_;
  wire [31:0] _29236_;
  wire [31:0] _29237_;
  wire [31:0] _29238_;
  wire [31:0] _29239_;
  wire [31:0] _29240_;
  wire [31:0] _29241_;
  wire [31:0] _29242_;
  wire [31:0] _29243_;
  wire [31:0] _29244_;
  wire [31:0] _29245_;
  wire [31:0] _29246_;
  wire [31:0] _29247_;
  wire [31:0] _29248_;
  wire [31:0] _29249_;
  wire [31:0] _29250_;
  wire [31:0] _29251_;
  wire [31:0] _29252_;
  wire [31:0] _29253_;
  wire [31:0] _29254_;
  wire [31:0] _29255_;
  wire [31:0] _29256_;
  wire [31:0] _29257_;
  wire [31:0] _29258_;
  wire [31:0] _29259_;
  wire [31:0] _29260_;
  wire [31:0] _29261_;
  wire [31:0] _29262_;
  wire [31:0] _29263_;
  wire [31:0] _29264_;
  wire [31:0] _29265_;
  wire [31:0] _29266_;
  wire [31:0] _29267_;
  wire [31:0] _29268_;
  wire [31:0] _29269_;
  wire [31:0] _29270_;
  wire [31:0] _29271_;
  wire [31:0] _29272_;
  wire [31:0] _29273_;
  wire [31:0] _29274_;
  wire [31:0] _29275_;
  wire [31:0] _29276_;
  wire [31:0] _29277_;
  wire [31:0] _29278_;
  wire [31:0] _29279_;
  wire [31:0] _29280_;
  wire [8:0] _29281_;
  wire [31:0] _29282_;
  wire [31:0] _29283_;
  wire [31:0] _29284_;
  wire [31:0] _29285_;
  wire [31:0] _29286_;
  wire [31:0] _29287_;
  wire [7:0] _29288_;
  wire [7:0] _29289_;
  wire [7:0] _29290_;
  wire [7:0] _29291_;
  wire [7:0] _29292_;
  wire [31:0] _29293_;
  wire [31:0] _29294_;
  wire [31:0] _29295_;
  wire [31:0] _29296_;
  wire [31:0] _29297_;
  wire [31:0] _29298_;
  wire [31:0] _29299_;
  wire [31:0] _29300_;
  wire [31:0] _29301_;
  wire [31:0] _29302_;
  wire [31:0] _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire [31:0] _29316_;
  wire [31:0] _29317_;
  wire [31:0] _29318_;
  wire [31:0] _29319_;
  wire [31:0] _29320_;
  wire [31:0] _29321_;
  wire [31:0] _29322_;
  wire [31:0] _29323_;
  wire [31:0] _29324_;
  wire [31:0] _29325_;
  wire [31:0] _29326_;
  wire [31:0] _29327_;
  wire [31:0] _29328_;
  wire [31:0] _29329_;
  wire [31:0] _29330_;
  wire [31:0] _29331_;
  wire [31:0] _29332_;
  wire [31:0] _29333_;
  wire [31:0] _29334_;
  wire [31:0] _29335_;
  wire [31:0] _29336_;
  wire [31:0] _29337_;
  wire [31:0] _29338_;
  wire [31:0] _29339_;
  wire [31:0] _29340_;
  wire [31:0] _29341_;
  wire [31:0] _29342_;
  wire [31:0] _29343_;
  wire [31:0] _29344_;
  wire [31:0] _29345_;
  wire [31:0] _29346_;
  wire [31:0] _29347_;
  wire [31:0] _29348_;
  wire [31:0] _29349_;
  wire [31:0] _29350_;
  wire [31:0] _29351_;
  wire [31:0] _29352_;
  wire [31:0] _29353_;
  wire [31:0] _29354_;
  wire [31:0] _29355_;
  wire [31:0] _29356_;
  wire [31:0] _29357_;
  wire [31:0] _29358_;
  wire [31:0] _29359_;
  wire [31:0] _29360_;
  wire [31:0] _29361_;
  wire [31:0] _29362_;
  wire [31:0] _29363_;
  wire [31:0] _29364_;
  wire [31:0] _29365_;
  wire [31:0] _29366_;
  wire [31:0] _29367_;
  wire [31:0] _29368_;
  wire [31:0] _29369_;
  wire [31:0] _29370_;
  wire [31:0] _29371_;
  wire [31:0] _29372_;
  wire [31:0] _29373_;
  wire [31:0] _29374_;
  wire [31:0] _29375_;
  wire [31:0] _29376_;
  wire [31:0] _29377_;
  wire [31:0] _29378_;
  wire [31:0] _29379_;
  wire [31:0] _29380_;
  wire [31:0] _29381_;
  wire [31:0] _29382_;
  wire [31:0] _29383_;
  wire [31:0] _29384_;
  wire [31:0] _29385_;
  wire [31:0] _29386_;
  wire [31:0] _29387_;
  wire [31:0] _29388_;
  wire [31:0] _29389_;
  wire [31:0] _29390_;
  wire [31:0] _29391_;
  wire [31:0] _29392_;
  wire [31:0] _29393_;
  wire [31:0] _29394_;
  wire [31:0] _29395_;
  wire [31:0] _29396_;
  wire [31:0] _29397_;
  wire [31:0] _29398_;
  wire [31:0] _29399_;
  wire [31:0] _29400_;
  wire [31:0] _29401_;
  wire [31:0] _29402_;
  wire [31:0] _29403_;
  wire [31:0] _29404_;
  wire [31:0] _29405_;
  wire [31:0] _29406_;
  wire [31:0] _29407_;
  wire [31:0] _29408_;
  wire [31:0] _29409_;
  wire [31:0] _29410_;
  wire [31:0] _29411_;
  wire [31:0] _29412_;
  wire [31:0] _29413_;
  wire [31:0] _29414_;
  wire [31:0] _29415_;
  wire [31:0] _29416_;
  wire [31:0] _29417_;
  wire [31:0] _29418_;
  wire [31:0] _29419_;
  wire [31:0] _29420_;
  wire [31:0] _29421_;
  wire [31:0] _29422_;
  wire [31:0] _29423_;
  wire [31:0] _29424_;
  wire [31:0] _29425_;
  wire [31:0] _29426_;
  wire [31:0] _29427_;
  wire [31:0] _29428_;
  wire [31:0] _29429_;
  wire [31:0] _29430_;
  wire [31:0] _29431_;
  wire [31:0] _29432_;
  wire [31:0] _29433_;
  wire [31:0] _29434_;
  wire [31:0] _29435_;
  wire [31:0] _29436_;
  wire [31:0] _29437_;
  wire [31:0] _29438_;
  wire [31:0] _29439_;
  wire [31:0] _29440_;
  wire [31:0] _29441_;
  wire [31:0] _29442_;
  wire [31:0] _29443_;
  wire [31:0] _29444_;
  wire [31:0] _29445_;
  wire [31:0] _29446_;
  wire [31:0] _29447_;
  wire [31:0] _29448_;
  wire [31:0] _29449_;
  wire [31:0] _29450_;
  wire [31:0] _29451_;
  wire [31:0] _29452_;
  wire RESETN_inv;
  wire RESETN_inv_buf;
  wire RST;
  wire _RESETN_inv_1;
  wire _RESETN_inv_2;
  wire [3:0] __delay_data_1000;
  wire [3:0] __delay_data_1001;
  wire [3:0] __delay_data_1002;
  wire [3:0] __delay_data_1003;
  wire [3:0] __delay_data_1004;
  wire [3:0] __delay_data_1005;
  wire [3:0] __delay_data_1006;
  wire [7:0] __delay_data_1007;
  wire [7:0] __delay_data_1008;
  wire [7:0] __delay_data_1009;
  wire [7:0] __delay_data_1010;
  wire [7:0] __delay_data_1011;
  wire [7:0] __delay_data_1012;
  wire __delay_data_1013;
  wire __delay_data_1014;
  wire __delay_data_1015;
  wire [7:0] __delay_data_1016;
  wire __delay_data_1017;
  wire __delay_data_1018;
  wire __delay_data_1019;
  wire [7:0] __delay_data_1020;
  wire __delay_data_1021;
  wire __delay_data_1022;
  wire __delay_data_1023;
  wire [7:0] __delay_data_1024;
  wire __delay_data_1025;
  wire __delay_data_1026;
  wire __delay_data_1027;
  wire __delay_data_1028;
  wire __delay_data_1029;
  wire __delay_data_1030;
  wire __delay_data_1031;
  wire [7:0] __delay_data_1032;
  wire __delay_data_1033;
  wire __delay_data_1034;
  wire __delay_data_1035;
  wire __delay_data_1036;
  wire __delay_data_1037;
  wire [7:0] __delay_data_1038;
  wire [7:0] __delay_data_1039;
  wire __delay_data_1040;
  wire __delay_data_1041;
  wire __delay_data_1042;
  wire __delay_data_1043;
  wire __delay_data_1044;
  wire __delay_data_1045;
  wire __delay_data_1046;
  wire [3:0] __delay_data_1047;
  wire [3:0] __delay_data_1048;
  wire [3:0] __delay_data_1049;
  wire [3:0] __delay_data_1050;
  wire [3:0] __delay_data_1051;
  wire [3:0] __delay_data_1052;
  wire [3:0] __delay_data_1053;
  wire [3:0] __delay_data_1054;
  wire [7:0] __delay_data_1055;
  wire [7:0] __delay_data_1056;
  wire [7:0] __delay_data_1057;
  wire [7:0] __delay_data_1058;
  wire [7:0] __delay_data_1059;
  wire [7:0] __delay_data_1060;
  wire __delay_data_1061;
  wire __delay_data_1062;
  wire __delay_data_1063;
  wire __delay_data_1064;
  wire __delay_data_1065;
  wire __delay_data_1066;
  wire __delay_data_1067;
  wire [7:0] __delay_data_1068;
  wire __delay_data_1069;
  wire __delay_data_1070;
  wire __delay_data_1071;
  wire __delay_data_1072;
  wire __delay_data_1073;
  wire [7:0] __delay_data_1074;
  wire __delay_data_1075;
  wire __delay_data_1076;
  wire __delay_data_1077;
  wire __delay_data_1078;
  wire __delay_data_1079;
  wire __delay_data_1080;
  wire __delay_data_1081;
  wire [3:0] __delay_data_1082;
  wire [3:0] __delay_data_1083;
  wire [3:0] __delay_data_1084;
  wire [3:0] __delay_data_1085;
  wire [3:0] __delay_data_1086;
  wire [3:0] __delay_data_1087;
  wire [3:0] __delay_data_1088;
  wire [3:0] __delay_data_1089;
  wire [7:0] __delay_data_1090;
  wire [7:0] __delay_data_1091;
  wire [7:0] __delay_data_1092;
  wire [7:0] __delay_data_1093;
  wire [7:0] __delay_data_1094;
  wire [7:0] __delay_data_1095;
  wire __delay_data_1096;
  wire __delay_data_1097;
  wire __delay_data_1098;
  wire __delay_data_1099;
  wire __delay_data_1100;
  wire __delay_data_1101;
  wire __delay_data_1102;
  wire [7:0] __delay_data_1103;
  wire __delay_data_1104;
  wire __delay_data_1105;
  wire __delay_data_1106;
  wire __delay_data_1107;
  wire __delay_data_1108;
  wire [7:0] __delay_data_1109;
  wire __delay_data_1110;
  wire __delay_data_1111;
  wire __delay_data_1112;
  wire __delay_data_1113;
  wire __delay_data_1114;
  wire __delay_data_1115;
  wire __delay_data_1116;
  wire [3:0] __delay_data_1117;
  wire [3:0] __delay_data_1118;
  wire [3:0] __delay_data_1119;
  wire [3:0] __delay_data_1120;
  wire [3:0] __delay_data_1121;
  wire [3:0] __delay_data_1122;
  wire [3:0] __delay_data_1123;
  wire [3:0] __delay_data_1124;
  wire [7:0] __delay_data_1125;
  wire [7:0] __delay_data_1126;
  wire [7:0] __delay_data_1127;
  wire [7:0] __delay_data_1128;
  wire [7:0] __delay_data_1129;
  wire [7:0] __delay_data_1130;
  wire __delay_data_1131;
  wire __delay_data_1132;
  wire __delay_data_1133;
  wire __delay_data_1134;
  wire __delay_data_1135;
  wire __delay_data_1136;
  wire __delay_data_1137;
  wire [7:0] __delay_data_1138;
  wire __delay_data_1139;
  wire __delay_data_1140;
  wire __delay_data_1141;
  wire __delay_data_1142;
  wire __delay_data_1143;
  wire [7:0] __delay_data_1144;
  wire __delay_data_1145;
  wire __delay_data_1146;
  wire __delay_data_1147;
  wire __delay_data_1148;
  wire __delay_data_1149;
  wire __delay_data_1150;
  wire __delay_data_1151;
  wire [3:0] __delay_data_1152;
  wire [3:0] __delay_data_1153;
  wire [3:0] __delay_data_1154;
  wire [3:0] __delay_data_1155;
  wire [3:0] __delay_data_1156;
  wire [3:0] __delay_data_1157;
  wire [3:0] __delay_data_1158;
  wire [3:0] __delay_data_1159;
  wire [7:0] __delay_data_1160;
  wire [7:0] __delay_data_1161;
  wire [7:0] __delay_data_1162;
  wire [7:0] __delay_data_1163;
  wire [7:0] __delay_data_1164;
  wire [7:0] __delay_data_1165;
  wire __delay_data_1166;
  wire __delay_data_1167;
  wire __delay_data_1168;
  wire __delay_data_1169;
  wire __delay_data_1170;
  wire __delay_data_1171;
  wire __delay_data_1172;
  wire __delay_data_1173;
  wire __delay_data_1174;
  wire __delay_data_1175;
  wire __delay_data_1176;
  wire __delay_data_1177;
  wire [7:0] __delay_data_1178;
  wire __delay_data_1179;
  wire __delay_data_1180;
  wire __delay_data_1181;
  wire __delay_data_1182;
  wire __delay_data_1183;
  wire __delay_data_1184;
  wire __delay_data_1185;
  wire [3:0] __delay_data_1186;
  wire [3:0] __delay_data_1187;
  wire [3:0] __delay_data_1188;
  wire [3:0] __delay_data_1189;
  wire [3:0] __delay_data_1190;
  wire [3:0] __delay_data_1191;
  wire [3:0] __delay_data_1192;
  wire [3:0] __delay_data_1193;
  wire [7:0] __delay_data_1194;
  wire [7:0] __delay_data_1195;
  wire [7:0] __delay_data_1196;
  wire [7:0] __delay_data_1197;
  wire [7:0] __delay_data_1198;
  wire [7:0] __delay_data_1199;
  wire __delay_data_1200;
  wire __delay_data_1201;
  wire __delay_data_1202;
  wire __delay_data_1203;
  wire __delay_data_1204;
  wire __delay_data_1205;
  wire __delay_data_1206;
  wire __delay_data_1207;
  wire __delay_data_1208;
  wire __delay_data_1209;
  wire __delay_data_1210;
  wire __delay_data_1211;
  wire [7:0] __delay_data_1212;
  wire __delay_data_1213;
  wire __delay_data_1214;
  wire __delay_data_1215;
  wire __delay_data_1216;
  wire __delay_data_1217;
  wire __delay_data_1218;
  wire __delay_data_1219;
  wire [3:0] __delay_data_1220;
  wire [3:0] __delay_data_1221;
  wire [3:0] __delay_data_1222;
  wire [3:0] __delay_data_1223;
  wire [3:0] __delay_data_1224;
  wire [3:0] __delay_data_1225;
  wire [3:0] __delay_data_1226;
  wire [3:0] __delay_data_1227;
  wire [7:0] __delay_data_1228;
  wire [7:0] __delay_data_1229;
  wire [7:0] __delay_data_1230;
  wire [7:0] __delay_data_1231;
  wire [7:0] __delay_data_1232;
  wire [7:0] __delay_data_1233;
  wire __delay_data_1234;
  wire __delay_data_1235;
  wire __delay_data_1236;
  wire __delay_data_1237;
  wire __delay_data_1238;
  wire __delay_data_1239;
  wire __delay_data_1240;
  wire __delay_data_1241;
  wire __delay_data_1242;
  wire __delay_data_1243;
  wire __delay_data_1244;
  wire __delay_data_1245;
  wire [7:0] __delay_data_1246;
  wire __delay_data_1247;
  wire __delay_data_1248;
  wire __delay_data_1249;
  wire __delay_data_1250;
  wire __delay_data_1251;
  wire __delay_data_1252;
  wire __delay_data_1253;
  wire [3:0] __delay_data_1254;
  wire [3:0] __delay_data_1255;
  wire [3:0] __delay_data_1256;
  wire [3:0] __delay_data_1257;
  wire [3:0] __delay_data_1258;
  wire [3:0] __delay_data_1259;
  wire [3:0] __delay_data_1260;
  wire [3:0] __delay_data_1261;
  wire [7:0] __delay_data_1262;
  wire [7:0] __delay_data_1263;
  wire [7:0] __delay_data_1264;
  wire [7:0] __delay_data_1265;
  wire [7:0] __delay_data_1266;
  wire [7:0] __delay_data_1267;
  wire __delay_data_1268;
  wire [7:0] __delay_data_1269;
  wire [7:0] __delay_data_1270;
  wire [7:0] __delay_data_1271;
  wire [7:0] __delay_data_1272;
  wire [7:0] __delay_data_1273;
  wire [7:0] __delay_data_1274;
  wire [7:0] __delay_data_1275;
  wire [7:0] __delay_data_1276;
  wire [7:0] __delay_data_1277;
  wire [7:0] __delay_data_1278;
  wire [7:0] __delay_data_1279;
  wire [7:0] __delay_data_1280;
  wire [7:0] __delay_data_1281;
  wire [7:0] __delay_data_1282;
  wire [7:0] __delay_data_1283;
  wire [7:0] __delay_data_1284;
  wire [7:0] __delay_data_1285;
  wire [7:0] __delay_data_1286;
  wire [7:0] __delay_data_1287;
  wire [7:0] __delay_data_1288;
  wire [5:0] __delay_data_1289;
  wire [5:0] __delay_data_1290;
  wire [5:0] __delay_data_1291;
  wire [5:0] __delay_data_1292;
  wire [5:0] __delay_data_1293;
  wire [5:0] __delay_data_1294;
  wire [5:0] __delay_data_1295;
  wire [5:0] __delay_data_1296;
  wire [5:0] __delay_data_1297;
  wire [5:0] __delay_data_1298;
  wire [5:0] __delay_data_1299;
  wire [5:0] __delay_data_1300;
  wire [5:0] __delay_data_1301;
  wire [5:0] __delay_data_1302;
  wire [5:0] __delay_data_1303;
  wire [5:0] __delay_data_1304;
  wire [5:0] __delay_data_1305;
  wire [5:0] __delay_data_1306;
  wire [5:0] __delay_data_1307;
  wire [5:0] __delay_data_1308;
  wire [5:0] __delay_data_1309;
  wire [5:0] __delay_data_1310;
  wire [7:0] __delay_data_1311;
  wire [7:0] __delay_data_1312;
  wire [7:0] __delay_data_1313;
  wire [7:0] __delay_data_1314;
  wire [7:0] __delay_data_1315;
  wire [7:0] __delay_data_1316;
  wire [7:0] __delay_data_1317;
  wire [7:0] __delay_data_1318;
  wire [7:0] __delay_data_1319;
  wire [7:0] __delay_data_1320;
  wire [7:0] __delay_data_1321;
  wire [7:0] __delay_data_1322;
  wire [7:0] __delay_data_1323;
  wire [7:0] __delay_data_1324;
  wire [7:0] __delay_data_1325;
  wire [7:0] __delay_data_1326;
  wire [7:0] __delay_data_1327;
  wire [7:0] __delay_data_1328;
  wire [7:0] __delay_data_1329;
  wire [7:0] __delay_data_1330;
  wire [7:0] __delay_data_1331;
  wire [7:0] __delay_data_1332;
  wire [7:0] __delay_data_1333;
  wire [7:0] __delay_data_1334;
  wire [7:0] __delay_data_1335;
  wire [7:0] __delay_data_1336;
  wire [7:0] __delay_data_1337;
  wire [7:0] __delay_data_1338;
  wire [3:0] __delay_data_1339;
  wire [7:0] __delay_data_1340;
  wire [7:0] __delay_data_1341;
  wire [7:0] __delay_data_1342;
  wire [7:0] __delay_data_1343;
  wire [7:0] __delay_data_1344;
  wire [7:0] __delay_data_1345;
  wire [7:0] __delay_data_1346;
  wire [7:0] __delay_data_1347;
  wire [7:0] __delay_data_1348;
  wire [7:0] __delay_data_1349;
  wire [7:0] __delay_data_1350;
  wire [7:0] __delay_data_1351;
  wire [7:0] __delay_data_1352;
  wire [7:0] __delay_data_1353;
  wire [7:0] __delay_data_1354;
  wire [7:0] __delay_data_1355;
  wire [7:0] __delay_data_1356;
  wire [7:0] __delay_data_1357;
  wire [7:0] __delay_data_1358;
  wire [7:0] __delay_data_1359;
  wire [7:0] __delay_data_1360;
  wire [7:0] __delay_data_1361;
  wire [7:0] __delay_data_1362;
  wire [7:0] __delay_data_1363;
  wire [7:0] __delay_data_1364;
  wire [7:0] __delay_data_1365;
  wire [7:0] __delay_data_1366;
  wire [7:0] __delay_data_1367;
  wire [7:0] __delay_data_1368;
  wire [7:0] __delay_data_1369;
  wire [7:0] __delay_data_1370;
  wire [7:0] __delay_data_1371;
  wire [7:0] __delay_data_1372;
  wire [7:0] __delay_data_1373;
  wire [7:0] __delay_data_1374;
  wire [7:0] __delay_data_1375;
  wire [7:0] __delay_data_1376;
  wire [7:0] __delay_data_1377;
  wire [7:0] __delay_data_1378;
  wire [7:0] __delay_data_1379;
  wire [7:0] __delay_data_1380;
  wire [7:0] __delay_data_1381;
  wire [7:0] __delay_data_1382;
  wire [7:0] __delay_data_1383;
  wire [7:0] __delay_data_1384;
  wire [7:0] __delay_data_1385;
  wire [7:0] __delay_data_1386;
  wire [7:0] __delay_data_1387;
  wire [7:0] __delay_data_1388;
  wire [7:0] __delay_data_1389;
  wire [7:0] __delay_data_1390;
  wire [7:0] __delay_data_1391;
  wire [7:0] __delay_data_1392;
  wire [7:0] __delay_data_1393;
  wire [7:0] __delay_data_1394;
  wire [7:0] __delay_data_1395;
  wire [7:0] __delay_data_1396;
  wire [7:0] __delay_data_1397;
  wire __delay_data_1398;
  wire __delay_data_1399;
  wire __delay_data_1400;
  wire __delay_data_1401;
  wire __delay_data_1402;
  wire __delay_data_1403;
  wire __delay_data_1404;
  wire __delay_data_1405;
  wire __delay_data_1406;
  wire __delay_data_1407;
  wire __delay_data_1408;
  wire __delay_data_1409;
  wire __delay_data_1410;
  wire [3:0] __delay_data_1411;
  wire [7:0] __delay_data_1412;
  wire [7:0] __delay_data_1413;
  wire [2:0] __delay_data_1414;
  wire [2:0] __delay_data_1415;
  wire [2:0] __delay_data_1416;
  wire [7:0] __delay_data_1417;
  wire __delay_data_1418;
  wire __delay_data_1419;
  wire __delay_data_1420;
  wire __delay_data_1421;
  wire __delay_data_1422;
  wire [3:0] __delay_data_1423;
  wire [3:0] __delay_data_1424;
  wire [3:0] __delay_data_1425;
  wire [3:0] __delay_data_1426;
  wire [7:0] __delay_data_1427;
  wire [7:0] __delay_data_1428;
  wire __delay_data_1429;
  wire [7:0] __delay_data_1430;
  wire [7:0] __delay_data_1431;
  wire [7:0] __delay_data_1432;
  wire [7:0] __delay_data_1433;
  wire [7:0] __delay_data_1434;
  wire [7:0] __delay_data_1435;
  wire [7:0] __delay_data_1436;
  wire [7:0] __delay_data_1437;
  wire [7:0] __delay_data_1438;
  wire [7:0] __delay_data_1439;
  wire [7:0] __delay_data_1440;
  wire [7:0] __delay_data_1441;
  wire [7:0] __delay_data_1442;
  wire [7:0] __delay_data_1443;
  wire [10:0] __delay_data_1444;
  wire [10:0] __delay_data_1445;
  wire [10:0] __delay_data_1446;
  wire [10:0] __delay_data_1447;
  wire [10:0] __delay_data_1448;
  wire [10:0] __delay_data_1449;
  wire [10:0] __delay_data_1450;
  wire [10:0] __delay_data_1451;
  wire [10:0] __delay_data_1452;
  wire [10:0] __delay_data_1453;
  wire [10:0] __delay_data_1454;
  wire [10:0] __delay_data_1455;
  wire [10:0] __delay_data_1456;
  wire [10:0] __delay_data_1457;
  wire [10:0] __delay_data_1458;
  wire [10:0] __delay_data_1459;
  wire [7:0] __delay_data_1460;
  wire [7:0] __delay_data_1461;
  wire [7:0] __delay_data_1462;
  wire [7:0] __delay_data_1463;
  wire [7:0] __delay_data_1464;
  wire [7:0] __delay_data_1465;
  wire [7:0] __delay_data_1466;
  wire [7:0] __delay_data_1467;
  wire [7:0] __delay_data_1468;
  wire [7:0] __delay_data_1469;
  wire [7:0] __delay_data_1470;
  wire [7:0] __delay_data_1471;
  wire [7:0] __delay_data_1472;
  wire [7:0] __delay_data_1473;
  wire [7:0] __delay_data_1474;
  wire [7:0] __delay_data_1475;
  wire [7:0] __delay_data_1476;
  wire [7:0] __delay_data_1477;
  wire [7:0] __delay_data_1478;
  wire [7:0] __delay_data_1479;
  wire [7:0] __delay_data_1480;
  wire [7:0] __delay_data_1481;
  wire [3:0] __delay_data_1482;
  wire [7:0] __delay_data_1483;
  wire [7:0] __delay_data_1484;
  wire [7:0] __delay_data_1485;
  wire [7:0] __delay_data_1486;
  wire [7:0] __delay_data_1487;
  wire [7:0] __delay_data_1488;
  wire [7:0] __delay_data_1489;
  wire [7:0] __delay_data_1490;
  wire [7:0] __delay_data_1491;
  wire [7:0] __delay_data_1492;
  wire [7:0] __delay_data_1493;
  wire [7:0] __delay_data_1494;
  wire [7:0] __delay_data_1495;
  wire [7:0] __delay_data_1496;
  wire [7:0] __delay_data_1497;
  wire [7:0] __delay_data_1498;
  wire [7:0] __delay_data_1499;
  wire [7:0] __delay_data_1500;
  wire [7:0] __delay_data_1501;
  wire [7:0] __delay_data_1502;
  wire [7:0] __delay_data_1503;
  wire [7:0] __delay_data_1504;
  wire [7:0] __delay_data_1505;
  wire [7:0] __delay_data_1506;
  wire [7:0] __delay_data_1507;
  wire [7:0] __delay_data_1508;
  wire [7:0] __delay_data_1509;
  wire [7:0] __delay_data_1510;
  wire [7:0] __delay_data_1511;
  wire [7:0] __delay_data_1512;
  wire [7:0] __delay_data_1513;
  wire [7:0] __delay_data_1514;
  wire [7:0] __delay_data_1515;
  wire [7:0] __delay_data_1516;
  wire [7:0] __delay_data_1517;
  wire [7:0] __delay_data_1518;
  wire [7:0] __delay_data_1519;
  wire [7:0] __delay_data_1520;
  wire [7:0] __delay_data_1521;
  wire [7:0] __delay_data_1522;
  wire [7:0] __delay_data_1523;
  wire [7:0] __delay_data_1524;
  wire [7:0] __delay_data_1525;
  wire [7:0] __delay_data_1526;
  wire [7:0] __delay_data_1527;
  wire [7:0] __delay_data_1528;
  wire __delay_data_1529;
  wire __delay_data_1530;
  wire __delay_data_1531;
  wire __delay_data_1532;
  wire __delay_data_1533;
  wire __delay_data_1534;
  wire __delay_data_1535;
  wire __delay_data_1536;
  wire __delay_data_1537;
  wire __delay_data_1538;
  wire __delay_data_1539;
  wire __delay_data_1540;
  wire __delay_data_1541;
  wire __delay_data_1542;
  wire __delay_data_1543;
  wire __delay_data_1544;
  wire __delay_data_1545;
  wire __delay_data_1546;
  wire __delay_data_1547;
  wire __delay_data_1548;
  wire __delay_data_1549;
  wire __delay_data_1550;
  wire __delay_data_1551;
  wire __delay_data_1552;
  wire __delay_data_1553;
  wire __delay_data_1554;
  wire __delay_data_1555;
  wire __delay_data_1556;
  wire __delay_data_1557;
  wire __delay_data_1558;
  wire __delay_data_1559;
  wire __delay_data_1560;
  wire __delay_data_1561;
  wire __delay_data_1562;
  wire __delay_data_1563;
  wire [7:0] __delay_data_1564;
  wire __delay_data_1565;
  wire __delay_data_1566;
  wire __delay_data_1567;
  wire __delay_data_1568;
  wire __delay_data_1569;
  wire __delay_data_1570;
  wire __delay_data_1571;
  wire __delay_data_1572;
  wire __delay_data_1573;
  wire __delay_data_1574;
  wire __delay_data_1575;
  wire __delay_data_1576;
  wire __delay_data_1577;
  wire __delay_data_1578;
  wire __delay_data_1579;
  wire __delay_data_1580;
  wire __delay_data_1581;
  wire __delay_data_1582;
  wire __delay_data_1583;
  wire __delay_data_1584;
  wire __delay_data_1585;
  wire __delay_data_1586;
  wire __delay_data_1587;
  wire __delay_data_1588;
  wire __delay_data_1589;
  wire __delay_data_1590;
  wire __delay_data_1591;
  wire __delay_data_1592;
  wire __delay_data_1593;
  wire __delay_data_1594;
  wire __delay_data_1595;
  wire __delay_data_1596;
  wire __delay_data_1597;
  wire __delay_data_1598;
  wire __delay_data_1599;
  wire __delay_data_1600;
  wire [7:0] __delay_data_1601;
  wire __delay_data_1602;
  wire __delay_data_1603;
  wire __delay_data_1604;
  wire __delay_data_1605;
  wire __delay_data_1606;
  wire __delay_data_1607;
  wire __delay_data_1608;
  wire __delay_data_1609;
  wire __delay_data_1610;
  wire __delay_data_1611;
  wire __delay_data_1612;
  wire __delay_data_1613;
  wire __delay_data_1614;
  wire __delay_data_1615;
  wire __delay_data_1616;
  wire __delay_data_593;
  wire [7:0] __delay_data_594;
  wire [7:0] __delay_data_595;
  wire [7:0] __delay_data_596;
  wire [3:0] __delay_data_597;
  wire [3:0] __delay_data_598;
  wire [3:0] __delay_data_599;
  wire [3:0] __delay_data_600;
  wire [3:0] __delay_data_601;
  wire [3:0] __delay_data_602;
  wire [3:0] __delay_data_603;
  wire [3:0] __delay_data_604;
  wire [3:0] __delay_data_605;
  wire [3:0] __delay_data_606;
  wire __delay_data_610;
  wire [7:0] __delay_data_611;
  wire [7:0] __delay_data_612;
  wire [7:0] __delay_data_613;
  wire [3:0] __delay_data_614;
  wire [3:0] __delay_data_615;
  wire [3:0] __delay_data_616;
  wire [3:0] __delay_data_617;
  wire [3:0] __delay_data_618;
  wire [3:0] __delay_data_619;
  wire [3:0] __delay_data_620;
  wire [3:0] __delay_data_621;
  wire [3:0] __delay_data_622;
  wire [3:0] __delay_data_623;
  wire __delay_data_627;
  wire [7:0] __delay_data_628;
  wire [7:0] __delay_data_629;
  wire [7:0] __delay_data_630;
  wire [3:0] __delay_data_631;
  wire [3:0] __delay_data_632;
  wire [3:0] __delay_data_633;
  wire [3:0] __delay_data_634;
  wire [3:0] __delay_data_635;
  wire [3:0] __delay_data_636;
  wire [3:0] __delay_data_637;
  wire [3:0] __delay_data_638;
  wire [3:0] __delay_data_639;
  wire [3:0] __delay_data_640;
  wire __delay_data_644;
  wire [7:0] __delay_data_645;
  wire [7:0] __delay_data_646;
  wire [7:0] __delay_data_647;
  wire [3:0] __delay_data_648;
  wire [3:0] __delay_data_649;
  wire [3:0] __delay_data_650;
  wire [3:0] __delay_data_651;
  wire [3:0] __delay_data_652;
  wire [3:0] __delay_data_653;
  wire [3:0] __delay_data_654;
  wire [3:0] __delay_data_655;
  wire [3:0] __delay_data_656;
  wire [3:0] __delay_data_657;
  wire __delay_data_661;
  wire [7:0] __delay_data_662;
  wire [7:0] __delay_data_663;
  wire [7:0] __delay_data_664;
  wire [3:0] __delay_data_665;
  wire [3:0] __delay_data_666;
  wire [3:0] __delay_data_667;
  wire [3:0] __delay_data_668;
  wire [3:0] __delay_data_669;
  wire [3:0] __delay_data_670;
  wire [3:0] __delay_data_671;
  wire [3:0] __delay_data_672;
  wire [3:0] __delay_data_673;
  wire [3:0] __delay_data_674;
  wire __delay_data_678;
  wire [7:0] __delay_data_679;
  wire [7:0] __delay_data_680;
  wire [7:0] __delay_data_681;
  wire [3:0] __delay_data_682;
  wire [3:0] __delay_data_683;
  wire [3:0] __delay_data_684;
  wire [3:0] __delay_data_685;
  wire [3:0] __delay_data_686;
  wire [3:0] __delay_data_687;
  wire [3:0] __delay_data_688;
  wire [3:0] __delay_data_689;
  wire [3:0] __delay_data_690;
  wire [3:0] __delay_data_691;
  wire __delay_data_695;
  wire [7:0] __delay_data_696;
  wire [7:0] __delay_data_697;
  wire [7:0] __delay_data_698;
  wire [3:0] __delay_data_699;
  wire [3:0] __delay_data_700;
  wire [3:0] __delay_data_701;
  wire [3:0] __delay_data_702;
  wire [3:0] __delay_data_703;
  wire [3:0] __delay_data_704;
  wire [3:0] __delay_data_705;
  wire [3:0] __delay_data_706;
  wire [3:0] __delay_data_707;
  wire [3:0] __delay_data_708;
  wire __delay_data_712;
  wire [7:0] __delay_data_713;
  wire [7:0] __delay_data_714;
  wire [7:0] __delay_data_715;
  wire [3:0] __delay_data_716;
  wire [3:0] __delay_data_717;
  wire [3:0] __delay_data_718;
  wire [3:0] __delay_data_719;
  wire [3:0] __delay_data_720;
  wire [3:0] __delay_data_721;
  wire [3:0] __delay_data_722;
  wire [3:0] __delay_data_723;
  wire [3:0] __delay_data_724;
  wire [3:0] __delay_data_725;
  wire __delay_data_729;
  wire [7:0] __delay_data_730;
  wire [7:0] __delay_data_731;
  wire [7:0] __delay_data_732;
  wire [3:0] __delay_data_733;
  wire [3:0] __delay_data_734;
  wire [3:0] __delay_data_735;
  wire [3:0] __delay_data_736;
  wire [3:0] __delay_data_737;
  wire [3:0] __delay_data_738;
  wire [3:0] __delay_data_739;
  wire [3:0] __delay_data_740;
  wire [3:0] __delay_data_741;
  wire [3:0] __delay_data_742;
  wire __delay_data_748;
  wire [31:0] __delay_data_749;
  wire [31:0] __delay_data_750;
  wire [5:0] __delay_data_751;
  wire [5:0] __delay_data_752;
  wire [5:0] __delay_data_753;
  wire [5:0] __delay_data_754;
  wire __delay_data_755;
  wire __delay_data_756;
  wire __delay_data_757;
  wire __delay_data_758;
  wire [5:0] __delay_data_764;
  wire [5:0] __delay_data_765;
  wire [5:0] __delay_data_766;
  wire [5:0] __delay_data_767;
  wire [39:0] __delay_data_768;
  wire __delay_data_769;
  wire [7:0] __delay_data_898;
  wire __delay_data_899;
  wire [7:0] __delay_data_900;
  wire [7:0] __delay_data_901;
  wire __delay_data_902;
  wire __delay_data_903;
  wire [7:0] __delay_data_904;
  wire [7:0] __delay_data_905;
  wire [7:0] __delay_data_906;
  wire [7:0] __delay_data_907;
  wire __delay_data_908;
  wire [7:0] __delay_data_909;
  wire [7:0] __delay_data_910;
  wire __delay_data_911;
  wire __delay_data_912;
  wire [7:0] __delay_data_913;
  wire [7:0] __delay_data_914;
  wire [7:0] __delay_data_915;
  wire [7:0] __delay_data_916;
  wire __delay_data_917;
  wire [7:0] __delay_data_918;
  wire [7:0] __delay_data_919;
  wire __delay_data_920;
  wire __delay_data_921;
  wire [7:0] __delay_data_922;
  wire [7:0] __delay_data_923;
  wire [7:0] __delay_data_924;
  wire __delay_data_925;
  wire __delay_data_926;
  wire __delay_data_927;
  wire __delay_data_928;
  wire __delay_data_929;
  wire __delay_data_930;
  wire __delay_data_931;
  wire [7:0] __delay_data_932;
  wire __delay_data_933;
  wire __delay_data_934;
  wire __delay_data_935;
  wire __delay_data_936;
  wire __delay_data_937;
  wire [7:0] __delay_data_938;
  wire [7:0] __delay_data_939;
  wire __delay_data_940;
  wire __delay_data_941;
  wire __delay_data_942;
  wire __delay_data_943;
  wire __delay_data_944;
  wire __delay_data_945;
  wire __delay_data_946;
  wire __delay_data_947;
  wire [3:0] __delay_data_948;
  wire [3:0] __delay_data_949;
  wire [3:0] __delay_data_950;
  wire [3:0] __delay_data_951;
  wire [3:0] __delay_data_952;
  wire [3:0] __delay_data_953;
  wire [3:0] __delay_data_954;
  wire [3:0] __delay_data_955;
  wire [7:0] __delay_data_956;
  wire [7:0] __delay_data_957;
  wire [7:0] __delay_data_958;
  wire [7:0] __delay_data_959;
  wire [7:0] __delay_data_960;
  wire [7:0] __delay_data_961;
  wire __delay_data_962;
  wire [7:0] __delay_data_963;
  wire __delay_data_964;
  wire __delay_data_965;
  wire [7:0] __delay_data_966;
  wire __delay_data_967;
  wire [7:0] __delay_data_968;
  wire __delay_data_969;
  wire __delay_data_970;
  wire [7:0] __delay_data_971;
  wire __delay_data_972;
  wire [7:0] __delay_data_973;
  wire __delay_data_974;
  wire __delay_data_975;
  wire [7:0] __delay_data_976;
  wire __delay_data_977;
  wire __delay_data_978;
  wire __delay_data_979;
  wire __delay_data_980;
  wire __delay_data_981;
  wire __delay_data_982;
  wire __delay_data_983;
  wire [7:0] __delay_data_984;
  wire __delay_data_985;
  wire __delay_data_986;
  wire __delay_data_987;
  wire __delay_data_988;
  wire __delay_data_989;
  wire [7:0] __delay_data_990;
  wire [7:0] __delay_data_991;
  wire __delay_data_992;
  wire __delay_data_993;
  wire __delay_data_994;
  wire __delay_data_995;
  wire __delay_data_996;
  wire __delay_data_997;
  wire __delay_data_998;
  wire [3:0] __delay_data_999;
  wire __maxi_read_fsm_cond_3_0_1;
  wire __maxi_read_fsm_cond_3_2_1;
  wire __maxi_read_fsm_cond_3_3_1;
  wire __maxi_read_fsm_cond_3_4_1;
  wire __maxi_read_fsm_cond_3_5_1;
  wire __maxi_read_fsm_cond_3_6_1;
  wire __maxi_read_fsm_cond_3_7_1;
  wire __maxi_read_fsm_cond_3_8_1;
  wire __maxi_read_fsm_cond_3_9_1;
  wire __maxi_read_fsm_cond_4_1_1;
  wire __maxi_write_fsm_cond_4_0_1;
  wire [11:0] __muladd_data_103;
  wire [11:0] __muladd_data_120;
  wire [11:0] __muladd_data_137;
  wire [11:0] __muladd_data_154;
  wire [11:0] __muladd_data_171;
  wire [11:0] __muladd_data_188;
  wire [11:0] __muladd_data_205;
  wire [11:0] __muladd_data_69;
  wire [11:0] __muladd_data_86;
  wire \__muladd_madd_103.CLK ;
  wire [7:0] \__muladd_madd_103.a ;
  wire [3:0] \__muladd_madd_103.b ;
  wire [11:0] \__muladd_madd_103.c ;
  wire [11:0] \__muladd_madd_103.d ;
  wire \__muladd_madd_103.madd.CLK ;
  wire [7:0] \__muladd_madd_103.madd._a ;
  wire [3:0] \__muladd_madd_103.madd._b ;
  wire [11:0] \__muladd_madd_103.madd._c ;
  wire [11:0] \__muladd_madd_103.madd._madd ;
  wire [11:0] \__muladd_madd_103.madd._mul ;
  wire [11:0] \__muladd_madd_103.madd._pipe_madd0 ;
  wire [11:0] \__muladd_madd_103.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_103.madd.a ;
  wire [3:0] \__muladd_madd_103.madd.b ;
  wire [11:0] \__muladd_madd_103.madd.c ;
  wire [11:0] \__muladd_madd_103.madd.d ;
  wire \__muladd_madd_103.madd.update ;
  wire \__muladd_madd_103.update ;
  wire \__muladd_madd_120.CLK ;
  wire [7:0] \__muladd_madd_120.a ;
  wire [3:0] \__muladd_madd_120.b ;
  wire [11:0] \__muladd_madd_120.c ;
  wire [11:0] \__muladd_madd_120.d ;
  wire \__muladd_madd_120.madd.CLK ;
  wire [7:0] \__muladd_madd_120.madd._a ;
  wire [3:0] \__muladd_madd_120.madd._b ;
  wire [11:0] \__muladd_madd_120.madd._c ;
  wire [11:0] \__muladd_madd_120.madd._madd ;
  wire [11:0] \__muladd_madd_120.madd._mul ;
  wire [11:0] \__muladd_madd_120.madd._pipe_madd0 ;
  wire [11:0] \__muladd_madd_120.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_120.madd.a ;
  wire [3:0] \__muladd_madd_120.madd.b ;
  wire [11:0] \__muladd_madd_120.madd.c ;
  wire [11:0] \__muladd_madd_120.madd.d ;
  wire \__muladd_madd_120.madd.update ;
  wire \__muladd_madd_120.update ;
  wire \__muladd_madd_137.CLK ;
  wire [7:0] \__muladd_madd_137.a ;
  wire [3:0] \__muladd_madd_137.b ;
  wire [11:0] \__muladd_madd_137.c ;
  wire [11:0] \__muladd_madd_137.d ;
  wire \__muladd_madd_137.madd.CLK ;
  wire [7:0] \__muladd_madd_137.madd._a ;
  wire [3:0] \__muladd_madd_137.madd._b ;
  wire [11:0] \__muladd_madd_137.madd._c ;
  wire [11:0] \__muladd_madd_137.madd._madd ;
  wire [11:0] \__muladd_madd_137.madd._mul ;
  wire [11:0] \__muladd_madd_137.madd._pipe_madd0 ;
  wire [11:0] \__muladd_madd_137.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_137.madd.a ;
  wire [3:0] \__muladd_madd_137.madd.b ;
  wire [11:0] \__muladd_madd_137.madd.c ;
  wire [11:0] \__muladd_madd_137.madd.d ;
  wire \__muladd_madd_137.madd.update ;
  wire \__muladd_madd_137.update ;
  wire \__muladd_madd_154.CLK ;
  wire [7:0] \__muladd_madd_154.a ;
  wire [3:0] \__muladd_madd_154.b ;
  wire [11:0] \__muladd_madd_154.c ;
  wire [11:0] \__muladd_madd_154.d ;
  wire \__muladd_madd_154.madd.CLK ;
  wire [7:0] \__muladd_madd_154.madd._a ;
  wire [3:0] \__muladd_madd_154.madd._b ;
  wire [11:0] \__muladd_madd_154.madd._c ;
  wire [11:0] \__muladd_madd_154.madd._madd ;
  wire [11:0] \__muladd_madd_154.madd._mul ;
  wire [11:0] \__muladd_madd_154.madd._pipe_madd0 ;
  wire [11:0] \__muladd_madd_154.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_154.madd.a ;
  wire [3:0] \__muladd_madd_154.madd.b ;
  wire [11:0] \__muladd_madd_154.madd.c ;
  wire [11:0] \__muladd_madd_154.madd.d ;
  wire \__muladd_madd_154.madd.update ;
  wire \__muladd_madd_154.update ;
  wire \__muladd_madd_171.CLK ;
  wire [7:0] \__muladd_madd_171.a ;
  wire [3:0] \__muladd_madd_171.b ;
  wire [11:0] \__muladd_madd_171.c ;
  wire [11:0] \__muladd_madd_171.d ;
  wire \__muladd_madd_171.madd.CLK ;
  wire [7:0] \__muladd_madd_171.madd._a ;
  wire [3:0] \__muladd_madd_171.madd._b ;
  wire [11:0] \__muladd_madd_171.madd._c ;
  wire [11:0] \__muladd_madd_171.madd._madd ;
  wire [11:0] \__muladd_madd_171.madd._mul ;
  wire [11:0] \__muladd_madd_171.madd._pipe_madd0 ;
  wire [11:0] \__muladd_madd_171.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_171.madd.a ;
  wire [3:0] \__muladd_madd_171.madd.b ;
  wire [11:0] \__muladd_madd_171.madd.c ;
  wire [11:0] \__muladd_madd_171.madd.d ;
  wire \__muladd_madd_171.madd.update ;
  wire \__muladd_madd_171.update ;
  wire \__muladd_madd_188.CLK ;
  wire [7:0] \__muladd_madd_188.a ;
  wire [3:0] \__muladd_madd_188.b ;
  wire [11:0] \__muladd_madd_188.c ;
  wire [11:0] \__muladd_madd_188.d ;
  wire \__muladd_madd_188.madd.CLK ;
  wire [7:0] \__muladd_madd_188.madd._a ;
  wire [3:0] \__muladd_madd_188.madd._b ;
  wire [11:0] \__muladd_madd_188.madd._c ;
  wire [11:0] \__muladd_madd_188.madd._madd ;
  wire [11:0] \__muladd_madd_188.madd._mul ;
  wire [11:0] \__muladd_madd_188.madd._pipe_madd0 ;
  wire [11:0] \__muladd_madd_188.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_188.madd.a ;
  wire [3:0] \__muladd_madd_188.madd.b ;
  wire [11:0] \__muladd_madd_188.madd.c ;
  wire [11:0] \__muladd_madd_188.madd.d ;
  wire \__muladd_madd_188.madd.update ;
  wire \__muladd_madd_188.update ;
  wire \__muladd_madd_205.CLK ;
  wire [7:0] \__muladd_madd_205.a ;
  wire [3:0] \__muladd_madd_205.b ;
  wire [11:0] \__muladd_madd_205.c ;
  wire [11:0] \__muladd_madd_205.d ;
  wire \__muladd_madd_205.madd.CLK ;
  wire [7:0] \__muladd_madd_205.madd._a ;
  wire [3:0] \__muladd_madd_205.madd._b ;
  wire [11:0] \__muladd_madd_205.madd._c ;
  wire [11:0] \__muladd_madd_205.madd._madd ;
  wire [11:0] \__muladd_madd_205.madd._mul ;
  wire [11:0] \__muladd_madd_205.madd._pipe_madd0 ;
  wire [11:0] \__muladd_madd_205.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_205.madd.a ;
  wire [3:0] \__muladd_madd_205.madd.b ;
  wire [11:0] \__muladd_madd_205.madd.c ;
  wire [11:0] \__muladd_madd_205.madd.d ;
  wire \__muladd_madd_205.madd.update ;
  wire \__muladd_madd_205.update ;
  wire \__muladd_madd_69.CLK ;
  wire [7:0] \__muladd_madd_69.a ;
  wire [3:0] \__muladd_madd_69.b ;
  wire [11:0] \__muladd_madd_69.c ;
  wire [11:0] \__muladd_madd_69.d ;
  wire \__muladd_madd_69.madd.CLK ;
  wire [7:0] \__muladd_madd_69.madd._a ;
  wire [3:0] \__muladd_madd_69.madd._b ;
  wire [11:0] \__muladd_madd_69.madd._c ;
  wire [11:0] \__muladd_madd_69.madd._madd ;
  wire [11:0] \__muladd_madd_69.madd._mul ;
  wire [11:0] \__muladd_madd_69.madd._pipe_madd0 ;
  wire [11:0] \__muladd_madd_69.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_69.madd.a ;
  wire [3:0] \__muladd_madd_69.madd.b ;
  wire [11:0] \__muladd_madd_69.madd.c ;
  wire [11:0] \__muladd_madd_69.madd.d ;
  wire \__muladd_madd_69.madd.update ;
  wire \__muladd_madd_69.update ;
  wire \__muladd_madd_86.CLK ;
  wire [7:0] \__muladd_madd_86.a ;
  wire [3:0] \__muladd_madd_86.b ;
  wire [11:0] \__muladd_madd_86.c ;
  wire [11:0] \__muladd_madd_86.d ;
  wire \__muladd_madd_86.madd.CLK ;
  wire [7:0] \__muladd_madd_86.madd._a ;
  wire [3:0] \__muladd_madd_86.madd._b ;
  wire [11:0] \__muladd_madd_86.madd._c ;
  wire [11:0] \__muladd_madd_86.madd._madd ;
  wire [11:0] \__muladd_madd_86.madd._mul ;
  wire [11:0] \__muladd_madd_86.madd._pipe_madd0 ;
  wire [11:0] \__muladd_madd_86.madd._pipe_madd1 ;
  wire [7:0] \__muladd_madd_86.madd.a ;
  wire [3:0] \__muladd_madd_86.madd.b ;
  wire [11:0] \__muladd_madd_86.madd.c ;
  wire [11:0] \__muladd_madd_86.madd.d ;
  wire \__muladd_madd_86.madd.update ;
  wire \__muladd_madd_86.update ;
  wire [11:0] __muladd_madd_odata_103;
  wire [11:0] __muladd_madd_odata_120;
  wire [11:0] __muladd_madd_odata_137;
  wire [11:0] __muladd_madd_odata_154;
  wire [11:0] __muladd_madd_odata_171;
  wire [11:0] __muladd_madd_odata_188;
  wire [11:0] __muladd_madd_odata_205;
  wire [11:0] __muladd_madd_odata_69;
  wire [11:0] __muladd_madd_odata_86;
  wire [11:0] __muladd_madd_odata_reg_103;
  wire [11:0] __muladd_madd_odata_reg_120;
  wire [11:0] __muladd_madd_odata_reg_137;
  wire [11:0] __muladd_madd_odata_reg_154;
  wire [11:0] __muladd_madd_odata_reg_171;
  wire [11:0] __muladd_madd_odata_reg_188;
  wire [11:0] __muladd_madd_odata_reg_205;
  wire [11:0] __muladd_madd_odata_reg_69;
  wire [11:0] __muladd_madd_odata_reg_86;
  wire __muladd_madd_update_103;
  wire __muladd_madd_update_120;
  wire __muladd_madd_update_137;
  wire __muladd_madd_update_154;
  wire __muladd_madd_update_171;
  wire __muladd_madd_update_188;
  wire __muladd_madd_update_205;
  wire __muladd_madd_update_69;
  wire __muladd_madd_update_86;
  wire [31:0] __plusn_data_34;
  wire [31:0] __plusn_data_35;
  wire [31:0] __plusn_data_36;
  wire [31:0] __plusn_data_37;
  wire __reduce_max_13_data_sink_wenable;
  wire [31:0] __reduce_max_13_fsm;
  wire __reduce_max_13_reduce_reset;
  wire __reduce_max_13_valid_sink_wenable;
  wire __reduce_max_13_x_idle;
  wire __reduce_max_13_x_source_ram_rvalid;
  wire __set_flag_1036_1;
  wire __set_flag_1036_2;
  wire __set_flag_1036_3;
  wire __set_flag_1036_4;
  wire __set_flag_1036_5;
  wire __set_flag_1036_6;
  wire __set_flag_1036_7;
  wire __set_flag_1036_8;
  wire __set_flag_1036_9;
  wire __set_flag_1224_1;
  wire __set_flag_1224_10;
  wire __set_flag_1224_11;
  wire __set_flag_1224_12;
  wire __set_flag_1224_13;
  wire __set_flag_1224_14;
  wire __set_flag_1224_15;
  wire __set_flag_1224_16;
  wire __set_flag_1224_17;
  wire __set_flag_1224_18;
  wire __set_flag_1224_19;
  wire __set_flag_1224_2;
  wire __set_flag_1224_20;
  wire __set_flag_1224_21;
  wire __set_flag_1224_22;
  wire __set_flag_1224_23;
  wire __set_flag_1224_24;
  wire __set_flag_1224_25;
  wire __set_flag_1224_26;
  wire __set_flag_1224_27;
  wire __set_flag_1224_28;
  wire __set_flag_1224_29;
  wire __set_flag_1224_3;
  wire __set_flag_1224_30;
  wire __set_flag_1224_31;
  wire __set_flag_1224_32;
  wire __set_flag_1224_33;
  wire __set_flag_1224_34;
  wire __set_flag_1224_35;
  wire __set_flag_1224_36;
  wire __set_flag_1224_37;
  wire __set_flag_1224_38;
  wire __set_flag_1224_39;
  wire __set_flag_1224_4;
  wire __set_flag_1224_40;
  wire __set_flag_1224_41;
  wire __set_flag_1224_5;
  wire __set_flag_1224_6;
  wire __set_flag_1224_7;
  wire __set_flag_1224_8;
  wire __set_flag_1224_9;
  wire __set_flag_710_1;
  wire __set_flag_710_10;
  wire __set_flag_710_11;
  wire __set_flag_710_12;
  wire __set_flag_710_13;
  wire __set_flag_710_14;
  wire __set_flag_710_15;
  wire __set_flag_710_16;
  wire __set_flag_710_17;
  wire __set_flag_710_18;
  wire __set_flag_710_19;
  wire __set_flag_710_2;
  wire __set_flag_710_20;
  wire __set_flag_710_21;
  wire __set_flag_710_22;
  wire __set_flag_710_23;
  wire __set_flag_710_24;
  wire __set_flag_710_25;
  wire __set_flag_710_26;
  wire __set_flag_710_27;
  wire __set_flag_710_28;
  wire __set_flag_710_29;
  wire __set_flag_710_3;
  wire __set_flag_710_30;
  wire __set_flag_710_31;
  wire __set_flag_710_32;
  wire __set_flag_710_33;
  wire __set_flag_710_34;
  wire __set_flag_710_35;
  wire __set_flag_710_36;
  wire __set_flag_710_37;
  wire __set_flag_710_38;
  wire __set_flag_710_39;
  wire __set_flag_710_4;
  wire __set_flag_710_40;
  wire __set_flag_710_41;
  wire __set_flag_710_42;
  wire __set_flag_710_43;
  wire __set_flag_710_44;
  wire __set_flag_710_45;
  wire __set_flag_710_5;
  wire __set_flag_710_6;
  wire __set_flag_710_7;
  wire __set_flag_710_8;
  wire __set_flag_710_9;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_1;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_10;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_11;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_12;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_13;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_14;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_15;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_16;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_17;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_18;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_19;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_2;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_20;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_21;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_22;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_23;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_24;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_25;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_26;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_27;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_28;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_29;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_3;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_30;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_31;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_32;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_33;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_34;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_35;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_36;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_37;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_38;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_39;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_4;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_40;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_41;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_42;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_43;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_44;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_45;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_5;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_6;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_7;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_8;
  wire [31:0] __stream_conv2d_16_sink_37_sink_offset_0_9;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_1;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_10;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_11;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_12;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_13;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_14;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_15;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_16;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_17;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_18;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_19;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_2;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_20;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_21;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_22;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_23;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_24;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_25;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_26;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_27;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_28;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_29;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_3;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_30;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_31;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_32;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_33;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_34;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_35;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_36;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_37;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_38;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_39;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_4;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_40;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_41;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_42;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_43;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_44;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_45;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_5;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_6;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_7;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_8;
  wire [32:0] __stream_conv2d_16_sink_37_sink_size_1_9;
  wire __stream_conv2d_16_start_1;
  wire __stream_conv2d_16_start_10;
  wire __stream_conv2d_16_start_11;
  wire __stream_conv2d_16_start_12;
  wire __stream_conv2d_16_start_13;
  wire __stream_conv2d_16_start_14;
  wire __stream_conv2d_16_start_15;
  wire __stream_conv2d_16_start_16;
  wire __stream_conv2d_16_start_17;
  wire __stream_conv2d_16_start_18;
  wire __stream_conv2d_16_start_19;
  wire __stream_conv2d_16_start_2;
  wire __stream_conv2d_16_start_20;
  wire __stream_conv2d_16_start_21;
  wire __stream_conv2d_16_start_22;
  wire __stream_conv2d_16_start_23;
  wire __stream_conv2d_16_start_24;
  wire __stream_conv2d_16_start_25;
  wire __stream_conv2d_16_start_26;
  wire __stream_conv2d_16_start_27;
  wire __stream_conv2d_16_start_28;
  wire __stream_conv2d_16_start_29;
  wire __stream_conv2d_16_start_3;
  wire __stream_conv2d_16_start_30;
  wire __stream_conv2d_16_start_31;
  wire __stream_conv2d_16_start_32;
  wire __stream_conv2d_16_start_33;
  wire __stream_conv2d_16_start_34;
  wire __stream_conv2d_16_start_35;
  wire __stream_conv2d_16_start_36;
  wire __stream_conv2d_16_start_37;
  wire __stream_conv2d_16_start_38;
  wire __stream_conv2d_16_start_39;
  wire __stream_conv2d_16_start_4;
  wire __stream_conv2d_16_start_40;
  wire __stream_conv2d_16_start_41;
  wire __stream_conv2d_16_start_42;
  wire __stream_conv2d_16_start_43;
  wire __stream_conv2d_16_start_44;
  wire __stream_conv2d_16_start_45;
  wire __stream_conv2d_16_start_46;
  wire __stream_conv2d_16_start_5;
  wire __stream_conv2d_16_start_6;
  wire __stream_conv2d_16_start_7;
  wire __stream_conv2d_16_start_8;
  wire __stream_conv2d_16_start_9;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_1;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_10;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_11;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_12;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_13;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_14;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_15;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_16;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_17;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_18;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_19;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_2;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_20;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_21;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_22;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_23;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_24;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_25;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_26;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_27;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_28;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_29;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_3;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_30;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_31;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_32;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_33;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_34;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_35;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_36;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_37;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_38;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_39;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_4;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_40;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_41;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_5;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_6;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_7;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_8;
  wire [31:0] __stream_matmul_29_sink_21_sink_offset_0_9;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_1;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_10;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_11;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_12;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_13;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_14;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_15;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_16;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_17;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_18;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_19;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_2;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_20;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_21;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_22;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_23;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_24;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_25;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_26;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_27;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_28;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_29;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_3;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_30;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_31;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_32;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_33;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_34;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_35;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_36;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_37;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_38;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_39;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_4;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_40;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_41;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_5;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_6;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_7;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_8;
  wire [32:0] __stream_matmul_29_sink_21_sink_size_1_9;
  wire __stream_matmul_29_start_1;
  wire __stream_matmul_29_start_10;
  wire __stream_matmul_29_start_11;
  wire __stream_matmul_29_start_12;
  wire __stream_matmul_29_start_13;
  wire __stream_matmul_29_start_14;
  wire __stream_matmul_29_start_15;
  wire __stream_matmul_29_start_16;
  wire __stream_matmul_29_start_17;
  wire __stream_matmul_29_start_18;
  wire __stream_matmul_29_start_19;
  wire __stream_matmul_29_start_2;
  wire __stream_matmul_29_start_20;
  wire __stream_matmul_29_start_21;
  wire __stream_matmul_29_start_22;
  wire __stream_matmul_29_start_23;
  wire __stream_matmul_29_start_24;
  wire __stream_matmul_29_start_25;
  wire __stream_matmul_29_start_26;
  wire __stream_matmul_29_start_27;
  wire __stream_matmul_29_start_28;
  wire __stream_matmul_29_start_29;
  wire __stream_matmul_29_start_3;
  wire __stream_matmul_29_start_30;
  wire __stream_matmul_29_start_31;
  wire __stream_matmul_29_start_32;
  wire __stream_matmul_29_start_33;
  wire __stream_matmul_29_start_34;
  wire __stream_matmul_29_start_35;
  wire __stream_matmul_29_start_36;
  wire __stream_matmul_29_start_37;
  wire __stream_matmul_29_start_38;
  wire __stream_matmul_29_start_39;
  wire __stream_matmul_29_start_4;
  wire __stream_matmul_29_start_40;
  wire __stream_matmul_29_start_41;
  wire __stream_matmul_29_start_42;
  wire __stream_matmul_29_start_5;
  wire __stream_matmul_29_start_6;
  wire __stream_matmul_29_start_7;
  wire __stream_matmul_29_start_8;
  wire __stream_matmul_29_start_9;
  wire [31:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_1;
  wire [31:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_2;
  wire [31:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_3;
  wire [31:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_4;
  wire [31:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_5;
  wire [31:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_6;
  wire [31:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_7;
  wire [31:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_8;
  wire [31:0] __stream_max_pool_serial_18_sink_3_sink_offset_0_9;
  wire [32:0] __stream_max_pool_serial_18_sink_3_sink_size_1_1;
  wire [32:0] __stream_max_pool_serial_18_sink_3_sink_size_1_2;
  wire [32:0] __stream_max_pool_serial_18_sink_3_sink_size_1_3;
  wire [32:0] __stream_max_pool_serial_18_sink_3_sink_size_1_4;
  wire [32:0] __stream_max_pool_serial_18_sink_3_sink_size_1_5;
  wire [32:0] __stream_max_pool_serial_18_sink_3_sink_size_1_6;
  wire [32:0] __stream_max_pool_serial_18_sink_3_sink_size_1_7;
  wire [32:0] __stream_max_pool_serial_18_sink_3_sink_size_1_8;
  wire [32:0] __stream_max_pool_serial_18_sink_3_sink_size_1_9;
  wire __stream_max_pool_serial_18_start_1;
  wire __stream_max_pool_serial_18_start_10;
  wire __stream_max_pool_serial_18_start_2;
  wire __stream_max_pool_serial_18_start_3;
  wire __stream_max_pool_serial_18_start_4;
  wire __stream_max_pool_serial_18_start_5;
  wire __stream_max_pool_serial_18_start_6;
  wire __stream_max_pool_serial_18_start_7;
  wire __stream_max_pool_serial_18_start_8;
  wire __stream_max_pool_serial_18_start_9;
  wire __stream_seq_14_cond_2_1;
  wire __stream_seq_14_cond_2_10;
  wire __stream_seq_14_cond_2_11;
  wire __stream_seq_14_cond_2_12;
  wire __stream_seq_14_cond_2_13;
  wire __stream_seq_14_cond_2_14;
  wire __stream_seq_14_cond_2_15;
  wire __stream_seq_14_cond_2_16;
  wire __stream_seq_14_cond_2_17;
  wire __stream_seq_14_cond_2_18;
  wire __stream_seq_14_cond_2_19;
  wire __stream_seq_14_cond_2_2;
  wire __stream_seq_14_cond_2_20;
  wire __stream_seq_14_cond_2_21;
  wire __stream_seq_14_cond_2_22;
  wire __stream_seq_14_cond_2_23;
  wire __stream_seq_14_cond_2_24;
  wire __stream_seq_14_cond_2_25;
  wire __stream_seq_14_cond_2_26;
  wire __stream_seq_14_cond_2_27;
  wire __stream_seq_14_cond_2_28;
  wire __stream_seq_14_cond_2_29;
  wire __stream_seq_14_cond_2_3;
  wire __stream_seq_14_cond_2_30;
  wire __stream_seq_14_cond_2_31;
  wire __stream_seq_14_cond_2_32;
  wire __stream_seq_14_cond_2_33;
  wire __stream_seq_14_cond_2_34;
  wire __stream_seq_14_cond_2_35;
  wire __stream_seq_14_cond_2_36;
  wire __stream_seq_14_cond_2_37;
  wire __stream_seq_14_cond_2_38;
  wire __stream_seq_14_cond_2_39;
  wire __stream_seq_14_cond_2_4;
  wire __stream_seq_14_cond_2_40;
  wire __stream_seq_14_cond_2_41;
  wire __stream_seq_14_cond_2_42;
  wire __stream_seq_14_cond_2_43;
  wire __stream_seq_14_cond_2_44;
  wire __stream_seq_14_cond_2_45;
  wire __stream_seq_14_cond_2_5;
  wire __stream_seq_14_cond_2_6;
  wire __stream_seq_14_cond_2_7;
  wire __stream_seq_14_cond_2_8;
  wire __stream_seq_14_cond_2_9;
  wire __stream_seq_15_cond_2_1;
  wire __stream_seq_15_cond_2_2;
  wire __stream_seq_15_cond_2_3;
  wire __stream_seq_15_cond_2_4;
  wire __stream_seq_15_cond_2_5;
  wire __stream_seq_15_cond_2_6;
  wire __stream_seq_15_cond_2_7;
  wire __stream_seq_15_cond_2_8;
  wire __stream_seq_15_cond_2_9;
  wire __stream_seq_16_cond_2_1;
  wire __stream_seq_16_cond_2_10;
  wire __stream_seq_16_cond_2_11;
  wire __stream_seq_16_cond_2_12;
  wire __stream_seq_16_cond_2_13;
  wire __stream_seq_16_cond_2_14;
  wire __stream_seq_16_cond_2_15;
  wire __stream_seq_16_cond_2_16;
  wire __stream_seq_16_cond_2_17;
  wire __stream_seq_16_cond_2_18;
  wire __stream_seq_16_cond_2_19;
  wire __stream_seq_16_cond_2_2;
  wire __stream_seq_16_cond_2_20;
  wire __stream_seq_16_cond_2_21;
  wire __stream_seq_16_cond_2_22;
  wire __stream_seq_16_cond_2_23;
  wire __stream_seq_16_cond_2_24;
  wire __stream_seq_16_cond_2_25;
  wire __stream_seq_16_cond_2_26;
  wire __stream_seq_16_cond_2_27;
  wire __stream_seq_16_cond_2_28;
  wire __stream_seq_16_cond_2_29;
  wire __stream_seq_16_cond_2_3;
  wire __stream_seq_16_cond_2_30;
  wire __stream_seq_16_cond_2_31;
  wire __stream_seq_16_cond_2_32;
  wire __stream_seq_16_cond_2_33;
  wire __stream_seq_16_cond_2_34;
  wire __stream_seq_16_cond_2_35;
  wire __stream_seq_16_cond_2_36;
  wire __stream_seq_16_cond_2_37;
  wire __stream_seq_16_cond_2_38;
  wire __stream_seq_16_cond_2_39;
  wire __stream_seq_16_cond_2_4;
  wire __stream_seq_16_cond_2_40;
  wire __stream_seq_16_cond_2_41;
  wire __stream_seq_16_cond_2_5;
  wire __stream_seq_16_cond_2_6;
  wire __stream_seq_16_cond_2_7;
  wire __stream_seq_16_cond_2_8;
  wire __stream_seq_16_cond_2_9;
  wire [11:0] __substreamoutput_data_608;
  wire [11:0] __substreamoutput_data_625;
  wire [11:0] __substreamoutput_data_642;
  wire [11:0] __substreamoutput_data_659;
  wire [11:0] __substreamoutput_data_676;
  wire [11:0] __substreamoutput_data_693;
  wire [11:0] __substreamoutput_data_710;
  wire [11:0] __substreamoutput_data_727;
  wire [11:0] __substreamoutput_data_744;
  wire [31:0] __substreamoutput_data_746;
  wire [31:0] __substreamoutput_data_760;
  wire __substreamoutput_data_761;
  wire [7:0] __substreamoutput_data_771;
  wire [7:0] __substreamoutput_data_793;
  wire __substreamoutput_data_794;
  wire [11:0] __substreamoutput_data_876;
  wire [31:0] __substreamoutput_data_878;
  wire [31:0] __substreamoutput_data_881;
  wire __substreamoutput_data_882;
  wire [7:0] __substreamoutput_data_886;
  wire __tmp_1000_1;
  wire [7:0] __tmp_1001_1;
  wire __tmp_1012_1;
  wire [7:0] __tmp_1013_1;
  wire [1:0] __tmp_1027_1;
  wire [1:0] __tmp_1027_2;
  wire __tmp_1035_1;
  wire __tmp_1040_1;
  wire __tmp_1040_2;
  wire __tmp_1040_3;
  wire __tmp_1040_4;
  wire __tmp_1040_5;
  wire __tmp_1042_1;
  wire __tmp_1042_2;
  wire __tmp_1042_3;
  wire __tmp_1042_4;
  wire __tmp_1042_5;
  wire __tmp_1042_6;
  wire __tmp_1042_7;
  wire __tmp_1042_8;
  wire __tmp_1042_9;
  wire __tmp_1044_1;
  wire __tmp_1044_2;
  wire __tmp_1044_3;
  wire __tmp_1044_4;
  wire __tmp_1044_5;
  wire __tmp_1044_6;
  wire __tmp_1044_7;
  wire __tmp_1046_1;
  wire __tmp_1046_2;
  wire __tmp_1046_3;
  wire __tmp_1046_4;
  wire __tmp_1046_5;
  wire __tmp_1046_6;
  wire __tmp_1046_7;
  wire __tmp_1048_1;
  wire __tmp_1050_1;
  wire __tmp_1050_2;
  wire __tmp_1050_3;
  wire __tmp_1050_4;
  wire __tmp_1050_5;
  wire __tmp_1052_1;
  wire __tmp_1052_2;
  wire __tmp_1052_3;
  wire __tmp_1052_4;
  wire __tmp_1054_1;
  wire __tmp_1054_2;
  wire __tmp_1054_3;
  wire __tmp_1054_4;
  wire __tmp_1056_1;
  wire __tmp_1056_2;
  wire __tmp_1056_3;
  wire __tmp_1056_4;
  wire __tmp_1056_5;
  wire __tmp_1058_1;
  wire __tmp_1058_2;
  wire __tmp_1058_3;
  wire __tmp_1058_4;
  wire __tmp_1058_5;
  wire __tmp_1060_1;
  wire __tmp_1060_2;
  wire __tmp_1060_3;
  wire __tmp_1060_4;
  wire __tmp_1060_5;
  wire __tmp_1062_1;
  wire __tmp_1062_10;
  wire __tmp_1062_2;
  wire __tmp_1062_3;
  wire __tmp_1062_4;
  wire __tmp_1062_5;
  wire __tmp_1062_6;
  wire __tmp_1062_7;
  wire __tmp_1062_8;
  wire __tmp_1062_9;
  wire __tmp_1064_1;
  wire __tmp_1064_10;
  wire __tmp_1064_2;
  wire __tmp_1064_3;
  wire __tmp_1064_4;
  wire __tmp_1064_5;
  wire __tmp_1064_6;
  wire __tmp_1064_7;
  wire __tmp_1064_8;
  wire __tmp_1064_9;
  wire __tmp_1066_1;
  wire __tmp_1066_10;
  wire __tmp_1066_2;
  wire __tmp_1066_3;
  wire __tmp_1066_4;
  wire __tmp_1066_5;
  wire __tmp_1066_6;
  wire __tmp_1066_7;
  wire __tmp_1066_8;
  wire __tmp_1066_9;
  wire __tmp_1068_1;
  wire __tmp_1068_10;
  wire __tmp_1068_2;
  wire __tmp_1068_3;
  wire __tmp_1068_4;
  wire __tmp_1068_5;
  wire __tmp_1068_6;
  wire __tmp_1068_7;
  wire __tmp_1068_8;
  wire __tmp_1068_9;
  wire __tmp_1070_1;
  wire __tmp_1070_2;
  wire __tmp_1070_3;
  wire __tmp_1070_4;
  wire __tmp_1070_5;
  wire __tmp_1070_6;
  wire __tmp_1077_1;
  wire [7:0] __tmp_1078_1;
  wire __tmp_1089_1;
  wire [7:0] __tmp_1090_1;
  wire __tmp_1101_1;
  wire [7:0] __tmp_1102_1;
  wire __tmp_1113_1;
  wire [7:0] __tmp_1114_1;
  wire [1:0] __tmp_1170_1;
  wire [1:0] __tmp_1170_2;
  wire __tmp_1178_1;
  wire [1:0] __tmp_1181_1;
  wire [1:0] __tmp_1181_2;
  wire __tmp_1189_1;
  wire [1:0] __tmp_1201_1;
  wire [1:0] __tmp_1201_2;
  wire __tmp_1209_1;
  wire [2:0] __tmp_1211_1;
  wire [2:0] __tmp_1211_2;
  wire __tmp_1223_1;
  wire __tmp_1227_1;
  wire __tmp_1227_2;
  wire __tmp_1227_3;
  wire __tmp_1227_4;
  wire __tmp_1227_5;
  wire __tmp_1229_1;
  wire __tmp_1229_2;
  wire __tmp_1229_3;
  wire __tmp_1229_4;
  wire __tmp_1229_5;
  wire __tmp_1229_6;
  wire __tmp_1229_7;
  wire __tmp_1229_8;
  wire __tmp_1231_1;
  wire __tmp_1231_2;
  wire __tmp_1231_3;
  wire __tmp_1231_4;
  wire __tmp_1231_5;
  wire __tmp_1231_6;
  wire __tmp_1231_7;
  wire __tmp_1231_8;
  wire __tmp_1233_1;
  wire __tmp_1233_2;
  wire __tmp_1233_3;
  wire __tmp_1233_4;
  wire __tmp_1233_5;
  wire __tmp_1233_6;
  wire __tmp_1233_7;
  wire __tmp_1233_8;
  wire __tmp_1235_1;
  wire __tmp_1235_10;
  wire __tmp_1235_11;
  wire __tmp_1235_12;
  wire __tmp_1235_13;
  wire __tmp_1235_14;
  wire __tmp_1235_15;
  wire __tmp_1235_16;
  wire __tmp_1235_17;
  wire __tmp_1235_18;
  wire __tmp_1235_2;
  wire __tmp_1235_3;
  wire __tmp_1235_4;
  wire __tmp_1235_5;
  wire __tmp_1235_6;
  wire __tmp_1235_7;
  wire __tmp_1235_8;
  wire __tmp_1235_9;
  wire __tmp_1237_1;
  wire __tmp_1237_10;
  wire __tmp_1237_11;
  wire __tmp_1237_12;
  wire __tmp_1237_13;
  wire __tmp_1237_14;
  wire __tmp_1237_15;
  wire __tmp_1237_16;
  wire __tmp_1237_17;
  wire __tmp_1237_18;
  wire __tmp_1237_19;
  wire __tmp_1237_2;
  wire __tmp_1237_20;
  wire __tmp_1237_21;
  wire __tmp_1237_22;
  wire __tmp_1237_3;
  wire __tmp_1237_4;
  wire __tmp_1237_5;
  wire __tmp_1237_6;
  wire __tmp_1237_7;
  wire __tmp_1237_8;
  wire __tmp_1237_9;
  wire __tmp_1239_1;
  wire __tmp_1239_10;
  wire __tmp_1239_11;
  wire __tmp_1239_12;
  wire __tmp_1239_13;
  wire __tmp_1239_14;
  wire __tmp_1239_15;
  wire __tmp_1239_16;
  wire __tmp_1239_17;
  wire __tmp_1239_18;
  wire __tmp_1239_19;
  wire __tmp_1239_2;
  wire __tmp_1239_20;
  wire __tmp_1239_3;
  wire __tmp_1239_4;
  wire __tmp_1239_5;
  wire __tmp_1239_6;
  wire __tmp_1239_7;
  wire __tmp_1239_8;
  wire __tmp_1239_9;
  wire __tmp_1241_1;
  wire __tmp_1241_10;
  wire __tmp_1241_11;
  wire __tmp_1241_12;
  wire __tmp_1241_13;
  wire __tmp_1241_14;
  wire __tmp_1241_15;
  wire __tmp_1241_16;
  wire __tmp_1241_17;
  wire __tmp_1241_18;
  wire __tmp_1241_19;
  wire __tmp_1241_2;
  wire __tmp_1241_20;
  wire __tmp_1241_3;
  wire __tmp_1241_4;
  wire __tmp_1241_5;
  wire __tmp_1241_6;
  wire __tmp_1241_7;
  wire __tmp_1241_8;
  wire __tmp_1241_9;
  wire __tmp_1243_1;
  wire __tmp_1243_10;
  wire __tmp_1243_11;
  wire __tmp_1243_12;
  wire __tmp_1243_13;
  wire __tmp_1243_14;
  wire __tmp_1243_15;
  wire __tmp_1243_16;
  wire __tmp_1243_17;
  wire __tmp_1243_18;
  wire __tmp_1243_19;
  wire __tmp_1243_2;
  wire __tmp_1243_20;
  wire __tmp_1243_3;
  wire __tmp_1243_4;
  wire __tmp_1243_5;
  wire __tmp_1243_6;
  wire __tmp_1243_7;
  wire __tmp_1243_8;
  wire __tmp_1243_9;
  wire __tmp_1245_1;
  wire __tmp_1245_10;
  wire __tmp_1245_11;
  wire __tmp_1245_12;
  wire __tmp_1245_13;
  wire __tmp_1245_14;
  wire __tmp_1245_15;
  wire __tmp_1245_16;
  wire __tmp_1245_17;
  wire __tmp_1245_18;
  wire __tmp_1245_19;
  wire __tmp_1245_2;
  wire __tmp_1245_20;
  wire __tmp_1245_21;
  wire __tmp_1245_22;
  wire __tmp_1245_23;
  wire __tmp_1245_24;
  wire __tmp_1245_25;
  wire __tmp_1245_26;
  wire __tmp_1245_27;
  wire __tmp_1245_28;
  wire __tmp_1245_3;
  wire __tmp_1245_4;
  wire __tmp_1245_5;
  wire __tmp_1245_6;
  wire __tmp_1245_7;
  wire __tmp_1245_8;
  wire __tmp_1245_9;
  wire __tmp_1247_1;
  wire __tmp_1247_10;
  wire __tmp_1247_11;
  wire __tmp_1247_12;
  wire __tmp_1247_13;
  wire __tmp_1247_14;
  wire __tmp_1247_15;
  wire __tmp_1247_16;
  wire __tmp_1247_17;
  wire __tmp_1247_18;
  wire __tmp_1247_19;
  wire __tmp_1247_2;
  wire __tmp_1247_20;
  wire __tmp_1247_21;
  wire __tmp_1247_22;
  wire __tmp_1247_23;
  wire __tmp_1247_24;
  wire __tmp_1247_25;
  wire __tmp_1247_26;
  wire __tmp_1247_27;
  wire __tmp_1247_28;
  wire __tmp_1247_3;
  wire __tmp_1247_4;
  wire __tmp_1247_5;
  wire __tmp_1247_6;
  wire __tmp_1247_7;
  wire __tmp_1247_8;
  wire __tmp_1247_9;
  wire __tmp_1249_1;
  wire __tmp_1249_10;
  wire __tmp_1249_11;
  wire __tmp_1249_12;
  wire __tmp_1249_13;
  wire __tmp_1249_14;
  wire __tmp_1249_15;
  wire __tmp_1249_16;
  wire __tmp_1249_17;
  wire __tmp_1249_18;
  wire __tmp_1249_19;
  wire __tmp_1249_2;
  wire __tmp_1249_20;
  wire __tmp_1249_21;
  wire __tmp_1249_22;
  wire __tmp_1249_23;
  wire __tmp_1249_24;
  wire __tmp_1249_25;
  wire __tmp_1249_26;
  wire __tmp_1249_27;
  wire __tmp_1249_28;
  wire __tmp_1249_3;
  wire __tmp_1249_4;
  wire __tmp_1249_5;
  wire __tmp_1249_6;
  wire __tmp_1249_7;
  wire __tmp_1249_8;
  wire __tmp_1249_9;
  wire __tmp_1251_1;
  wire __tmp_1253_1;
  wire __tmp_1253_2;
  wire __tmp_1253_3;
  wire __tmp_1253_4;
  wire __tmp_1253_5;
  wire __tmp_1255_1;
  wire __tmp_1255_2;
  wire __tmp_1255_3;
  wire __tmp_1255_4;
  wire __tmp_1255_5;
  wire __tmp_1257_1;
  wire __tmp_1257_2;
  wire __tmp_1257_3;
  wire __tmp_1257_4;
  wire __tmp_1257_5;
  wire __tmp_1259_1;
  wire __tmp_1259_10;
  wire __tmp_1259_11;
  wire __tmp_1259_12;
  wire __tmp_1259_2;
  wire __tmp_1259_3;
  wire __tmp_1259_4;
  wire __tmp_1259_5;
  wire __tmp_1259_6;
  wire __tmp_1259_7;
  wire __tmp_1259_8;
  wire __tmp_1259_9;
  wire __tmp_1261_1;
  wire __tmp_1261_10;
  wire __tmp_1261_11;
  wire __tmp_1261_12;
  wire __tmp_1261_2;
  wire __tmp_1261_3;
  wire __tmp_1261_4;
  wire __tmp_1261_5;
  wire __tmp_1261_6;
  wire __tmp_1261_7;
  wire __tmp_1261_8;
  wire __tmp_1261_9;
  wire __tmp_1263_1;
  wire __tmp_1263_10;
  wire __tmp_1263_11;
  wire __tmp_1263_12;
  wire __tmp_1263_2;
  wire __tmp_1263_3;
  wire __tmp_1263_4;
  wire __tmp_1263_5;
  wire __tmp_1263_6;
  wire __tmp_1263_7;
  wire __tmp_1263_8;
  wire __tmp_1263_9;
  wire __tmp_1265_1;
  wire __tmp_1265_10;
  wire __tmp_1265_11;
  wire __tmp_1265_12;
  wire __tmp_1265_13;
  wire __tmp_1265_14;
  wire __tmp_1265_15;
  wire __tmp_1265_2;
  wire __tmp_1265_3;
  wire __tmp_1265_4;
  wire __tmp_1265_5;
  wire __tmp_1265_6;
  wire __tmp_1265_7;
  wire __tmp_1265_8;
  wire __tmp_1265_9;
  wire __tmp_1267_1;
  wire __tmp_1267_2;
  wire __tmp_1267_3;
  wire __tmp_1267_4;
  wire __tmp_1269_1;
  wire __tmp_1269_2;
  wire __tmp_1269_3;
  wire __tmp_1269_4;
  wire __tmp_1271_1;
  wire __tmp_1271_2;
  wire __tmp_1271_3;
  wire __tmp_1271_4;
  wire __tmp_1273_1;
  wire __tmp_1273_10;
  wire __tmp_1273_11;
  wire __tmp_1273_12;
  wire __tmp_1273_13;
  wire __tmp_1273_14;
  wire __tmp_1273_15;
  wire __tmp_1273_16;
  wire __tmp_1273_17;
  wire __tmp_1273_18;
  wire __tmp_1273_2;
  wire __tmp_1273_3;
  wire __tmp_1273_4;
  wire __tmp_1273_5;
  wire __tmp_1273_6;
  wire __tmp_1273_7;
  wire __tmp_1273_8;
  wire __tmp_1273_9;
  wire __tmp_1275_1;
  wire __tmp_1275_10;
  wire __tmp_1275_11;
  wire __tmp_1275_12;
  wire __tmp_1275_13;
  wire __tmp_1275_14;
  wire __tmp_1275_15;
  wire __tmp_1275_16;
  wire __tmp_1275_17;
  wire __tmp_1275_2;
  wire __tmp_1275_3;
  wire __tmp_1275_4;
  wire __tmp_1275_5;
  wire __tmp_1275_6;
  wire __tmp_1275_7;
  wire __tmp_1275_8;
  wire __tmp_1275_9;
  wire __tmp_1277_1;
  wire __tmp_1277_10;
  wire __tmp_1277_11;
  wire __tmp_1277_12;
  wire __tmp_1277_13;
  wire __tmp_1277_14;
  wire __tmp_1277_15;
  wire __tmp_1277_16;
  wire __tmp_1277_17;
  wire __tmp_1277_2;
  wire __tmp_1277_3;
  wire __tmp_1277_4;
  wire __tmp_1277_5;
  wire __tmp_1277_6;
  wire __tmp_1277_7;
  wire __tmp_1277_8;
  wire __tmp_1277_9;
  wire __tmp_1279_1;
  wire __tmp_1279_10;
  wire __tmp_1279_11;
  wire __tmp_1279_12;
  wire __tmp_1279_13;
  wire __tmp_1279_14;
  wire __tmp_1279_15;
  wire __tmp_1279_16;
  wire __tmp_1279_17;
  wire __tmp_1279_2;
  wire __tmp_1279_3;
  wire __tmp_1279_4;
  wire __tmp_1279_5;
  wire __tmp_1279_6;
  wire __tmp_1279_7;
  wire __tmp_1279_8;
  wire __tmp_1279_9;
  wire __tmp_1281_1;
  wire __tmp_1281_2;
  wire __tmp_1281_3;
  wire __tmp_1281_4;
  wire __tmp_1281_5;
  wire __tmp_1281_6;
  wire __tmp_1281_7;
  wire __tmp_1281_8;
  wire __tmp_1281_9;
  wire __tmp_1283_1;
  wire __tmp_1283_2;
  wire __tmp_1283_3;
  wire __tmp_1283_4;
  wire __tmp_1283_5;
  wire __tmp_1283_6;
  wire __tmp_1283_7;
  wire __tmp_1283_8;
  wire __tmp_1283_9;
  wire __tmp_1285_1;
  wire __tmp_1285_2;
  wire __tmp_1285_3;
  wire __tmp_1285_4;
  wire __tmp_1285_5;
  wire __tmp_1285_6;
  wire __tmp_1285_7;
  wire __tmp_1285_8;
  wire __tmp_1285_9;
  wire __tmp_1287_1;
  wire __tmp_1287_10;
  wire __tmp_1287_11;
  wire __tmp_1287_12;
  wire __tmp_1287_13;
  wire __tmp_1287_14;
  wire __tmp_1287_15;
  wire __tmp_1287_16;
  wire __tmp_1287_17;
  wire __tmp_1287_18;
  wire __tmp_1287_19;
  wire __tmp_1287_2;
  wire __tmp_1287_20;
  wire __tmp_1287_21;
  wire __tmp_1287_22;
  wire __tmp_1287_23;
  wire __tmp_1287_24;
  wire __tmp_1287_25;
  wire __tmp_1287_3;
  wire __tmp_1287_4;
  wire __tmp_1287_5;
  wire __tmp_1287_6;
  wire __tmp_1287_7;
  wire __tmp_1287_8;
  wire __tmp_1287_9;
  wire __tmp_1289_1;
  wire __tmp_1289_10;
  wire __tmp_1289_11;
  wire __tmp_1289_12;
  wire __tmp_1289_13;
  wire __tmp_1289_14;
  wire __tmp_1289_15;
  wire __tmp_1289_16;
  wire __tmp_1289_17;
  wire __tmp_1289_18;
  wire __tmp_1289_19;
  wire __tmp_1289_2;
  wire __tmp_1289_20;
  wire __tmp_1289_21;
  wire __tmp_1289_22;
  wire __tmp_1289_23;
  wire __tmp_1289_24;
  wire __tmp_1289_25;
  wire __tmp_1289_3;
  wire __tmp_1289_4;
  wire __tmp_1289_5;
  wire __tmp_1289_6;
  wire __tmp_1289_7;
  wire __tmp_1289_8;
  wire __tmp_1289_9;
  wire __tmp_1291_1;
  wire __tmp_1291_10;
  wire __tmp_1291_11;
  wire __tmp_1291_12;
  wire __tmp_1291_13;
  wire __tmp_1291_14;
  wire __tmp_1291_15;
  wire __tmp_1291_16;
  wire __tmp_1291_17;
  wire __tmp_1291_18;
  wire __tmp_1291_19;
  wire __tmp_1291_2;
  wire __tmp_1291_20;
  wire __tmp_1291_21;
  wire __tmp_1291_22;
  wire __tmp_1291_23;
  wire __tmp_1291_24;
  wire __tmp_1291_25;
  wire __tmp_1291_3;
  wire __tmp_1291_4;
  wire __tmp_1291_5;
  wire __tmp_1291_6;
  wire __tmp_1291_7;
  wire __tmp_1291_8;
  wire __tmp_1291_9;
  wire __tmp_1293_1;
  wire __tmp_1293_10;
  wire __tmp_1293_11;
  wire __tmp_1293_12;
  wire __tmp_1293_2;
  wire __tmp_1293_3;
  wire __tmp_1293_4;
  wire __tmp_1293_5;
  wire __tmp_1293_6;
  wire __tmp_1293_7;
  wire __tmp_1293_8;
  wire __tmp_1293_9;
  wire __tmp_1295_1;
  wire __tmp_1295_10;
  wire __tmp_1295_11;
  wire __tmp_1295_12;
  wire __tmp_1295_2;
  wire __tmp_1295_3;
  wire __tmp_1295_4;
  wire __tmp_1295_5;
  wire __tmp_1295_6;
  wire __tmp_1295_7;
  wire __tmp_1295_8;
  wire __tmp_1295_9;
  wire __tmp_1297_1;
  wire __tmp_1297_10;
  wire __tmp_1297_11;
  wire __tmp_1297_12;
  wire __tmp_1297_2;
  wire __tmp_1297_3;
  wire __tmp_1297_4;
  wire __tmp_1297_5;
  wire __tmp_1297_6;
  wire __tmp_1297_7;
  wire __tmp_1297_8;
  wire __tmp_1297_9;
  wire __tmp_1299_1;
  wire __tmp_1299_10;
  wire __tmp_1299_11;
  wire __tmp_1299_12;
  wire __tmp_1299_13;
  wire __tmp_1299_14;
  wire __tmp_1299_15;
  wire __tmp_1299_16;
  wire __tmp_1299_17;
  wire __tmp_1299_18;
  wire __tmp_1299_19;
  wire __tmp_1299_2;
  wire __tmp_1299_20;
  wire __tmp_1299_21;
  wire __tmp_1299_22;
  wire __tmp_1299_23;
  wire __tmp_1299_24;
  wire __tmp_1299_25;
  wire __tmp_1299_26;
  wire __tmp_1299_27;
  wire __tmp_1299_28;
  wire __tmp_1299_29;
  wire __tmp_1299_3;
  wire __tmp_1299_30;
  wire __tmp_1299_31;
  wire __tmp_1299_32;
  wire __tmp_1299_33;
  wire __tmp_1299_34;
  wire __tmp_1299_35;
  wire __tmp_1299_36;
  wire __tmp_1299_37;
  wire __tmp_1299_38;
  wire __tmp_1299_39;
  wire __tmp_1299_4;
  wire __tmp_1299_40;
  wire __tmp_1299_41;
  wire __tmp_1299_42;
  wire __tmp_1299_5;
  wire __tmp_1299_6;
  wire __tmp_1299_7;
  wire __tmp_1299_8;
  wire __tmp_1299_9;
  wire __tmp_1301_1;
  wire __tmp_1301_10;
  wire __tmp_1301_11;
  wire __tmp_1301_12;
  wire __tmp_1301_13;
  wire __tmp_1301_14;
  wire __tmp_1301_15;
  wire __tmp_1301_16;
  wire __tmp_1301_17;
  wire __tmp_1301_18;
  wire __tmp_1301_19;
  wire __tmp_1301_2;
  wire __tmp_1301_20;
  wire __tmp_1301_21;
  wire __tmp_1301_22;
  wire __tmp_1301_23;
  wire __tmp_1301_24;
  wire __tmp_1301_25;
  wire __tmp_1301_26;
  wire __tmp_1301_27;
  wire __tmp_1301_28;
  wire __tmp_1301_29;
  wire __tmp_1301_3;
  wire __tmp_1301_30;
  wire __tmp_1301_31;
  wire __tmp_1301_32;
  wire __tmp_1301_33;
  wire __tmp_1301_34;
  wire __tmp_1301_35;
  wire __tmp_1301_36;
  wire __tmp_1301_37;
  wire __tmp_1301_38;
  wire __tmp_1301_39;
  wire __tmp_1301_4;
  wire __tmp_1301_40;
  wire __tmp_1301_41;
  wire __tmp_1301_42;
  wire __tmp_1301_5;
  wire __tmp_1301_6;
  wire __tmp_1301_7;
  wire __tmp_1301_8;
  wire __tmp_1301_9;
  wire __tmp_1303_1;
  wire __tmp_1303_10;
  wire __tmp_1303_11;
  wire __tmp_1303_12;
  wire __tmp_1303_13;
  wire __tmp_1303_14;
  wire __tmp_1303_15;
  wire __tmp_1303_16;
  wire __tmp_1303_17;
  wire __tmp_1303_18;
  wire __tmp_1303_19;
  wire __tmp_1303_2;
  wire __tmp_1303_20;
  wire __tmp_1303_21;
  wire __tmp_1303_22;
  wire __tmp_1303_23;
  wire __tmp_1303_24;
  wire __tmp_1303_25;
  wire __tmp_1303_26;
  wire __tmp_1303_27;
  wire __tmp_1303_28;
  wire __tmp_1303_29;
  wire __tmp_1303_3;
  wire __tmp_1303_30;
  wire __tmp_1303_31;
  wire __tmp_1303_32;
  wire __tmp_1303_33;
  wire __tmp_1303_34;
  wire __tmp_1303_35;
  wire __tmp_1303_36;
  wire __tmp_1303_37;
  wire __tmp_1303_38;
  wire __tmp_1303_39;
  wire __tmp_1303_4;
  wire __tmp_1303_40;
  wire __tmp_1303_41;
  wire __tmp_1303_42;
  wire __tmp_1303_5;
  wire __tmp_1303_6;
  wire __tmp_1303_7;
  wire __tmp_1303_8;
  wire __tmp_1303_9;
  wire __tmp_1305_1;
  wire __tmp_1305_10;
  wire __tmp_1305_11;
  wire __tmp_1305_12;
  wire __tmp_1305_13;
  wire __tmp_1305_14;
  wire __tmp_1305_15;
  wire __tmp_1305_16;
  wire __tmp_1305_17;
  wire __tmp_1305_18;
  wire __tmp_1305_19;
  wire __tmp_1305_2;
  wire __tmp_1305_20;
  wire __tmp_1305_21;
  wire __tmp_1305_22;
  wire __tmp_1305_23;
  wire __tmp_1305_24;
  wire __tmp_1305_25;
  wire __tmp_1305_26;
  wire __tmp_1305_27;
  wire __tmp_1305_28;
  wire __tmp_1305_29;
  wire __tmp_1305_3;
  wire __tmp_1305_30;
  wire __tmp_1305_31;
  wire __tmp_1305_32;
  wire __tmp_1305_33;
  wire __tmp_1305_34;
  wire __tmp_1305_35;
  wire __tmp_1305_36;
  wire __tmp_1305_37;
  wire __tmp_1305_38;
  wire __tmp_1305_39;
  wire __tmp_1305_4;
  wire __tmp_1305_40;
  wire __tmp_1305_41;
  wire __tmp_1305_42;
  wire __tmp_1305_5;
  wire __tmp_1305_6;
  wire __tmp_1305_7;
  wire __tmp_1305_8;
  wire __tmp_1305_9;
  wire __tmp_1307_1;
  wire __tmp_1307_10;
  wire __tmp_1307_11;
  wire __tmp_1307_12;
  wire __tmp_1307_13;
  wire __tmp_1307_14;
  wire __tmp_1307_15;
  wire __tmp_1307_16;
  wire __tmp_1307_17;
  wire __tmp_1307_18;
  wire __tmp_1307_19;
  wire __tmp_1307_2;
  wire __tmp_1307_20;
  wire __tmp_1307_21;
  wire __tmp_1307_22;
  wire __tmp_1307_23;
  wire __tmp_1307_24;
  wire __tmp_1307_25;
  wire __tmp_1307_26;
  wire __tmp_1307_27;
  wire __tmp_1307_28;
  wire __tmp_1307_29;
  wire __tmp_1307_3;
  wire __tmp_1307_30;
  wire __tmp_1307_31;
  wire __tmp_1307_32;
  wire __tmp_1307_33;
  wire __tmp_1307_34;
  wire __tmp_1307_35;
  wire __tmp_1307_36;
  wire __tmp_1307_37;
  wire __tmp_1307_38;
  wire __tmp_1307_4;
  wire __tmp_1307_5;
  wire __tmp_1307_6;
  wire __tmp_1307_7;
  wire __tmp_1307_8;
  wire __tmp_1307_9;
  wire __tmp_1314_1;
  wire [7:0] __tmp_1315_1;
  wire __tmp_1326_1;
  wire [7:0] __tmp_1327_1;
  wire __tmp_1338_1;
  wire [7:0] __tmp_1339_1;
  wire __tmp_1350_1;
  wire [7:0] __tmp_1351_1;
  wire [1:0] __tmp_464_1;
  wire [1:0] __tmp_464_2;
  wire __tmp_472_1;
  wire [1:0] __tmp_475_1;
  wire [1:0] __tmp_475_2;
  wire __tmp_483_1;
  wire [1:0] __tmp_495_1;
  wire [1:0] __tmp_495_2;
  wire __tmp_503_1;
  wire [1:0] __tmp_505_1;
  wire [1:0] __tmp_505_2;
  wire __tmp_513_1;
  wire [1:0] __tmp_515_1;
  wire [1:0] __tmp_515_2;
  wire __tmp_523_1;
  wire [1:0] __tmp_525_1;
  wire [1:0] __tmp_525_2;
  wire __tmp_533_1;
  wire [1:0] __tmp_535_1;
  wire [1:0] __tmp_535_2;
  wire __tmp_543_1;
  wire [1:0] __tmp_545_1;
  wire [1:0] __tmp_545_2;
  wire __tmp_553_1;
  wire [1:0] __tmp_555_1;
  wire [1:0] __tmp_555_2;
  wire __tmp_563_1;
  wire [1:0] __tmp_565_1;
  wire [1:0] __tmp_565_2;
  wire __tmp_573_1;
  wire [1:0] __tmp_575_1;
  wire [1:0] __tmp_575_2;
  wire __tmp_583_1;
  wire [2:0] __tmp_585_1;
  wire [2:0] __tmp_585_2;
  wire __tmp_597_1;
  wire [2:0] __tmp_599_1;
  wire [2:0] __tmp_599_2;
  wire __tmp_611_1;
  wire [2:0] __tmp_613_1;
  wire [2:0] __tmp_613_2;
  wire __tmp_625_1;
  wire [2:0] __tmp_627_1;
  wire [2:0] __tmp_627_2;
  wire __tmp_639_1;
  wire [2:0] __tmp_641_1;
  wire [2:0] __tmp_641_2;
  wire __tmp_653_1;
  wire [2:0] __tmp_655_1;
  wire [2:0] __tmp_655_2;
  wire __tmp_667_1;
  wire [2:0] __tmp_669_1;
  wire [2:0] __tmp_669_2;
  wire __tmp_681_1;
  wire [2:0] __tmp_683_1;
  wire [2:0] __tmp_683_2;
  wire __tmp_695_1;
  wire [2:0] __tmp_697_1;
  wire [2:0] __tmp_697_2;
  wire __tmp_709_1;
  wire __tmp_713_1;
  wire __tmp_713_2;
  wire __tmp_713_3;
  wire __tmp_713_4;
  wire __tmp_713_5;
  wire __tmp_715_1;
  wire __tmp_715_10;
  wire __tmp_715_11;
  wire __tmp_715_12;
  wire __tmp_715_2;
  wire __tmp_715_3;
  wire __tmp_715_4;
  wire __tmp_715_5;
  wire __tmp_715_6;
  wire __tmp_715_7;
  wire __tmp_715_8;
  wire __tmp_715_9;
  wire __tmp_717_1;
  wire __tmp_717_10;
  wire __tmp_717_11;
  wire __tmp_717_12;
  wire __tmp_717_2;
  wire __tmp_717_3;
  wire __tmp_717_4;
  wire __tmp_717_5;
  wire __tmp_717_6;
  wire __tmp_717_7;
  wire __tmp_717_8;
  wire __tmp_717_9;
  wire __tmp_719_1;
  wire __tmp_719_10;
  wire __tmp_719_11;
  wire __tmp_719_12;
  wire __tmp_719_2;
  wire __tmp_719_3;
  wire __tmp_719_4;
  wire __tmp_719_5;
  wire __tmp_719_6;
  wire __tmp_719_7;
  wire __tmp_719_8;
  wire __tmp_719_9;
  wire __tmp_721_1;
  wire __tmp_721_10;
  wire __tmp_721_11;
  wire __tmp_721_12;
  wire __tmp_721_2;
  wire __tmp_721_3;
  wire __tmp_721_4;
  wire __tmp_721_5;
  wire __tmp_721_6;
  wire __tmp_721_7;
  wire __tmp_721_8;
  wire __tmp_721_9;
  wire __tmp_723_1;
  wire __tmp_723_10;
  wire __tmp_723_11;
  wire __tmp_723_12;
  wire __tmp_723_2;
  wire __tmp_723_3;
  wire __tmp_723_4;
  wire __tmp_723_5;
  wire __tmp_723_6;
  wire __tmp_723_7;
  wire __tmp_723_8;
  wire __tmp_723_9;
  wire __tmp_725_1;
  wire __tmp_725_10;
  wire __tmp_725_11;
  wire __tmp_725_12;
  wire __tmp_725_2;
  wire __tmp_725_3;
  wire __tmp_725_4;
  wire __tmp_725_5;
  wire __tmp_725_6;
  wire __tmp_725_7;
  wire __tmp_725_8;
  wire __tmp_725_9;
  wire __tmp_727_1;
  wire __tmp_727_10;
  wire __tmp_727_11;
  wire __tmp_727_12;
  wire __tmp_727_2;
  wire __tmp_727_3;
  wire __tmp_727_4;
  wire __tmp_727_5;
  wire __tmp_727_6;
  wire __tmp_727_7;
  wire __tmp_727_8;
  wire __tmp_727_9;
  wire __tmp_729_1;
  wire __tmp_729_10;
  wire __tmp_729_11;
  wire __tmp_729_12;
  wire __tmp_729_2;
  wire __tmp_729_3;
  wire __tmp_729_4;
  wire __tmp_729_5;
  wire __tmp_729_6;
  wire __tmp_729_7;
  wire __tmp_729_8;
  wire __tmp_729_9;
  wire __tmp_731_1;
  wire __tmp_731_10;
  wire __tmp_731_11;
  wire __tmp_731_12;
  wire __tmp_731_2;
  wire __tmp_731_3;
  wire __tmp_731_4;
  wire __tmp_731_5;
  wire __tmp_731_6;
  wire __tmp_731_7;
  wire __tmp_731_8;
  wire __tmp_731_9;
  wire __tmp_733_1;
  wire __tmp_733_10;
  wire __tmp_733_11;
  wire __tmp_733_12;
  wire __tmp_733_2;
  wire __tmp_733_3;
  wire __tmp_733_4;
  wire __tmp_733_5;
  wire __tmp_733_6;
  wire __tmp_733_7;
  wire __tmp_733_8;
  wire __tmp_733_9;
  wire __tmp_735_1;
  wire __tmp_735_10;
  wire __tmp_735_11;
  wire __tmp_735_12;
  wire __tmp_735_2;
  wire __tmp_735_3;
  wire __tmp_735_4;
  wire __tmp_735_5;
  wire __tmp_735_6;
  wire __tmp_735_7;
  wire __tmp_735_8;
  wire __tmp_735_9;
  wire __tmp_737_1;
  wire __tmp_737_10;
  wire __tmp_737_11;
  wire __tmp_737_12;
  wire __tmp_737_2;
  wire __tmp_737_3;
  wire __tmp_737_4;
  wire __tmp_737_5;
  wire __tmp_737_6;
  wire __tmp_737_7;
  wire __tmp_737_8;
  wire __tmp_737_9;
  wire __tmp_739_1;
  wire __tmp_739_10;
  wire __tmp_739_11;
  wire __tmp_739_12;
  wire __tmp_739_2;
  wire __tmp_739_3;
  wire __tmp_739_4;
  wire __tmp_739_5;
  wire __tmp_739_6;
  wire __tmp_739_7;
  wire __tmp_739_8;
  wire __tmp_739_9;
  wire __tmp_741_1;
  wire __tmp_741_10;
  wire __tmp_741_11;
  wire __tmp_741_12;
  wire __tmp_741_2;
  wire __tmp_741_3;
  wire __tmp_741_4;
  wire __tmp_741_5;
  wire __tmp_741_6;
  wire __tmp_741_7;
  wire __tmp_741_8;
  wire __tmp_741_9;
  wire __tmp_743_1;
  wire __tmp_743_10;
  wire __tmp_743_11;
  wire __tmp_743_12;
  wire __tmp_743_2;
  wire __tmp_743_3;
  wire __tmp_743_4;
  wire __tmp_743_5;
  wire __tmp_743_6;
  wire __tmp_743_7;
  wire __tmp_743_8;
  wire __tmp_743_9;
  wire __tmp_745_1;
  wire __tmp_745_10;
  wire __tmp_745_11;
  wire __tmp_745_12;
  wire __tmp_745_2;
  wire __tmp_745_3;
  wire __tmp_745_4;
  wire __tmp_745_5;
  wire __tmp_745_6;
  wire __tmp_745_7;
  wire __tmp_745_8;
  wire __tmp_745_9;
  wire __tmp_747_1;
  wire __tmp_747_10;
  wire __tmp_747_11;
  wire __tmp_747_12;
  wire __tmp_747_2;
  wire __tmp_747_3;
  wire __tmp_747_4;
  wire __tmp_747_5;
  wire __tmp_747_6;
  wire __tmp_747_7;
  wire __tmp_747_8;
  wire __tmp_747_9;
  wire __tmp_749_1;
  wire __tmp_749_10;
  wire __tmp_749_11;
  wire __tmp_749_12;
  wire __tmp_749_2;
  wire __tmp_749_3;
  wire __tmp_749_4;
  wire __tmp_749_5;
  wire __tmp_749_6;
  wire __tmp_749_7;
  wire __tmp_749_8;
  wire __tmp_749_9;
  wire __tmp_751_1;
  wire __tmp_751_10;
  wire __tmp_751_11;
  wire __tmp_751_12;
  wire __tmp_751_2;
  wire __tmp_751_3;
  wire __tmp_751_4;
  wire __tmp_751_5;
  wire __tmp_751_6;
  wire __tmp_751_7;
  wire __tmp_751_8;
  wire __tmp_751_9;
  wire __tmp_753_1;
  wire __tmp_753_10;
  wire __tmp_753_11;
  wire __tmp_753_12;
  wire __tmp_753_2;
  wire __tmp_753_3;
  wire __tmp_753_4;
  wire __tmp_753_5;
  wire __tmp_753_6;
  wire __tmp_753_7;
  wire __tmp_753_8;
  wire __tmp_753_9;
  wire __tmp_755_1;
  wire __tmp_755_10;
  wire __tmp_755_11;
  wire __tmp_755_12;
  wire __tmp_755_2;
  wire __tmp_755_3;
  wire __tmp_755_4;
  wire __tmp_755_5;
  wire __tmp_755_6;
  wire __tmp_755_7;
  wire __tmp_755_8;
  wire __tmp_755_9;
  wire __tmp_757_1;
  wire __tmp_757_10;
  wire __tmp_757_11;
  wire __tmp_757_12;
  wire __tmp_757_2;
  wire __tmp_757_3;
  wire __tmp_757_4;
  wire __tmp_757_5;
  wire __tmp_757_6;
  wire __tmp_757_7;
  wire __tmp_757_8;
  wire __tmp_757_9;
  wire __tmp_759_1;
  wire __tmp_759_10;
  wire __tmp_759_11;
  wire __tmp_759_12;
  wire __tmp_759_2;
  wire __tmp_759_3;
  wire __tmp_759_4;
  wire __tmp_759_5;
  wire __tmp_759_6;
  wire __tmp_759_7;
  wire __tmp_759_8;
  wire __tmp_759_9;
  wire __tmp_761_1;
  wire __tmp_761_10;
  wire __tmp_761_11;
  wire __tmp_761_12;
  wire __tmp_761_2;
  wire __tmp_761_3;
  wire __tmp_761_4;
  wire __tmp_761_5;
  wire __tmp_761_6;
  wire __tmp_761_7;
  wire __tmp_761_8;
  wire __tmp_761_9;
  wire __tmp_763_1;
  wire __tmp_763_10;
  wire __tmp_763_11;
  wire __tmp_763_12;
  wire __tmp_763_2;
  wire __tmp_763_3;
  wire __tmp_763_4;
  wire __tmp_763_5;
  wire __tmp_763_6;
  wire __tmp_763_7;
  wire __tmp_763_8;
  wire __tmp_763_9;
  wire __tmp_765_1;
  wire __tmp_765_10;
  wire __tmp_765_11;
  wire __tmp_765_12;
  wire __tmp_765_2;
  wire __tmp_765_3;
  wire __tmp_765_4;
  wire __tmp_765_5;
  wire __tmp_765_6;
  wire __tmp_765_7;
  wire __tmp_765_8;
  wire __tmp_765_9;
  wire __tmp_767_1;
  wire __tmp_767_10;
  wire __tmp_767_11;
  wire __tmp_767_12;
  wire __tmp_767_2;
  wire __tmp_767_3;
  wire __tmp_767_4;
  wire __tmp_767_5;
  wire __tmp_767_6;
  wire __tmp_767_7;
  wire __tmp_767_8;
  wire __tmp_767_9;
  wire __tmp_769_1;
  wire __tmp_769_10;
  wire __tmp_769_11;
  wire __tmp_769_12;
  wire __tmp_769_13;
  wire __tmp_769_14;
  wire __tmp_769_15;
  wire __tmp_769_16;
  wire __tmp_769_17;
  wire __tmp_769_18;
  wire __tmp_769_19;
  wire __tmp_769_2;
  wire __tmp_769_20;
  wire __tmp_769_21;
  wire __tmp_769_22;
  wire __tmp_769_3;
  wire __tmp_769_4;
  wire __tmp_769_5;
  wire __tmp_769_6;
  wire __tmp_769_7;
  wire __tmp_769_8;
  wire __tmp_769_9;
  wire __tmp_771_1;
  wire __tmp_771_10;
  wire __tmp_771_11;
  wire __tmp_771_12;
  wire __tmp_771_13;
  wire __tmp_771_14;
  wire __tmp_771_15;
  wire __tmp_771_16;
  wire __tmp_771_17;
  wire __tmp_771_18;
  wire __tmp_771_19;
  wire __tmp_771_2;
  wire __tmp_771_20;
  wire __tmp_771_21;
  wire __tmp_771_22;
  wire __tmp_771_3;
  wire __tmp_771_4;
  wire __tmp_771_5;
  wire __tmp_771_6;
  wire __tmp_771_7;
  wire __tmp_771_8;
  wire __tmp_771_9;
  wire __tmp_773_1;
  wire __tmp_773_10;
  wire __tmp_773_11;
  wire __tmp_773_12;
  wire __tmp_773_13;
  wire __tmp_773_14;
  wire __tmp_773_15;
  wire __tmp_773_16;
  wire __tmp_773_17;
  wire __tmp_773_18;
  wire __tmp_773_19;
  wire __tmp_773_2;
  wire __tmp_773_20;
  wire __tmp_773_21;
  wire __tmp_773_22;
  wire __tmp_773_3;
  wire __tmp_773_4;
  wire __tmp_773_5;
  wire __tmp_773_6;
  wire __tmp_773_7;
  wire __tmp_773_8;
  wire __tmp_773_9;
  wire __tmp_775_1;
  wire __tmp_775_10;
  wire __tmp_775_11;
  wire __tmp_775_12;
  wire __tmp_775_13;
  wire __tmp_775_14;
  wire __tmp_775_15;
  wire __tmp_775_16;
  wire __tmp_775_17;
  wire __tmp_775_18;
  wire __tmp_775_19;
  wire __tmp_775_2;
  wire __tmp_775_20;
  wire __tmp_775_21;
  wire __tmp_775_22;
  wire __tmp_775_3;
  wire __tmp_775_4;
  wire __tmp_775_5;
  wire __tmp_775_6;
  wire __tmp_775_7;
  wire __tmp_775_8;
  wire __tmp_775_9;
  wire __tmp_777_1;
  wire __tmp_777_10;
  wire __tmp_777_11;
  wire __tmp_777_12;
  wire __tmp_777_13;
  wire __tmp_777_14;
  wire __tmp_777_15;
  wire __tmp_777_16;
  wire __tmp_777_17;
  wire __tmp_777_18;
  wire __tmp_777_19;
  wire __tmp_777_2;
  wire __tmp_777_20;
  wire __tmp_777_21;
  wire __tmp_777_22;
  wire __tmp_777_3;
  wire __tmp_777_4;
  wire __tmp_777_5;
  wire __tmp_777_6;
  wire __tmp_777_7;
  wire __tmp_777_8;
  wire __tmp_777_9;
  wire __tmp_779_1;
  wire __tmp_779_10;
  wire __tmp_779_11;
  wire __tmp_779_12;
  wire __tmp_779_13;
  wire __tmp_779_14;
  wire __tmp_779_15;
  wire __tmp_779_16;
  wire __tmp_779_17;
  wire __tmp_779_18;
  wire __tmp_779_19;
  wire __tmp_779_2;
  wire __tmp_779_20;
  wire __tmp_779_21;
  wire __tmp_779_22;
  wire __tmp_779_3;
  wire __tmp_779_4;
  wire __tmp_779_5;
  wire __tmp_779_6;
  wire __tmp_779_7;
  wire __tmp_779_8;
  wire __tmp_779_9;
  wire __tmp_781_1;
  wire __tmp_781_10;
  wire __tmp_781_11;
  wire __tmp_781_12;
  wire __tmp_781_13;
  wire __tmp_781_14;
  wire __tmp_781_15;
  wire __tmp_781_16;
  wire __tmp_781_17;
  wire __tmp_781_18;
  wire __tmp_781_19;
  wire __tmp_781_2;
  wire __tmp_781_20;
  wire __tmp_781_21;
  wire __tmp_781_22;
  wire __tmp_781_3;
  wire __tmp_781_4;
  wire __tmp_781_5;
  wire __tmp_781_6;
  wire __tmp_781_7;
  wire __tmp_781_8;
  wire __tmp_781_9;
  wire __tmp_783_1;
  wire __tmp_783_10;
  wire __tmp_783_11;
  wire __tmp_783_12;
  wire __tmp_783_13;
  wire __tmp_783_14;
  wire __tmp_783_15;
  wire __tmp_783_16;
  wire __tmp_783_17;
  wire __tmp_783_18;
  wire __tmp_783_19;
  wire __tmp_783_2;
  wire __tmp_783_20;
  wire __tmp_783_21;
  wire __tmp_783_22;
  wire __tmp_783_3;
  wire __tmp_783_4;
  wire __tmp_783_5;
  wire __tmp_783_6;
  wire __tmp_783_7;
  wire __tmp_783_8;
  wire __tmp_783_9;
  wire __tmp_785_1;
  wire __tmp_785_10;
  wire __tmp_785_11;
  wire __tmp_785_12;
  wire __tmp_785_13;
  wire __tmp_785_14;
  wire __tmp_785_15;
  wire __tmp_785_16;
  wire __tmp_785_17;
  wire __tmp_785_18;
  wire __tmp_785_19;
  wire __tmp_785_2;
  wire __tmp_785_20;
  wire __tmp_785_21;
  wire __tmp_785_22;
  wire __tmp_785_3;
  wire __tmp_785_4;
  wire __tmp_785_5;
  wire __tmp_785_6;
  wire __tmp_785_7;
  wire __tmp_785_8;
  wire __tmp_785_9;
  wire __tmp_787_1;
  wire __tmp_787_10;
  wire __tmp_787_11;
  wire __tmp_787_12;
  wire __tmp_787_13;
  wire __tmp_787_14;
  wire __tmp_787_15;
  wire __tmp_787_16;
  wire __tmp_787_17;
  wire __tmp_787_18;
  wire __tmp_787_19;
  wire __tmp_787_2;
  wire __tmp_787_20;
  wire __tmp_787_21;
  wire __tmp_787_22;
  wire __tmp_787_23;
  wire __tmp_787_24;
  wire __tmp_787_25;
  wire __tmp_787_26;
  wire __tmp_787_27;
  wire __tmp_787_28;
  wire __tmp_787_3;
  wire __tmp_787_4;
  wire __tmp_787_5;
  wire __tmp_787_6;
  wire __tmp_787_7;
  wire __tmp_787_8;
  wire __tmp_787_9;
  wire __tmp_789_1;
  wire __tmp_789_10;
  wire __tmp_789_11;
  wire __tmp_789_12;
  wire __tmp_789_13;
  wire __tmp_789_14;
  wire __tmp_789_15;
  wire __tmp_789_16;
  wire __tmp_789_17;
  wire __tmp_789_18;
  wire __tmp_789_19;
  wire __tmp_789_2;
  wire __tmp_789_20;
  wire __tmp_789_21;
  wire __tmp_789_22;
  wire __tmp_789_23;
  wire __tmp_789_24;
  wire __tmp_789_25;
  wire __tmp_789_26;
  wire __tmp_789_3;
  wire __tmp_789_4;
  wire __tmp_789_5;
  wire __tmp_789_6;
  wire __tmp_789_7;
  wire __tmp_789_8;
  wire __tmp_789_9;
  wire __tmp_791_1;
  wire __tmp_791_10;
  wire __tmp_791_11;
  wire __tmp_791_12;
  wire __tmp_791_13;
  wire __tmp_791_14;
  wire __tmp_791_15;
  wire __tmp_791_16;
  wire __tmp_791_17;
  wire __tmp_791_18;
  wire __tmp_791_19;
  wire __tmp_791_2;
  wire __tmp_791_20;
  wire __tmp_791_21;
  wire __tmp_791_22;
  wire __tmp_791_23;
  wire __tmp_791_24;
  wire __tmp_791_25;
  wire __tmp_791_26;
  wire __tmp_791_3;
  wire __tmp_791_4;
  wire __tmp_791_5;
  wire __tmp_791_6;
  wire __tmp_791_7;
  wire __tmp_791_8;
  wire __tmp_791_9;
  wire __tmp_793_1;
  wire __tmp_793_10;
  wire __tmp_793_11;
  wire __tmp_793_12;
  wire __tmp_793_13;
  wire __tmp_793_14;
  wire __tmp_793_15;
  wire __tmp_793_16;
  wire __tmp_793_17;
  wire __tmp_793_18;
  wire __tmp_793_19;
  wire __tmp_793_2;
  wire __tmp_793_20;
  wire __tmp_793_21;
  wire __tmp_793_22;
  wire __tmp_793_23;
  wire __tmp_793_24;
  wire __tmp_793_25;
  wire __tmp_793_26;
  wire __tmp_793_3;
  wire __tmp_793_4;
  wire __tmp_793_5;
  wire __tmp_793_6;
  wire __tmp_793_7;
  wire __tmp_793_8;
  wire __tmp_793_9;
  wire __tmp_795_1;
  wire __tmp_795_10;
  wire __tmp_795_11;
  wire __tmp_795_12;
  wire __tmp_795_13;
  wire __tmp_795_14;
  wire __tmp_795_15;
  wire __tmp_795_16;
  wire __tmp_795_17;
  wire __tmp_795_18;
  wire __tmp_795_19;
  wire __tmp_795_2;
  wire __tmp_795_20;
  wire __tmp_795_21;
  wire __tmp_795_22;
  wire __tmp_795_23;
  wire __tmp_795_24;
  wire __tmp_795_25;
  wire __tmp_795_26;
  wire __tmp_795_27;
  wire __tmp_795_28;
  wire __tmp_795_29;
  wire __tmp_795_3;
  wire __tmp_795_30;
  wire __tmp_795_31;
  wire __tmp_795_32;
  wire __tmp_795_33;
  wire __tmp_795_34;
  wire __tmp_795_4;
  wire __tmp_795_5;
  wire __tmp_795_6;
  wire __tmp_795_7;
  wire __tmp_795_8;
  wire __tmp_795_9;
  wire __tmp_797_1;
  wire __tmp_797_10;
  wire __tmp_797_11;
  wire __tmp_797_12;
  wire __tmp_797_13;
  wire __tmp_797_14;
  wire __tmp_797_15;
  wire __tmp_797_16;
  wire __tmp_797_17;
  wire __tmp_797_18;
  wire __tmp_797_19;
  wire __tmp_797_2;
  wire __tmp_797_20;
  wire __tmp_797_21;
  wire __tmp_797_22;
  wire __tmp_797_23;
  wire __tmp_797_24;
  wire __tmp_797_25;
  wire __tmp_797_26;
  wire __tmp_797_27;
  wire __tmp_797_28;
  wire __tmp_797_29;
  wire __tmp_797_3;
  wire __tmp_797_30;
  wire __tmp_797_31;
  wire __tmp_797_32;
  wire __tmp_797_33;
  wire __tmp_797_34;
  wire __tmp_797_4;
  wire __tmp_797_5;
  wire __tmp_797_6;
  wire __tmp_797_7;
  wire __tmp_797_8;
  wire __tmp_797_9;
  wire __tmp_799_1;
  wire __tmp_799_10;
  wire __tmp_799_11;
  wire __tmp_799_12;
  wire __tmp_799_13;
  wire __tmp_799_14;
  wire __tmp_799_15;
  wire __tmp_799_16;
  wire __tmp_799_17;
  wire __tmp_799_18;
  wire __tmp_799_19;
  wire __tmp_799_2;
  wire __tmp_799_20;
  wire __tmp_799_21;
  wire __tmp_799_22;
  wire __tmp_799_23;
  wire __tmp_799_24;
  wire __tmp_799_25;
  wire __tmp_799_26;
  wire __tmp_799_27;
  wire __tmp_799_28;
  wire __tmp_799_29;
  wire __tmp_799_3;
  wire __tmp_799_30;
  wire __tmp_799_31;
  wire __tmp_799_32;
  wire __tmp_799_33;
  wire __tmp_799_34;
  wire __tmp_799_4;
  wire __tmp_799_5;
  wire __tmp_799_6;
  wire __tmp_799_7;
  wire __tmp_799_8;
  wire __tmp_799_9;
  wire __tmp_801_1;
  wire __tmp_803_1;
  wire __tmp_803_2;
  wire __tmp_803_3;
  wire __tmp_803_4;
  wire __tmp_803_5;
  wire __tmp_803_6;
  wire __tmp_803_7;
  wire __tmp_803_8;
  wire __tmp_803_9;
  wire __tmp_805_1;
  wire __tmp_805_2;
  wire __tmp_805_3;
  wire __tmp_805_4;
  wire __tmp_805_5;
  wire __tmp_805_6;
  wire __tmp_805_7;
  wire __tmp_805_8;
  wire __tmp_805_9;
  wire __tmp_807_1;
  wire __tmp_807_2;
  wire __tmp_807_3;
  wire __tmp_807_4;
  wire __tmp_807_5;
  wire __tmp_807_6;
  wire __tmp_807_7;
  wire __tmp_807_8;
  wire __tmp_807_9;
  wire __tmp_809_1;
  wire __tmp_809_10;
  wire __tmp_809_11;
  wire __tmp_809_12;
  wire __tmp_809_2;
  wire __tmp_809_3;
  wire __tmp_809_4;
  wire __tmp_809_5;
  wire __tmp_809_6;
  wire __tmp_809_7;
  wire __tmp_809_8;
  wire __tmp_809_9;
  wire __tmp_811_1;
  wire __tmp_811_10;
  wire __tmp_811_11;
  wire __tmp_811_12;
  wire __tmp_811_2;
  wire __tmp_811_3;
  wire __tmp_811_4;
  wire __tmp_811_5;
  wire __tmp_811_6;
  wire __tmp_811_7;
  wire __tmp_811_8;
  wire __tmp_811_9;
  wire __tmp_813_1;
  wire __tmp_813_10;
  wire __tmp_813_11;
  wire __tmp_813_12;
  wire __tmp_813_2;
  wire __tmp_813_3;
  wire __tmp_813_4;
  wire __tmp_813_5;
  wire __tmp_813_6;
  wire __tmp_813_7;
  wire __tmp_813_8;
  wire __tmp_813_9;
  wire __tmp_815_1;
  wire __tmp_815_2;
  wire __tmp_815_3;
  wire __tmp_815_4;
  wire __tmp_815_5;
  wire __tmp_815_6;
  wire __tmp_815_7;
  wire __tmp_815_8;
  wire __tmp_815_9;
  wire __tmp_817_1;
  wire __tmp_817_2;
  wire __tmp_817_3;
  wire __tmp_817_4;
  wire __tmp_817_5;
  wire __tmp_817_6;
  wire __tmp_817_7;
  wire __tmp_817_8;
  wire __tmp_817_9;
  wire __tmp_819_1;
  wire __tmp_819_2;
  wire __tmp_819_3;
  wire __tmp_819_4;
  wire __tmp_819_5;
  wire __tmp_819_6;
  wire __tmp_819_7;
  wire __tmp_819_8;
  wire __tmp_819_9;
  wire __tmp_821_1;
  wire __tmp_821_10;
  wire __tmp_821_11;
  wire __tmp_821_12;
  wire __tmp_821_2;
  wire __tmp_821_3;
  wire __tmp_821_4;
  wire __tmp_821_5;
  wire __tmp_821_6;
  wire __tmp_821_7;
  wire __tmp_821_8;
  wire __tmp_821_9;
  wire __tmp_823_1;
  wire __tmp_823_10;
  wire __tmp_823_11;
  wire __tmp_823_12;
  wire __tmp_823_2;
  wire __tmp_823_3;
  wire __tmp_823_4;
  wire __tmp_823_5;
  wire __tmp_823_6;
  wire __tmp_823_7;
  wire __tmp_823_8;
  wire __tmp_823_9;
  wire __tmp_825_1;
  wire __tmp_825_10;
  wire __tmp_825_11;
  wire __tmp_825_12;
  wire __tmp_825_2;
  wire __tmp_825_3;
  wire __tmp_825_4;
  wire __tmp_825_5;
  wire __tmp_825_6;
  wire __tmp_825_7;
  wire __tmp_825_8;
  wire __tmp_825_9;
  wire __tmp_827_1;
  wire __tmp_827_2;
  wire __tmp_827_3;
  wire __tmp_827_4;
  wire __tmp_827_5;
  wire __tmp_827_6;
  wire __tmp_827_7;
  wire __tmp_827_8;
  wire __tmp_827_9;
  wire __tmp_829_1;
  wire __tmp_829_2;
  wire __tmp_829_3;
  wire __tmp_829_4;
  wire __tmp_829_5;
  wire __tmp_829_6;
  wire __tmp_829_7;
  wire __tmp_829_8;
  wire __tmp_829_9;
  wire __tmp_831_1;
  wire __tmp_831_2;
  wire __tmp_831_3;
  wire __tmp_831_4;
  wire __tmp_831_5;
  wire __tmp_831_6;
  wire __tmp_831_7;
  wire __tmp_831_8;
  wire __tmp_831_9;
  wire __tmp_833_1;
  wire __tmp_833_10;
  wire __tmp_833_11;
  wire __tmp_833_12;
  wire __tmp_833_2;
  wire __tmp_833_3;
  wire __tmp_833_4;
  wire __tmp_833_5;
  wire __tmp_833_6;
  wire __tmp_833_7;
  wire __tmp_833_8;
  wire __tmp_833_9;
  wire __tmp_835_1;
  wire __tmp_835_10;
  wire __tmp_835_11;
  wire __tmp_835_12;
  wire __tmp_835_2;
  wire __tmp_835_3;
  wire __tmp_835_4;
  wire __tmp_835_5;
  wire __tmp_835_6;
  wire __tmp_835_7;
  wire __tmp_835_8;
  wire __tmp_835_9;
  wire __tmp_837_1;
  wire __tmp_837_10;
  wire __tmp_837_11;
  wire __tmp_837_12;
  wire __tmp_837_2;
  wire __tmp_837_3;
  wire __tmp_837_4;
  wire __tmp_837_5;
  wire __tmp_837_6;
  wire __tmp_837_7;
  wire __tmp_837_8;
  wire __tmp_837_9;
  wire __tmp_839_1;
  wire __tmp_839_2;
  wire __tmp_839_3;
  wire __tmp_839_4;
  wire __tmp_839_5;
  wire __tmp_839_6;
  wire __tmp_839_7;
  wire __tmp_839_8;
  wire __tmp_839_9;
  wire __tmp_841_1;
  wire __tmp_841_2;
  wire __tmp_841_3;
  wire __tmp_841_4;
  wire __tmp_841_5;
  wire __tmp_841_6;
  wire __tmp_841_7;
  wire __tmp_841_8;
  wire __tmp_841_9;
  wire __tmp_843_1;
  wire __tmp_843_2;
  wire __tmp_843_3;
  wire __tmp_843_4;
  wire __tmp_843_5;
  wire __tmp_843_6;
  wire __tmp_843_7;
  wire __tmp_843_8;
  wire __tmp_843_9;
  wire __tmp_845_1;
  wire __tmp_845_10;
  wire __tmp_845_11;
  wire __tmp_845_12;
  wire __tmp_845_2;
  wire __tmp_845_3;
  wire __tmp_845_4;
  wire __tmp_845_5;
  wire __tmp_845_6;
  wire __tmp_845_7;
  wire __tmp_845_8;
  wire __tmp_845_9;
  wire __tmp_847_1;
  wire __tmp_847_10;
  wire __tmp_847_11;
  wire __tmp_847_12;
  wire __tmp_847_2;
  wire __tmp_847_3;
  wire __tmp_847_4;
  wire __tmp_847_5;
  wire __tmp_847_6;
  wire __tmp_847_7;
  wire __tmp_847_8;
  wire __tmp_847_9;
  wire __tmp_849_1;
  wire __tmp_849_10;
  wire __tmp_849_11;
  wire __tmp_849_12;
  wire __tmp_849_2;
  wire __tmp_849_3;
  wire __tmp_849_4;
  wire __tmp_849_5;
  wire __tmp_849_6;
  wire __tmp_849_7;
  wire __tmp_849_8;
  wire __tmp_849_9;
  wire __tmp_851_1;
  wire __tmp_851_2;
  wire __tmp_851_3;
  wire __tmp_851_4;
  wire __tmp_851_5;
  wire __tmp_851_6;
  wire __tmp_851_7;
  wire __tmp_851_8;
  wire __tmp_851_9;
  wire __tmp_853_1;
  wire __tmp_853_2;
  wire __tmp_853_3;
  wire __tmp_853_4;
  wire __tmp_853_5;
  wire __tmp_853_6;
  wire __tmp_853_7;
  wire __tmp_853_8;
  wire __tmp_853_9;
  wire __tmp_855_1;
  wire __tmp_855_2;
  wire __tmp_855_3;
  wire __tmp_855_4;
  wire __tmp_855_5;
  wire __tmp_855_6;
  wire __tmp_855_7;
  wire __tmp_855_8;
  wire __tmp_855_9;
  wire __tmp_857_1;
  wire __tmp_857_10;
  wire __tmp_857_11;
  wire __tmp_857_12;
  wire __tmp_857_2;
  wire __tmp_857_3;
  wire __tmp_857_4;
  wire __tmp_857_5;
  wire __tmp_857_6;
  wire __tmp_857_7;
  wire __tmp_857_8;
  wire __tmp_857_9;
  wire __tmp_859_1;
  wire __tmp_859_10;
  wire __tmp_859_11;
  wire __tmp_859_12;
  wire __tmp_859_2;
  wire __tmp_859_3;
  wire __tmp_859_4;
  wire __tmp_859_5;
  wire __tmp_859_6;
  wire __tmp_859_7;
  wire __tmp_859_8;
  wire __tmp_859_9;
  wire __tmp_861_1;
  wire __tmp_861_10;
  wire __tmp_861_11;
  wire __tmp_861_12;
  wire __tmp_861_2;
  wire __tmp_861_3;
  wire __tmp_861_4;
  wire __tmp_861_5;
  wire __tmp_861_6;
  wire __tmp_861_7;
  wire __tmp_861_8;
  wire __tmp_861_9;
  wire __tmp_863_1;
  wire __tmp_863_2;
  wire __tmp_863_3;
  wire __tmp_863_4;
  wire __tmp_863_5;
  wire __tmp_863_6;
  wire __tmp_863_7;
  wire __tmp_863_8;
  wire __tmp_863_9;
  wire __tmp_865_1;
  wire __tmp_865_2;
  wire __tmp_865_3;
  wire __tmp_865_4;
  wire __tmp_865_5;
  wire __tmp_865_6;
  wire __tmp_865_7;
  wire __tmp_865_8;
  wire __tmp_865_9;
  wire __tmp_867_1;
  wire __tmp_867_2;
  wire __tmp_867_3;
  wire __tmp_867_4;
  wire __tmp_867_5;
  wire __tmp_867_6;
  wire __tmp_867_7;
  wire __tmp_867_8;
  wire __tmp_867_9;
  wire __tmp_869_1;
  wire __tmp_869_10;
  wire __tmp_869_11;
  wire __tmp_869_12;
  wire __tmp_869_2;
  wire __tmp_869_3;
  wire __tmp_869_4;
  wire __tmp_869_5;
  wire __tmp_869_6;
  wire __tmp_869_7;
  wire __tmp_869_8;
  wire __tmp_869_9;
  wire __tmp_871_1;
  wire __tmp_871_10;
  wire __tmp_871_11;
  wire __tmp_871_12;
  wire __tmp_871_2;
  wire __tmp_871_3;
  wire __tmp_871_4;
  wire __tmp_871_5;
  wire __tmp_871_6;
  wire __tmp_871_7;
  wire __tmp_871_8;
  wire __tmp_871_9;
  wire __tmp_873_1;
  wire __tmp_873_10;
  wire __tmp_873_11;
  wire __tmp_873_12;
  wire __tmp_873_2;
  wire __tmp_873_3;
  wire __tmp_873_4;
  wire __tmp_873_5;
  wire __tmp_873_6;
  wire __tmp_873_7;
  wire __tmp_873_8;
  wire __tmp_873_9;
  wire __tmp_875_1;
  wire __tmp_875_2;
  wire __tmp_875_3;
  wire __tmp_875_4;
  wire __tmp_875_5;
  wire __tmp_875_6;
  wire __tmp_875_7;
  wire __tmp_875_8;
  wire __tmp_875_9;
  wire __tmp_877_1;
  wire __tmp_877_2;
  wire __tmp_877_3;
  wire __tmp_877_4;
  wire __tmp_877_5;
  wire __tmp_877_6;
  wire __tmp_877_7;
  wire __tmp_877_8;
  wire __tmp_877_9;
  wire __tmp_879_1;
  wire __tmp_879_2;
  wire __tmp_879_3;
  wire __tmp_879_4;
  wire __tmp_879_5;
  wire __tmp_879_6;
  wire __tmp_879_7;
  wire __tmp_879_8;
  wire __tmp_879_9;
  wire __tmp_881_1;
  wire __tmp_881_10;
  wire __tmp_881_11;
  wire __tmp_881_12;
  wire __tmp_881_2;
  wire __tmp_881_3;
  wire __tmp_881_4;
  wire __tmp_881_5;
  wire __tmp_881_6;
  wire __tmp_881_7;
  wire __tmp_881_8;
  wire __tmp_881_9;
  wire __tmp_883_1;
  wire __tmp_883_10;
  wire __tmp_883_11;
  wire __tmp_883_12;
  wire __tmp_883_2;
  wire __tmp_883_3;
  wire __tmp_883_4;
  wire __tmp_883_5;
  wire __tmp_883_6;
  wire __tmp_883_7;
  wire __tmp_883_8;
  wire __tmp_883_9;
  wire __tmp_885_1;
  wire __tmp_885_10;
  wire __tmp_885_11;
  wire __tmp_885_12;
  wire __tmp_885_2;
  wire __tmp_885_3;
  wire __tmp_885_4;
  wire __tmp_885_5;
  wire __tmp_885_6;
  wire __tmp_885_7;
  wire __tmp_885_8;
  wire __tmp_885_9;
  wire __tmp_887_1;
  wire __tmp_887_2;
  wire __tmp_887_3;
  wire __tmp_887_4;
  wire __tmp_887_5;
  wire __tmp_887_6;
  wire __tmp_887_7;
  wire __tmp_887_8;
  wire __tmp_887_9;
  wire __tmp_889_1;
  wire __tmp_889_2;
  wire __tmp_889_3;
  wire __tmp_889_4;
  wire __tmp_889_5;
  wire __tmp_889_6;
  wire __tmp_889_7;
  wire __tmp_889_8;
  wire __tmp_889_9;
  wire __tmp_891_1;
  wire __tmp_891_2;
  wire __tmp_891_3;
  wire __tmp_891_4;
  wire __tmp_891_5;
  wire __tmp_891_6;
  wire __tmp_891_7;
  wire __tmp_891_8;
  wire __tmp_891_9;
  wire __tmp_893_1;
  wire __tmp_893_10;
  wire __tmp_893_11;
  wire __tmp_893_12;
  wire __tmp_893_2;
  wire __tmp_893_3;
  wire __tmp_893_4;
  wire __tmp_893_5;
  wire __tmp_893_6;
  wire __tmp_893_7;
  wire __tmp_893_8;
  wire __tmp_893_9;
  wire __tmp_895_1;
  wire __tmp_895_10;
  wire __tmp_895_11;
  wire __tmp_895_12;
  wire __tmp_895_2;
  wire __tmp_895_3;
  wire __tmp_895_4;
  wire __tmp_895_5;
  wire __tmp_895_6;
  wire __tmp_895_7;
  wire __tmp_895_8;
  wire __tmp_895_9;
  wire __tmp_897_1;
  wire __tmp_897_10;
  wire __tmp_897_11;
  wire __tmp_897_12;
  wire __tmp_897_2;
  wire __tmp_897_3;
  wire __tmp_897_4;
  wire __tmp_897_5;
  wire __tmp_897_6;
  wire __tmp_897_7;
  wire __tmp_897_8;
  wire __tmp_897_9;
  wire __tmp_899_1;
  wire __tmp_899_2;
  wire __tmp_899_3;
  wire __tmp_899_4;
  wire __tmp_899_5;
  wire __tmp_899_6;
  wire __tmp_899_7;
  wire __tmp_899_8;
  wire __tmp_899_9;
  wire __tmp_901_1;
  wire __tmp_901_2;
  wire __tmp_901_3;
  wire __tmp_901_4;
  wire __tmp_901_5;
  wire __tmp_901_6;
  wire __tmp_901_7;
  wire __tmp_901_8;
  wire __tmp_901_9;
  wire __tmp_903_1;
  wire __tmp_903_2;
  wire __tmp_903_3;
  wire __tmp_903_4;
  wire __tmp_903_5;
  wire __tmp_903_6;
  wire __tmp_903_7;
  wire __tmp_903_8;
  wire __tmp_903_9;
  wire __tmp_905_1;
  wire __tmp_905_10;
  wire __tmp_905_11;
  wire __tmp_905_12;
  wire __tmp_905_2;
  wire __tmp_905_3;
  wire __tmp_905_4;
  wire __tmp_905_5;
  wire __tmp_905_6;
  wire __tmp_905_7;
  wire __tmp_905_8;
  wire __tmp_905_9;
  wire __tmp_907_1;
  wire __tmp_907_10;
  wire __tmp_907_11;
  wire __tmp_907_12;
  wire __tmp_907_2;
  wire __tmp_907_3;
  wire __tmp_907_4;
  wire __tmp_907_5;
  wire __tmp_907_6;
  wire __tmp_907_7;
  wire __tmp_907_8;
  wire __tmp_907_9;
  wire __tmp_909_1;
  wire __tmp_909_10;
  wire __tmp_909_11;
  wire __tmp_909_12;
  wire __tmp_909_2;
  wire __tmp_909_3;
  wire __tmp_909_4;
  wire __tmp_909_5;
  wire __tmp_909_6;
  wire __tmp_909_7;
  wire __tmp_909_8;
  wire __tmp_909_9;
  wire __tmp_911_1;
  wire __tmp_911_10;
  wire __tmp_911_11;
  wire __tmp_911_12;
  wire __tmp_911_13;
  wire __tmp_911_14;
  wire __tmp_911_15;
  wire __tmp_911_16;
  wire __tmp_911_17;
  wire __tmp_911_18;
  wire __tmp_911_19;
  wire __tmp_911_2;
  wire __tmp_911_3;
  wire __tmp_911_4;
  wire __tmp_911_5;
  wire __tmp_911_6;
  wire __tmp_911_7;
  wire __tmp_911_8;
  wire __tmp_911_9;
  wire __tmp_913_1;
  wire __tmp_913_10;
  wire __tmp_913_11;
  wire __tmp_913_12;
  wire __tmp_913_13;
  wire __tmp_913_14;
  wire __tmp_913_15;
  wire __tmp_913_16;
  wire __tmp_913_17;
  wire __tmp_913_18;
  wire __tmp_913_19;
  wire __tmp_913_2;
  wire __tmp_913_3;
  wire __tmp_913_4;
  wire __tmp_913_5;
  wire __tmp_913_6;
  wire __tmp_913_7;
  wire __tmp_913_8;
  wire __tmp_913_9;
  wire __tmp_915_1;
  wire __tmp_915_10;
  wire __tmp_915_11;
  wire __tmp_915_12;
  wire __tmp_915_13;
  wire __tmp_915_14;
  wire __tmp_915_15;
  wire __tmp_915_16;
  wire __tmp_915_17;
  wire __tmp_915_18;
  wire __tmp_915_19;
  wire __tmp_915_2;
  wire __tmp_915_3;
  wire __tmp_915_4;
  wire __tmp_915_5;
  wire __tmp_915_6;
  wire __tmp_915_7;
  wire __tmp_915_8;
  wire __tmp_915_9;
  wire __tmp_917_1;
  wire __tmp_917_10;
  wire __tmp_917_11;
  wire __tmp_917_12;
  wire __tmp_917_13;
  wire __tmp_917_14;
  wire __tmp_917_15;
  wire __tmp_917_16;
  wire __tmp_917_17;
  wire __tmp_917_18;
  wire __tmp_917_19;
  wire __tmp_917_2;
  wire __tmp_917_3;
  wire __tmp_917_4;
  wire __tmp_917_5;
  wire __tmp_917_6;
  wire __tmp_917_7;
  wire __tmp_917_8;
  wire __tmp_917_9;
  wire __tmp_919_1;
  wire __tmp_919_10;
  wire __tmp_919_11;
  wire __tmp_919_12;
  wire __tmp_919_13;
  wire __tmp_919_14;
  wire __tmp_919_15;
  wire __tmp_919_16;
  wire __tmp_919_17;
  wire __tmp_919_18;
  wire __tmp_919_19;
  wire __tmp_919_2;
  wire __tmp_919_3;
  wire __tmp_919_4;
  wire __tmp_919_5;
  wire __tmp_919_6;
  wire __tmp_919_7;
  wire __tmp_919_8;
  wire __tmp_919_9;
  wire __tmp_921_1;
  wire __tmp_921_10;
  wire __tmp_921_11;
  wire __tmp_921_12;
  wire __tmp_921_13;
  wire __tmp_921_14;
  wire __tmp_921_15;
  wire __tmp_921_16;
  wire __tmp_921_17;
  wire __tmp_921_18;
  wire __tmp_921_19;
  wire __tmp_921_2;
  wire __tmp_921_3;
  wire __tmp_921_4;
  wire __tmp_921_5;
  wire __tmp_921_6;
  wire __tmp_921_7;
  wire __tmp_921_8;
  wire __tmp_921_9;
  wire __tmp_923_1;
  wire __tmp_923_10;
  wire __tmp_923_11;
  wire __tmp_923_12;
  wire __tmp_923_13;
  wire __tmp_923_14;
  wire __tmp_923_15;
  wire __tmp_923_16;
  wire __tmp_923_17;
  wire __tmp_923_18;
  wire __tmp_923_19;
  wire __tmp_923_2;
  wire __tmp_923_3;
  wire __tmp_923_4;
  wire __tmp_923_5;
  wire __tmp_923_6;
  wire __tmp_923_7;
  wire __tmp_923_8;
  wire __tmp_923_9;
  wire __tmp_925_1;
  wire __tmp_925_10;
  wire __tmp_925_11;
  wire __tmp_925_12;
  wire __tmp_925_13;
  wire __tmp_925_14;
  wire __tmp_925_15;
  wire __tmp_925_16;
  wire __tmp_925_17;
  wire __tmp_925_18;
  wire __tmp_925_19;
  wire __tmp_925_2;
  wire __tmp_925_3;
  wire __tmp_925_4;
  wire __tmp_925_5;
  wire __tmp_925_6;
  wire __tmp_925_7;
  wire __tmp_925_8;
  wire __tmp_925_9;
  wire __tmp_927_1;
  wire __tmp_927_10;
  wire __tmp_927_11;
  wire __tmp_927_12;
  wire __tmp_927_13;
  wire __tmp_927_14;
  wire __tmp_927_15;
  wire __tmp_927_16;
  wire __tmp_927_17;
  wire __tmp_927_18;
  wire __tmp_927_19;
  wire __tmp_927_2;
  wire __tmp_927_3;
  wire __tmp_927_4;
  wire __tmp_927_5;
  wire __tmp_927_6;
  wire __tmp_927_7;
  wire __tmp_927_8;
  wire __tmp_927_9;
  wire __tmp_929_1;
  wire __tmp_929_2;
  wire __tmp_929_3;
  wire __tmp_929_4;
  wire __tmp_929_5;
  wire __tmp_929_6;
  wire __tmp_931_1;
  wire __tmp_931_2;
  wire __tmp_931_3;
  wire __tmp_931_4;
  wire __tmp_931_5;
  wire __tmp_931_6;
  wire __tmp_933_1;
  wire __tmp_933_2;
  wire __tmp_933_3;
  wire __tmp_933_4;
  wire __tmp_933_5;
  wire __tmp_933_6;
  wire __tmp_935_1;
  wire __tmp_935_10;
  wire __tmp_935_11;
  wire __tmp_935_12;
  wire __tmp_935_13;
  wire __tmp_935_14;
  wire __tmp_935_15;
  wire __tmp_935_16;
  wire __tmp_935_17;
  wire __tmp_935_18;
  wire __tmp_935_19;
  wire __tmp_935_2;
  wire __tmp_935_20;
  wire __tmp_935_21;
  wire __tmp_935_22;
  wire __tmp_935_23;
  wire __tmp_935_24;
  wire __tmp_935_3;
  wire __tmp_935_4;
  wire __tmp_935_5;
  wire __tmp_935_6;
  wire __tmp_935_7;
  wire __tmp_935_8;
  wire __tmp_935_9;
  wire __tmp_937_1;
  wire __tmp_937_10;
  wire __tmp_937_11;
  wire __tmp_937_12;
  wire __tmp_937_13;
  wire __tmp_937_14;
  wire __tmp_937_15;
  wire __tmp_937_16;
  wire __tmp_937_17;
  wire __tmp_937_18;
  wire __tmp_937_19;
  wire __tmp_937_2;
  wire __tmp_937_20;
  wire __tmp_937_21;
  wire __tmp_937_22;
  wire __tmp_937_23;
  wire __tmp_937_3;
  wire __tmp_937_4;
  wire __tmp_937_5;
  wire __tmp_937_6;
  wire __tmp_937_7;
  wire __tmp_937_8;
  wire __tmp_937_9;
  wire __tmp_939_1;
  wire __tmp_939_10;
  wire __tmp_939_11;
  wire __tmp_939_12;
  wire __tmp_939_13;
  wire __tmp_939_14;
  wire __tmp_939_15;
  wire __tmp_939_16;
  wire __tmp_939_17;
  wire __tmp_939_18;
  wire __tmp_939_19;
  wire __tmp_939_2;
  wire __tmp_939_20;
  wire __tmp_939_21;
  wire __tmp_939_22;
  wire __tmp_939_23;
  wire __tmp_939_3;
  wire __tmp_939_4;
  wire __tmp_939_5;
  wire __tmp_939_6;
  wire __tmp_939_7;
  wire __tmp_939_8;
  wire __tmp_939_9;
  wire __tmp_941_1;
  wire __tmp_941_10;
  wire __tmp_941_11;
  wire __tmp_941_12;
  wire __tmp_941_13;
  wire __tmp_941_14;
  wire __tmp_941_15;
  wire __tmp_941_16;
  wire __tmp_941_17;
  wire __tmp_941_18;
  wire __tmp_941_19;
  wire __tmp_941_2;
  wire __tmp_941_20;
  wire __tmp_941_21;
  wire __tmp_941_22;
  wire __tmp_941_23;
  wire __tmp_941_3;
  wire __tmp_941_4;
  wire __tmp_941_5;
  wire __tmp_941_6;
  wire __tmp_941_7;
  wire __tmp_941_8;
  wire __tmp_941_9;
  wire __tmp_943_1;
  wire __tmp_943_2;
  wire __tmp_943_3;
  wire __tmp_943_4;
  wire __tmp_943_5;
  wire __tmp_943_6;
  wire __tmp_943_7;
  wire __tmp_943_8;
  wire __tmp_943_9;
  wire __tmp_945_1;
  wire __tmp_945_2;
  wire __tmp_945_3;
  wire __tmp_945_4;
  wire __tmp_945_5;
  wire __tmp_945_6;
  wire __tmp_945_7;
  wire __tmp_945_8;
  wire __tmp_945_9;
  wire __tmp_947_1;
  wire __tmp_947_2;
  wire __tmp_947_3;
  wire __tmp_947_4;
  wire __tmp_947_5;
  wire __tmp_947_6;
  wire __tmp_947_7;
  wire __tmp_947_8;
  wire __tmp_947_9;
  wire __tmp_949_1;
  wire __tmp_949_10;
  wire __tmp_949_11;
  wire __tmp_949_12;
  wire __tmp_949_13;
  wire __tmp_949_14;
  wire __tmp_949_15;
  wire __tmp_949_16;
  wire __tmp_949_17;
  wire __tmp_949_18;
  wire __tmp_949_19;
  wire __tmp_949_2;
  wire __tmp_949_20;
  wire __tmp_949_21;
  wire __tmp_949_22;
  wire __tmp_949_23;
  wire __tmp_949_24;
  wire __tmp_949_25;
  wire __tmp_949_26;
  wire __tmp_949_27;
  wire __tmp_949_28;
  wire __tmp_949_29;
  wire __tmp_949_3;
  wire __tmp_949_30;
  wire __tmp_949_31;
  wire __tmp_949_4;
  wire __tmp_949_5;
  wire __tmp_949_6;
  wire __tmp_949_7;
  wire __tmp_949_8;
  wire __tmp_949_9;
  wire __tmp_951_1;
  wire __tmp_951_10;
  wire __tmp_951_11;
  wire __tmp_951_12;
  wire __tmp_951_13;
  wire __tmp_951_14;
  wire __tmp_951_15;
  wire __tmp_951_16;
  wire __tmp_951_17;
  wire __tmp_951_18;
  wire __tmp_951_19;
  wire __tmp_951_2;
  wire __tmp_951_20;
  wire __tmp_951_21;
  wire __tmp_951_22;
  wire __tmp_951_23;
  wire __tmp_951_24;
  wire __tmp_951_25;
  wire __tmp_951_26;
  wire __tmp_951_27;
  wire __tmp_951_28;
  wire __tmp_951_29;
  wire __tmp_951_3;
  wire __tmp_951_30;
  wire __tmp_951_31;
  wire __tmp_951_4;
  wire __tmp_951_5;
  wire __tmp_951_6;
  wire __tmp_951_7;
  wire __tmp_951_8;
  wire __tmp_951_9;
  wire __tmp_953_1;
  wire __tmp_953_10;
  wire __tmp_953_11;
  wire __tmp_953_12;
  wire __tmp_953_13;
  wire __tmp_953_14;
  wire __tmp_953_15;
  wire __tmp_953_16;
  wire __tmp_953_17;
  wire __tmp_953_18;
  wire __tmp_953_19;
  wire __tmp_953_2;
  wire __tmp_953_20;
  wire __tmp_953_21;
  wire __tmp_953_22;
  wire __tmp_953_23;
  wire __tmp_953_24;
  wire __tmp_953_25;
  wire __tmp_953_26;
  wire __tmp_953_27;
  wire __tmp_953_28;
  wire __tmp_953_29;
  wire __tmp_953_3;
  wire __tmp_953_30;
  wire __tmp_953_31;
  wire __tmp_953_4;
  wire __tmp_953_5;
  wire __tmp_953_6;
  wire __tmp_953_7;
  wire __tmp_953_8;
  wire __tmp_953_9;
  wire __tmp_955_1;
  wire __tmp_955_10;
  wire __tmp_955_11;
  wire __tmp_955_12;
  wire __tmp_955_2;
  wire __tmp_955_3;
  wire __tmp_955_4;
  wire __tmp_955_5;
  wire __tmp_955_6;
  wire __tmp_955_7;
  wire __tmp_955_8;
  wire __tmp_955_9;
  wire __tmp_957_1;
  wire __tmp_957_10;
  wire __tmp_957_11;
  wire __tmp_957_12;
  wire __tmp_957_2;
  wire __tmp_957_3;
  wire __tmp_957_4;
  wire __tmp_957_5;
  wire __tmp_957_6;
  wire __tmp_957_7;
  wire __tmp_957_8;
  wire __tmp_957_9;
  wire __tmp_959_1;
  wire __tmp_959_10;
  wire __tmp_959_11;
  wire __tmp_959_12;
  wire __tmp_959_2;
  wire __tmp_959_3;
  wire __tmp_959_4;
  wire __tmp_959_5;
  wire __tmp_959_6;
  wire __tmp_959_7;
  wire __tmp_959_8;
  wire __tmp_959_9;
  wire __tmp_961_1;
  wire __tmp_961_10;
  wire __tmp_961_11;
  wire __tmp_961_12;
  wire __tmp_961_13;
  wire __tmp_961_14;
  wire __tmp_961_15;
  wire __tmp_961_16;
  wire __tmp_961_17;
  wire __tmp_961_18;
  wire __tmp_961_19;
  wire __tmp_961_2;
  wire __tmp_961_20;
  wire __tmp_961_21;
  wire __tmp_961_22;
  wire __tmp_961_23;
  wire __tmp_961_24;
  wire __tmp_961_25;
  wire __tmp_961_26;
  wire __tmp_961_27;
  wire __tmp_961_28;
  wire __tmp_961_29;
  wire __tmp_961_3;
  wire __tmp_961_30;
  wire __tmp_961_31;
  wire __tmp_961_32;
  wire __tmp_961_33;
  wire __tmp_961_34;
  wire __tmp_961_35;
  wire __tmp_961_36;
  wire __tmp_961_37;
  wire __tmp_961_38;
  wire __tmp_961_39;
  wire __tmp_961_4;
  wire __tmp_961_40;
  wire __tmp_961_41;
  wire __tmp_961_42;
  wire __tmp_961_43;
  wire __tmp_961_44;
  wire __tmp_961_45;
  wire __tmp_961_46;
  wire __tmp_961_5;
  wire __tmp_961_6;
  wire __tmp_961_7;
  wire __tmp_961_8;
  wire __tmp_961_9;
  wire __tmp_963_1;
  wire __tmp_963_10;
  wire __tmp_963_11;
  wire __tmp_963_12;
  wire __tmp_963_13;
  wire __tmp_963_14;
  wire __tmp_963_15;
  wire __tmp_963_16;
  wire __tmp_963_17;
  wire __tmp_963_18;
  wire __tmp_963_19;
  wire __tmp_963_2;
  wire __tmp_963_20;
  wire __tmp_963_21;
  wire __tmp_963_22;
  wire __tmp_963_23;
  wire __tmp_963_24;
  wire __tmp_963_25;
  wire __tmp_963_26;
  wire __tmp_963_27;
  wire __tmp_963_28;
  wire __tmp_963_29;
  wire __tmp_963_3;
  wire __tmp_963_30;
  wire __tmp_963_31;
  wire __tmp_963_32;
  wire __tmp_963_33;
  wire __tmp_963_34;
  wire __tmp_963_35;
  wire __tmp_963_36;
  wire __tmp_963_37;
  wire __tmp_963_38;
  wire __tmp_963_39;
  wire __tmp_963_4;
  wire __tmp_963_40;
  wire __tmp_963_41;
  wire __tmp_963_42;
  wire __tmp_963_43;
  wire __tmp_963_44;
  wire __tmp_963_45;
  wire __tmp_963_46;
  wire __tmp_963_5;
  wire __tmp_963_6;
  wire __tmp_963_7;
  wire __tmp_963_8;
  wire __tmp_963_9;
  wire __tmp_965_1;
  wire __tmp_965_10;
  wire __tmp_965_11;
  wire __tmp_965_12;
  wire __tmp_965_13;
  wire __tmp_965_14;
  wire __tmp_965_15;
  wire __tmp_965_16;
  wire __tmp_965_17;
  wire __tmp_965_18;
  wire __tmp_965_19;
  wire __tmp_965_2;
  wire __tmp_965_20;
  wire __tmp_965_21;
  wire __tmp_965_22;
  wire __tmp_965_23;
  wire __tmp_965_24;
  wire __tmp_965_25;
  wire __tmp_965_26;
  wire __tmp_965_27;
  wire __tmp_965_28;
  wire __tmp_965_29;
  wire __tmp_965_3;
  wire __tmp_965_30;
  wire __tmp_965_31;
  wire __tmp_965_32;
  wire __tmp_965_33;
  wire __tmp_965_34;
  wire __tmp_965_35;
  wire __tmp_965_36;
  wire __tmp_965_37;
  wire __tmp_965_38;
  wire __tmp_965_39;
  wire __tmp_965_4;
  wire __tmp_965_40;
  wire __tmp_965_41;
  wire __tmp_965_42;
  wire __tmp_965_43;
  wire __tmp_965_44;
  wire __tmp_965_45;
  wire __tmp_965_46;
  wire __tmp_965_5;
  wire __tmp_965_6;
  wire __tmp_965_7;
  wire __tmp_965_8;
  wire __tmp_965_9;
  wire __tmp_967_1;
  wire __tmp_967_10;
  wire __tmp_967_11;
  wire __tmp_967_12;
  wire __tmp_967_13;
  wire __tmp_967_14;
  wire __tmp_967_15;
  wire __tmp_967_16;
  wire __tmp_967_17;
  wire __tmp_967_18;
  wire __tmp_967_19;
  wire __tmp_967_2;
  wire __tmp_967_20;
  wire __tmp_967_21;
  wire __tmp_967_22;
  wire __tmp_967_23;
  wire __tmp_967_24;
  wire __tmp_967_25;
  wire __tmp_967_26;
  wire __tmp_967_27;
  wire __tmp_967_28;
  wire __tmp_967_29;
  wire __tmp_967_3;
  wire __tmp_967_30;
  wire __tmp_967_31;
  wire __tmp_967_32;
  wire __tmp_967_33;
  wire __tmp_967_34;
  wire __tmp_967_35;
  wire __tmp_967_36;
  wire __tmp_967_37;
  wire __tmp_967_38;
  wire __tmp_967_39;
  wire __tmp_967_4;
  wire __tmp_967_40;
  wire __tmp_967_41;
  wire __tmp_967_42;
  wire __tmp_967_43;
  wire __tmp_967_44;
  wire __tmp_967_45;
  wire __tmp_967_46;
  wire __tmp_967_5;
  wire __tmp_967_6;
  wire __tmp_967_7;
  wire __tmp_967_8;
  wire __tmp_967_9;
  wire __tmp_969_1;
  wire __tmp_969_10;
  wire __tmp_969_11;
  wire __tmp_969_12;
  wire __tmp_969_13;
  wire __tmp_969_14;
  wire __tmp_969_15;
  wire __tmp_969_16;
  wire __tmp_969_17;
  wire __tmp_969_18;
  wire __tmp_969_19;
  wire __tmp_969_2;
  wire __tmp_969_20;
  wire __tmp_969_21;
  wire __tmp_969_22;
  wire __tmp_969_23;
  wire __tmp_969_24;
  wire __tmp_969_25;
  wire __tmp_969_26;
  wire __tmp_969_27;
  wire __tmp_969_28;
  wire __tmp_969_29;
  wire __tmp_969_3;
  wire __tmp_969_30;
  wire __tmp_969_31;
  wire __tmp_969_32;
  wire __tmp_969_33;
  wire __tmp_969_34;
  wire __tmp_969_35;
  wire __tmp_969_36;
  wire __tmp_969_37;
  wire __tmp_969_38;
  wire __tmp_969_39;
  wire __tmp_969_4;
  wire __tmp_969_40;
  wire __tmp_969_41;
  wire __tmp_969_42;
  wire __tmp_969_5;
  wire __tmp_969_6;
  wire __tmp_969_7;
  wire __tmp_969_8;
  wire __tmp_969_9;
  wire __tmp_976_1;
  wire [7:0] __tmp_977_1;
  wire __tmp_988_1;
  wire [7:0] __tmp_989_1;
  wire [31:0] __variable_wdata_0;
  wire [5:0] __variable_wdata_1;
  wire [7:0] __variable_wdata_105;
  wire [3:0] __variable_wdata_106;
  wire [3:0] __variable_wdata_107;
  wire [7:0] __variable_wdata_122;
  wire [3:0] __variable_wdata_123;
  wire [3:0] __variable_wdata_124;
  wire [7:0] __variable_wdata_139;
  wire [3:0] __variable_wdata_140;
  wire [3:0] __variable_wdata_141;
  wire [7:0] __variable_wdata_156;
  wire [3:0] __variable_wdata_157;
  wire [3:0] __variable_wdata_158;
  wire [7:0] __variable_wdata_173;
  wire [3:0] __variable_wdata_174;
  wire [3:0] __variable_wdata_175;
  wire [7:0] __variable_wdata_190;
  wire [3:0] __variable_wdata_191;
  wire [3:0] __variable_wdata_192;
  wire [31:0] __variable_wdata_2;
  wire [7:0] __variable_wdata_207;
  wire [7:0] __variable_wdata_208;
  wire [5:0] __variable_wdata_214;
  wire [1:0] __variable_wdata_215;
  wire [1:0] __variable_wdata_216;
  wire [8:0] __variable_wdata_217;
  wire [31:0] __variable_wdata_22;
  wire [7:0] __variable_wdata_230;
  wire [7:0] __variable_wdata_237;
  wire [31:0] __variable_wdata_24;
  wire [7:0] __variable_wdata_244;
  wire [31:0] __variable_wdata_25;
  wire [7:0] __variable_wdata_251;
  wire [7:0] __variable_wdata_258;
  wire [31:0] __variable_wdata_26;
  wire __variable_wdata_264;
  wire __variable_wdata_265;
  wire [3:0] __variable_wdata_266;
  wire [7:0] __variable_wdata_268;
  wire [7:0] __variable_wdata_269;
  wire [31:0] __variable_wdata_27;
  wire [7:0] __variable_wdata_270;
  wire [7:0] __variable_wdata_271;
  wire [7:0] __variable_wdata_272;
  wire [7:0] __variable_wdata_273;
  wire [7:0] __variable_wdata_274;
  wire [7:0] __variable_wdata_275;
  wire [7:0] __variable_wdata_276;
  wire [31:0] __variable_wdata_28;
  wire [31:0] __variable_wdata_29;
  wire [31:0] __variable_wdata_30;
  wire [31:0] __variable_wdata_31;
  wire [31:0] __variable_wdata_32;
  wire [31:0] __variable_wdata_38;
  wire [7:0] __variable_wdata_39;
  wire [5:0] __variable_wdata_40;
  wire [3:0] __variable_wdata_502;
  wire [3:0] __variable_wdata_503;
  wire [3:0] __variable_wdata_504;
  wire [3:0] __variable_wdata_505;
  wire [3:0] __variable_wdata_506;
  wire [3:0] __variable_wdata_507;
  wire [3:0] __variable_wdata_508;
  wire [3:0] __variable_wdata_509;
  wire [3:0] __variable_wdata_510;
  wire [7:0] __variable_wdata_54;
  wire [3:0] __variable_wdata_55;
  wire [3:0] __variable_wdata_56;
  wire [7:0] __variable_wdata_71;
  wire [3:0] __variable_wdata_72;
  wire [3:0] __variable_wdata_73;
  wire [2:0] __variable_wdata_777;
  wire [7:0] __variable_wdata_778;
  wire [3:0] __variable_wdata_779;
  wire [10:0] __variable_wdata_796;
  wire __variable_wdata_797;
  wire __variable_wdata_798;
  wire __variable_wdata_799;
  wire [7:0] __variable_wdata_812;
  wire [7:0] __variable_wdata_819;
  wire [7:0] __variable_wdata_826;
  wire [7:0] __variable_wdata_833;
  wire [7:0] __variable_wdata_840;
  wire __variable_wdata_846;
  wire __variable_wdata_847;
  wire [3:0] __variable_wdata_848;
  wire [1:0] __variable_wdata_849;
  wire [7:0] __variable_wdata_850;
  wire [3:0] __variable_wdata_864;
  wire [7:0] __variable_wdata_88;
  wire [3:0] __variable_wdata_89;
  wire [3:0] __variable_wdata_90;
  wire [31:0] _acc_0_fsm;
  wire _acc_0_reduce_reset;
  wire _acc_0_rshift_idle;
  wire _acc_0_rshift_source_ram_rvalid;
  wire _acc_0_sum_sink_wenable;
  wire _acc_0_valid_sink_wenable;
  wire _acc_0_x_idle;
  wire _acc_0_x_source_ram_rvalid;
  wire [31:0] _add_tree_1_fsm;
  wire _add_tree_1_sum_sink_wenable;
  wire _add_tree_1_var0_idle;
  wire _add_tree_1_var0_source_ram_rvalid;
  wire [31:0] _add_tree_2_fsm;
  wire _add_tree_2_sum_sink_wenable;
  wire _add_tree_2_var0_idle;
  wire _add_tree_2_var0_source_ram_rvalid;
  wire _add_tree_2_var1_idle;
  wire _add_tree_2_var1_source_ram_rvalid;
  wire _add_tree_2_var2_idle;
  wire _add_tree_2_var2_source_ram_rvalid;
  wire _add_tree_2_var3_idle;
  wire _add_tree_2_var3_source_ram_rvalid;
  wire _add_tree_2_var4_idle;
  wire _add_tree_2_var4_source_ram_rvalid;
  wire _add_tree_2_var5_idle;
  wire _add_tree_2_var5_source_ram_rvalid;
  wire _add_tree_2_var6_idle;
  wire _add_tree_2_var6_source_ram_rvalid;
  wire _add_tree_2_var7_idle;
  wire _add_tree_2_var7_source_ram_rvalid;
  wire _add_tree_2_var8_idle;
  wire _add_tree_2_var8_source_ram_rvalid;
  wire [31:0] _cast_data_23;
  wire [31:0] _cast_src_23;
  wire [11:0] _cond_data_101;
  wire [11:0] _cond_data_118;
  wire [31:0] _cond_data_13;
  wire [11:0] _cond_data_135;
  wire [11:0] _cond_data_152;
  wire [11:0] _cond_data_169;
  wire [11:0] _cond_data_186;
  wire [11:0] _cond_data_203;
  wire [7:0] _cond_data_235;
  wire [7:0] _cond_data_242;
  wire [7:0] _cond_data_249;
  wire [7:0] _cond_data_256;
  wire [7:0] _cond_data_263;
  wire [7:0] _cond_data_279;
  wire [7:0] _cond_data_283;
  wire [7:0] _cond_data_286;
  wire [7:0] _cond_data_289;
  wire [7:0] _cond_data_293;
  wire [7:0] _cond_data_296;
  wire [7:0] _cond_data_299;
  wire [7:0] _cond_data_303;
  wire [7:0] _cond_data_306;
  wire [7:0] _cond_data_309;
  wire [7:0] _cond_data_313;
  wire [7:0] _cond_data_316;
  wire [7:0] _cond_data_319;
  wire [7:0] _cond_data_323;
  wire [7:0] _cond_data_326;
  wire [7:0] _cond_data_329;
  wire [7:0] _cond_data_333;
  wire [7:0] _cond_data_336;
  wire [7:0] _cond_data_339;
  wire [7:0] _cond_data_343;
  wire [7:0] _cond_data_346;
  wire [7:0] _cond_data_349;
  wire [7:0] _cond_data_353;
  wire [7:0] _cond_data_356;
  wire [7:0] _cond_data_359;
  wire [7:0] _cond_data_363;
  wire [7:0] _cond_data_366;
  wire [7:0] _cond_data_369;
  wire [7:0] _cond_data_373;
  wire [7:0] _cond_data_376;
  wire [7:0] _cond_data_379;
  wire [7:0] _cond_data_383;
  wire [7:0] _cond_data_386;
  wire [7:0] _cond_data_389;
  wire [7:0] _cond_data_393;
  wire [7:0] _cond_data_396;
  wire [7:0] _cond_data_399;
  wire [7:0] _cond_data_403;
  wire [7:0] _cond_data_406;
  wire [7:0] _cond_data_409;
  wire [7:0] _cond_data_413;
  wire [7:0] _cond_data_416;
  wire [7:0] _cond_data_419;
  wire [7:0] _cond_data_423;
  wire [7:0] _cond_data_426;
  wire [7:0] _cond_data_429;
  wire [7:0] _cond_data_433;
  wire [7:0] _cond_data_436;
  wire [7:0] _cond_data_439;
  wire [7:0] _cond_data_443;
  wire [7:0] _cond_data_446;
  wire [7:0] _cond_data_449;
  wire [39:0] _cond_data_45;
  wire [7:0] _cond_data_453;
  wire [7:0] _cond_data_456;
  wire [39:0] _cond_data_49;
  wire [7:0] _cond_data_53;
  wire [7:0] _cond_data_575;
  wire [7:0] _cond_data_577;
  wire [7:0] _cond_data_579;
  wire [7:0] _cond_data_581;
  wire [7:0] _cond_data_583;
  wire [7:0] _cond_data_585;
  wire [7:0] _cond_data_587;
  wire [7:0] _cond_data_589;
  wire [7:0] _cond_data_591;
  wire [11:0] _cond_data_67;
  wire [7:0] _cond_data_775;
  wire [8:0] _cond_data_791;
  wire [7:0] _cond_data_817;
  wire [7:0] _cond_data_824;
  wire [7:0] _cond_data_831;
  wire [7:0] _cond_data_838;
  wire [11:0] _cond_data_84;
  wire [7:0] _cond_data_845;
  wire [7:0] _cond_data_853;
  wire [7:0] _cond_data_857;
  wire [7:0] _cond_data_873;
  wire [7:0] _cond_data_890;
  wire [7:0] _cond_data_893;
  wire [7:0] _cond_data_896;
  wire _control_conv2d_16_cond_14_2_1;
  wire _control_conv2d_16_cond_15_3_1;
  wire _control_conv2d_16_cond_23_4_1;
  wire _control_conv2d_16_cond_24_5_1;
  wire _control_conv2d_16_cond_30_6_1;
  wire _control_conv2d_16_cond_31_7_1;
  wire _control_conv2d_16_cond_37_8_1;
  wire _control_conv2d_16_cond_38_9_1;
  wire _control_conv2d_16_cond_3_0_1;
  wire _control_conv2d_16_cond_48_10_1;
  wire _control_conv2d_16_cond_8_1_1;
  wire _control_matmul_29_cond_14_2_1;
  wire _control_matmul_29_cond_22_3_1;
  wire _control_matmul_29_cond_32_4_1;
  wire _control_matmul_29_cond_3_0_1;
  wire _control_matmul_29_cond_8_1_1;
  wire _control_max_pool_serial_18_cond_11_1_1;
  wire _control_max_pool_serial_18_cond_19_2_1;
  wire _control_max_pool_serial_18_cond_5_0_1;
  wire [31:0] _counter_count_782;
  wire [31:0] _counter_data_782;
  wire [31:0] _d1__maxi_read_fsm;
  wire [31:0] _d1__maxi_write_fsm;
  wire [31:0] _d1_control_conv2d_16;
  wire [31:0] _d1_control_matmul_29;
  wire [31:0] _d1_control_max_pool_serial_18;
  wire [31:0] _dataflow_cat_data_107;
  wire [31:0] _dataflow_cat_data_167;
  wire [31:0] _dataflow_cat_data_98;
  wire [31:0] _dataflow_cat_odata_107;
  wire [31:0] _dataflow_cat_odata_167;
  wire [31:0] _dataflow_cat_odata_98;
  wire _dataflow_cat_ovalid_107;
  wire _dataflow_cat_ovalid_167;
  wire _dataflow_cat_ovalid_98;
  wire _dataflow_cat_valid_107;
  wire _dataflow_cat_valid_167;
  wire _dataflow_cat_valid_98;
  wire [7:0] _dataflow_slice_data_111;
  wire [7:0] _dataflow_slice_data_114;
  wire [7:0] _dataflow_slice_data_117;
  wire [7:0] _dataflow_slice_data_12;
  wire [7:0] _dataflow_slice_data_120;
  wire [3:0] _dataflow_slice_data_124;
  wire [3:0] _dataflow_slice_data_127;
  wire [3:0] _dataflow_slice_data_130;
  wire [3:0] _dataflow_slice_data_133;
  wire [3:0] _dataflow_slice_data_136;
  wire [3:0] _dataflow_slice_data_139;
  wire [3:0] _dataflow_slice_data_142;
  wire [3:0] _dataflow_slice_data_145;
  wire [7:0] _dataflow_slice_data_149;
  wire [7:0] _dataflow_slice_data_152;
  wire [7:0] _dataflow_slice_data_155;
  wire [7:0] _dataflow_slice_data_158;
  wire [7:0] _dataflow_slice_data_16;
  wire [7:0] _dataflow_slice_data_19;
  wire [7:0] _dataflow_slice_data_22;
  wire [7:0] _dataflow_slice_data_25;
  wire [3:0] _dataflow_slice_data_29;
  wire [7:0] _dataflow_slice_data_3;
  wire [3:0] _dataflow_slice_data_32;
  wire [3:0] _dataflow_slice_data_35;
  wire [3:0] _dataflow_slice_data_38;
  wire [3:0] _dataflow_slice_data_41;
  wire [3:0] _dataflow_slice_data_44;
  wire [3:0] _dataflow_slice_data_47;
  wire [3:0] _dataflow_slice_data_50;
  wire [7:0] _dataflow_slice_data_54;
  wire [7:0] _dataflow_slice_data_57;
  wire [7:0] _dataflow_slice_data_6;
  wire [7:0] _dataflow_slice_data_60;
  wire [7:0] _dataflow_slice_data_63;
  wire [7:0] _dataflow_slice_data_67;
  wire [7:0] _dataflow_slice_data_70;
  wire [7:0] _dataflow_slice_data_73;
  wire [7:0] _dataflow_slice_data_76;
  wire [7:0] _dataflow_slice_data_80;
  wire [7:0] _dataflow_slice_data_83;
  wire [7:0] _dataflow_slice_data_86;
  wire [7:0] _dataflow_slice_data_89;
  wire [7:0] _dataflow_slice_data_9;
  wire [7:0] _dataflow_slice_odata_111;
  wire [7:0] _dataflow_slice_odata_114;
  wire [7:0] _dataflow_slice_odata_117;
  wire [7:0] _dataflow_slice_odata_12;
  wire [7:0] _dataflow_slice_odata_120;
  wire [3:0] _dataflow_slice_odata_124;
  wire [3:0] _dataflow_slice_odata_127;
  wire [3:0] _dataflow_slice_odata_130;
  wire [3:0] _dataflow_slice_odata_133;
  wire [3:0] _dataflow_slice_odata_136;
  wire [3:0] _dataflow_slice_odata_139;
  wire [3:0] _dataflow_slice_odata_142;
  wire [3:0] _dataflow_slice_odata_145;
  wire [7:0] _dataflow_slice_odata_149;
  wire [7:0] _dataflow_slice_odata_152;
  wire [7:0] _dataflow_slice_odata_155;
  wire [7:0] _dataflow_slice_odata_158;
  wire [7:0] _dataflow_slice_odata_16;
  wire [7:0] _dataflow_slice_odata_19;
  wire [7:0] _dataflow_slice_odata_22;
  wire [7:0] _dataflow_slice_odata_25;
  wire [3:0] _dataflow_slice_odata_29;
  wire [7:0] _dataflow_slice_odata_3;
  wire [3:0] _dataflow_slice_odata_32;
  wire [3:0] _dataflow_slice_odata_35;
  wire [3:0] _dataflow_slice_odata_38;
  wire [3:0] _dataflow_slice_odata_41;
  wire [3:0] _dataflow_slice_odata_44;
  wire [3:0] _dataflow_slice_odata_47;
  wire [3:0] _dataflow_slice_odata_50;
  wire [7:0] _dataflow_slice_odata_54;
  wire [7:0] _dataflow_slice_odata_57;
  wire [7:0] _dataflow_slice_odata_6;
  wire [7:0] _dataflow_slice_odata_60;
  wire [7:0] _dataflow_slice_odata_63;
  wire [7:0] _dataflow_slice_odata_67;
  wire [7:0] _dataflow_slice_odata_70;
  wire [7:0] _dataflow_slice_odata_73;
  wire [7:0] _dataflow_slice_odata_76;
  wire [7:0] _dataflow_slice_odata_80;
  wire [7:0] _dataflow_slice_odata_83;
  wire [7:0] _dataflow_slice_odata_86;
  wire [7:0] _dataflow_slice_odata_89;
  wire [7:0] _dataflow_slice_odata_9;
  wire _dataflow_slice_ovalid_111;
  wire _dataflow_slice_ovalid_114;
  wire _dataflow_slice_ovalid_117;
  wire _dataflow_slice_ovalid_12;
  wire _dataflow_slice_ovalid_120;
  wire _dataflow_slice_ovalid_124;
  wire _dataflow_slice_ovalid_127;
  wire _dataflow_slice_ovalid_130;
  wire _dataflow_slice_ovalid_133;
  wire _dataflow_slice_ovalid_136;
  wire _dataflow_slice_ovalid_139;
  wire _dataflow_slice_ovalid_142;
  wire _dataflow_slice_ovalid_145;
  wire _dataflow_slice_ovalid_149;
  wire _dataflow_slice_ovalid_152;
  wire _dataflow_slice_ovalid_155;
  wire _dataflow_slice_ovalid_158;
  wire _dataflow_slice_ovalid_16;
  wire _dataflow_slice_ovalid_19;
  wire _dataflow_slice_ovalid_22;
  wire _dataflow_slice_ovalid_25;
  wire _dataflow_slice_ovalid_29;
  wire _dataflow_slice_ovalid_3;
  wire _dataflow_slice_ovalid_32;
  wire _dataflow_slice_ovalid_35;
  wire _dataflow_slice_ovalid_38;
  wire _dataflow_slice_ovalid_41;
  wire _dataflow_slice_ovalid_44;
  wire _dataflow_slice_ovalid_47;
  wire _dataflow_slice_ovalid_50;
  wire _dataflow_slice_ovalid_54;
  wire _dataflow_slice_ovalid_57;
  wire _dataflow_slice_ovalid_6;
  wire _dataflow_slice_ovalid_60;
  wire _dataflow_slice_ovalid_63;
  wire _dataflow_slice_ovalid_67;
  wire _dataflow_slice_ovalid_70;
  wire _dataflow_slice_ovalid_73;
  wire _dataflow_slice_ovalid_76;
  wire _dataflow_slice_ovalid_80;
  wire _dataflow_slice_ovalid_83;
  wire _dataflow_slice_ovalid_86;
  wire _dataflow_slice_ovalid_89;
  wire _dataflow_slice_ovalid_9;
  wire _dataflow_slice_valid_111;
  wire _dataflow_slice_valid_114;
  wire _dataflow_slice_valid_117;
  wire _dataflow_slice_valid_12;
  wire _dataflow_slice_valid_120;
  wire _dataflow_slice_valid_124;
  wire _dataflow_slice_valid_127;
  wire _dataflow_slice_valid_130;
  wire _dataflow_slice_valid_133;
  wire _dataflow_slice_valid_136;
  wire _dataflow_slice_valid_139;
  wire _dataflow_slice_valid_142;
  wire _dataflow_slice_valid_145;
  wire _dataflow_slice_valid_149;
  wire _dataflow_slice_valid_152;
  wire _dataflow_slice_valid_155;
  wire _dataflow_slice_valid_158;
  wire _dataflow_slice_valid_16;
  wire _dataflow_slice_valid_19;
  wire _dataflow_slice_valid_22;
  wire _dataflow_slice_valid_25;
  wire _dataflow_slice_valid_29;
  wire _dataflow_slice_valid_3;
  wire _dataflow_slice_valid_32;
  wire _dataflow_slice_valid_35;
  wire _dataflow_slice_valid_38;
  wire _dataflow_slice_valid_41;
  wire _dataflow_slice_valid_44;
  wire _dataflow_slice_valid_47;
  wire _dataflow_slice_valid_50;
  wire _dataflow_slice_valid_54;
  wire _dataflow_slice_valid_57;
  wire _dataflow_slice_valid_6;
  wire _dataflow_slice_valid_60;
  wire _dataflow_slice_valid_63;
  wire _dataflow_slice_valid_67;
  wire _dataflow_slice_valid_70;
  wire _dataflow_slice_valid_73;
  wire _dataflow_slice_valid_76;
  wire _dataflow_slice_valid_80;
  wire _dataflow_slice_valid_83;
  wire _dataflow_slice_valid_86;
  wire _dataflow_slice_valid_89;
  wire _dataflow_slice_valid_9;
  wire _eq_data_277;
  wire _eq_data_281;
  wire _eq_data_284;
  wire _eq_data_287;
  wire _eq_data_291;
  wire _eq_data_294;
  wire _eq_data_297;
  wire _eq_data_301;
  wire _eq_data_304;
  wire _eq_data_307;
  wire _eq_data_311;
  wire _eq_data_314;
  wire _eq_data_317;
  wire _eq_data_321;
  wire _eq_data_324;
  wire _eq_data_327;
  wire _eq_data_331;
  wire _eq_data_334;
  wire _eq_data_337;
  wire _eq_data_341;
  wire _eq_data_344;
  wire _eq_data_347;
  wire _eq_data_351;
  wire _eq_data_354;
  wire _eq_data_357;
  wire _eq_data_361;
  wire _eq_data_364;
  wire _eq_data_367;
  wire _eq_data_371;
  wire _eq_data_374;
  wire _eq_data_377;
  wire _eq_data_381;
  wire _eq_data_384;
  wire _eq_data_387;
  wire _eq_data_391;
  wire _eq_data_394;
  wire _eq_data_397;
  wire _eq_data_401;
  wire _eq_data_404;
  wire _eq_data_407;
  wire _eq_data_411;
  wire _eq_data_414;
  wire _eq_data_417;
  wire _eq_data_421;
  wire _eq_data_424;
  wire _eq_data_427;
  wire _eq_data_431;
  wire _eq_data_434;
  wire _eq_data_437;
  wire _eq_data_441;
  wire _eq_data_444;
  wire _eq_data_447;
  wire _eq_data_451;
  wire _eq_data_454;
  wire _eq_data_851;
  wire _eq_data_855;
  wire _eq_data_891;
  wire _eq_data_894;
  wire _greatereq_data_51;
  wire _greaterthan_data_108;
  wire _greaterthan_data_125;
  wire _greaterthan_data_142;
  wire _greaterthan_data_159;
  wire _greaterthan_data_176;
  wire _greaterthan_data_193;
  wire _greaterthan_data_3;
  wire _greaterthan_data_43;
  wire _greaterthan_data_57;
  wire _greaterthan_data_74;
  wire _greaterthan_data_773;
  wire _greaterthan_data_888;
  wire _greaterthan_data_91;
  wire _lessthan_data_47;
  wire _maxi_cond_0_1;
  wire _maxi_cond_1_1;
  wire _maxi_cond_2_1;
  wire _maxi_cond_3_1;
  wire _maxi_cond_4_1;
  wire [31:0] _maxi_global_base_addr;
  wire [31:0] _maxi_ram_w4_l8192_id0_1_read_global_addr;
  wire [31:0] _maxi_ram_w4_l8192_id0_1_read_local_addr;
  wire [31:0] _maxi_ram_w4_l8192_id0_1_read_local_stride;
  wire [7:0] _maxi_ram_w4_l8192_id0_1_read_op_sel;
  wire [32:0] _maxi_ram_w4_l8192_id0_1_read_size;
  wire _maxi_ram_w4_l8192_id0_1_read_start;
  wire [31:0] _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_global_addr;
  wire [31:0] _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_addr;
  wire [31:0] _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_stride;
  wire [7:0] _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_op_sel;
  wire [32:0] _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_size;
  wire _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id0_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id0_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id0_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id0_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id0_1_read_size;
  wire _maxi_ram_w8_l2048_id0_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id0_1_write_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id0_1_write_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id0_1_write_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id0_1_write_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id0_1_write_size;
  wire _maxi_ram_w8_l2048_id0_1_write_start;
  wire [31:0] _maxi_ram_w8_l2048_id11_1_write_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id11_1_write_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id11_1_write_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id11_1_write_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id11_1_write_size;
  wire _maxi_ram_w8_l2048_id11_1_write_start;
  wire [31:0] _maxi_ram_w8_l2048_id1_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id1_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id1_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id1_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id1_1_read_size;
  wire _maxi_ram_w8_l2048_id1_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id1_1_write_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id1_1_write_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id1_1_write_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id1_1_write_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id1_1_write_size;
  wire _maxi_ram_w8_l2048_id1_1_write_start;
  wire [31:0] _maxi_ram_w8_l2048_id2_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id2_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id2_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id2_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id2_1_read_size;
  wire _maxi_ram_w8_l2048_id2_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_size;
  wire _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id3_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id3_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id3_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id3_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id3_1_read_size;
  wire _maxi_ram_w8_l2048_id3_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_size;
  wire _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start;
  wire [31:0] _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_global_addr;
  wire [31:0] _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_addr;
  wire [31:0] _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_stride;
  wire [7:0] _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_op_sel;
  wire [32:0] _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_size;
  wire _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start;
  wire [31:0] _maxi_read_cur_global_addr;
  wire [32:0] _maxi_read_cur_size;
  wire [31:0] _maxi_read_fsm;
  wire [31:0] _maxi_read_global_addr;
  wire _maxi_read_idle;
  wire [31:0] _maxi_read_local_addr;
  wire [31:0] _maxi_read_local_stride;
  wire [7:0] _maxi_read_op_sel;
  wire [32:0] _maxi_read_rest_size;
  wire [32:0] _maxi_read_size;
  wire _maxi_read_start;
  wire [31:0] _maxi_write_cur_global_addr;
  wire [32:0] _maxi_write_cur_size;
  wire _maxi_write_data_done;
  wire [31:0] _maxi_write_fsm;
  wire [31:0] _maxi_write_global_addr;
  wire _maxi_write_idle;
  wire [31:0] _maxi_write_local_addr;
  wire [31:0] _maxi_write_local_stride;
  wire [7:0] _maxi_write_op_sel;
  wire [32:0] _maxi_write_rest_size;
  wire [32:0] _maxi_write_size;
  wire _maxi_write_start;
  wire [3:0] _minus_data_110;
  wire [3:0] _minus_data_127;
  wire [3:0] _minus_data_144;
  wire [3:0] _minus_data_161;
  wire [3:0] _minus_data_178;
  wire [3:0] _minus_data_195;
  wire [5:0] _minus_data_5;
  wire [3:0] _minus_data_59;
  wire [3:0] _minus_data_76;
  wire [3:0] _minus_data_93;
  wire [31:0] _mul_10_fsm;
  wire _mul_10_rshift_idle;
  wire _mul_10_rshift_source_ram_rvalid;
  wire _mul_10_x_idle;
  wire _mul_10_x_source_ram_rvalid;
  wire _mul_10_y_idle;
  wire _mul_10_y_source_ram_rvalid;
  wire _mul_10_z_sink_wenable;
  wire [31:0] _mul_11_fsm;
  wire _mul_11_rshift_idle;
  wire _mul_11_rshift_source_ram_rvalid;
  wire _mul_11_x_idle;
  wire _mul_11_x_source_ram_rvalid;
  wire _mul_11_y_idle;
  wire _mul_11_y_source_ram_rvalid;
  wire _mul_11_z_sink_wenable;
  wire [31:0] _mul_12_fsm;
  wire _mul_12_rshift_idle;
  wire _mul_12_rshift_source_ram_rvalid;
  wire _mul_12_x_idle;
  wire _mul_12_x_source_ram_rvalid;
  wire _mul_12_y_idle;
  wire _mul_12_y_source_ram_rvalid;
  wire _mul_12_z_sink_wenable;
  wire [31:0] _mul_4_fsm;
  wire _mul_4_rshift_idle;
  wire _mul_4_rshift_source_ram_rvalid;
  wire _mul_4_x_idle;
  wire _mul_4_x_source_ram_rvalid;
  wire _mul_4_y_idle;
  wire _mul_4_y_source_ram_rvalid;
  wire _mul_4_z_sink_wenable;
  wire [31:0] _mul_5_fsm;
  wire _mul_5_rshift_idle;
  wire _mul_5_rshift_source_ram_rvalid;
  wire _mul_5_x_idle;
  wire _mul_5_x_source_ram_rvalid;
  wire _mul_5_y_idle;
  wire _mul_5_y_source_ram_rvalid;
  wire _mul_5_z_sink_wenable;
  wire [31:0] _mul_6_fsm;
  wire _mul_6_rshift_idle;
  wire _mul_6_rshift_source_ram_rvalid;
  wire _mul_6_x_idle;
  wire _mul_6_x_source_ram_rvalid;
  wire _mul_6_y_idle;
  wire _mul_6_y_source_ram_rvalid;
  wire _mul_6_z_sink_wenable;
  wire [31:0] _mul_7_fsm;
  wire _mul_7_rshift_idle;
  wire _mul_7_rshift_source_ram_rvalid;
  wire _mul_7_x_idle;
  wire _mul_7_x_source_ram_rvalid;
  wire _mul_7_y_idle;
  wire _mul_7_y_source_ram_rvalid;
  wire _mul_7_z_sink_wenable;
  wire [31:0] _mul_8_fsm;
  wire _mul_8_rshift_idle;
  wire _mul_8_rshift_source_ram_rvalid;
  wire _mul_8_x_idle;
  wire _mul_8_x_source_ram_rvalid;
  wire _mul_8_y_idle;
  wire _mul_8_y_source_ram_rvalid;
  wire _mul_8_z_sink_wenable;
  wire [31:0] _mul_9_fsm;
  wire _mul_9_rshift_idle;
  wire _mul_9_rshift_source_ram_rvalid;
  wire _mul_9_x_idle;
  wire _mul_9_x_source_ram_rvalid;
  wire _mul_9_y_idle;
  wire _mul_9_y_source_ram_rvalid;
  wire _mul_9_z_sink_wenable;
  wire [31:0] _mul_rshift_clip_3_fsm;
  wire _mul_rshift_clip_3_rshift_idle;
  wire _mul_rshift_clip_3_rshift_source_ram_rvalid;
  wire _mul_rshift_clip_3_x_idle;
  wire _mul_rshift_clip_3_x_source_ram_rvalid;
  wire _mul_rshift_clip_3_y_idle;
  wire _mul_rshift_clip_3_y_source_ram_rvalid;
  wire _mul_rshift_clip_3_z_sink_wenable;
  wire [31:0] _plus_data_20;
  wire [7:0] _plus_data_607;
  wire [7:0] _plus_data_624;
  wire [7:0] _plus_data_641;
  wire [7:0] _plus_data_658;
  wire [7:0] _plus_data_675;
  wire [7:0] _plus_data_692;
  wire [7:0] _plus_data_709;
  wire [7:0] _plus_data_726;
  wire [7:0] _plus_data_743;
  wire [7:0] _plus_data_759;
  wire [31:0] _plus_data_762;
  wire [7:0] _plus_data_770;
  wire [7:0] _plus_data_875;
  wire [7:0] _plus_data_880;
  wire [31:0] _plus_data_883;
  wire [7:0] _plus_data_885;
  wire _pointer_data_556;
  wire _pointer_data_558;
  wire _pointer_data_560;
  wire _pointer_data_562;
  wire _pointer_data_564;
  wire _pointer_data_566;
  wire _pointer_data_568;
  wire _pointer_data_570;
  wire _pointer_data_572;
  wire _pointer_data_784;
  wire _pointer_data_870;
  wire [32:0] _pulse_count_19;
  wire [8:0] _pulse_count_213;
  wire _pulse_data_19;
  wire _pulse_data_213;
  wire _ram_w4_l8192_id0_0_cond_0_1;
  wire _ram_w4_l8192_id0_0_cond_1_1;
  wire _ram_w4_l8192_id0_0_cond_2_1;
  wire _ram_w4_l8192_id0_0_cond_3_1;
  wire _ram_w4_l8192_id0_0_cond_4_1;
  wire _ram_w4_l8192_id0_0_cond_5_1;
  wire _ram_w4_l8192_id0_0_cond_6_1;
  wire _ram_w4_l8192_id0_1_cond_0_1;
  wire _ram_w4_l8192_id0_1_cond_1_1;
  wire _ram_w4_l8192_id0_1_cond_2_1;
  wire _ram_w4_l8192_id0_1_cond_3_1;
  wire _ram_w4_l8192_id0_1_cond_4_1;
  wire _ram_w4_l8192_id0_1_cond_5_1;
  wire _ram_w4_l8192_id0_1_cond_6_1;
  wire _ram_w4_l8192_id0_2_cond_0_1;
  wire _ram_w4_l8192_id0_2_cond_1_1;
  wire _ram_w4_l8192_id0_2_cond_2_1;
  wire _ram_w4_l8192_id0_2_cond_3_1;
  wire _ram_w4_l8192_id0_2_cond_4_1;
  wire _ram_w4_l8192_id0_2_cond_5_1;
  wire _ram_w4_l8192_id0_2_cond_6_1;
  wire _ram_w4_l8192_id0_3_cond_0_1;
  wire _ram_w4_l8192_id0_3_cond_1_1;
  wire _ram_w4_l8192_id0_3_cond_2_1;
  wire _ram_w4_l8192_id0_3_cond_3_1;
  wire _ram_w4_l8192_id0_3_cond_4_1;
  wire _ram_w4_l8192_id0_3_cond_5_1;
  wire _ram_w4_l8192_id0_3_cond_6_1;
  wire _ram_w4_l8192_id0_4_cond_0_1;
  wire _ram_w4_l8192_id0_4_cond_1_1;
  wire _ram_w4_l8192_id0_4_cond_2_1;
  wire _ram_w4_l8192_id0_4_cond_3_1;
  wire _ram_w4_l8192_id0_4_cond_4_1;
  wire _ram_w4_l8192_id0_4_cond_5_1;
  wire _ram_w4_l8192_id0_4_cond_6_1;
  wire _ram_w4_l8192_id0_5_cond_0_1;
  wire _ram_w4_l8192_id0_5_cond_1_1;
  wire _ram_w4_l8192_id0_5_cond_2_1;
  wire _ram_w4_l8192_id0_5_cond_3_1;
  wire _ram_w4_l8192_id0_5_cond_4_1;
  wire _ram_w4_l8192_id0_5_cond_5_1;
  wire _ram_w4_l8192_id0_5_cond_6_1;
  wire _ram_w4_l8192_id0_6_cond_0_1;
  wire _ram_w4_l8192_id0_6_cond_1_1;
  wire _ram_w4_l8192_id0_6_cond_2_1;
  wire _ram_w4_l8192_id0_6_cond_3_1;
  wire _ram_w4_l8192_id0_6_cond_4_1;
  wire _ram_w4_l8192_id0_6_cond_5_1;
  wire _ram_w4_l8192_id0_6_cond_6_1;
  wire _ram_w4_l8192_id0_7_cond_0_1;
  wire _ram_w4_l8192_id0_7_cond_1_1;
  wire _ram_w4_l8192_id0_7_cond_2_1;
  wire _ram_w4_l8192_id0_7_cond_3_1;
  wire _ram_w4_l8192_id0_7_cond_4_1;
  wire _ram_w4_l8192_id0_7_cond_5_1;
  wire _ram_w4_l8192_id0_7_cond_6_1;
  wire _ram_w4_l8192_id1_0_cond_0_1;
  wire _ram_w4_l8192_id1_0_cond_1_1;
  wire _ram_w4_l8192_id1_0_cond_2_1;
  wire _ram_w4_l8192_id1_1_cond_0_1;
  wire _ram_w4_l8192_id1_1_cond_1_1;
  wire _ram_w4_l8192_id1_1_cond_2_1;
  wire _ram_w4_l8192_id1_2_cond_0_1;
  wire _ram_w4_l8192_id1_2_cond_1_1;
  wire _ram_w4_l8192_id1_2_cond_2_1;
  wire _ram_w4_l8192_id1_3_cond_0_1;
  wire _ram_w4_l8192_id1_3_cond_1_1;
  wire _ram_w4_l8192_id1_3_cond_2_1;
  wire _ram_w4_l8192_id1_4_cond_0_1;
  wire _ram_w4_l8192_id1_4_cond_1_1;
  wire _ram_w4_l8192_id1_4_cond_2_1;
  wire _ram_w4_l8192_id1_5_cond_0_1;
  wire _ram_w4_l8192_id1_5_cond_1_1;
  wire _ram_w4_l8192_id1_5_cond_2_1;
  wire _ram_w4_l8192_id1_6_cond_0_1;
  wire _ram_w4_l8192_id1_6_cond_1_1;
  wire _ram_w4_l8192_id1_6_cond_2_1;
  wire _ram_w4_l8192_id1_7_cond_0_1;
  wire _ram_w4_l8192_id1_7_cond_1_1;
  wire _ram_w4_l8192_id1_7_cond_2_1;
  wire _ram_w4_l8192_id2_0_cond_0_1;
  wire _ram_w4_l8192_id2_0_cond_1_1;
  wire _ram_w4_l8192_id2_0_cond_2_1;
  wire _ram_w4_l8192_id2_1_cond_0_1;
  wire _ram_w4_l8192_id2_1_cond_1_1;
  wire _ram_w4_l8192_id2_1_cond_2_1;
  wire _ram_w4_l8192_id2_2_cond_0_1;
  wire _ram_w4_l8192_id2_2_cond_1_1;
  wire _ram_w4_l8192_id2_2_cond_2_1;
  wire _ram_w4_l8192_id2_3_cond_0_1;
  wire _ram_w4_l8192_id2_3_cond_1_1;
  wire _ram_w4_l8192_id2_3_cond_2_1;
  wire _ram_w4_l8192_id2_4_cond_0_1;
  wire _ram_w4_l8192_id2_4_cond_1_1;
  wire _ram_w4_l8192_id2_4_cond_2_1;
  wire _ram_w4_l8192_id2_5_cond_0_1;
  wire _ram_w4_l8192_id2_5_cond_1_1;
  wire _ram_w4_l8192_id2_5_cond_2_1;
  wire _ram_w4_l8192_id2_6_cond_0_1;
  wire _ram_w4_l8192_id2_6_cond_1_1;
  wire _ram_w4_l8192_id2_6_cond_2_1;
  wire _ram_w4_l8192_id2_7_cond_0_1;
  wire _ram_w4_l8192_id2_7_cond_1_1;
  wire _ram_w4_l8192_id2_7_cond_2_1;
  wire _ram_w4_l8192_id3_0_cond_0_1;
  wire _ram_w4_l8192_id3_0_cond_1_1;
  wire _ram_w4_l8192_id3_0_cond_2_1;
  wire _ram_w4_l8192_id3_1_cond_0_1;
  wire _ram_w4_l8192_id3_1_cond_1_1;
  wire _ram_w4_l8192_id3_1_cond_2_1;
  wire _ram_w4_l8192_id3_2_cond_0_1;
  wire _ram_w4_l8192_id3_2_cond_1_1;
  wire _ram_w4_l8192_id3_2_cond_2_1;
  wire _ram_w4_l8192_id3_3_cond_0_1;
  wire _ram_w4_l8192_id3_3_cond_1_1;
  wire _ram_w4_l8192_id3_3_cond_2_1;
  wire _ram_w4_l8192_id3_4_cond_0_1;
  wire _ram_w4_l8192_id3_4_cond_1_1;
  wire _ram_w4_l8192_id3_4_cond_2_1;
  wire _ram_w4_l8192_id3_5_cond_0_1;
  wire _ram_w4_l8192_id3_5_cond_1_1;
  wire _ram_w4_l8192_id3_5_cond_2_1;
  wire _ram_w4_l8192_id3_6_cond_0_1;
  wire _ram_w4_l8192_id3_6_cond_1_1;
  wire _ram_w4_l8192_id3_6_cond_2_1;
  wire _ram_w4_l8192_id3_7_cond_0_1;
  wire _ram_w4_l8192_id3_7_cond_1_1;
  wire _ram_w4_l8192_id3_7_cond_2_1;
  wire _ram_w4_l8192_id4_0_cond_0_1;
  wire _ram_w4_l8192_id4_0_cond_1_1;
  wire _ram_w4_l8192_id4_0_cond_2_1;
  wire _ram_w4_l8192_id4_1_cond_0_1;
  wire _ram_w4_l8192_id4_1_cond_1_1;
  wire _ram_w4_l8192_id4_1_cond_2_1;
  wire _ram_w4_l8192_id4_2_cond_0_1;
  wire _ram_w4_l8192_id4_2_cond_1_1;
  wire _ram_w4_l8192_id4_2_cond_2_1;
  wire _ram_w4_l8192_id4_3_cond_0_1;
  wire _ram_w4_l8192_id4_3_cond_1_1;
  wire _ram_w4_l8192_id4_3_cond_2_1;
  wire _ram_w4_l8192_id4_4_cond_0_1;
  wire _ram_w4_l8192_id4_4_cond_1_1;
  wire _ram_w4_l8192_id4_4_cond_2_1;
  wire _ram_w4_l8192_id4_5_cond_0_1;
  wire _ram_w4_l8192_id4_5_cond_1_1;
  wire _ram_w4_l8192_id4_5_cond_2_1;
  wire _ram_w4_l8192_id4_6_cond_0_1;
  wire _ram_w4_l8192_id4_6_cond_1_1;
  wire _ram_w4_l8192_id4_6_cond_2_1;
  wire _ram_w4_l8192_id4_7_cond_0_1;
  wire _ram_w4_l8192_id4_7_cond_1_1;
  wire _ram_w4_l8192_id4_7_cond_2_1;
  wire _ram_w4_l8192_id5_0_cond_0_1;
  wire _ram_w4_l8192_id5_0_cond_1_1;
  wire _ram_w4_l8192_id5_0_cond_2_1;
  wire _ram_w4_l8192_id5_1_cond_0_1;
  wire _ram_w4_l8192_id5_1_cond_1_1;
  wire _ram_w4_l8192_id5_1_cond_2_1;
  wire _ram_w4_l8192_id5_2_cond_0_1;
  wire _ram_w4_l8192_id5_2_cond_1_1;
  wire _ram_w4_l8192_id5_2_cond_2_1;
  wire _ram_w4_l8192_id5_3_cond_0_1;
  wire _ram_w4_l8192_id5_3_cond_1_1;
  wire _ram_w4_l8192_id5_3_cond_2_1;
  wire _ram_w4_l8192_id5_4_cond_0_1;
  wire _ram_w4_l8192_id5_4_cond_1_1;
  wire _ram_w4_l8192_id5_4_cond_2_1;
  wire _ram_w4_l8192_id5_5_cond_0_1;
  wire _ram_w4_l8192_id5_5_cond_1_1;
  wire _ram_w4_l8192_id5_5_cond_2_1;
  wire _ram_w4_l8192_id5_6_cond_0_1;
  wire _ram_w4_l8192_id5_6_cond_1_1;
  wire _ram_w4_l8192_id5_6_cond_2_1;
  wire _ram_w4_l8192_id5_7_cond_0_1;
  wire _ram_w4_l8192_id5_7_cond_1_1;
  wire _ram_w4_l8192_id5_7_cond_2_1;
  wire _ram_w4_l8192_id6_0_cond_0_1;
  wire _ram_w4_l8192_id6_0_cond_1_1;
  wire _ram_w4_l8192_id6_0_cond_2_1;
  wire _ram_w4_l8192_id6_1_cond_0_1;
  wire _ram_w4_l8192_id6_1_cond_1_1;
  wire _ram_w4_l8192_id6_1_cond_2_1;
  wire _ram_w4_l8192_id6_2_cond_0_1;
  wire _ram_w4_l8192_id6_2_cond_1_1;
  wire _ram_w4_l8192_id6_2_cond_2_1;
  wire _ram_w4_l8192_id6_3_cond_0_1;
  wire _ram_w4_l8192_id6_3_cond_1_1;
  wire _ram_w4_l8192_id6_3_cond_2_1;
  wire _ram_w4_l8192_id6_4_cond_0_1;
  wire _ram_w4_l8192_id6_4_cond_1_1;
  wire _ram_w4_l8192_id6_4_cond_2_1;
  wire _ram_w4_l8192_id6_5_cond_0_1;
  wire _ram_w4_l8192_id6_5_cond_1_1;
  wire _ram_w4_l8192_id6_5_cond_2_1;
  wire _ram_w4_l8192_id6_6_cond_0_1;
  wire _ram_w4_l8192_id6_6_cond_1_1;
  wire _ram_w4_l8192_id6_6_cond_2_1;
  wire _ram_w4_l8192_id6_7_cond_0_1;
  wire _ram_w4_l8192_id6_7_cond_1_1;
  wire _ram_w4_l8192_id6_7_cond_2_1;
  wire _ram_w4_l8192_id7_0_cond_0_1;
  wire _ram_w4_l8192_id7_0_cond_1_1;
  wire _ram_w4_l8192_id7_0_cond_2_1;
  wire _ram_w4_l8192_id7_1_cond_0_1;
  wire _ram_w4_l8192_id7_1_cond_1_1;
  wire _ram_w4_l8192_id7_1_cond_2_1;
  wire _ram_w4_l8192_id7_2_cond_0_1;
  wire _ram_w4_l8192_id7_2_cond_1_1;
  wire _ram_w4_l8192_id7_2_cond_2_1;
  wire _ram_w4_l8192_id7_3_cond_0_1;
  wire _ram_w4_l8192_id7_3_cond_1_1;
  wire _ram_w4_l8192_id7_3_cond_2_1;
  wire _ram_w4_l8192_id7_4_cond_0_1;
  wire _ram_w4_l8192_id7_4_cond_1_1;
  wire _ram_w4_l8192_id7_4_cond_2_1;
  wire _ram_w4_l8192_id7_5_cond_0_1;
  wire _ram_w4_l8192_id7_5_cond_1_1;
  wire _ram_w4_l8192_id7_5_cond_2_1;
  wire _ram_w4_l8192_id7_6_cond_0_1;
  wire _ram_w4_l8192_id7_6_cond_1_1;
  wire _ram_w4_l8192_id7_6_cond_2_1;
  wire _ram_w4_l8192_id7_7_cond_0_1;
  wire _ram_w4_l8192_id7_7_cond_1_1;
  wire _ram_w4_l8192_id7_7_cond_2_1;
  wire _ram_w4_l8192_id8_0_cond_0_1;
  wire _ram_w4_l8192_id8_0_cond_1_1;
  wire _ram_w4_l8192_id8_0_cond_2_1;
  wire _ram_w4_l8192_id8_1_cond_0_1;
  wire _ram_w4_l8192_id8_1_cond_1_1;
  wire _ram_w4_l8192_id8_1_cond_2_1;
  wire _ram_w4_l8192_id8_2_cond_0_1;
  wire _ram_w4_l8192_id8_2_cond_1_1;
  wire _ram_w4_l8192_id8_2_cond_2_1;
  wire _ram_w4_l8192_id8_3_cond_0_1;
  wire _ram_w4_l8192_id8_3_cond_1_1;
  wire _ram_w4_l8192_id8_3_cond_2_1;
  wire _ram_w4_l8192_id8_4_cond_0_1;
  wire _ram_w4_l8192_id8_4_cond_1_1;
  wire _ram_w4_l8192_id8_4_cond_2_1;
  wire _ram_w4_l8192_id8_5_cond_0_1;
  wire _ram_w4_l8192_id8_5_cond_1_1;
  wire _ram_w4_l8192_id8_5_cond_2_1;
  wire _ram_w4_l8192_id8_6_cond_0_1;
  wire _ram_w4_l8192_id8_6_cond_1_1;
  wire _ram_w4_l8192_id8_6_cond_2_1;
  wire _ram_w4_l8192_id8_7_cond_0_1;
  wire _ram_w4_l8192_id8_7_cond_1_1;
  wire _ram_w4_l8192_id8_7_cond_2_1;
  wire _ram_w8_l2048_id0_0_cond_0_1;
  wire _ram_w8_l2048_id0_0_cond_1_1;
  wire _ram_w8_l2048_id0_0_cond_2_1;
  wire _ram_w8_l2048_id0_0_cond_3_1;
  wire _ram_w8_l2048_id0_0_cond_4_1;
  wire _ram_w8_l2048_id0_0_cond_5_1;
  wire _ram_w8_l2048_id0_1_cond_0_1;
  wire _ram_w8_l2048_id0_1_cond_1_1;
  wire _ram_w8_l2048_id0_1_cond_2_1;
  wire _ram_w8_l2048_id0_1_cond_3_1;
  wire _ram_w8_l2048_id0_1_cond_4_1;
  wire _ram_w8_l2048_id0_1_cond_5_1;
  wire _ram_w8_l2048_id0_2_cond_0_1;
  wire _ram_w8_l2048_id0_2_cond_1_1;
  wire _ram_w8_l2048_id0_2_cond_2_1;
  wire _ram_w8_l2048_id0_2_cond_3_1;
  wire _ram_w8_l2048_id0_2_cond_4_1;
  wire _ram_w8_l2048_id0_2_cond_5_1;
  wire _ram_w8_l2048_id0_3_cond_0_1;
  wire _ram_w8_l2048_id0_3_cond_1_1;
  wire _ram_w8_l2048_id0_3_cond_2_1;
  wire _ram_w8_l2048_id0_3_cond_3_1;
  wire _ram_w8_l2048_id0_3_cond_4_1;
  wire _ram_w8_l2048_id0_3_cond_5_1;
  wire _ram_w8_l2048_id10_0_cond_0_1;
  wire _ram_w8_l2048_id10_0_cond_1_1;
  wire _ram_w8_l2048_id10_0_cond_2_1;
  wire _ram_w8_l2048_id10_1_cond_0_1;
  wire _ram_w8_l2048_id10_1_cond_1_1;
  wire _ram_w8_l2048_id10_1_cond_2_1;
  wire _ram_w8_l2048_id10_2_cond_0_1;
  wire _ram_w8_l2048_id10_2_cond_1_1;
  wire _ram_w8_l2048_id10_2_cond_2_1;
  wire _ram_w8_l2048_id10_3_cond_0_1;
  wire _ram_w8_l2048_id10_3_cond_1_1;
  wire _ram_w8_l2048_id10_3_cond_2_1;
  wire _ram_w8_l2048_id11_0_cond_0_1;
  wire _ram_w8_l2048_id11_1_cond_0_1;
  wire _ram_w8_l2048_id11_2_cond_0_1;
  wire _ram_w8_l2048_id11_3_cond_0_1;
  wire _ram_w8_l2048_id1_0_cond_0_1;
  wire _ram_w8_l2048_id1_0_cond_1_1;
  wire _ram_w8_l2048_id1_0_cond_2_1;
  wire _ram_w8_l2048_id1_0_cond_3_1;
  wire _ram_w8_l2048_id1_0_cond_4_1;
  wire _ram_w8_l2048_id1_0_cond_5_1;
  wire _ram_w8_l2048_id1_1_cond_0_1;
  wire _ram_w8_l2048_id1_1_cond_1_1;
  wire _ram_w8_l2048_id1_1_cond_2_1;
  wire _ram_w8_l2048_id1_1_cond_3_1;
  wire _ram_w8_l2048_id1_1_cond_4_1;
  wire _ram_w8_l2048_id1_1_cond_5_1;
  wire _ram_w8_l2048_id1_2_cond_0_1;
  wire _ram_w8_l2048_id1_2_cond_1_1;
  wire _ram_w8_l2048_id1_2_cond_2_1;
  wire _ram_w8_l2048_id1_2_cond_3_1;
  wire _ram_w8_l2048_id1_2_cond_4_1;
  wire _ram_w8_l2048_id1_2_cond_5_1;
  wire _ram_w8_l2048_id1_3_cond_0_1;
  wire _ram_w8_l2048_id1_3_cond_1_1;
  wire _ram_w8_l2048_id1_3_cond_2_1;
  wire _ram_w8_l2048_id1_3_cond_3_1;
  wire _ram_w8_l2048_id1_3_cond_4_1;
  wire _ram_w8_l2048_id1_3_cond_5_1;
  wire _ram_w8_l2048_id2_0_cond_0_1;
  wire _ram_w8_l2048_id2_0_cond_1_1;
  wire _ram_w8_l2048_id2_0_cond_2_1;
  wire _ram_w8_l2048_id2_0_cond_3_1;
  wire _ram_w8_l2048_id2_0_cond_4_1;
  wire _ram_w8_l2048_id2_0_cond_5_1;
  wire _ram_w8_l2048_id2_0_cond_6_1;
  wire _ram_w8_l2048_id2_1_cond_0_1;
  wire _ram_w8_l2048_id2_1_cond_1_1;
  wire _ram_w8_l2048_id2_1_cond_2_1;
  wire _ram_w8_l2048_id2_1_cond_3_1;
  wire _ram_w8_l2048_id2_1_cond_4_1;
  wire _ram_w8_l2048_id2_1_cond_5_1;
  wire _ram_w8_l2048_id2_1_cond_6_1;
  wire _ram_w8_l2048_id2_2_cond_0_1;
  wire _ram_w8_l2048_id2_2_cond_1_1;
  wire _ram_w8_l2048_id2_2_cond_2_1;
  wire _ram_w8_l2048_id2_2_cond_3_1;
  wire _ram_w8_l2048_id2_2_cond_4_1;
  wire _ram_w8_l2048_id2_2_cond_5_1;
  wire _ram_w8_l2048_id2_2_cond_6_1;
  wire _ram_w8_l2048_id2_3_cond_0_1;
  wire _ram_w8_l2048_id2_3_cond_1_1;
  wire _ram_w8_l2048_id2_3_cond_2_1;
  wire _ram_w8_l2048_id2_3_cond_3_1;
  wire _ram_w8_l2048_id2_3_cond_4_1;
  wire _ram_w8_l2048_id2_3_cond_5_1;
  wire _ram_w8_l2048_id2_3_cond_6_1;
  wire _ram_w8_l2048_id3_0_cond_0_1;
  wire _ram_w8_l2048_id3_0_cond_1_1;
  wire _ram_w8_l2048_id3_0_cond_2_1;
  wire _ram_w8_l2048_id3_0_cond_3_1;
  wire _ram_w8_l2048_id3_0_cond_4_1;
  wire _ram_w8_l2048_id3_0_cond_5_1;
  wire _ram_w8_l2048_id3_1_cond_0_1;
  wire _ram_w8_l2048_id3_1_cond_1_1;
  wire _ram_w8_l2048_id3_1_cond_2_1;
  wire _ram_w8_l2048_id3_1_cond_3_1;
  wire _ram_w8_l2048_id3_1_cond_4_1;
  wire _ram_w8_l2048_id3_1_cond_5_1;
  wire _ram_w8_l2048_id3_2_cond_0_1;
  wire _ram_w8_l2048_id3_2_cond_1_1;
  wire _ram_w8_l2048_id3_2_cond_2_1;
  wire _ram_w8_l2048_id3_2_cond_3_1;
  wire _ram_w8_l2048_id3_2_cond_4_1;
  wire _ram_w8_l2048_id3_2_cond_5_1;
  wire _ram_w8_l2048_id3_3_cond_0_1;
  wire _ram_w8_l2048_id3_3_cond_1_1;
  wire _ram_w8_l2048_id3_3_cond_2_1;
  wire _ram_w8_l2048_id3_3_cond_3_1;
  wire _ram_w8_l2048_id3_3_cond_4_1;
  wire _ram_w8_l2048_id3_3_cond_5_1;
  wire _ram_w8_l2048_id4_0_cond_0_1;
  wire _ram_w8_l2048_id4_0_cond_1_1;
  wire _ram_w8_l2048_id4_0_cond_2_1;
  wire _ram_w8_l2048_id4_1_cond_0_1;
  wire _ram_w8_l2048_id4_1_cond_1_1;
  wire _ram_w8_l2048_id4_1_cond_2_1;
  wire _ram_w8_l2048_id4_2_cond_0_1;
  wire _ram_w8_l2048_id4_2_cond_1_1;
  wire _ram_w8_l2048_id4_2_cond_2_1;
  wire _ram_w8_l2048_id4_3_cond_0_1;
  wire _ram_w8_l2048_id4_3_cond_1_1;
  wire _ram_w8_l2048_id4_3_cond_2_1;
  wire _ram_w8_l2048_id5_0_cond_0_1;
  wire _ram_w8_l2048_id5_0_cond_1_1;
  wire _ram_w8_l2048_id5_0_cond_2_1;
  wire _ram_w8_l2048_id5_0_cond_3_1;
  wire _ram_w8_l2048_id5_1_cond_0_1;
  wire _ram_w8_l2048_id5_1_cond_1_1;
  wire _ram_w8_l2048_id5_1_cond_2_1;
  wire _ram_w8_l2048_id5_1_cond_3_1;
  wire _ram_w8_l2048_id5_2_cond_0_1;
  wire _ram_w8_l2048_id5_2_cond_1_1;
  wire _ram_w8_l2048_id5_2_cond_2_1;
  wire _ram_w8_l2048_id5_2_cond_3_1;
  wire _ram_w8_l2048_id5_3_cond_0_1;
  wire _ram_w8_l2048_id5_3_cond_1_1;
  wire _ram_w8_l2048_id5_3_cond_2_1;
  wire _ram_w8_l2048_id5_3_cond_3_1;
  wire _ram_w8_l2048_id6_0_cond_0_1;
  wire _ram_w8_l2048_id6_0_cond_1_1;
  wire _ram_w8_l2048_id6_0_cond_2_1;
  wire _ram_w8_l2048_id6_1_cond_0_1;
  wire _ram_w8_l2048_id6_1_cond_1_1;
  wire _ram_w8_l2048_id6_1_cond_2_1;
  wire _ram_w8_l2048_id6_2_cond_0_1;
  wire _ram_w8_l2048_id6_2_cond_1_1;
  wire _ram_w8_l2048_id6_2_cond_2_1;
  wire _ram_w8_l2048_id6_3_cond_0_1;
  wire _ram_w8_l2048_id6_3_cond_1_1;
  wire _ram_w8_l2048_id6_3_cond_2_1;
  wire _ram_w8_l2048_id7_0_cond_0_1;
  wire _ram_w8_l2048_id7_0_cond_1_1;
  wire _ram_w8_l2048_id7_0_cond_2_1;
  wire _ram_w8_l2048_id7_1_cond_0_1;
  wire _ram_w8_l2048_id7_1_cond_1_1;
  wire _ram_w8_l2048_id7_1_cond_2_1;
  wire _ram_w8_l2048_id7_2_cond_0_1;
  wire _ram_w8_l2048_id7_2_cond_1_1;
  wire _ram_w8_l2048_id7_2_cond_2_1;
  wire _ram_w8_l2048_id7_3_cond_0_1;
  wire _ram_w8_l2048_id7_3_cond_1_1;
  wire _ram_w8_l2048_id7_3_cond_2_1;
  wire _ram_w8_l2048_id8_0_cond_0_1;
  wire _ram_w8_l2048_id8_0_cond_1_1;
  wire _ram_w8_l2048_id8_0_cond_2_1;
  wire _ram_w8_l2048_id8_0_cond_3_1;
  wire _ram_w8_l2048_id8_1_cond_0_1;
  wire _ram_w8_l2048_id8_1_cond_1_1;
  wire _ram_w8_l2048_id8_1_cond_2_1;
  wire _ram_w8_l2048_id8_1_cond_3_1;
  wire _ram_w8_l2048_id8_2_cond_0_1;
  wire _ram_w8_l2048_id8_2_cond_1_1;
  wire _ram_w8_l2048_id8_2_cond_2_1;
  wire _ram_w8_l2048_id8_2_cond_3_1;
  wire _ram_w8_l2048_id8_3_cond_0_1;
  wire _ram_w8_l2048_id8_3_cond_1_1;
  wire _ram_w8_l2048_id8_3_cond_2_1;
  wire _ram_w8_l2048_id8_3_cond_3_1;
  wire _ram_w8_l2048_id9_0_cond_0_1;
  wire _ram_w8_l2048_id9_0_cond_1_1;
  wire _ram_w8_l2048_id9_0_cond_2_1;
  wire _ram_w8_l2048_id9_1_cond_0_1;
  wire _ram_w8_l2048_id9_1_cond_1_1;
  wire _ram_w8_l2048_id9_1_cond_2_1;
  wire _ram_w8_l2048_id9_2_cond_0_1;
  wire _ram_w8_l2048_id9_2_cond_1_1;
  wire _ram_w8_l2048_id9_2_cond_2_1;
  wire _ram_w8_l2048_id9_3_cond_0_1;
  wire _ram_w8_l2048_id9_3_cond_1_1;
  wire _ram_w8_l2048_id9_3_cond_2_1;
  wire [7:0] _reduce_max_13_data_data;
  wire [7:0] _reduce_max_13_size_data;
  wire _reduce_max_13_valid_data;
  wire [7:0] _reduce_max_13_x_data;
  wire [32:0] _reduceadd_count_17;
  wire [31:0] _reduceadd_data_17;
  wire [8:0] _reducemax_count_211;
  wire [7:0] _reducemax_data_211;
  wire [7:0] _reinterpretcast_data_234;
  wire [7:0] _reinterpretcast_data_241;
  wire [7:0] _reinterpretcast_data_248;
  wire [7:0] _reinterpretcast_data_255;
  wire [7:0] _reinterpretcast_data_262;
  wire [7:0] _reinterpretcast_data_493;
  wire [7:0] _reinterpretcast_data_494;
  wire [7:0] _reinterpretcast_data_495;
  wire [7:0] _reinterpretcast_data_496;
  wire [7:0] _reinterpretcast_data_497;
  wire [7:0] _reinterpretcast_data_498;
  wire [7:0] _reinterpretcast_data_499;
  wire [7:0] _reinterpretcast_data_500;
  wire [7:0] _reinterpretcast_data_501;
  wire [3:0] _reinterpretcast_data_547;
  wire [3:0] _reinterpretcast_data_548;
  wire [3:0] _reinterpretcast_data_549;
  wire [3:0] _reinterpretcast_data_550;
  wire [3:0] _reinterpretcast_data_551;
  wire [3:0] _reinterpretcast_data_552;
  wire [3:0] _reinterpretcast_data_553;
  wire [3:0] _reinterpretcast_data_554;
  wire [3:0] _reinterpretcast_data_555;
  wire [7:0] _reinterpretcast_data_776;
  wire [7:0] _reinterpretcast_data_789;
  wire [7:0] _reinterpretcast_data_795;
  wire [7:0] _reinterpretcast_data_816;
  wire [7:0] _reinterpretcast_data_823;
  wire [7:0] _reinterpretcast_data_830;
  wire [7:0] _reinterpretcast_data_837;
  wire [7:0] _reinterpretcast_data_844;
  wire [7:0] _reinterpretcast_data_863;
  wire [3:0] _reinterpretcast_data_869;
  wire [7:0] _reinterpretcast_data_897;
  wire [7:0] _reinterpretcast_src_234;
  wire [7:0] _reinterpretcast_src_241;
  wire [7:0] _reinterpretcast_src_248;
  wire [7:0] _reinterpretcast_src_255;
  wire [7:0] _reinterpretcast_src_262;
  wire [7:0] _reinterpretcast_src_493;
  wire [7:0] _reinterpretcast_src_494;
  wire [7:0] _reinterpretcast_src_495;
  wire [7:0] _reinterpretcast_src_496;
  wire [7:0] _reinterpretcast_src_497;
  wire [7:0] _reinterpretcast_src_498;
  wire [7:0] _reinterpretcast_src_499;
  wire [7:0] _reinterpretcast_src_500;
  wire [7:0] _reinterpretcast_src_501;
  wire [3:0] _reinterpretcast_src_547;
  wire [3:0] _reinterpretcast_src_548;
  wire [3:0] _reinterpretcast_src_549;
  wire [3:0] _reinterpretcast_src_550;
  wire [3:0] _reinterpretcast_src_551;
  wire [3:0] _reinterpretcast_src_552;
  wire [3:0] _reinterpretcast_src_553;
  wire [3:0] _reinterpretcast_src_554;
  wire [3:0] _reinterpretcast_src_555;
  wire [7:0] _reinterpretcast_src_776;
  wire [7:0] _reinterpretcast_src_789;
  wire [7:0] _reinterpretcast_src_795;
  wire [7:0] _reinterpretcast_src_816;
  wire [7:0] _reinterpretcast_src_823;
  wire [7:0] _reinterpretcast_src_830;
  wire [7:0] _reinterpretcast_src_837;
  wire [7:0] _reinterpretcast_src_844;
  wire [7:0] _reinterpretcast_src_863;
  wire [3:0] _reinterpretcast_src_869;
  wire [7:0] _reinterpretcast_src_897;
  wire _rst_logic_1;
  wire _rst_logic_2;
  wire _saxi_cond_0_1;
  wire _saxi_flag_0;
  wire _saxi_flag_1;
  wire _saxi_flag_10;
  wire _saxi_flag_11;
  wire _saxi_flag_12;
  wire _saxi_flag_13;
  wire _saxi_flag_2;
  wire _saxi_flag_3;
  wire _saxi_flag_4;
  wire _saxi_flag_5;
  wire _saxi_flag_6;
  wire _saxi_flag_7;
  wire _saxi_flag_8;
  wire _saxi_flag_9;
  wire [31:0] _saxi_register_0;
  wire [31:0] _saxi_register_1;
  wire [31:0] _saxi_register_10;
  wire [31:0] _saxi_register_11;
  wire [31:0] _saxi_register_12;
  wire [31:0] _saxi_register_13;
  wire [31:0] _saxi_register_2;
  wire [31:0] _saxi_register_3;
  wire [31:0] _saxi_register_4;
  wire [31:0] _saxi_register_5;
  wire [31:0] _saxi_register_6;
  wire [31:0] _saxi_register_7;
  wire [31:0] _saxi_register_8;
  wire [31:0] _saxi_register_9;
  wire [31:0] _saxi_register_fsm;
  wire [31:0] _saxi_resetval_0;
  wire [31:0] _saxi_resetval_1;
  wire [31:0] _saxi_resetval_10;
  wire [31:0] _saxi_resetval_11;
  wire [31:0] _saxi_resetval_12;
  wire [31:0] _saxi_resetval_13;
  wire [31:0] _saxi_resetval_2;
  wire [31:0] _saxi_resetval_3;
  wire [31:0] _saxi_resetval_4;
  wire [31:0] _saxi_resetval_5;
  wire [31:0] _saxi_resetval_6;
  wire [31:0] _saxi_resetval_7;
  wire [31:0] _saxi_resetval_8;
  wire [31:0] _saxi_resetval_9;
  wire _set_flag_1024;
  wire _set_flag_1025;
  wire _set_flag_1026;
  wire _set_flag_1036;
  wire _set_flag_1038;
  wire _set_flag_1163;
  wire _set_flag_1164;
  wire _set_flag_1165;
  wire _set_flag_1166;
  wire _set_flag_1167;
  wire _set_flag_1168;
  wire _set_flag_1169;
  wire _set_flag_1179;
  wire _set_flag_1180;
  wire _set_flag_1190;
  wire _set_flag_1191;
  wire _set_flag_1192;
  wire _set_flag_1193;
  wire _set_flag_1194;
  wire _set_flag_1195;
  wire _set_flag_1196;
  wire _set_flag_1197;
  wire _set_flag_1198;
  wire _set_flag_1199;
  wire _set_flag_1200;
  wire _set_flag_1210;
  wire _set_flag_1224;
  wire _set_flag_457;
  wire _set_flag_458;
  wire _set_flag_459;
  wire _set_flag_460;
  wire _set_flag_461;
  wire _set_flag_462;
  wire _set_flag_463;
  wire _set_flag_473;
  wire _set_flag_474;
  wire _set_flag_484;
  wire _set_flag_485;
  wire _set_flag_486;
  wire _set_flag_487;
  wire _set_flag_488;
  wire _set_flag_489;
  wire _set_flag_490;
  wire _set_flag_491;
  wire _set_flag_492;
  wire _set_flag_493;
  wire _set_flag_494;
  wire _set_flag_504;
  wire _set_flag_514;
  wire _set_flag_524;
  wire _set_flag_534;
  wire _set_flag_544;
  wire _set_flag_554;
  wire _set_flag_564;
  wire _set_flag_574;
  wire _set_flag_584;
  wire _set_flag_598;
  wire _set_flag_612;
  wire _set_flag_626;
  wire _set_flag_640;
  wire _set_flag_654;
  wire _set_flag_668;
  wire _set_flag_682;
  wire _set_flag_696;
  wire _set_flag_710;
  wire [7:0] _slice_data_233;
  wire [7:0] _slice_data_240;
  wire [7:0] _slice_data_247;
  wire [7:0] _slice_data_254;
  wire [7:0] _slice_data_261;
  wire [7:0] _slice_data_815;
  wire [7:0] _slice_data_822;
  wire [7:0] _slice_data_829;
  wire [7:0] _slice_data_836;
  wire [7:0] _slice_data_843;
  wire [17:0] _sll_data_112;
  wire [17:0] _sll_data_129;
  wire [17:0] _sll_data_146;
  wire [17:0] _sll_data_163;
  wire [17:0] _sll_data_180;
  wire [17:0] _sll_data_197;
  wire [17:0] _sll_data_61;
  wire [65:0] _sll_data_7;
  wire [17:0] _sll_data_78;
  wire [17:0] _sll_data_95;
  wire [32:0] _source_stream_conv2d_16_source_19_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_19_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_19_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_19_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_19_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_19_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_19_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_19_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_19_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_19_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_19_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_19_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_19_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_19_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_19_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_19_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_19_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_19_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_19_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_19_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_19_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_19_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_19_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_19_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_20_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_20_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_20_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_20_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_20_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_20_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_20_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_20_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_20_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_20_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_20_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_20_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_20_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_20_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_20_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_20_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_20_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_20_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_20_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_20_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_20_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_20_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_20_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_20_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_21_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_21_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_21_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_21_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_21_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_21_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_21_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_21_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_21_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_21_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_21_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_21_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_21_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_21_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_21_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_21_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_21_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_21_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_21_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_21_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_21_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_21_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_21_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_21_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_22_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_22_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_22_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_22_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_22_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_22_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_22_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_22_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_22_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_22_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_22_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_22_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_22_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_22_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_22_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_22_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_22_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_22_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_22_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_22_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_22_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_22_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_22_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_22_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_23_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_23_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_23_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_23_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_23_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_23_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_23_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_23_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_23_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_23_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_23_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_23_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_23_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_23_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_23_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_23_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_23_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_23_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_23_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_23_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_23_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_23_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_23_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_23_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_24_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_24_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_24_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_24_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_24_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_24_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_24_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_24_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_24_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_24_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_24_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_24_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_24_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_24_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_24_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_24_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_24_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_24_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_24_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_24_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_24_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_24_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_24_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_24_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_25_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_25_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_25_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_25_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_25_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_25_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_25_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_25_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_25_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_25_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_25_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_25_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_25_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_25_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_25_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_25_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_25_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_25_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_25_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_25_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_25_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_25_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_25_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_25_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_26_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_26_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_26_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_26_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_26_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_26_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_26_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_26_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_26_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_26_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_26_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_26_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_26_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_26_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_26_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_26_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_26_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_26_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_26_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_26_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_26_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_26_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_26_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_26_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_27_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_27_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_27_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_27_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_27_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_27_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_27_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_27_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_27_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_27_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_27_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_27_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_27_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_27_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_27_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_27_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_27_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_27_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_27_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_27_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_27_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_27_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_27_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_27_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_28_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_28_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_28_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_28_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_28_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_28_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_28_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_28_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_28_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_28_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_28_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_28_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_28_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_28_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_28_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_28_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_28_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_28_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_28_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_28_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_28_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_28_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_28_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_28_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_29_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_29_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_29_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_29_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_29_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_29_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_29_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_29_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_29_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_29_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_29_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_29_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_29_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_29_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_29_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_29_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_29_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_29_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_29_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_29_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_29_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_29_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_29_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_29_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_30_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_30_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_30_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_30_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_30_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_30_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_30_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_30_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_30_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_30_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_30_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_30_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_30_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_30_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_30_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_30_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_30_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_30_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_30_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_30_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_30_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_30_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_30_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_30_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_31_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_31_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_31_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_31_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_31_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_31_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_31_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_31_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_31_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_31_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_31_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_31_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_31_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_31_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_31_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_31_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_31_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_31_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_31_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_31_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_31_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_31_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_31_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_31_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_32_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_32_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_32_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_32_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_32_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_32_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_32_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_32_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_32_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_32_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_32_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_32_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_32_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_32_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_32_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_32_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_32_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_32_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_32_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_32_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_32_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_32_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_32_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_32_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_33_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_33_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_33_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_33_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_33_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_33_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_33_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_33_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_33_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_33_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_33_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_33_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_33_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_33_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_33_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_33_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_33_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_33_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_33_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_33_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_33_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_33_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_33_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_33_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_34_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_34_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_34_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_34_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_34_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_34_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_34_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_34_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_34_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_34_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_34_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_34_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_34_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_34_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_34_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_34_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_34_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_34_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_34_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_34_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_34_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_34_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_34_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_34_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_35_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_35_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_35_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_35_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_35_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_35_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_35_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_35_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_35_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_35_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_35_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_35_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_35_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_35_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_35_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_35_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_35_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_35_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_35_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_35_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_35_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_35_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_35_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_35_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_36_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_36_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_36_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_36_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_36_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_36_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_36_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_36_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_36_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_36_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_36_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_36_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_36_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_36_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_36_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_36_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_36_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_36_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_36_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_36_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_36_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_36_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_36_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_36_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_6_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_6_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_6_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_6_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_6_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_6_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_6_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_6_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_6_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_6_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_6_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_6_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_6_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_6_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_6_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_6_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_6_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_6_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_6_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_6_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_6_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_6_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_6_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_6_pat_stride_buf_3;
  wire [32:0] _source_stream_conv2d_16_source_8_pat_count_0;
  wire [32:0] _source_stream_conv2d_16_source_8_pat_count_1;
  wire [32:0] _source_stream_conv2d_16_source_8_pat_count_2;
  wire [32:0] _source_stream_conv2d_16_source_8_pat_count_3;
  wire [31:0] _source_stream_conv2d_16_source_8_pat_cur_offset_0;
  wire [31:0] _source_stream_conv2d_16_source_8_pat_cur_offset_1;
  wire [31:0] _source_stream_conv2d_16_source_8_pat_cur_offset_2;
  wire [31:0] _source_stream_conv2d_16_source_8_pat_cur_offset_3;
  wire [32:0] _source_stream_conv2d_16_source_8_pat_size_0;
  wire [32:0] _source_stream_conv2d_16_source_8_pat_size_1;
  wire [32:0] _source_stream_conv2d_16_source_8_pat_size_2;
  wire [32:0] _source_stream_conv2d_16_source_8_pat_size_3;
  wire [32:0] _source_stream_conv2d_16_source_8_pat_size_buf_0;
  wire [32:0] _source_stream_conv2d_16_source_8_pat_size_buf_1;
  wire [32:0] _source_stream_conv2d_16_source_8_pat_size_buf_2;
  wire [32:0] _source_stream_conv2d_16_source_8_pat_size_buf_3;
  wire [31:0] _source_stream_conv2d_16_source_8_pat_stride_0;
  wire [31:0] _source_stream_conv2d_16_source_8_pat_stride_1;
  wire [31:0] _source_stream_conv2d_16_source_8_pat_stride_2;
  wire [31:0] _source_stream_conv2d_16_source_8_pat_stride_3;
  wire [31:0] _source_stream_conv2d_16_source_8_pat_stride_buf_0;
  wire [31:0] _source_stream_conv2d_16_source_8_pat_stride_buf_1;
  wire [31:0] _source_stream_conv2d_16_source_8_pat_stride_buf_2;
  wire [31:0] _source_stream_conv2d_16_source_8_pat_stride_buf_3;
  wire [32:0] _source_stream_matmul_29_source_19_pat_count_0;
  wire [32:0] _source_stream_matmul_29_source_19_pat_count_1;
  wire [32:0] _source_stream_matmul_29_source_19_pat_count_2;
  wire [32:0] _source_stream_matmul_29_source_19_pat_count_3;
  wire [31:0] _source_stream_matmul_29_source_19_pat_cur_offset_0;
  wire [31:0] _source_stream_matmul_29_source_19_pat_cur_offset_1;
  wire [31:0] _source_stream_matmul_29_source_19_pat_cur_offset_2;
  wire [31:0] _source_stream_matmul_29_source_19_pat_cur_offset_3;
  wire [32:0] _source_stream_matmul_29_source_19_pat_size_0;
  wire [32:0] _source_stream_matmul_29_source_19_pat_size_1;
  wire [32:0] _source_stream_matmul_29_source_19_pat_size_2;
  wire [32:0] _source_stream_matmul_29_source_19_pat_size_3;
  wire [32:0] _source_stream_matmul_29_source_19_pat_size_buf_0;
  wire [32:0] _source_stream_matmul_29_source_19_pat_size_buf_1;
  wire [32:0] _source_stream_matmul_29_source_19_pat_size_buf_2;
  wire [32:0] _source_stream_matmul_29_source_19_pat_size_buf_3;
  wire [31:0] _source_stream_matmul_29_source_19_pat_stride_0;
  wire [31:0] _source_stream_matmul_29_source_19_pat_stride_1;
  wire [31:0] _source_stream_matmul_29_source_19_pat_stride_2;
  wire [31:0] _source_stream_matmul_29_source_19_pat_stride_3;
  wire [31:0] _source_stream_matmul_29_source_19_pat_stride_buf_0;
  wire [31:0] _source_stream_matmul_29_source_19_pat_stride_buf_1;
  wire [31:0] _source_stream_matmul_29_source_19_pat_stride_buf_2;
  wire [31:0] _source_stream_matmul_29_source_19_pat_stride_buf_3;
  wire [32:0] _source_stream_matmul_29_source_20_pat_count_0;
  wire [32:0] _source_stream_matmul_29_source_20_pat_count_1;
  wire [32:0] _source_stream_matmul_29_source_20_pat_count_2;
  wire [32:0] _source_stream_matmul_29_source_20_pat_count_3;
  wire [31:0] _source_stream_matmul_29_source_20_pat_cur_offset_0;
  wire [31:0] _source_stream_matmul_29_source_20_pat_cur_offset_1;
  wire [31:0] _source_stream_matmul_29_source_20_pat_cur_offset_2;
  wire [31:0] _source_stream_matmul_29_source_20_pat_cur_offset_3;
  wire [32:0] _source_stream_matmul_29_source_20_pat_size_0;
  wire [32:0] _source_stream_matmul_29_source_20_pat_size_1;
  wire [32:0] _source_stream_matmul_29_source_20_pat_size_2;
  wire [32:0] _source_stream_matmul_29_source_20_pat_size_3;
  wire [32:0] _source_stream_matmul_29_source_20_pat_size_buf_0;
  wire [32:0] _source_stream_matmul_29_source_20_pat_size_buf_1;
  wire [32:0] _source_stream_matmul_29_source_20_pat_size_buf_2;
  wire [32:0] _source_stream_matmul_29_source_20_pat_size_buf_3;
  wire [31:0] _source_stream_matmul_29_source_20_pat_stride_0;
  wire [31:0] _source_stream_matmul_29_source_20_pat_stride_1;
  wire [31:0] _source_stream_matmul_29_source_20_pat_stride_2;
  wire [31:0] _source_stream_matmul_29_source_20_pat_stride_3;
  wire [31:0] _source_stream_matmul_29_source_20_pat_stride_buf_0;
  wire [31:0] _source_stream_matmul_29_source_20_pat_stride_buf_1;
  wire [31:0] _source_stream_matmul_29_source_20_pat_stride_buf_2;
  wire [31:0] _source_stream_matmul_29_source_20_pat_stride_buf_3;
  wire [32:0] _source_stream_matmul_29_source_6_pat_count_0;
  wire [32:0] _source_stream_matmul_29_source_6_pat_count_1;
  wire [32:0] _source_stream_matmul_29_source_6_pat_count_2;
  wire [32:0] _source_stream_matmul_29_source_6_pat_count_3;
  wire [31:0] _source_stream_matmul_29_source_6_pat_cur_offset_0;
  wire [31:0] _source_stream_matmul_29_source_6_pat_cur_offset_1;
  wire [31:0] _source_stream_matmul_29_source_6_pat_cur_offset_2;
  wire [31:0] _source_stream_matmul_29_source_6_pat_cur_offset_3;
  wire [32:0] _source_stream_matmul_29_source_6_pat_size_0;
  wire [32:0] _source_stream_matmul_29_source_6_pat_size_1;
  wire [32:0] _source_stream_matmul_29_source_6_pat_size_2;
  wire [32:0] _source_stream_matmul_29_source_6_pat_size_3;
  wire [32:0] _source_stream_matmul_29_source_6_pat_size_buf_0;
  wire [32:0] _source_stream_matmul_29_source_6_pat_size_buf_1;
  wire [32:0] _source_stream_matmul_29_source_6_pat_size_buf_2;
  wire [32:0] _source_stream_matmul_29_source_6_pat_size_buf_3;
  wire [31:0] _source_stream_matmul_29_source_6_pat_stride_0;
  wire [31:0] _source_stream_matmul_29_source_6_pat_stride_1;
  wire [31:0] _source_stream_matmul_29_source_6_pat_stride_2;
  wire [31:0] _source_stream_matmul_29_source_6_pat_stride_3;
  wire [31:0] _source_stream_matmul_29_source_6_pat_stride_buf_0;
  wire [31:0] _source_stream_matmul_29_source_6_pat_stride_buf_1;
  wire [31:0] _source_stream_matmul_29_source_6_pat_stride_buf_2;
  wire [31:0] _source_stream_matmul_29_source_6_pat_stride_buf_3;
  wire [32:0] _source_stream_matmul_29_source_8_pat_count_0;
  wire [32:0] _source_stream_matmul_29_source_8_pat_count_1;
  wire [32:0] _source_stream_matmul_29_source_8_pat_count_2;
  wire [32:0] _source_stream_matmul_29_source_8_pat_count_3;
  wire [31:0] _source_stream_matmul_29_source_8_pat_cur_offset_0;
  wire [31:0] _source_stream_matmul_29_source_8_pat_cur_offset_1;
  wire [31:0] _source_stream_matmul_29_source_8_pat_cur_offset_2;
  wire [31:0] _source_stream_matmul_29_source_8_pat_cur_offset_3;
  wire [32:0] _source_stream_matmul_29_source_8_pat_size_0;
  wire [32:0] _source_stream_matmul_29_source_8_pat_size_1;
  wire [32:0] _source_stream_matmul_29_source_8_pat_size_2;
  wire [32:0] _source_stream_matmul_29_source_8_pat_size_3;
  wire [32:0] _source_stream_matmul_29_source_8_pat_size_buf_0;
  wire [32:0] _source_stream_matmul_29_source_8_pat_size_buf_1;
  wire [32:0] _source_stream_matmul_29_source_8_pat_size_buf_2;
  wire [32:0] _source_stream_matmul_29_source_8_pat_size_buf_3;
  wire [31:0] _source_stream_matmul_29_source_8_pat_stride_0;
  wire [31:0] _source_stream_matmul_29_source_8_pat_stride_1;
  wire [31:0] _source_stream_matmul_29_source_8_pat_stride_2;
  wire [31:0] _source_stream_matmul_29_source_8_pat_stride_3;
  wire [31:0] _source_stream_matmul_29_source_8_pat_stride_buf_0;
  wire [31:0] _source_stream_matmul_29_source_8_pat_stride_buf_1;
  wire [31:0] _source_stream_matmul_29_source_8_pat_stride_buf_2;
  wire [31:0] _source_stream_matmul_29_source_8_pat_stride_buf_3;
  wire [32:0] _source_stream_max_pool_serial_18_source_1_pat_count_0;
  wire [32:0] _source_stream_max_pool_serial_18_source_1_pat_count_1;
  wire [32:0] _source_stream_max_pool_serial_18_source_1_pat_count_2;
  wire [32:0] _source_stream_max_pool_serial_18_source_1_pat_count_3;
  wire [31:0] _source_stream_max_pool_serial_18_source_1_pat_cur_offset_0;
  wire [31:0] _source_stream_max_pool_serial_18_source_1_pat_cur_offset_1;
  wire [31:0] _source_stream_max_pool_serial_18_source_1_pat_cur_offset_2;
  wire [31:0] _source_stream_max_pool_serial_18_source_1_pat_cur_offset_3;
  wire [32:0] _source_stream_max_pool_serial_18_source_1_pat_size_0;
  wire [32:0] _source_stream_max_pool_serial_18_source_1_pat_size_1;
  wire [32:0] _source_stream_max_pool_serial_18_source_1_pat_size_2;
  wire [32:0] _source_stream_max_pool_serial_18_source_1_pat_size_3;
  wire [32:0] _source_stream_max_pool_serial_18_source_1_pat_size_buf_0;
  wire [32:0] _source_stream_max_pool_serial_18_source_1_pat_size_buf_1;
  wire [32:0] _source_stream_max_pool_serial_18_source_1_pat_size_buf_2;
  wire [32:0] _source_stream_max_pool_serial_18_source_1_pat_size_buf_3;
  wire [31:0] _source_stream_max_pool_serial_18_source_1_pat_stride_0;
  wire [31:0] _source_stream_max_pool_serial_18_source_1_pat_stride_1;
  wire [31:0] _source_stream_max_pool_serial_18_source_1_pat_stride_2;
  wire [31:0] _source_stream_max_pool_serial_18_source_1_pat_stride_3;
  wire [31:0] _source_stream_max_pool_serial_18_source_1_pat_stride_buf_0;
  wire [31:0] _source_stream_max_pool_serial_18_source_1_pat_stride_buf_1;
  wire [31:0] _source_stream_max_pool_serial_18_source_1_pat_stride_buf_2;
  wire [31:0] _source_stream_max_pool_serial_18_source_1_pat_stride_buf_3;
  wire [11:0] _sra_data_104;
  wire [11:0] _sra_data_121;
  wire [11:0] _sra_data_138;
  wire [11:0] _sra_data_155;
  wire [11:0] _sra_data_172;
  wire [11:0] _sra_data_189;
  wire [11:0] _sra_data_206;
  wire [31:0] _sra_data_21;
  wire [39:0] _sra_data_42;
  wire [11:0] _sra_data_70;
  wire [11:0] _sra_data_87;
  wire [5:0] _stream_conv2d_16_constant_0_next_constant_data;
  wire _stream_conv2d_16_constant_15_next_constant_data;
  wire _stream_conv2d_16_constant_16_next_constant_data;
  wire [3:0] _stream_conv2d_16_constant_17_next_constant_data;
  wire [1:0] _stream_conv2d_16_constant_1_next_constant_data;
  wire [1:0] _stream_conv2d_16_constant_2_next_constant_data;
  wire [8:0] _stream_conv2d_16_constant_3_next_constant_data;
  wire _stream_conv2d_16_done;
  wire _stream_conv2d_16_end_flag;
  wire [31:0] _stream_conv2d_16_fsm;
  wire [32:0] _stream_conv2d_16_sink_37_sink_count;
  wire [31:0] _stream_conv2d_16_sink_37_sink_fsm_20;
  wire [2:0] _stream_conv2d_16_sink_37_sink_mode;
  wire [31:0] _stream_conv2d_16_sink_37_sink_offset;
  wire [7:0] _stream_conv2d_16_sink_37_sink_ram_sel;
  wire [32:0] _stream_conv2d_16_sink_37_sink_size;
  wire [31:0] _stream_conv2d_16_sink_37_sink_stride;
  wire [31:0] _stream_conv2d_16_sink_37_sink_stride_buf;
  wire [31:0] _stream_conv2d_16_sink_37_sink_waddr;
  wire [7:0] _stream_conv2d_16_sink_37_sink_wdata;
  wire _stream_conv2d_16_sink_37_sink_wenable;
  wire _stream_conv2d_16_sink_38_sink_wenable;
  wire _stream_conv2d_16_source_10_idle;
  wire [7:0] _stream_conv2d_16_source_10_source_empty_data;
  wire _stream_conv2d_16_source_10_source_ram_rvalid;
  wire _stream_conv2d_16_source_12_idle;
  wire [7:0] _stream_conv2d_16_source_12_source_empty_data;
  wire _stream_conv2d_16_source_12_source_ram_rvalid;
  wire _stream_conv2d_16_source_14_idle;
  wire [7:0] _stream_conv2d_16_source_14_source_empty_data;
  wire _stream_conv2d_16_source_14_source_ram_rvalid;
  wire _stream_conv2d_16_source_19_idle;
  wire [2:0] _stream_conv2d_16_source_19_source_mode;
  wire [31:0] _stream_conv2d_16_source_19_source_offset;
  wire [31:0] _stream_conv2d_16_source_19_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_19_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_19_source_pat_fsm_2;
  wire [31:0] _stream_conv2d_16_source_19_source_ram_raddr;
  wire [7:0] _stream_conv2d_16_source_19_source_ram_rdata;
  wire _stream_conv2d_16_source_19_source_ram_renable;
  wire _stream_conv2d_16_source_19_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_19_source_ram_sel;
  wire _stream_conv2d_16_source_20_idle;
  wire [2:0] _stream_conv2d_16_source_20_source_mode;
  wire [31:0] _stream_conv2d_16_source_20_source_offset;
  wire [31:0] _stream_conv2d_16_source_20_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_20_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_20_source_pat_fsm_3;
  wire [31:0] _stream_conv2d_16_source_20_source_ram_raddr;
  wire [7:0] _stream_conv2d_16_source_20_source_ram_rdata;
  wire _stream_conv2d_16_source_20_source_ram_renable;
  wire _stream_conv2d_16_source_20_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_20_source_ram_sel;
  wire _stream_conv2d_16_source_21_idle;
  wire [2:0] _stream_conv2d_16_source_21_source_mode;
  wire [31:0] _stream_conv2d_16_source_21_source_offset;
  wire [31:0] _stream_conv2d_16_source_21_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_21_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_21_source_pat_fsm_4;
  wire [31:0] _stream_conv2d_16_source_21_source_ram_raddr;
  wire [7:0] _stream_conv2d_16_source_21_source_ram_rdata;
  wire _stream_conv2d_16_source_21_source_ram_renable;
  wire _stream_conv2d_16_source_21_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_21_source_ram_sel;
  wire _stream_conv2d_16_source_22_idle;
  wire [2:0] _stream_conv2d_16_source_22_source_mode;
  wire [31:0] _stream_conv2d_16_source_22_source_offset;
  wire [31:0] _stream_conv2d_16_source_22_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_22_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_22_source_pat_fsm_5;
  wire [31:0] _stream_conv2d_16_source_22_source_ram_raddr;
  wire [7:0] _stream_conv2d_16_source_22_source_ram_rdata;
  wire _stream_conv2d_16_source_22_source_ram_renable;
  wire _stream_conv2d_16_source_22_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_22_source_ram_sel;
  wire _stream_conv2d_16_source_23_idle;
  wire [2:0] _stream_conv2d_16_source_23_source_mode;
  wire [31:0] _stream_conv2d_16_source_23_source_offset;
  wire [31:0] _stream_conv2d_16_source_23_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_23_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_23_source_pat_fsm_6;
  wire [31:0] _stream_conv2d_16_source_23_source_ram_raddr;
  wire [7:0] _stream_conv2d_16_source_23_source_ram_rdata;
  wire _stream_conv2d_16_source_23_source_ram_renable;
  wire _stream_conv2d_16_source_23_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_23_source_ram_sel;
  wire _stream_conv2d_16_source_24_idle;
  wire [2:0] _stream_conv2d_16_source_24_source_mode;
  wire [31:0] _stream_conv2d_16_source_24_source_offset;
  wire [31:0] _stream_conv2d_16_source_24_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_24_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_24_source_pat_fsm_7;
  wire [31:0] _stream_conv2d_16_source_24_source_ram_raddr;
  wire [7:0] _stream_conv2d_16_source_24_source_ram_rdata;
  wire _stream_conv2d_16_source_24_source_ram_renable;
  wire _stream_conv2d_16_source_24_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_24_source_ram_sel;
  wire _stream_conv2d_16_source_25_idle;
  wire [2:0] _stream_conv2d_16_source_25_source_mode;
  wire [31:0] _stream_conv2d_16_source_25_source_offset;
  wire [31:0] _stream_conv2d_16_source_25_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_25_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_25_source_pat_fsm_8;
  wire [31:0] _stream_conv2d_16_source_25_source_ram_raddr;
  wire [7:0] _stream_conv2d_16_source_25_source_ram_rdata;
  wire _stream_conv2d_16_source_25_source_ram_renable;
  wire _stream_conv2d_16_source_25_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_25_source_ram_sel;
  wire _stream_conv2d_16_source_26_idle;
  wire [2:0] _stream_conv2d_16_source_26_source_mode;
  wire [31:0] _stream_conv2d_16_source_26_source_offset;
  wire [31:0] _stream_conv2d_16_source_26_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_26_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_26_source_pat_fsm_9;
  wire [31:0] _stream_conv2d_16_source_26_source_ram_raddr;
  wire [7:0] _stream_conv2d_16_source_26_source_ram_rdata;
  wire _stream_conv2d_16_source_26_source_ram_renable;
  wire _stream_conv2d_16_source_26_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_26_source_ram_sel;
  wire _stream_conv2d_16_source_27_idle;
  wire [2:0] _stream_conv2d_16_source_27_source_mode;
  wire [31:0] _stream_conv2d_16_source_27_source_offset;
  wire [31:0] _stream_conv2d_16_source_27_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_27_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_27_source_pat_fsm_10;
  wire [31:0] _stream_conv2d_16_source_27_source_ram_raddr;
  wire [7:0] _stream_conv2d_16_source_27_source_ram_rdata;
  wire _stream_conv2d_16_source_27_source_ram_renable;
  wire _stream_conv2d_16_source_27_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_27_source_ram_sel;
  wire _stream_conv2d_16_source_28_idle;
  wire [2:0] _stream_conv2d_16_source_28_source_mode;
  wire [31:0] _stream_conv2d_16_source_28_source_offset;
  wire [31:0] _stream_conv2d_16_source_28_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_28_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_28_source_pat_fsm_11;
  wire [31:0] _stream_conv2d_16_source_28_source_ram_raddr;
  wire [3:0] _stream_conv2d_16_source_28_source_ram_rdata;
  wire _stream_conv2d_16_source_28_source_ram_renable;
  wire _stream_conv2d_16_source_28_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_28_source_ram_sel;
  wire _stream_conv2d_16_source_29_idle;
  wire [2:0] _stream_conv2d_16_source_29_source_mode;
  wire [31:0] _stream_conv2d_16_source_29_source_offset;
  wire [31:0] _stream_conv2d_16_source_29_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_29_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_29_source_pat_fsm_12;
  wire [31:0] _stream_conv2d_16_source_29_source_ram_raddr;
  wire [3:0] _stream_conv2d_16_source_29_source_ram_rdata;
  wire _stream_conv2d_16_source_29_source_ram_renable;
  wire _stream_conv2d_16_source_29_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_29_source_ram_sel;
  wire _stream_conv2d_16_source_30_idle;
  wire [2:0] _stream_conv2d_16_source_30_source_mode;
  wire [31:0] _stream_conv2d_16_source_30_source_offset;
  wire [31:0] _stream_conv2d_16_source_30_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_30_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_30_source_pat_fsm_13;
  wire [31:0] _stream_conv2d_16_source_30_source_ram_raddr;
  wire [3:0] _stream_conv2d_16_source_30_source_ram_rdata;
  wire _stream_conv2d_16_source_30_source_ram_renable;
  wire _stream_conv2d_16_source_30_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_30_source_ram_sel;
  wire _stream_conv2d_16_source_31_idle;
  wire [2:0] _stream_conv2d_16_source_31_source_mode;
  wire [31:0] _stream_conv2d_16_source_31_source_offset;
  wire [31:0] _stream_conv2d_16_source_31_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_31_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_31_source_pat_fsm_14;
  wire [31:0] _stream_conv2d_16_source_31_source_ram_raddr;
  wire [3:0] _stream_conv2d_16_source_31_source_ram_rdata;
  wire _stream_conv2d_16_source_31_source_ram_renable;
  wire _stream_conv2d_16_source_31_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_31_source_ram_sel;
  wire _stream_conv2d_16_source_32_idle;
  wire [2:0] _stream_conv2d_16_source_32_source_mode;
  wire [31:0] _stream_conv2d_16_source_32_source_offset;
  wire [31:0] _stream_conv2d_16_source_32_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_32_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_32_source_pat_fsm_15;
  wire [31:0] _stream_conv2d_16_source_32_source_ram_raddr;
  wire [3:0] _stream_conv2d_16_source_32_source_ram_rdata;
  wire _stream_conv2d_16_source_32_source_ram_renable;
  wire _stream_conv2d_16_source_32_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_32_source_ram_sel;
  wire _stream_conv2d_16_source_33_idle;
  wire [2:0] _stream_conv2d_16_source_33_source_mode;
  wire [31:0] _stream_conv2d_16_source_33_source_offset;
  wire [31:0] _stream_conv2d_16_source_33_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_33_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_33_source_pat_fsm_16;
  wire [31:0] _stream_conv2d_16_source_33_source_ram_raddr;
  wire [3:0] _stream_conv2d_16_source_33_source_ram_rdata;
  wire _stream_conv2d_16_source_33_source_ram_renable;
  wire _stream_conv2d_16_source_33_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_33_source_ram_sel;
  wire _stream_conv2d_16_source_34_idle;
  wire [2:0] _stream_conv2d_16_source_34_source_mode;
  wire [31:0] _stream_conv2d_16_source_34_source_offset;
  wire [31:0] _stream_conv2d_16_source_34_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_34_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_34_source_pat_fsm_17;
  wire [31:0] _stream_conv2d_16_source_34_source_ram_raddr;
  wire [3:0] _stream_conv2d_16_source_34_source_ram_rdata;
  wire _stream_conv2d_16_source_34_source_ram_renable;
  wire _stream_conv2d_16_source_34_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_34_source_ram_sel;
  wire _stream_conv2d_16_source_35_idle;
  wire [2:0] _stream_conv2d_16_source_35_source_mode;
  wire [31:0] _stream_conv2d_16_source_35_source_offset;
  wire [31:0] _stream_conv2d_16_source_35_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_35_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_35_source_pat_fsm_18;
  wire [31:0] _stream_conv2d_16_source_35_source_ram_raddr;
  wire [3:0] _stream_conv2d_16_source_35_source_ram_rdata;
  wire _stream_conv2d_16_source_35_source_ram_renable;
  wire _stream_conv2d_16_source_35_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_35_source_ram_sel;
  wire _stream_conv2d_16_source_36_idle;
  wire [2:0] _stream_conv2d_16_source_36_source_mode;
  wire [31:0] _stream_conv2d_16_source_36_source_offset;
  wire [31:0] _stream_conv2d_16_source_36_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_36_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_36_source_pat_fsm_19;
  wire [31:0] _stream_conv2d_16_source_36_source_ram_raddr;
  wire [3:0] _stream_conv2d_16_source_36_source_ram_rdata;
  wire _stream_conv2d_16_source_36_source_ram_renable;
  wire _stream_conv2d_16_source_36_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_36_source_ram_sel;
  wire _stream_conv2d_16_source_6_idle;
  wire [2:0] _stream_conv2d_16_source_6_source_mode;
  wire [31:0] _stream_conv2d_16_source_6_source_offset;
  wire [31:0] _stream_conv2d_16_source_6_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_6_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_6_source_pat_fsm_0;
  wire [31:0] _stream_conv2d_16_source_6_source_ram_raddr;
  wire [7:0] _stream_conv2d_16_source_6_source_ram_rdata;
  wire _stream_conv2d_16_source_6_source_ram_renable;
  wire _stream_conv2d_16_source_6_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_6_source_ram_sel;
  wire _stream_conv2d_16_source_8_idle;
  wire [2:0] _stream_conv2d_16_source_8_source_mode;
  wire [31:0] _stream_conv2d_16_source_8_source_offset;
  wire [31:0] _stream_conv2d_16_source_8_source_offset_buf;
  wire [31:0] _stream_conv2d_16_source_8_source_pat_all_offset;
  wire [31:0] _stream_conv2d_16_source_8_source_pat_fsm_1;
  wire [31:0] _stream_conv2d_16_source_8_source_ram_raddr;
  wire [7:0] _stream_conv2d_16_source_8_source_ram_rdata;
  wire _stream_conv2d_16_source_8_source_ram_renable;
  wire _stream_conv2d_16_source_8_source_ram_rvalid;
  wire [7:0] _stream_conv2d_16_source_8_source_ram_sel;
  wire _stream_conv2d_16_source_busy;
  wire _stream_conv2d_16_start;
  wire _stream_conv2d_16_start_flag;
  wire _stream_conv2d_16_term_sink;
  wire [10:0] _stream_matmul_29_constant_0_next_constant_data;
  wire _stream_matmul_29_constant_15_next_constant_data;
  wire _stream_matmul_29_constant_16_next_constant_data;
  wire [3:0] _stream_matmul_29_constant_17_next_constant_data;
  wire [1:0] _stream_matmul_29_constant_18_next_constant_data;
  wire _stream_matmul_29_constant_1_next_constant_data;
  wire _stream_matmul_29_constant_2_next_constant_data;
  wire _stream_matmul_29_constant_3_next_constant_data;
  wire _stream_matmul_29_done;
  wire _stream_matmul_29_end_flag;
  wire [31:0] _stream_matmul_29_fsm;
  wire [32:0] _stream_matmul_29_sink_21_sink_count;
  wire [31:0] _stream_matmul_29_sink_21_sink_fsm_4;
  wire [2:0] _stream_matmul_29_sink_21_sink_mode;
  wire [31:0] _stream_matmul_29_sink_21_sink_offset;
  wire [7:0] _stream_matmul_29_sink_21_sink_ram_sel;
  wire [32:0] _stream_matmul_29_sink_21_sink_size;
  wire [31:0] _stream_matmul_29_sink_21_sink_stride;
  wire [31:0] _stream_matmul_29_sink_21_sink_stride_buf;
  wire [31:0] _stream_matmul_29_sink_21_sink_waddr;
  wire [7:0] _stream_matmul_29_sink_21_sink_wdata;
  wire _stream_matmul_29_sink_21_sink_wenable;
  wire _stream_matmul_29_sink_22_sink_wenable;
  wire _stream_matmul_29_source_10_idle;
  wire [7:0] _stream_matmul_29_source_10_source_empty_data;
  wire _stream_matmul_29_source_10_source_ram_rvalid;
  wire _stream_matmul_29_source_12_idle;
  wire [7:0] _stream_matmul_29_source_12_source_empty_data;
  wire _stream_matmul_29_source_12_source_ram_rvalid;
  wire _stream_matmul_29_source_14_idle;
  wire [7:0] _stream_matmul_29_source_14_source_empty_data;
  wire _stream_matmul_29_source_14_source_ram_rvalid;
  wire _stream_matmul_29_source_19_idle;
  wire [2:0] _stream_matmul_29_source_19_source_mode;
  wire [31:0] _stream_matmul_29_source_19_source_offset;
  wire [31:0] _stream_matmul_29_source_19_source_offset_buf;
  wire [31:0] _stream_matmul_29_source_19_source_pat_all_offset;
  wire [31:0] _stream_matmul_29_source_19_source_pat_fsm_2;
  wire [31:0] _stream_matmul_29_source_19_source_ram_raddr;
  wire [7:0] _stream_matmul_29_source_19_source_ram_rdata;
  wire _stream_matmul_29_source_19_source_ram_renable;
  wire _stream_matmul_29_source_19_source_ram_rvalid;
  wire [7:0] _stream_matmul_29_source_19_source_ram_sel;
  wire _stream_matmul_29_source_20_idle;
  wire [2:0] _stream_matmul_29_source_20_source_mode;
  wire [31:0] _stream_matmul_29_source_20_source_offset;
  wire [31:0] _stream_matmul_29_source_20_source_offset_buf;
  wire [31:0] _stream_matmul_29_source_20_source_pat_all_offset;
  wire [31:0] _stream_matmul_29_source_20_source_pat_fsm_3;
  wire [31:0] _stream_matmul_29_source_20_source_ram_raddr;
  wire [3:0] _stream_matmul_29_source_20_source_ram_rdata;
  wire _stream_matmul_29_source_20_source_ram_renable;
  wire _stream_matmul_29_source_20_source_ram_rvalid;
  wire [7:0] _stream_matmul_29_source_20_source_ram_sel;
  wire _stream_matmul_29_source_6_idle;
  wire [2:0] _stream_matmul_29_source_6_source_mode;
  wire [31:0] _stream_matmul_29_source_6_source_offset;
  wire [31:0] _stream_matmul_29_source_6_source_offset_buf;
  wire [31:0] _stream_matmul_29_source_6_source_pat_all_offset;
  wire [31:0] _stream_matmul_29_source_6_source_pat_fsm_0;
  wire [31:0] _stream_matmul_29_source_6_source_ram_raddr;
  wire [7:0] _stream_matmul_29_source_6_source_ram_rdata;
  wire _stream_matmul_29_source_6_source_ram_renable;
  wire _stream_matmul_29_source_6_source_ram_rvalid;
  wire [7:0] _stream_matmul_29_source_6_source_ram_sel;
  wire _stream_matmul_29_source_8_idle;
  wire [2:0] _stream_matmul_29_source_8_source_mode;
  wire [31:0] _stream_matmul_29_source_8_source_offset;
  wire [31:0] _stream_matmul_29_source_8_source_offset_buf;
  wire [31:0] _stream_matmul_29_source_8_source_pat_all_offset;
  wire [31:0] _stream_matmul_29_source_8_source_pat_fsm_1;
  wire [31:0] _stream_matmul_29_source_8_source_ram_raddr;
  wire [7:0] _stream_matmul_29_source_8_source_ram_rdata;
  wire _stream_matmul_29_source_8_source_ram_renable;
  wire _stream_matmul_29_source_8_source_ram_rvalid;
  wire [7:0] _stream_matmul_29_source_8_source_ram_sel;
  wire _stream_matmul_29_source_busy;
  wire _stream_matmul_29_start;
  wire _stream_matmul_29_start_flag;
  wire _stream_matmul_29_term_sink;
  wire [2:0] _stream_max_pool_serial_18_constant_0_next_constant_data;
  wire [3:0] _stream_max_pool_serial_18_constant_2_next_constant_data;
  wire _stream_max_pool_serial_18_done;
  wire _stream_max_pool_serial_18_end_flag;
  wire [31:0] _stream_max_pool_serial_18_fsm;
  wire _stream_max_pool_serial_18_reduce_reset;
  wire [32:0] _stream_max_pool_serial_18_sink_3_sink_count;
  wire [31:0] _stream_max_pool_serial_18_sink_3_sink_fsm_1;
  wire [2:0] _stream_max_pool_serial_18_sink_3_sink_mode;
  wire [31:0] _stream_max_pool_serial_18_sink_3_sink_offset;
  wire [7:0] _stream_max_pool_serial_18_sink_3_sink_ram_sel;
  wire [32:0] _stream_max_pool_serial_18_sink_3_sink_size;
  wire [31:0] _stream_max_pool_serial_18_sink_3_sink_stride;
  wire [31:0] _stream_max_pool_serial_18_sink_3_sink_stride_buf;
  wire [31:0] _stream_max_pool_serial_18_sink_3_sink_waddr;
  wire [7:0] _stream_max_pool_serial_18_sink_3_sink_wdata;
  wire _stream_max_pool_serial_18_sink_3_sink_wenable;
  wire _stream_max_pool_serial_18_sink_4_sink_wenable;
  wire _stream_max_pool_serial_18_source_1_idle;
  wire [2:0] _stream_max_pool_serial_18_source_1_source_mode;
  wire [31:0] _stream_max_pool_serial_18_source_1_source_offset;
  wire [31:0] _stream_max_pool_serial_18_source_1_source_offset_buf;
  wire [31:0] _stream_max_pool_serial_18_source_1_source_pat_all_offset;
  wire [31:0] _stream_max_pool_serial_18_source_1_source_pat_fsm_0;
  wire [31:0] _stream_max_pool_serial_18_source_1_source_ram_raddr;
  wire [7:0] _stream_max_pool_serial_18_source_1_source_ram_rdata;
  wire _stream_max_pool_serial_18_source_1_source_ram_renable;
  wire _stream_max_pool_serial_18_source_1_source_ram_rvalid;
  wire [7:0] _stream_max_pool_serial_18_source_1_source_ram_sel;
  wire _stream_max_pool_serial_18_source_busy;
  wire _stream_max_pool_serial_18_start;
  wire _stream_max_pool_serial_18_start_flag;
  wire _stream_max_pool_serial_18_term_sink;
  wire _substream__reduce_max_13_size_data_cond_792_43;
  wire _substream__reduce_max_13_x_data_cond_792_42;
  wire _substream_acc_0_rshift_data_cond_747_37;
  wire _substream_acc_0_rshift_data_cond_879_49;
  wire _substream_acc_0_size_data_cond_747_38;
  wire _substream_acc_0_size_data_cond_879_50;
  wire _substream_acc_0_x_data_cond_747_36;
  wire _substream_acc_0_x_data_cond_879_48;
  wire _substream_add_tree_1_var0_data_cond_877_47;
  wire _substream_add_tree_2_var0_data_cond_745_27;
  wire _substream_add_tree_2_var1_data_cond_745_28;
  wire _substream_add_tree_2_var2_data_cond_745_29;
  wire _substream_add_tree_2_var3_data_cond_745_30;
  wire _substream_add_tree_2_var4_data_cond_745_31;
  wire _substream_add_tree_2_var5_data_cond_745_32;
  wire _substream_add_tree_2_var6_data_cond_745_33;
  wire _substream_add_tree_2_var7_data_cond_745_34;
  wire _substream_add_tree_2_var8_data_cond_745_35;
  wire _substream_mul_10_rshift_data_cond_694_20;
  wire _substream_mul_10_x_data_cond_694_18;
  wire _substream_mul_10_y_data_cond_694_19;
  wire _substream_mul_11_rshift_data_cond_711_23;
  wire _substream_mul_11_x_data_cond_711_21;
  wire _substream_mul_11_y_data_cond_711_22;
  wire _substream_mul_12_rshift_data_cond_728_26;
  wire _substream_mul_12_x_data_cond_728_24;
  wire _substream_mul_12_y_data_cond_728_25;
  wire _substream_mul_4_rshift_data_cond_592_2;
  wire _substream_mul_4_rshift_data_cond_874_46;
  wire _substream_mul_4_x_data_cond_592_0;
  wire _substream_mul_4_x_data_cond_874_44;
  wire _substream_mul_4_y_data_cond_592_1;
  wire _substream_mul_4_y_data_cond_874_45;
  wire _substream_mul_5_rshift_data_cond_609_5;
  wire _substream_mul_5_x_data_cond_609_3;
  wire _substream_mul_5_y_data_cond_609_4;
  wire _substream_mul_6_rshift_data_cond_626_8;
  wire _substream_mul_6_x_data_cond_626_6;
  wire _substream_mul_6_y_data_cond_626_7;
  wire _substream_mul_7_rshift_data_cond_643_11;
  wire _substream_mul_7_x_data_cond_643_9;
  wire _substream_mul_7_y_data_cond_643_10;
  wire _substream_mul_8_rshift_data_cond_660_14;
  wire _substream_mul_8_x_data_cond_660_12;
  wire _substream_mul_8_y_data_cond_660_13;
  wire _substream_mul_9_rshift_data_cond_677_17;
  wire _substream_mul_9_x_data_cond_677_15;
  wire _substream_mul_9_y_data_cond_677_16;
  wire _substream_mul_rshift_clip_3_rshift_data_cond_763_41;
  wire _substream_mul_rshift_clip_3_rshift_data_cond_884_53;
  wire _substream_mul_rshift_clip_3_x_data_cond_763_39;
  wire _substream_mul_rshift_clip_3_x_data_cond_884_51;
  wire _substream_mul_rshift_clip_3_y_data_cond_763_40;
  wire _substream_mul_rshift_clip_3_y_data_cond_884_52;
  wire [39:0] _times_data_41;
  wire \_times_mul_41.CLK ;
  wire [31:0] \_times_mul_41.a ;
  wire [7:0] \_times_mul_41.b ;
  wire [39:0] \_times_mul_41.c ;
  wire \_times_mul_41.mult.CLK ;
  wire [31:0] \_times_mul_41.mult._a ;
  wire [7:0] \_times_mul_41.mult._b ;
  wire [39:0] \_times_mul_41.mult._mul ;
  wire [39:0] \_times_mul_41.mult._pipe_mul0 ;
  wire [39:0] \_times_mul_41.mult._pipe_mul1 ;
  wire [31:0] \_times_mul_41.mult.a ;
  wire [7:0] \_times_mul_41.mult.b ;
  wire [39:0] \_times_mul_41.mult.c ;
  wire \_times_mul_41.mult.update ;
  wire \_times_mul_41.update ;
  wire [39:0] _times_mul_odata_41;
  wire [39:0] _times_mul_odata_reg_41;
  wire _times_mul_update_41;
  wire [5:0] _tmp_0;
  wire _tmp_1;
  wire [10:0] _tmp_100;
  wire _tmp_1000;
  wire [7:0] _tmp_1001;
  wire _tmp_1002;
  wire _tmp_1003;
  wire _tmp_1004;
  wire _tmp_1005;
  wire [33:0] _tmp_1006;
  wire _tmp_1007;
  wire [33:0] _tmp_101;
  wire _tmp_1010;
  wire _tmp_1012;
  wire [7:0] _tmp_1013;
  wire _tmp_1014;
  wire _tmp_1015;
  wire _tmp_1016;
  wire _tmp_1017;
  wire [33:0] _tmp_1018;
  wire [8:0] _tmp_1019;
  wire _tmp_102;
  wire _tmp_1020;
  wire [1:0] _tmp_1027;
  wire [9:0] _tmp_103;
  wire [7:0] _tmp_1032;
  wire _tmp_1035;
  wire [1:0] _tmp_1037;
  wire [9:0] _tmp_104;
  wire _tmp_1040;
  wire _tmp_1042;
  wire _tmp_1044;
  wire _tmp_1046;
  wire _tmp_1048;
  wire [9:0] _tmp_105;
  wire _tmp_1050;
  wire _tmp_1052;
  wire _tmp_1054;
  wire _tmp_1056;
  wire _tmp_1058;
  wire [9:0] _tmp_106;
  wire _tmp_1060;
  wire _tmp_1062;
  wire _tmp_1064;
  wire _tmp_1066;
  wire _tmp_1068;
  wire [9:0] _tmp_107;
  wire _tmp_1070;
  wire _tmp_1072;
  wire _tmp_1075;
  wire _tmp_1077;
  wire [7:0] _tmp_1078;
  wire _tmp_1079;
  wire [9:0] _tmp_108;
  wire _tmp_1080;
  wire _tmp_1081;
  wire _tmp_1082;
  wire [33:0] _tmp_1083;
  wire _tmp_1084;
  wire _tmp_1087;
  wire _tmp_1089;
  wire [9:0] _tmp_109;
  wire [7:0] _tmp_1090;
  wire _tmp_1091;
  wire _tmp_1092;
  wire _tmp_1093;
  wire _tmp_1094;
  wire [33:0] _tmp_1095;
  wire _tmp_1096;
  wire _tmp_1099;
  wire [9:0] _tmp_110;
  wire _tmp_1101;
  wire [7:0] _tmp_1102;
  wire _tmp_1103;
  wire _tmp_1104;
  wire _tmp_1105;
  wire _tmp_1106;
  wire [33:0] _tmp_1107;
  wire _tmp_1108;
  wire [9:0] _tmp_111;
  wire _tmp_1111;
  wire _tmp_1113;
  wire [7:0] _tmp_1114;
  wire _tmp_1115;
  wire _tmp_1116;
  wire _tmp_1117;
  wire _tmp_1118;
  wire [33:0] _tmp_1119;
  wire [9:0] _tmp_112;
  wire _tmp_1120;
  wire [33:0] _tmp_1124;
  wire _tmp_1125;
  wire [33:0] _tmp_1126;
  wire _tmp_1127;
  wire [33:0] _tmp_1128;
  wire _tmp_1129;
  wire [9:0] _tmp_113;
  wire [33:0] _tmp_1130;
  wire _tmp_1131;
  wire [33:0] _tmp_1136;
  wire _tmp_1137;
  wire [33:0] _tmp_1138;
  wire _tmp_1139;
  wire [9:0] _tmp_114;
  wire [33:0] _tmp_1140;
  wire _tmp_1141;
  wire [33:0] _tmp_1142;
  wire _tmp_1143;
  wire [33:0] _tmp_1144;
  wire _tmp_1145;
  wire [33:0] _tmp_1146;
  wire _tmp_1147;
  wire [33:0] _tmp_1148;
  wire _tmp_1149;
  wire [9:0] _tmp_115;
  wire [33:0] _tmp_1150;
  wire _tmp_1151;
  wire [33:0] _tmp_1155;
  wire _tmp_1156;
  wire [33:0] _tmp_1157;
  wire _tmp_1158;
  wire [33:0] _tmp_1159;
  wire [9:0] _tmp_116;
  wire _tmp_1160;
  wire [33:0] _tmp_1161;
  wire _tmp_1162;
  wire [9:0] _tmp_117;
  wire [1:0] _tmp_1170;
  wire [7:0] _tmp_1175;
  wire _tmp_1178;
  wire [9:0] _tmp_118;
  wire [1:0] _tmp_1181;
  wire [7:0] _tmp_1186;
  wire _tmp_1189;
  wire [9:0] _tmp_119;
  wire [33:0] _tmp_12;
  wire [9:0] _tmp_120;
  wire [1:0] _tmp_1201;
  wire [7:0] _tmp_1206;
  wire _tmp_1209;
  wire [9:0] _tmp_121;
  wire [2:0] _tmp_1211;
  wire [9:0] _tmp_122;
  wire [3:0] _tmp_1220;
  wire _tmp_1223;
  wire [1:0] _tmp_1225;
  wire _tmp_1227;
  wire _tmp_1229;
  wire [9:0] _tmp_123;
  wire _tmp_1231;
  wire _tmp_1233;
  wire _tmp_1235;
  wire _tmp_1237;
  wire _tmp_1239;
  wire [9:0] _tmp_124;
  wire _tmp_1241;
  wire _tmp_1243;
  wire _tmp_1245;
  wire _tmp_1247;
  wire _tmp_1249;
  wire [9:0] _tmp_125;
  wire _tmp_1251;
  wire _tmp_1253;
  wire _tmp_1255;
  wire _tmp_1257;
  wire _tmp_1259;
  wire [9:0] _tmp_126;
  wire _tmp_1261;
  wire _tmp_1263;
  wire _tmp_1265;
  wire _tmp_1267;
  wire _tmp_1269;
  wire [9:0] _tmp_127;
  wire _tmp_1271;
  wire _tmp_1273;
  wire _tmp_1275;
  wire _tmp_1277;
  wire _tmp_1279;
  wire [9:0] _tmp_128;
  wire _tmp_1281;
  wire _tmp_1283;
  wire _tmp_1285;
  wire _tmp_1287;
  wire _tmp_1289;
  wire [9:0] _tmp_129;
  wire _tmp_1291;
  wire _tmp_1293;
  wire _tmp_1295;
  wire _tmp_1297;
  wire _tmp_1299;
  wire _tmp_13;
  wire [3:0] _tmp_130;
  wire _tmp_1301;
  wire _tmp_1303;
  wire _tmp_1305;
  wire _tmp_1307;
  wire _tmp_1309;
  wire [10:0] _tmp_131;
  wire _tmp_1312;
  wire _tmp_1314;
  wire [7:0] _tmp_1315;
  wire _tmp_1316;
  wire _tmp_1317;
  wire _tmp_1318;
  wire _tmp_1319;
  wire [33:0] _tmp_132;
  wire [33:0] _tmp_1320;
  wire _tmp_1321;
  wire _tmp_1324;
  wire _tmp_1326;
  wire [7:0] _tmp_1327;
  wire _tmp_1328;
  wire _tmp_1329;
  wire _tmp_133;
  wire _tmp_1330;
  wire _tmp_1331;
  wire [33:0] _tmp_1332;
  wire _tmp_1333;
  wire _tmp_1336;
  wire _tmp_1338;
  wire [7:0] _tmp_1339;
  wire [9:0] _tmp_134;
  wire _tmp_1340;
  wire _tmp_1341;
  wire _tmp_1342;
  wire _tmp_1343;
  wire [33:0] _tmp_1344;
  wire _tmp_1345;
  wire _tmp_1348;
  wire [9:0] _tmp_135;
  wire _tmp_1350;
  wire [7:0] _tmp_1351;
  wire _tmp_1352;
  wire _tmp_1353;
  wire _tmp_1354;
  wire _tmp_1355;
  wire [33:0] _tmp_1356;
  wire _tmp_1357;
  wire [9:0] _tmp_136;
  wire [9:0] _tmp_137;
  wire [9:0] _tmp_138;
  wire [9:0] _tmp_139;
  wire [33:0] _tmp_14;
  wire [9:0] _tmp_140;
  wire [9:0] _tmp_141;
  wire [9:0] _tmp_142;
  wire [9:0] _tmp_143;
  wire [9:0] _tmp_144;
  wire [9:0] _tmp_145;
  wire [9:0] _tmp_146;
  wire [9:0] _tmp_147;
  wire [9:0] _tmp_148;
  wire [9:0] _tmp_149;
  wire _tmp_15;
  wire [9:0] _tmp_150;
  wire [9:0] _tmp_151;
  wire [9:0] _tmp_152;
  wire [9:0] _tmp_153;
  wire [9:0] _tmp_154;
  wire [9:0] _tmp_155;
  wire [9:0] _tmp_156;
  wire [9:0] _tmp_157;
  wire [9:0] _tmp_158;
  wire [9:0] _tmp_159;
  wire [33:0] _tmp_16;
  wire [9:0] _tmp_160;
  wire [3:0] _tmp_161;
  wire [10:0] _tmp_162;
  wire [33:0] _tmp_163;
  wire _tmp_164;
  wire [9:0] _tmp_165;
  wire [9:0] _tmp_166;
  wire [9:0] _tmp_167;
  wire [9:0] _tmp_168;
  wire [9:0] _tmp_169;
  wire _tmp_17;
  wire [9:0] _tmp_170;
  wire [9:0] _tmp_171;
  wire [9:0] _tmp_172;
  wire [9:0] _tmp_173;
  wire [9:0] _tmp_174;
  wire [9:0] _tmp_175;
  wire [9:0] _tmp_176;
  wire [9:0] _tmp_177;
  wire [9:0] _tmp_178;
  wire [9:0] _tmp_179;
  wire [33:0] _tmp_18;
  wire [9:0] _tmp_180;
  wire [9:0] _tmp_181;
  wire [9:0] _tmp_182;
  wire [9:0] _tmp_183;
  wire [9:0] _tmp_184;
  wire [9:0] _tmp_185;
  wire [9:0] _tmp_186;
  wire [9:0] _tmp_187;
  wire [9:0] _tmp_188;
  wire [9:0] _tmp_189;
  wire _tmp_19;
  wire [9:0] _tmp_190;
  wire [9:0] _tmp_191;
  wire [3:0] _tmp_192;
  wire [10:0] _tmp_193;
  wire [33:0] _tmp_194;
  wire _tmp_195;
  wire [9:0] _tmp_196;
  wire [9:0] _tmp_197;
  wire [9:0] _tmp_198;
  wire [9:0] _tmp_199;
  wire _tmp_2;
  wire [8:0] _tmp_20;
  wire [9:0] _tmp_200;
  wire [9:0] _tmp_201;
  wire [9:0] _tmp_202;
  wire [9:0] _tmp_203;
  wire [9:0] _tmp_204;
  wire [9:0] _tmp_205;
  wire [9:0] _tmp_206;
  wire [9:0] _tmp_207;
  wire [9:0] _tmp_208;
  wire [9:0] _tmp_209;
  wire [9:0] _tmp_210;
  wire [9:0] _tmp_211;
  wire [9:0] _tmp_212;
  wire [9:0] _tmp_213;
  wire [9:0] _tmp_214;
  wire [9:0] _tmp_215;
  wire [9:0] _tmp_216;
  wire [9:0] _tmp_217;
  wire [9:0] _tmp_218;
  wire [9:0] _tmp_219;
  wire [9:0] _tmp_220;
  wire [9:0] _tmp_221;
  wire [9:0] _tmp_222;
  wire [3:0] _tmp_223;
  wire [10:0] _tmp_224;
  wire [33:0] _tmp_225;
  wire _tmp_226;
  wire [9:0] _tmp_227;
  wire [9:0] _tmp_228;
  wire [9:0] _tmp_229;
  wire [9:0] _tmp_230;
  wire [9:0] _tmp_231;
  wire [9:0] _tmp_232;
  wire [9:0] _tmp_233;
  wire [9:0] _tmp_234;
  wire [9:0] _tmp_235;
  wire [9:0] _tmp_236;
  wire [9:0] _tmp_237;
  wire [9:0] _tmp_238;
  wire [9:0] _tmp_239;
  wire [9:0] _tmp_240;
  wire [9:0] _tmp_241;
  wire [9:0] _tmp_242;
  wire [9:0] _tmp_243;
  wire [9:0] _tmp_244;
  wire [9:0] _tmp_245;
  wire [9:0] _tmp_246;
  wire [9:0] _tmp_247;
  wire [9:0] _tmp_248;
  wire [9:0] _tmp_249;
  wire [33:0] _tmp_25;
  wire [9:0] _tmp_250;
  wire [9:0] _tmp_251;
  wire [9:0] _tmp_252;
  wire [9:0] _tmp_253;
  wire [3:0] _tmp_254;
  wire [10:0] _tmp_255;
  wire [33:0] _tmp_256;
  wire _tmp_257;
  wire [9:0] _tmp_258;
  wire [9:0] _tmp_259;
  wire _tmp_26;
  wire [9:0] _tmp_260;
  wire [9:0] _tmp_261;
  wire [9:0] _tmp_262;
  wire [9:0] _tmp_263;
  wire [9:0] _tmp_264;
  wire [9:0] _tmp_265;
  wire [9:0] _tmp_266;
  wire [9:0] _tmp_267;
  wire [9:0] _tmp_268;
  wire [9:0] _tmp_269;
  wire [33:0] _tmp_27;
  wire [9:0] _tmp_270;
  wire [9:0] _tmp_271;
  wire [9:0] _tmp_272;
  wire [9:0] _tmp_273;
  wire [9:0] _tmp_274;
  wire [9:0] _tmp_275;
  wire [9:0] _tmp_276;
  wire [9:0] _tmp_277;
  wire [9:0] _tmp_278;
  wire [9:0] _tmp_279;
  wire _tmp_28;
  wire [9:0] _tmp_280;
  wire [9:0] _tmp_281;
  wire [9:0] _tmp_282;
  wire [9:0] _tmp_283;
  wire [9:0] _tmp_284;
  wire [3:0] _tmp_285;
  wire [33:0] _tmp_29;
  wire [9:0] _tmp_291;
  wire [33:0] _tmp_292;
  wire _tmp_293;
  wire [8:0] _tmp_294;
  wire [8:0] _tmp_295;
  wire [8:0] _tmp_296;
  wire [8:0] _tmp_297;
  wire [8:0] _tmp_298;
  wire [8:0] _tmp_299;
  wire _tmp_3;
  wire _tmp_30;
  wire [8:0] _tmp_300;
  wire [8:0] _tmp_301;
  wire [8:0] _tmp_302;
  wire [1:0] _tmp_303;
  wire [9:0] _tmp_304;
  wire [33:0] _tmp_305;
  wire _tmp_306;
  wire [8:0] _tmp_307;
  wire [8:0] _tmp_308;
  wire [8:0] _tmp_309;
  wire [33:0] _tmp_31;
  wire [8:0] _tmp_310;
  wire [8:0] _tmp_311;
  wire [8:0] _tmp_312;
  wire [8:0] _tmp_313;
  wire [8:0] _tmp_314;
  wire [8:0] _tmp_315;
  wire [1:0] _tmp_316;
  wire [9:0] _tmp_317;
  wire [33:0] _tmp_318;
  wire _tmp_319;
  wire _tmp_32;
  wire [8:0] _tmp_320;
  wire [8:0] _tmp_321;
  wire [8:0] _tmp_322;
  wire [8:0] _tmp_323;
  wire [8:0] _tmp_324;
  wire [8:0] _tmp_325;
  wire [8:0] _tmp_326;
  wire [8:0] _tmp_327;
  wire [8:0] _tmp_328;
  wire [1:0] _tmp_329;
  wire [9:0] _tmp_330;
  wire [33:0] _tmp_331;
  wire _tmp_332;
  wire [8:0] _tmp_333;
  wire [8:0] _tmp_334;
  wire [8:0] _tmp_335;
  wire [8:0] _tmp_336;
  wire [8:0] _tmp_337;
  wire [8:0] _tmp_338;
  wire [8:0] _tmp_339;
  wire [8:0] _tmp_340;
  wire [8:0] _tmp_341;
  wire [1:0] _tmp_342;
  wire [9:0] _tmp_348;
  wire [33:0] _tmp_349;
  wire _tmp_350;
  wire [8:0] _tmp_351;
  wire [8:0] _tmp_352;
  wire [8:0] _tmp_353;
  wire [8:0] _tmp_354;
  wire [8:0] _tmp_355;
  wire [8:0] _tmp_356;
  wire [8:0] _tmp_357;
  wire [8:0] _tmp_358;
  wire [8:0] _tmp_359;
  wire [1:0] _tmp_360;
  wire [9:0] _tmp_361;
  wire [33:0] _tmp_362;
  wire _tmp_363;
  wire [8:0] _tmp_364;
  wire [8:0] _tmp_365;
  wire [8:0] _tmp_366;
  wire [8:0] _tmp_367;
  wire [8:0] _tmp_368;
  wire [8:0] _tmp_369;
  wire [8:0] _tmp_370;
  wire [8:0] _tmp_371;
  wire [8:0] _tmp_372;
  wire [1:0] _tmp_373;
  wire [9:0] _tmp_374;
  wire [33:0] _tmp_375;
  wire _tmp_376;
  wire [8:0] _tmp_377;
  wire [8:0] _tmp_378;
  wire [8:0] _tmp_379;
  wire [10:0] _tmp_38;
  wire [8:0] _tmp_380;
  wire [8:0] _tmp_381;
  wire [8:0] _tmp_382;
  wire [8:0] _tmp_383;
  wire [8:0] _tmp_384;
  wire [8:0] _tmp_385;
  wire [1:0] _tmp_386;
  wire [9:0] _tmp_387;
  wire [33:0] _tmp_388;
  wire _tmp_389;
  wire [33:0] _tmp_39;
  wire [8:0] _tmp_390;
  wire [8:0] _tmp_391;
  wire [8:0] _tmp_392;
  wire [8:0] _tmp_393;
  wire [8:0] _tmp_394;
  wire [8:0] _tmp_395;
  wire [8:0] _tmp_396;
  wire [8:0] _tmp_397;
  wire [8:0] _tmp_398;
  wire [1:0] _tmp_399;
  wire _tmp_4;
  wire _tmp_40;
  wire [9:0] _tmp_405;
  wire [33:0] _tmp_406;
  wire _tmp_407;
  wire [8:0] _tmp_408;
  wire [8:0] _tmp_409;
  wire [9:0] _tmp_41;
  wire [8:0] _tmp_410;
  wire [8:0] _tmp_411;
  wire [8:0] _tmp_412;
  wire [8:0] _tmp_413;
  wire [8:0] _tmp_414;
  wire [8:0] _tmp_415;
  wire [8:0] _tmp_416;
  wire [1:0] _tmp_417;
  wire [9:0] _tmp_418;
  wire [33:0] _tmp_419;
  wire [9:0] _tmp_42;
  wire _tmp_420;
  wire [8:0] _tmp_421;
  wire [8:0] _tmp_422;
  wire [8:0] _tmp_423;
  wire [8:0] _tmp_424;
  wire [8:0] _tmp_425;
  wire [8:0] _tmp_426;
  wire [8:0] _tmp_427;
  wire [8:0] _tmp_428;
  wire [8:0] _tmp_429;
  wire [9:0] _tmp_43;
  wire [1:0] _tmp_430;
  wire [9:0] _tmp_431;
  wire [33:0] _tmp_432;
  wire _tmp_433;
  wire [8:0] _tmp_434;
  wire [8:0] _tmp_435;
  wire [8:0] _tmp_436;
  wire [8:0] _tmp_437;
  wire [8:0] _tmp_438;
  wire [8:0] _tmp_439;
  wire [9:0] _tmp_44;
  wire [8:0] _tmp_440;
  wire [8:0] _tmp_441;
  wire [8:0] _tmp_442;
  wire [1:0] _tmp_443;
  wire [9:0] _tmp_444;
  wire [33:0] _tmp_445;
  wire _tmp_446;
  wire [8:0] _tmp_447;
  wire [8:0] _tmp_448;
  wire [8:0] _tmp_449;
  wire [9:0] _tmp_45;
  wire [8:0] _tmp_450;
  wire [8:0] _tmp_451;
  wire [8:0] _tmp_452;
  wire [8:0] _tmp_453;
  wire [8:0] _tmp_454;
  wire [8:0] _tmp_455;
  wire [1:0] _tmp_456;
  wire [9:0] _tmp_46;
  wire [1:0] _tmp_464;
  wire [7:0] _tmp_469;
  wire [9:0] _tmp_47;
  wire _tmp_472;
  wire [1:0] _tmp_475;
  wire [9:0] _tmp_48;
  wire [7:0] _tmp_480;
  wire _tmp_483;
  wire [9:0] _tmp_49;
  wire [1:0] _tmp_495;
  wire [3:0] _tmp_5;
  wire [9:0] _tmp_50;
  wire [7:0] _tmp_500;
  wire _tmp_503;
  wire [1:0] _tmp_505;
  wire [9:0] _tmp_51;
  wire [7:0] _tmp_510;
  wire _tmp_513;
  wire [1:0] _tmp_515;
  wire [9:0] _tmp_52;
  wire [7:0] _tmp_520;
  wire _tmp_523;
  wire [1:0] _tmp_525;
  wire [9:0] _tmp_53;
  wire [7:0] _tmp_530;
  wire _tmp_533;
  wire [1:0] _tmp_535;
  wire [9:0] _tmp_54;
  wire [7:0] _tmp_540;
  wire _tmp_543;
  wire [1:0] _tmp_545;
  wire [9:0] _tmp_55;
  wire [7:0] _tmp_550;
  wire _tmp_553;
  wire [1:0] _tmp_555;
  wire [9:0] _tmp_56;
  wire [7:0] _tmp_560;
  wire _tmp_563;
  wire [1:0] _tmp_565;
  wire [9:0] _tmp_57;
  wire [7:0] _tmp_570;
  wire _tmp_573;
  wire [1:0] _tmp_575;
  wire [9:0] _tmp_58;
  wire [7:0] _tmp_580;
  wire _tmp_583;
  wire [2:0] _tmp_585;
  wire [9:0] _tmp_59;
  wire [3:0] _tmp_594;
  wire _tmp_597;
  wire [2:0] _tmp_599;
  wire [31:0] _tmp_6;
  wire [9:0] _tmp_60;
  wire [3:0] _tmp_608;
  wire [9:0] _tmp_61;
  wire _tmp_611;
  wire [2:0] _tmp_613;
  wire [9:0] _tmp_62;
  wire [3:0] _tmp_622;
  wire _tmp_625;
  wire [2:0] _tmp_627;
  wire [9:0] _tmp_63;
  wire [3:0] _tmp_636;
  wire _tmp_639;
  wire [9:0] _tmp_64;
  wire [2:0] _tmp_641;
  wire [9:0] _tmp_65;
  wire [3:0] _tmp_650;
  wire _tmp_653;
  wire [2:0] _tmp_655;
  wire [9:0] _tmp_66;
  wire [3:0] _tmp_664;
  wire _tmp_667;
  wire [2:0] _tmp_669;
  wire [9:0] _tmp_67;
  wire [3:0] _tmp_678;
  wire [3:0] _tmp_68;
  wire _tmp_681;
  wire [2:0] _tmp_683;
  wire [10:0] _tmp_69;
  wire [3:0] _tmp_692;
  wire _tmp_695;
  wire [2:0] _tmp_697;
  wire _tmp_7;
  wire [33:0] _tmp_70;
  wire [3:0] _tmp_706;
  wire _tmp_709;
  wire _tmp_71;
  wire [1:0] _tmp_711;
  wire _tmp_713;
  wire _tmp_715;
  wire _tmp_717;
  wire _tmp_719;
  wire [9:0] _tmp_72;
  wire _tmp_721;
  wire _tmp_723;
  wire _tmp_725;
  wire _tmp_727;
  wire _tmp_729;
  wire [9:0] _tmp_73;
  wire _tmp_731;
  wire _tmp_733;
  wire _tmp_735;
  wire _tmp_737;
  wire _tmp_739;
  wire [9:0] _tmp_74;
  wire _tmp_741;
  wire _tmp_743;
  wire _tmp_745;
  wire _tmp_747;
  wire _tmp_749;
  wire [9:0] _tmp_75;
  wire _tmp_751;
  wire _tmp_753;
  wire _tmp_755;
  wire _tmp_757;
  wire _tmp_759;
  wire [9:0] _tmp_76;
  wire _tmp_761;
  wire _tmp_763;
  wire _tmp_765;
  wire _tmp_767;
  wire _tmp_769;
  wire [9:0] _tmp_77;
  wire _tmp_771;
  wire _tmp_773;
  wire _tmp_775;
  wire _tmp_777;
  wire _tmp_779;
  wire [9:0] _tmp_78;
  wire _tmp_781;
  wire _tmp_783;
  wire _tmp_785;
  wire _tmp_787;
  wire _tmp_789;
  wire [9:0] _tmp_79;
  wire _tmp_791;
  wire _tmp_793;
  wire _tmp_795;
  wire _tmp_797;
  wire _tmp_799;
  wire [31:0] _tmp_8;
  wire [9:0] _tmp_80;
  wire _tmp_801;
  wire _tmp_803;
  wire _tmp_805;
  wire _tmp_807;
  wire _tmp_809;
  wire [9:0] _tmp_81;
  wire _tmp_811;
  wire _tmp_813;
  wire _tmp_815;
  wire _tmp_817;
  wire _tmp_819;
  wire [9:0] _tmp_82;
  wire _tmp_821;
  wire _tmp_823;
  wire _tmp_825;
  wire _tmp_827;
  wire _tmp_829;
  wire [9:0] _tmp_83;
  wire _tmp_831;
  wire _tmp_833;
  wire _tmp_835;
  wire _tmp_837;
  wire _tmp_839;
  wire [9:0] _tmp_84;
  wire _tmp_841;
  wire _tmp_843;
  wire _tmp_845;
  wire _tmp_847;
  wire _tmp_849;
  wire [9:0] _tmp_85;
  wire _tmp_851;
  wire _tmp_853;
  wire _tmp_855;
  wire _tmp_857;
  wire _tmp_859;
  wire [9:0] _tmp_86;
  wire _tmp_861;
  wire _tmp_863;
  wire _tmp_865;
  wire _tmp_867;
  wire _tmp_869;
  wire [9:0] _tmp_87;
  wire _tmp_871;
  wire _tmp_873;
  wire _tmp_875;
  wire _tmp_877;
  wire _tmp_879;
  wire [9:0] _tmp_88;
  wire _tmp_881;
  wire _tmp_883;
  wire _tmp_885;
  wire _tmp_887;
  wire _tmp_889;
  wire [9:0] _tmp_89;
  wire _tmp_891;
  wire _tmp_893;
  wire _tmp_895;
  wire _tmp_897;
  wire _tmp_899;
  wire [9:0] _tmp_90;
  wire _tmp_901;
  wire _tmp_903;
  wire _tmp_905;
  wire _tmp_907;
  wire _tmp_909;
  wire [9:0] _tmp_91;
  wire _tmp_911;
  wire _tmp_913;
  wire _tmp_915;
  wire _tmp_917;
  wire _tmp_919;
  wire [9:0] _tmp_92;
  wire _tmp_921;
  wire _tmp_923;
  wire _tmp_925;
  wire _tmp_927;
  wire _tmp_929;
  wire [9:0] _tmp_93;
  wire _tmp_931;
  wire _tmp_933;
  wire _tmp_935;
  wire _tmp_937;
  wire _tmp_939;
  wire [9:0] _tmp_94;
  wire _tmp_941;
  wire _tmp_943;
  wire _tmp_945;
  wire _tmp_947;
  wire _tmp_949;
  wire [9:0] _tmp_95;
  wire _tmp_951;
  wire _tmp_953;
  wire _tmp_955;
  wire _tmp_957;
  wire _tmp_959;
  wire [9:0] _tmp_96;
  wire _tmp_961;
  wire _tmp_963;
  wire _tmp_965;
  wire _tmp_967;
  wire _tmp_969;
  wire [9:0] _tmp_97;
  wire _tmp_971;
  wire _tmp_974;
  wire _tmp_976;
  wire [7:0] _tmp_977;
  wire _tmp_978;
  wire _tmp_979;
  wire [9:0] _tmp_98;
  wire _tmp_980;
  wire _tmp_981;
  wire [33:0] _tmp_982;
  wire _tmp_983;
  wire _tmp_986;
  wire _tmp_988;
  wire [7:0] _tmp_989;
  wire [3:0] _tmp_99;
  wire _tmp_990;
  wire _tmp_991;
  wire _tmp_992;
  wire _tmp_993;
  wire [33:0] _tmp_994;
  wire _tmp_995;
  wire _tmp_998;
  wire [31:0] _wdata_10;
  wire [31:0] _wdata_1122;
  wire [31:0] _wdata_1134;
  wire [31:0] _wdata_1153;
  wire [31:0] _wdata_23;
  wire [31:0] _wdata_289;
  wire [31:0] _wdata_346;
  wire [31:0] _wdata_36;
  wire [31:0] _wdata_403;
  wire _wvalid_11;
  wire _wvalid_1123;
  wire _wvalid_1135;
  wire _wvalid_1154;
  wire _wvalid_24;
  wire _wvalid_290;
  wire _wvalid_347;
  wire _wvalid_37;
  wire _wvalid_404;
  wire [5:0] acc_0_rshift_data;
  wire [31:0] acc_0_size_data;
  wire [31:0] acc_0_sum_data;
  wire acc_0_valid_data;
  wire [31:0] acc_0_x_data;
  wire [31:0] add_tree_1_sum_data;
  wire [31:0] add_tree_1_var0_data;
  wire [31:0] add_tree_2_sum_data;
  wire [31:0] add_tree_2_var0_data;
  wire [31:0] add_tree_2_var1_data;
  wire [31:0] add_tree_2_var2_data;
  wire [31:0] add_tree_2_var3_data;
  wire [31:0] add_tree_2_var4_data;
  wire [31:0] add_tree_2_var5_data;
  wire [31:0] add_tree_2_var6_data;
  wire [31:0] add_tree_2_var7_data;
  wire [31:0] add_tree_2_var8_data;
  wire axim_flag_1021;
  wire axim_flag_1022;
  wire axim_flag_1023;
  wire axim_flag_1071;
  wire axim_flag_1121;
  wire axim_flag_1132;
  wire axim_flag_1133;
  wire axim_flag_1152;
  wire axim_flag_1308;
  wire axim_flag_21;
  wire axim_flag_22;
  wire axim_flag_288;
  wire axim_flag_345;
  wire axim_flag_35;
  wire axim_flag_402;
  wire axim_flag_9;
  wire axim_flag_970;
  wire [31:0] control_conv2d_16;
  wire [31:0] control_matmul_29;
  wire [31:0] control_max_pool_serial_18;
  wire [31:0] conv2d_16_act_base_offset;
  wire [31:0] conv2d_16_act_base_offset_bat;
  wire [31:0] conv2d_16_act_base_offset_row;
  wire [31:0] conv2d_16_act_page_comp_offset_0;
  wire [31:0] conv2d_16_act_page_comp_offset_1;
  wire [31:0] conv2d_16_act_page_comp_offset_2;
  wire [31:0] conv2d_16_act_page_comp_offset_buf_0;
  wire [31:0] conv2d_16_act_page_comp_offset_buf_1;
  wire [31:0] conv2d_16_act_page_comp_offset_buf_2;
  wire [31:0] conv2d_16_act_page_dma_offset_0;
  wire [31:0] conv2d_16_act_page_dma_offset_1;
  wire [31:0] conv2d_16_act_page_dma_offset_2;
  wire [31:0] conv2d_16_arg_objaddr_0;
  wire [31:0] conv2d_16_arg_objaddr_1;
  wire [31:0] conv2d_16_arg_objaddr_2;
  wire [31:0] conv2d_16_arg_objaddr_3;
  wire [31:0] conv2d_16_bat_count;
  wire [31:0] conv2d_16_col_count;
  wire [1:0] conv2d_16_col_select;
  wire [31:0] conv2d_16_comp_fsm;
  wire [1:0] conv2d_16_control_param_index;
  wire conv2d_16_dma_flag_0;
  wire conv2d_16_dma_flag_1;
  wire conv2d_16_dma_flag_2;
  wire conv2d_16_dma_out_mask_0;
  wire conv2d_16_dma_pad_mask_0;
  wire conv2d_16_dma_pad_mask_1;
  wire conv2d_16_dma_pad_mask_2;
  wire [31:0] conv2d_16_filter_base_offset;
  wire [31:0] conv2d_16_filter_page_comp_offset;
  wire [31:0] conv2d_16_filter_page_comp_offset_buf;
  wire [31:0] conv2d_16_filter_page_dma_offset;
  wire [31:0] conv2d_16_mux_act_gaddr_0;
  wire [31:0] conv2d_16_mux_act_gaddr_1;
  wire [31:0] conv2d_16_mux_act_gaddr_2;
  wire conv2d_16_mux_dma_flag_0;
  wire conv2d_16_mux_dma_flag_1;
  wire conv2d_16_mux_dma_flag_2;
  wire conv2d_16_mux_dma_pad_mask_0;
  wire conv2d_16_mux_dma_pad_mask_1;
  wire conv2d_16_mux_dma_pad_mask_2;
  wire conv2d_16_mux_next_dma_flag_0;
  wire conv2d_16_mux_next_dma_flag_1;
  wire conv2d_16_mux_next_dma_flag_2;
  wire [31:0] conv2d_16_next_out_write_size;
  wire [31:0] conv2d_16_next_stream_num_ops;
  wire [31:0] conv2d_16_objaddr;
  wire [31:0] conv2d_16_och_count;
  wire [31:0] conv2d_16_och_count_buf;
  wire [31:0] conv2d_16_out_base_offset;
  wire [31:0] conv2d_16_out_base_offset_bat;
  wire [31:0] conv2d_16_out_base_offset_col;
  wire [31:0] conv2d_16_out_base_offset_och;
  wire [31:0] conv2d_16_out_base_offset_row;
  wire [31:0] conv2d_16_out_base_offset_val;
  wire [31:0] conv2d_16_out_laddr_offset;
  wire conv2d_16_out_page;
  wire [31:0] conv2d_16_out_page_comp_offset;
  wire [31:0] conv2d_16_out_page_comp_offset_buf;
  wire [31:0] conv2d_16_out_page_dma_offset;
  wire [31:0] conv2d_16_out_ram_select;
  wire [31:0] conv2d_16_out_row_count;
  wire [31:0] conv2d_16_prev_bat_count;
  wire [31:0] conv2d_16_prev_och_count;
  wire [31:0] conv2d_16_prev_row_count;
  wire [1:0] conv2d_16_prev_row_select;
  wire [31:0] conv2d_16_row_count;
  wire [31:0] conv2d_16_row_count_buf;
  wire [1:0] conv2d_16_row_select;
  wire [1:0] conv2d_16_row_select_buf;
  wire conv2d_16_skip_comp;
  wire conv2d_16_skip_read_act;
  wire conv2d_16_skip_read_filter;
  wire conv2d_16_skip_write_out;
  wire [31:0] conv2d_16_stream_act_local_0;
  wire [31:0] conv2d_16_stream_act_local_1;
  wire [31:0] conv2d_16_stream_act_local_2;
  wire [31:0] conv2d_16_stream_act_local_3;
  wire [31:0] conv2d_16_stream_act_local_4;
  wire [31:0] conv2d_16_stream_act_local_5;
  wire [31:0] conv2d_16_stream_act_local_6;
  wire [31:0] conv2d_16_stream_act_local_7;
  wire [31:0] conv2d_16_stream_act_local_8;
  wire [31:0] conv2d_16_stream_out_local;
  wire [31:0] conv2d_16_stream_out_local_col;
  wire [31:0] conv2d_16_stream_out_local_val;
  wire conv2d_16_stream_pad_mask_0_0;
  wire conv2d_16_stream_pad_mask_0_1;
  wire conv2d_16_stream_pad_mask_0_2;
  wire conv2d_16_stream_pad_mask_1_0;
  wire conv2d_16_stream_pad_mask_1_1;
  wire conv2d_16_stream_pad_mask_1_2;
  wire conv2d_16_stream_pad_mask_2_0;
  wire conv2d_16_stream_pad_mask_2_1;
  wire conv2d_16_stream_pad_mask_2_2;
  wire [8:0] conv2d_16_stream_pad_masks;
  wire [31:0] conv2d_16_sync_comp_count;
  wire [31:0] conv2d_16_sync_out_count;
  wire conv2d_16_update_act;
  wire conv2d_16_update_filter;
  wire cparam_conv2d_16_act_func_index;
  wire [5:0] cparam_conv2d_16_act_num_col;
  wire [5:0] cparam_conv2d_16_act_num_row;
  wire [31:0] cparam_conv2d_16_act_offset_values_0;
  wire [31:0] cparam_conv2d_16_act_offset_values_1;
  wire [31:0] cparam_conv2d_16_act_offset_values_2;
  wire [5:0] cparam_conv2d_16_act_read_block;
  wire [8:0] cparam_conv2d_16_act_read_size;
  wire [6:0] cparam_conv2d_16_act_read_step;
  wire [8:0] cparam_conv2d_16_act_row_step;
  wire [6:0] cparam_conv2d_16_bias_num;
  wire cparam_conv2d_16_bias_scala;
  wire [1:0] cparam_conv2d_16_col_select_initval;
  wire cparam_conv2d_16_cshamt_mul_value;
  wire [3:0] cparam_conv2d_16_cshamt_out_value;
  wire cparam_conv2d_16_cshamt_sum_value;
  wire cparam_conv2d_16_data_stationary;
  wire cparam_conv2d_16_dma_flag_conds_0;
  wire cparam_conv2d_16_dma_flag_conds_1;
  wire cparam_conv2d_16_dma_flag_conds_2;
  wire [13:0] cparam_conv2d_16_filter_base_step;
  wire [1:0] cparam_conv2d_16_filter_num_col_minus_stride_col_mod;
  wire [5:0] cparam_conv2d_16_filter_read_block;
  wire [14:0] cparam_conv2d_16_filter_read_size;
  wire [11:0] cparam_conv2d_16_filter_read_step;
  wire cparam_conv2d_16_inc_act_laddr_conds_0;
  wire cparam_conv2d_16_inc_act_laddr_conds_1;
  wire cparam_conv2d_16_inc_act_laddr_conds_10;
  wire cparam_conv2d_16_inc_act_laddr_conds_11;
  wire cparam_conv2d_16_inc_act_laddr_conds_12;
  wire cparam_conv2d_16_inc_act_laddr_conds_13;
  wire cparam_conv2d_16_inc_act_laddr_conds_14;
  wire cparam_conv2d_16_inc_act_laddr_conds_15;
  wire cparam_conv2d_16_inc_act_laddr_conds_16;
  wire cparam_conv2d_16_inc_act_laddr_conds_17;
  wire cparam_conv2d_16_inc_act_laddr_conds_18;
  wire cparam_conv2d_16_inc_act_laddr_conds_19;
  wire cparam_conv2d_16_inc_act_laddr_conds_2;
  wire cparam_conv2d_16_inc_act_laddr_conds_20;
  wire cparam_conv2d_16_inc_act_laddr_conds_21;
  wire cparam_conv2d_16_inc_act_laddr_conds_22;
  wire cparam_conv2d_16_inc_act_laddr_conds_23;
  wire cparam_conv2d_16_inc_act_laddr_conds_24;
  wire cparam_conv2d_16_inc_act_laddr_conds_25;
  wire cparam_conv2d_16_inc_act_laddr_conds_26;
  wire cparam_conv2d_16_inc_act_laddr_conds_3;
  wire cparam_conv2d_16_inc_act_laddr_conds_4;
  wire cparam_conv2d_16_inc_act_laddr_conds_5;
  wire cparam_conv2d_16_inc_act_laddr_conds_6;
  wire cparam_conv2d_16_inc_act_laddr_conds_7;
  wire cparam_conv2d_16_inc_act_laddr_conds_8;
  wire cparam_conv2d_16_inc_act_laddr_conds_9;
  wire [5:0] cparam_conv2d_16_inc_act_laddr_large;
  wire cparam_conv2d_16_inc_act_laddr_small;
  wire [6:0] cparam_conv2d_16_inc_out_laddr_col;
  wire [5:0] cparam_conv2d_16_inc_sync_out;
  wire cparam_conv2d_16_inc_sync_out_res;
  wire cparam_conv2d_16_keep_filter;
  wire cparam_conv2d_16_keep_input;
  wire cparam_conv2d_16_max_bat_count;
  wire [4:0] cparam_conv2d_16_max_col_count;
  wire cparam_conv2d_16_max_och_count;
  wire [4:0] cparam_conv2d_16_max_row_count;
  wire [7:0] cparam_conv2d_16_och_count_step;
  wire [6:0] cparam_conv2d_16_out_col_step;
  wire [5:0] cparam_conv2d_16_out_num_col;
  wire [5:0] cparam_conv2d_16_out_num_row;
  wire [6:0] cparam_conv2d_16_out_och_step;
  wire cparam_conv2d_16_out_offset_values_0;
  wire [9:0] cparam_conv2d_16_out_row_step;
  wire [9:0] cparam_conv2d_16_out_write_size;
  wire [9:0] cparam_conv2d_16_out_write_size_res;
  wire cparam_conv2d_16_pad_col_left;
  wire cparam_conv2d_16_pad_row_top;
  wire cparam_conv2d_16_scale_num;
  wire cparam_conv2d_16_scale_scala;
  wire cparam_conv2d_16_stream_act_local_large_flags_0;
  wire cparam_conv2d_16_stream_act_local_large_flags_1;
  wire cparam_conv2d_16_stream_act_local_large_flags_2;
  wire [6:0] cparam_conv2d_16_stream_act_local_large_offset;
  wire cparam_conv2d_16_stream_act_local_small_flags_0;
  wire cparam_conv2d_16_stream_act_local_small_flags_1;
  wire cparam_conv2d_16_stream_act_local_small_flags_2;
  wire cparam_conv2d_16_stream_act_local_small_offset;
  wire [5:0] cparam_conv2d_16_stream_aligned_reduce_size;
  wire [6:0] cparam_conv2d_16_stream_num_ops;
  wire [6:0] cparam_conv2d_16_stream_num_ops_res;
  wire cparam_conv2d_16_stream_omit_mask;
  wire [5:0] cparam_conv2d_16_stream_reduce_size;
  wire cparam_conv2d_16_stride_col_mod_filter_num;
  wire cparam_conv2d_16_stride_col_par_col;
  wire cparam_conv2d_16_stride_row_par_row;
  wire cparam_conv2d_16_vshamt_mul_num;
  wire cparam_conv2d_16_vshamt_mul_scala;
  wire cparam_conv2d_16_vshamt_out_num;
  wire cparam_conv2d_16_vshamt_out_scala;
  wire cparam_conv2d_16_vshamt_sum_num;
  wire cparam_conv2d_16_vshamt_sum_scala;
  wire [10:0] cparam_matmul_29_act_bat_step;
  wire cparam_matmul_29_act_func_index;
  wire cparam_matmul_29_act_num_col;
  wire cparam_matmul_29_act_num_row;
  wire [31:0] cparam_matmul_29_act_offset_values_0;
  wire [10:0] cparam_matmul_29_act_read_size;
  wire [10:0] cparam_matmul_29_act_read_step;
  wire [10:0] cparam_matmul_29_act_row_step;
  wire [8:0] cparam_matmul_29_bias_num;
  wire cparam_matmul_29_bias_scala;
  wire cparam_matmul_29_col_select_initval;
  wire cparam_matmul_29_cshamt_mul_value;
  wire [3:0] cparam_matmul_29_cshamt_out_value;
  wire cparam_matmul_29_cshamt_sum_value;
  wire cparam_matmul_29_data_stationary;
  wire cparam_matmul_29_dma_flag_conds_0;
  wire [11:0] cparam_matmul_29_filter_base_step;
  wire cparam_matmul_29_filter_num_col_minus_stride_col_mod;
  wire [12:0] cparam_matmul_29_filter_read_size;
  wire [12:0] cparam_matmul_29_filter_read_step;
  wire cparam_matmul_29_inc_act_laddr_conds_0;
  wire [10:0] cparam_matmul_29_inc_act_laddr_large;
  wire [10:0] cparam_matmul_29_inc_act_laddr_small;
  wire [8:0] cparam_matmul_29_inc_out_laddr_col;
  wire cparam_matmul_29_inc_sync_out;
  wire cparam_matmul_29_inc_sync_out_res;
  wire cparam_matmul_29_keep_filter;
  wire cparam_matmul_29_keep_input;
  wire cparam_matmul_29_max_bat_count;
  wire cparam_matmul_29_max_col_count;
  wire [7:0] cparam_matmul_29_max_och_count;
  wire cparam_matmul_29_max_row_count;
  wire [5:0] cparam_matmul_29_och_count_step;
  wire [8:0] cparam_matmul_29_out_bat_step;
  wire [8:0] cparam_matmul_29_out_col_step;
  wire cparam_matmul_29_out_num_col;
  wire cparam_matmul_29_out_num_row;
  wire [4:0] cparam_matmul_29_out_och_step;
  wire cparam_matmul_29_out_offset_values_0;
  wire [8:0] cparam_matmul_29_out_row_step;
  wire [4:0] cparam_matmul_29_out_write_size;
  wire [4:0] cparam_matmul_29_out_write_size_res;
  wire cparam_matmul_29_pad_col_left;
  wire cparam_matmul_29_pad_row_top;
  wire cparam_matmul_29_scale_num;
  wire cparam_matmul_29_scale_scala;
  wire cparam_matmul_29_stream_act_local_large_flags_0;
  wire cparam_matmul_29_stream_act_local_large_offset;
  wire cparam_matmul_29_stream_act_local_small_flags_0;
  wire cparam_matmul_29_stream_act_local_small_offset;
  wire [10:0] cparam_matmul_29_stream_aligned_reduce_size;
  wire [4:0] cparam_matmul_29_stream_num_ops;
  wire [4:0] cparam_matmul_29_stream_num_ops_res;
  wire cparam_matmul_29_stream_omit_mask;
  wire [10:0] cparam_matmul_29_stream_reduce_size;
  wire cparam_matmul_29_stride_col_mod_filter_num;
  wire cparam_matmul_29_stride_col_par_col;
  wire cparam_matmul_29_stride_row_par_row;
  wire cparam_matmul_29_vshamt_mul_num;
  wire cparam_matmul_29_vshamt_mul_scala;
  wire cparam_matmul_29_vshamt_out_num;
  wire cparam_matmul_29_vshamt_out_scala;
  wire cparam_matmul_29_vshamt_sum_num;
  wire cparam_matmul_29_vshamt_sum_scala;
  wire [5:0] cparam_max_pool_serial_18_act_num_col;
  wire [5:0] cparam_max_pool_serial_18_act_num_row;
  wire [31:0] cparam_max_pool_serial_18_act_offset_values_0;
  wire [31:0] cparam_max_pool_serial_18_act_offset_values_1;
  wire [6:0] cparam_max_pool_serial_18_act_read_block;
  wire [9:0] cparam_max_pool_serial_18_act_read_size;
  wire [10:0] cparam_max_pool_serial_18_act_row_step;
  wire cparam_max_pool_serial_18_col_select_initval;
  wire [7:0] cparam_max_pool_serial_18_inc_act_laddr;
  wire [6:0] cparam_max_pool_serial_18_inc_out_laddr;
  wire [1:0] cparam_max_pool_serial_18_ksize_col_minus_stride_col_mod;
  wire cparam_max_pool_serial_18_local_pad_offset;
  wire cparam_max_pool_serial_18_max_bat_count;
  wire [4:0] cparam_max_pool_serial_18_max_col_count;
  wire [4:0] cparam_max_pool_serial_18_max_row_count;
  wire [8:0] cparam_max_pool_serial_18_out_row_step;
  wire [8:0] cparam_max_pool_serial_18_out_write_size;
  wire cparam_max_pool_serial_18_pad_col_left;
  wire cparam_max_pool_serial_18_pad_row_top;
  wire [6:0] cparam_max_pool_serial_18_stream_size;
  wire [1:0] cparam_max_pool_serial_18_stride_col;
  wire cparam_max_pool_serial_18_stride_col_mod_ksize;
  wire [1:0] cparam_max_pool_serial_18_stride_row;
  wire [31:0] main_fsm;
  wire [31:0] matmul_29_act_base_offset;
  wire [31:0] matmul_29_act_base_offset_bat;
  wire [31:0] matmul_29_act_base_offset_row;
  wire [31:0] matmul_29_act_page_comp_offset_0;
  wire [31:0] matmul_29_act_page_comp_offset_buf_0;
  wire [31:0] matmul_29_act_page_dma_offset_0;
  wire [31:0] matmul_29_arg_objaddr_0;
  wire [31:0] matmul_29_arg_objaddr_1;
  wire [31:0] matmul_29_arg_objaddr_2;
  wire [31:0] matmul_29_arg_objaddr_3;
  wire [31:0] matmul_29_bat_count;
  wire [31:0] matmul_29_col_count;
  wire matmul_29_col_select;
  wire [31:0] matmul_29_comp_fsm;
  wire [1:0] matmul_29_control_param_index;
  wire matmul_29_dma_flag_0;
  wire matmul_29_dma_out_mask_0;
  wire matmul_29_dma_pad_mask_0;
  wire [31:0] matmul_29_filter_base_offset;
  wire [31:0] matmul_29_filter_page_comp_offset;
  wire [31:0] matmul_29_filter_page_comp_offset_buf;
  wire [31:0] matmul_29_filter_page_dma_offset;
  wire [31:0] matmul_29_mux_act_gaddr_0;
  wire matmul_29_mux_dma_flag_0;
  wire matmul_29_mux_dma_pad_mask_0;
  wire [31:0] matmul_29_next_out_write_size;
  wire [31:0] matmul_29_next_stream_num_ops;
  wire [31:0] matmul_29_objaddr;
  wire [31:0] matmul_29_och_count;
  wire [31:0] matmul_29_och_count_buf;
  wire [31:0] matmul_29_out_base_offset;
  wire [31:0] matmul_29_out_base_offset_bat;
  wire [31:0] matmul_29_out_base_offset_col;
  wire [31:0] matmul_29_out_base_offset_och;
  wire [31:0] matmul_29_out_base_offset_row;
  wire [31:0] matmul_29_out_base_offset_val;
  wire [31:0] matmul_29_out_laddr_offset;
  wire matmul_29_out_page;
  wire [31:0] matmul_29_out_page_comp_offset;
  wire [31:0] matmul_29_out_page_comp_offset_buf;
  wire [31:0] matmul_29_out_page_dma_offset;
  wire [31:0] matmul_29_out_ram_select;
  wire [31:0] matmul_29_out_row_count;
  wire [31:0] matmul_29_prev_bat_count;
  wire [31:0] matmul_29_prev_och_count;
  wire [31:0] matmul_29_prev_row_count;
  wire matmul_29_prev_row_select;
  wire [31:0] matmul_29_row_count;
  wire [31:0] matmul_29_row_count_buf;
  wire matmul_29_row_select;
  wire matmul_29_row_select_buf;
  wire matmul_29_skip_comp;
  wire matmul_29_skip_read_act;
  wire matmul_29_skip_read_filter;
  wire matmul_29_skip_write_out;
  wire [31:0] matmul_29_stream_act_local_0;
  wire [31:0] matmul_29_stream_out_local;
  wire [31:0] matmul_29_stream_out_local_col;
  wire [31:0] matmul_29_stream_out_local_val;
  wire matmul_29_stream_pad_mask_0_0;
  wire matmul_29_stream_pad_masks;
  wire [31:0] matmul_29_sync_comp_count;
  wire [31:0] matmul_29_sync_out_count;
  wire matmul_29_update_act;
  wire matmul_29_update_filter;
  wire [31:0] max_pool_serial_18_act_base_offset;
  wire [31:0] max_pool_serial_18_act_base_offset_bat;
  wire [31:0] max_pool_serial_18_act_base_offset_row;
  wire max_pool_serial_18_act_page;
  wire [31:0] max_pool_serial_18_act_page_comp_offset;
  wire [31:0] max_pool_serial_18_act_page_comp_offset_buf;
  wire [31:0] max_pool_serial_18_act_page_dma_offset;
  wire [31:0] max_pool_serial_18_arg_objaddr_0;
  wire [31:0] max_pool_serial_18_bat_count;
  wire [31:0] max_pool_serial_18_col_count;
  wire [31:0] max_pool_serial_18_comp_count;
  wire [31:0] max_pool_serial_18_comp_fsm;
  wire [1:0] max_pool_serial_18_control_param_index;
  wire max_pool_serial_18_dma_pad_mask_0;
  wire max_pool_serial_18_dma_pad_mask_1;
  wire [31:0] max_pool_serial_18_objaddr;
  wire [31:0] max_pool_serial_18_out_base_offset;
  wire [31:0] max_pool_serial_18_out_base_offset_bat;
  wire [31:0] max_pool_serial_18_out_base_offset_row;
  wire [31:0] max_pool_serial_18_out_count;
  wire max_pool_serial_18_out_page;
  wire [31:0] max_pool_serial_18_out_page_comp_offset;
  wire [31:0] max_pool_serial_18_out_page_comp_offset_buf;
  wire [31:0] max_pool_serial_18_out_page_dma_offset;
  wire [31:0] max_pool_serial_18_prev_bat_count;
  wire [31:0] max_pool_serial_18_prev_row_count;
  wire [31:0] max_pool_serial_18_row_count;
  wire [31:0] max_pool_serial_18_row_count_buf;
  wire max_pool_serial_18_skip_comp;
  wire max_pool_serial_18_skip_read_act;
  wire max_pool_serial_18_skip_write_out;
  wire [31:0] max_pool_serial_18_stream_act_local;
  wire [31:0] max_pool_serial_18_stream_out_local;
  wire max_pool_serial_18_stream_pad_mask_0_0;
  wire max_pool_serial_18_stream_pad_mask_0_1;
  wire max_pool_serial_18_stream_pad_mask_1_0;
  wire max_pool_serial_18_stream_pad_mask_1_1;
  wire [3:0] max_pool_serial_18_stream_pad_masks;
  wire [3:0] mul_10_rshift_data;
  wire [7:0] mul_10_x_data;
  wire [3:0] mul_10_y_data;
  wire [11:0] mul_10_z_data;
  wire [3:0] mul_11_rshift_data;
  wire [7:0] mul_11_x_data;
  wire [3:0] mul_11_y_data;
  wire [11:0] mul_11_z_data;
  wire [3:0] mul_12_rshift_data;
  wire [7:0] mul_12_x_data;
  wire [3:0] mul_12_y_data;
  wire [11:0] mul_12_z_data;
  wire [3:0] mul_4_rshift_data;
  wire [7:0] mul_4_x_data;
  wire [3:0] mul_4_y_data;
  wire [11:0] mul_4_z_data;
  wire [3:0] mul_5_rshift_data;
  wire [7:0] mul_5_x_data;
  wire [3:0] mul_5_y_data;
  wire [11:0] mul_5_z_data;
  wire [3:0] mul_6_rshift_data;
  wire [7:0] mul_6_x_data;
  wire [3:0] mul_6_y_data;
  wire [11:0] mul_6_z_data;
  wire [3:0] mul_7_rshift_data;
  wire [7:0] mul_7_x_data;
  wire [3:0] mul_7_y_data;
  wire [11:0] mul_7_z_data;
  wire [3:0] mul_8_rshift_data;
  wire [7:0] mul_8_x_data;
  wire [3:0] mul_8_y_data;
  wire [11:0] mul_8_z_data;
  wire [3:0] mul_9_rshift_data;
  wire [7:0] mul_9_x_data;
  wire [3:0] mul_9_y_data;
  wire [11:0] mul_9_z_data;
  wire [5:0] mul_rshift_clip_3_rshift_data;
  wire [31:0] mul_rshift_clip_3_x_data;
  wire [7:0] mul_rshift_clip_3_y_data;
  wire [7:0] mul_rshift_clip_3_z_data;
  wire [9:0] ram_w4_l8192_id0_0_0_addr;
  wire [3:0] ram_w4_l8192_id0_0_0_rdata;
  wire [3:0] ram_w4_l8192_id0_0_0_wdata;
  wire ram_w4_l8192_id0_0_0_wenable;
  wire [9:0] ram_w4_l8192_id0_0_1_addr;
  wire [3:0] ram_w4_l8192_id0_0_1_rdata;
  wire [3:0] ram_w4_l8192_id0_0_1_wdata;
  wire ram_w4_l8192_id0_0_1_wenable;
  wire [9:0] ram_w4_l8192_id0_1_0_addr;
  wire [3:0] ram_w4_l8192_id0_1_0_rdata;
  wire [3:0] ram_w4_l8192_id0_1_0_wdata;
  wire ram_w4_l8192_id0_1_0_wenable;
  wire [9:0] ram_w4_l8192_id0_1_1_addr;
  wire [3:0] ram_w4_l8192_id0_1_1_rdata;
  wire [3:0] ram_w4_l8192_id0_1_1_wdata;
  wire ram_w4_l8192_id0_1_1_wenable;
  wire [9:0] ram_w4_l8192_id0_2_0_addr;
  wire [3:0] ram_w4_l8192_id0_2_0_rdata;
  wire [3:0] ram_w4_l8192_id0_2_0_wdata;
  wire ram_w4_l8192_id0_2_0_wenable;
  wire [9:0] ram_w4_l8192_id0_2_1_addr;
  wire [3:0] ram_w4_l8192_id0_2_1_rdata;
  wire [3:0] ram_w4_l8192_id0_2_1_wdata;
  wire ram_w4_l8192_id0_2_1_wenable;
  wire [9:0] ram_w4_l8192_id0_3_0_addr;
  wire [3:0] ram_w4_l8192_id0_3_0_rdata;
  wire [3:0] ram_w4_l8192_id0_3_0_wdata;
  wire ram_w4_l8192_id0_3_0_wenable;
  wire [9:0] ram_w4_l8192_id0_3_1_addr;
  wire [3:0] ram_w4_l8192_id0_3_1_rdata;
  wire [3:0] ram_w4_l8192_id0_3_1_wdata;
  wire ram_w4_l8192_id0_3_1_wenable;
  wire [9:0] ram_w4_l8192_id0_4_0_addr;
  wire [3:0] ram_w4_l8192_id0_4_0_rdata;
  wire [3:0] ram_w4_l8192_id0_4_0_wdata;
  wire ram_w4_l8192_id0_4_0_wenable;
  wire [9:0] ram_w4_l8192_id0_4_1_addr;
  wire [3:0] ram_w4_l8192_id0_4_1_rdata;
  wire [3:0] ram_w4_l8192_id0_4_1_wdata;
  wire ram_w4_l8192_id0_4_1_wenable;
  wire [9:0] ram_w4_l8192_id0_5_0_addr;
  wire [3:0] ram_w4_l8192_id0_5_0_rdata;
  wire [3:0] ram_w4_l8192_id0_5_0_wdata;
  wire ram_w4_l8192_id0_5_0_wenable;
  wire [9:0] ram_w4_l8192_id0_5_1_addr;
  wire [3:0] ram_w4_l8192_id0_5_1_rdata;
  wire [3:0] ram_w4_l8192_id0_5_1_wdata;
  wire ram_w4_l8192_id0_5_1_wenable;
  wire [9:0] ram_w4_l8192_id0_6_0_addr;
  wire [3:0] ram_w4_l8192_id0_6_0_rdata;
  wire [3:0] ram_w4_l8192_id0_6_0_wdata;
  wire ram_w4_l8192_id0_6_0_wenable;
  wire [9:0] ram_w4_l8192_id0_6_1_addr;
  wire [3:0] ram_w4_l8192_id0_6_1_rdata;
  wire [3:0] ram_w4_l8192_id0_6_1_wdata;
  wire ram_w4_l8192_id0_6_1_wenable;
  wire [9:0] ram_w4_l8192_id0_7_0_addr;
  wire [3:0] ram_w4_l8192_id0_7_0_rdata;
  wire [3:0] ram_w4_l8192_id0_7_0_wdata;
  wire ram_w4_l8192_id0_7_0_wenable;
  wire [9:0] ram_w4_l8192_id0_7_1_addr;
  wire [3:0] ram_w4_l8192_id0_7_1_rdata;
  wire [3:0] ram_w4_l8192_id0_7_1_wdata;
  wire ram_w4_l8192_id0_7_1_wenable;
  wire [9:0] ram_w4_l8192_id1_0_0_addr;
  wire [3:0] ram_w4_l8192_id1_0_0_rdata;
  wire [3:0] ram_w4_l8192_id1_0_0_wdata;
  wire ram_w4_l8192_id1_0_0_wenable;
  wire [9:0] ram_w4_l8192_id1_0_1_addr;
  wire [3:0] ram_w4_l8192_id1_0_1_rdata;
  wire [3:0] ram_w4_l8192_id1_0_1_wdata;
  wire ram_w4_l8192_id1_0_1_wenable;
  wire [9:0] ram_w4_l8192_id1_1_0_addr;
  wire [3:0] ram_w4_l8192_id1_1_0_rdata;
  wire [3:0] ram_w4_l8192_id1_1_0_wdata;
  wire ram_w4_l8192_id1_1_0_wenable;
  wire [9:0] ram_w4_l8192_id1_1_1_addr;
  wire [3:0] ram_w4_l8192_id1_1_1_rdata;
  wire [3:0] ram_w4_l8192_id1_1_1_wdata;
  wire ram_w4_l8192_id1_1_1_wenable;
  wire [9:0] ram_w4_l8192_id1_2_0_addr;
  wire [3:0] ram_w4_l8192_id1_2_0_rdata;
  wire [3:0] ram_w4_l8192_id1_2_0_wdata;
  wire ram_w4_l8192_id1_2_0_wenable;
  wire [9:0] ram_w4_l8192_id1_2_1_addr;
  wire [3:0] ram_w4_l8192_id1_2_1_rdata;
  wire [3:0] ram_w4_l8192_id1_2_1_wdata;
  wire ram_w4_l8192_id1_2_1_wenable;
  wire [9:0] ram_w4_l8192_id1_3_0_addr;
  wire [3:0] ram_w4_l8192_id1_3_0_rdata;
  wire [3:0] ram_w4_l8192_id1_3_0_wdata;
  wire ram_w4_l8192_id1_3_0_wenable;
  wire [9:0] ram_w4_l8192_id1_3_1_addr;
  wire [3:0] ram_w4_l8192_id1_3_1_rdata;
  wire [3:0] ram_w4_l8192_id1_3_1_wdata;
  wire ram_w4_l8192_id1_3_1_wenable;
  wire [9:0] ram_w4_l8192_id1_4_0_addr;
  wire [3:0] ram_w4_l8192_id1_4_0_rdata;
  wire [3:0] ram_w4_l8192_id1_4_0_wdata;
  wire ram_w4_l8192_id1_4_0_wenable;
  wire [9:0] ram_w4_l8192_id1_4_1_addr;
  wire [3:0] ram_w4_l8192_id1_4_1_rdata;
  wire [3:0] ram_w4_l8192_id1_4_1_wdata;
  wire ram_w4_l8192_id1_4_1_wenable;
  wire [9:0] ram_w4_l8192_id1_5_0_addr;
  wire [3:0] ram_w4_l8192_id1_5_0_rdata;
  wire [3:0] ram_w4_l8192_id1_5_0_wdata;
  wire ram_w4_l8192_id1_5_0_wenable;
  wire [9:0] ram_w4_l8192_id1_5_1_addr;
  wire [3:0] ram_w4_l8192_id1_5_1_rdata;
  wire [3:0] ram_w4_l8192_id1_5_1_wdata;
  wire ram_w4_l8192_id1_5_1_wenable;
  wire [9:0] ram_w4_l8192_id1_6_0_addr;
  wire [3:0] ram_w4_l8192_id1_6_0_rdata;
  wire [3:0] ram_w4_l8192_id1_6_0_wdata;
  wire ram_w4_l8192_id1_6_0_wenable;
  wire [9:0] ram_w4_l8192_id1_6_1_addr;
  wire [3:0] ram_w4_l8192_id1_6_1_rdata;
  wire [3:0] ram_w4_l8192_id1_6_1_wdata;
  wire ram_w4_l8192_id1_6_1_wenable;
  wire [9:0] ram_w4_l8192_id1_7_0_addr;
  wire [3:0] ram_w4_l8192_id1_7_0_rdata;
  wire [3:0] ram_w4_l8192_id1_7_0_wdata;
  wire ram_w4_l8192_id1_7_0_wenable;
  wire [9:0] ram_w4_l8192_id1_7_1_addr;
  wire [3:0] ram_w4_l8192_id1_7_1_rdata;
  wire [3:0] ram_w4_l8192_id1_7_1_wdata;
  wire ram_w4_l8192_id1_7_1_wenable;
  wire [9:0] ram_w4_l8192_id2_0_0_addr;
  wire [3:0] ram_w4_l8192_id2_0_0_rdata;
  wire [3:0] ram_w4_l8192_id2_0_0_wdata;
  wire ram_w4_l8192_id2_0_0_wenable;
  wire [9:0] ram_w4_l8192_id2_0_1_addr;
  wire [3:0] ram_w4_l8192_id2_0_1_rdata;
  wire [3:0] ram_w4_l8192_id2_0_1_wdata;
  wire ram_w4_l8192_id2_0_1_wenable;
  wire [9:0] ram_w4_l8192_id2_1_0_addr;
  wire [3:0] ram_w4_l8192_id2_1_0_rdata;
  wire [3:0] ram_w4_l8192_id2_1_0_wdata;
  wire ram_w4_l8192_id2_1_0_wenable;
  wire [9:0] ram_w4_l8192_id2_1_1_addr;
  wire [3:0] ram_w4_l8192_id2_1_1_rdata;
  wire [3:0] ram_w4_l8192_id2_1_1_wdata;
  wire ram_w4_l8192_id2_1_1_wenable;
  wire [9:0] ram_w4_l8192_id2_2_0_addr;
  wire [3:0] ram_w4_l8192_id2_2_0_rdata;
  wire [3:0] ram_w4_l8192_id2_2_0_wdata;
  wire ram_w4_l8192_id2_2_0_wenable;
  wire [9:0] ram_w4_l8192_id2_2_1_addr;
  wire [3:0] ram_w4_l8192_id2_2_1_rdata;
  wire [3:0] ram_w4_l8192_id2_2_1_wdata;
  wire ram_w4_l8192_id2_2_1_wenable;
  wire [9:0] ram_w4_l8192_id2_3_0_addr;
  wire [3:0] ram_w4_l8192_id2_3_0_rdata;
  wire [3:0] ram_w4_l8192_id2_3_0_wdata;
  wire ram_w4_l8192_id2_3_0_wenable;
  wire [9:0] ram_w4_l8192_id2_3_1_addr;
  wire [3:0] ram_w4_l8192_id2_3_1_rdata;
  wire [3:0] ram_w4_l8192_id2_3_1_wdata;
  wire ram_w4_l8192_id2_3_1_wenable;
  wire [9:0] ram_w4_l8192_id2_4_0_addr;
  wire [3:0] ram_w4_l8192_id2_4_0_rdata;
  wire [3:0] ram_w4_l8192_id2_4_0_wdata;
  wire ram_w4_l8192_id2_4_0_wenable;
  wire [9:0] ram_w4_l8192_id2_4_1_addr;
  wire [3:0] ram_w4_l8192_id2_4_1_rdata;
  wire [3:0] ram_w4_l8192_id2_4_1_wdata;
  wire ram_w4_l8192_id2_4_1_wenable;
  wire [9:0] ram_w4_l8192_id2_5_0_addr;
  wire [3:0] ram_w4_l8192_id2_5_0_rdata;
  wire [3:0] ram_w4_l8192_id2_5_0_wdata;
  wire ram_w4_l8192_id2_5_0_wenable;
  wire [9:0] ram_w4_l8192_id2_5_1_addr;
  wire [3:0] ram_w4_l8192_id2_5_1_rdata;
  wire [3:0] ram_w4_l8192_id2_5_1_wdata;
  wire ram_w4_l8192_id2_5_1_wenable;
  wire [9:0] ram_w4_l8192_id2_6_0_addr;
  wire [3:0] ram_w4_l8192_id2_6_0_rdata;
  wire [3:0] ram_w4_l8192_id2_6_0_wdata;
  wire ram_w4_l8192_id2_6_0_wenable;
  wire [9:0] ram_w4_l8192_id2_6_1_addr;
  wire [3:0] ram_w4_l8192_id2_6_1_rdata;
  wire [3:0] ram_w4_l8192_id2_6_1_wdata;
  wire ram_w4_l8192_id2_6_1_wenable;
  wire [9:0] ram_w4_l8192_id2_7_0_addr;
  wire [3:0] ram_w4_l8192_id2_7_0_rdata;
  wire [3:0] ram_w4_l8192_id2_7_0_wdata;
  wire ram_w4_l8192_id2_7_0_wenable;
  wire [9:0] ram_w4_l8192_id2_7_1_addr;
  wire [3:0] ram_w4_l8192_id2_7_1_rdata;
  wire [3:0] ram_w4_l8192_id2_7_1_wdata;
  wire ram_w4_l8192_id2_7_1_wenable;
  wire [9:0] ram_w4_l8192_id3_0_0_addr;
  wire [3:0] ram_w4_l8192_id3_0_0_rdata;
  wire [3:0] ram_w4_l8192_id3_0_0_wdata;
  wire ram_w4_l8192_id3_0_0_wenable;
  wire [9:0] ram_w4_l8192_id3_0_1_addr;
  wire [3:0] ram_w4_l8192_id3_0_1_rdata;
  wire [3:0] ram_w4_l8192_id3_0_1_wdata;
  wire ram_w4_l8192_id3_0_1_wenable;
  wire [9:0] ram_w4_l8192_id3_1_0_addr;
  wire [3:0] ram_w4_l8192_id3_1_0_rdata;
  wire [3:0] ram_w4_l8192_id3_1_0_wdata;
  wire ram_w4_l8192_id3_1_0_wenable;
  wire [9:0] ram_w4_l8192_id3_1_1_addr;
  wire [3:0] ram_w4_l8192_id3_1_1_rdata;
  wire [3:0] ram_w4_l8192_id3_1_1_wdata;
  wire ram_w4_l8192_id3_1_1_wenable;
  wire [9:0] ram_w4_l8192_id3_2_0_addr;
  wire [3:0] ram_w4_l8192_id3_2_0_rdata;
  wire [3:0] ram_w4_l8192_id3_2_0_wdata;
  wire ram_w4_l8192_id3_2_0_wenable;
  wire [9:0] ram_w4_l8192_id3_2_1_addr;
  wire [3:0] ram_w4_l8192_id3_2_1_rdata;
  wire [3:0] ram_w4_l8192_id3_2_1_wdata;
  wire ram_w4_l8192_id3_2_1_wenable;
  wire [9:0] ram_w4_l8192_id3_3_0_addr;
  wire [3:0] ram_w4_l8192_id3_3_0_rdata;
  wire [3:0] ram_w4_l8192_id3_3_0_wdata;
  wire ram_w4_l8192_id3_3_0_wenable;
  wire [9:0] ram_w4_l8192_id3_3_1_addr;
  wire [3:0] ram_w4_l8192_id3_3_1_rdata;
  wire [3:0] ram_w4_l8192_id3_3_1_wdata;
  wire ram_w4_l8192_id3_3_1_wenable;
  wire [9:0] ram_w4_l8192_id3_4_0_addr;
  wire [3:0] ram_w4_l8192_id3_4_0_rdata;
  wire [3:0] ram_w4_l8192_id3_4_0_wdata;
  wire ram_w4_l8192_id3_4_0_wenable;
  wire [9:0] ram_w4_l8192_id3_4_1_addr;
  wire [3:0] ram_w4_l8192_id3_4_1_rdata;
  wire [3:0] ram_w4_l8192_id3_4_1_wdata;
  wire ram_w4_l8192_id3_4_1_wenable;
  wire [9:0] ram_w4_l8192_id3_5_0_addr;
  wire [3:0] ram_w4_l8192_id3_5_0_rdata;
  wire [3:0] ram_w4_l8192_id3_5_0_wdata;
  wire ram_w4_l8192_id3_5_0_wenable;
  wire [9:0] ram_w4_l8192_id3_5_1_addr;
  wire [3:0] ram_w4_l8192_id3_5_1_rdata;
  wire [3:0] ram_w4_l8192_id3_5_1_wdata;
  wire ram_w4_l8192_id3_5_1_wenable;
  wire [9:0] ram_w4_l8192_id3_6_0_addr;
  wire [3:0] ram_w4_l8192_id3_6_0_rdata;
  wire [3:0] ram_w4_l8192_id3_6_0_wdata;
  wire ram_w4_l8192_id3_6_0_wenable;
  wire [9:0] ram_w4_l8192_id3_6_1_addr;
  wire [3:0] ram_w4_l8192_id3_6_1_rdata;
  wire [3:0] ram_w4_l8192_id3_6_1_wdata;
  wire ram_w4_l8192_id3_6_1_wenable;
  wire [9:0] ram_w4_l8192_id3_7_0_addr;
  wire [3:0] ram_w4_l8192_id3_7_0_rdata;
  wire [3:0] ram_w4_l8192_id3_7_0_wdata;
  wire ram_w4_l8192_id3_7_0_wenable;
  wire [9:0] ram_w4_l8192_id3_7_1_addr;
  wire [3:0] ram_w4_l8192_id3_7_1_rdata;
  wire [3:0] ram_w4_l8192_id3_7_1_wdata;
  wire ram_w4_l8192_id3_7_1_wenable;
  wire [9:0] ram_w4_l8192_id4_0_0_addr;
  wire [3:0] ram_w4_l8192_id4_0_0_rdata;
  wire [3:0] ram_w4_l8192_id4_0_0_wdata;
  wire ram_w4_l8192_id4_0_0_wenable;
  wire [9:0] ram_w4_l8192_id4_0_1_addr;
  wire [3:0] ram_w4_l8192_id4_0_1_rdata;
  wire [3:0] ram_w4_l8192_id4_0_1_wdata;
  wire ram_w4_l8192_id4_0_1_wenable;
  wire [9:0] ram_w4_l8192_id4_1_0_addr;
  wire [3:0] ram_w4_l8192_id4_1_0_rdata;
  wire [3:0] ram_w4_l8192_id4_1_0_wdata;
  wire ram_w4_l8192_id4_1_0_wenable;
  wire [9:0] ram_w4_l8192_id4_1_1_addr;
  wire [3:0] ram_w4_l8192_id4_1_1_rdata;
  wire [3:0] ram_w4_l8192_id4_1_1_wdata;
  wire ram_w4_l8192_id4_1_1_wenable;
  wire [9:0] ram_w4_l8192_id4_2_0_addr;
  wire [3:0] ram_w4_l8192_id4_2_0_rdata;
  wire [3:0] ram_w4_l8192_id4_2_0_wdata;
  wire ram_w4_l8192_id4_2_0_wenable;
  wire [9:0] ram_w4_l8192_id4_2_1_addr;
  wire [3:0] ram_w4_l8192_id4_2_1_rdata;
  wire [3:0] ram_w4_l8192_id4_2_1_wdata;
  wire ram_w4_l8192_id4_2_1_wenable;
  wire [9:0] ram_w4_l8192_id4_3_0_addr;
  wire [3:0] ram_w4_l8192_id4_3_0_rdata;
  wire [3:0] ram_w4_l8192_id4_3_0_wdata;
  wire ram_w4_l8192_id4_3_0_wenable;
  wire [9:0] ram_w4_l8192_id4_3_1_addr;
  wire [3:0] ram_w4_l8192_id4_3_1_rdata;
  wire [3:0] ram_w4_l8192_id4_3_1_wdata;
  wire ram_w4_l8192_id4_3_1_wenable;
  wire [9:0] ram_w4_l8192_id4_4_0_addr;
  wire [3:0] ram_w4_l8192_id4_4_0_rdata;
  wire [3:0] ram_w4_l8192_id4_4_0_wdata;
  wire ram_w4_l8192_id4_4_0_wenable;
  wire [9:0] ram_w4_l8192_id4_4_1_addr;
  wire [3:0] ram_w4_l8192_id4_4_1_rdata;
  wire [3:0] ram_w4_l8192_id4_4_1_wdata;
  wire ram_w4_l8192_id4_4_1_wenable;
  wire [9:0] ram_w4_l8192_id4_5_0_addr;
  wire [3:0] ram_w4_l8192_id4_5_0_rdata;
  wire [3:0] ram_w4_l8192_id4_5_0_wdata;
  wire ram_w4_l8192_id4_5_0_wenable;
  wire [9:0] ram_w4_l8192_id4_5_1_addr;
  wire [3:0] ram_w4_l8192_id4_5_1_rdata;
  wire [3:0] ram_w4_l8192_id4_5_1_wdata;
  wire ram_w4_l8192_id4_5_1_wenable;
  wire [9:0] ram_w4_l8192_id4_6_0_addr;
  wire [3:0] ram_w4_l8192_id4_6_0_rdata;
  wire [3:0] ram_w4_l8192_id4_6_0_wdata;
  wire ram_w4_l8192_id4_6_0_wenable;
  wire [9:0] ram_w4_l8192_id4_6_1_addr;
  wire [3:0] ram_w4_l8192_id4_6_1_rdata;
  wire [3:0] ram_w4_l8192_id4_6_1_wdata;
  wire ram_w4_l8192_id4_6_1_wenable;
  wire [9:0] ram_w4_l8192_id4_7_0_addr;
  wire [3:0] ram_w4_l8192_id4_7_0_rdata;
  wire [3:0] ram_w4_l8192_id4_7_0_wdata;
  wire ram_w4_l8192_id4_7_0_wenable;
  wire [9:0] ram_w4_l8192_id4_7_1_addr;
  wire [3:0] ram_w4_l8192_id4_7_1_rdata;
  wire [3:0] ram_w4_l8192_id4_7_1_wdata;
  wire ram_w4_l8192_id4_7_1_wenable;
  wire [9:0] ram_w4_l8192_id5_0_0_addr;
  wire [3:0] ram_w4_l8192_id5_0_0_rdata;
  wire [3:0] ram_w4_l8192_id5_0_0_wdata;
  wire ram_w4_l8192_id5_0_0_wenable;
  wire [9:0] ram_w4_l8192_id5_0_1_addr;
  wire [3:0] ram_w4_l8192_id5_0_1_rdata;
  wire [3:0] ram_w4_l8192_id5_0_1_wdata;
  wire ram_w4_l8192_id5_0_1_wenable;
  wire [9:0] ram_w4_l8192_id5_1_0_addr;
  wire [3:0] ram_w4_l8192_id5_1_0_rdata;
  wire [3:0] ram_w4_l8192_id5_1_0_wdata;
  wire ram_w4_l8192_id5_1_0_wenable;
  wire [9:0] ram_w4_l8192_id5_1_1_addr;
  wire [3:0] ram_w4_l8192_id5_1_1_rdata;
  wire [3:0] ram_w4_l8192_id5_1_1_wdata;
  wire ram_w4_l8192_id5_1_1_wenable;
  wire [9:0] ram_w4_l8192_id5_2_0_addr;
  wire [3:0] ram_w4_l8192_id5_2_0_rdata;
  wire [3:0] ram_w4_l8192_id5_2_0_wdata;
  wire ram_w4_l8192_id5_2_0_wenable;
  wire [9:0] ram_w4_l8192_id5_2_1_addr;
  wire [3:0] ram_w4_l8192_id5_2_1_rdata;
  wire [3:0] ram_w4_l8192_id5_2_1_wdata;
  wire ram_w4_l8192_id5_2_1_wenable;
  wire [9:0] ram_w4_l8192_id5_3_0_addr;
  wire [3:0] ram_w4_l8192_id5_3_0_rdata;
  wire [3:0] ram_w4_l8192_id5_3_0_wdata;
  wire ram_w4_l8192_id5_3_0_wenable;
  wire [9:0] ram_w4_l8192_id5_3_1_addr;
  wire [3:0] ram_w4_l8192_id5_3_1_rdata;
  wire [3:0] ram_w4_l8192_id5_3_1_wdata;
  wire ram_w4_l8192_id5_3_1_wenable;
  wire [9:0] ram_w4_l8192_id5_4_0_addr;
  wire [3:0] ram_w4_l8192_id5_4_0_rdata;
  wire [3:0] ram_w4_l8192_id5_4_0_wdata;
  wire ram_w4_l8192_id5_4_0_wenable;
  wire [9:0] ram_w4_l8192_id5_4_1_addr;
  wire [3:0] ram_w4_l8192_id5_4_1_rdata;
  wire [3:0] ram_w4_l8192_id5_4_1_wdata;
  wire ram_w4_l8192_id5_4_1_wenable;
  wire [9:0] ram_w4_l8192_id5_5_0_addr;
  wire [3:0] ram_w4_l8192_id5_5_0_rdata;
  wire [3:0] ram_w4_l8192_id5_5_0_wdata;
  wire ram_w4_l8192_id5_5_0_wenable;
  wire [9:0] ram_w4_l8192_id5_5_1_addr;
  wire [3:0] ram_w4_l8192_id5_5_1_rdata;
  wire [3:0] ram_w4_l8192_id5_5_1_wdata;
  wire ram_w4_l8192_id5_5_1_wenable;
  wire [9:0] ram_w4_l8192_id5_6_0_addr;
  wire [3:0] ram_w4_l8192_id5_6_0_rdata;
  wire [3:0] ram_w4_l8192_id5_6_0_wdata;
  wire ram_w4_l8192_id5_6_0_wenable;
  wire [9:0] ram_w4_l8192_id5_6_1_addr;
  wire [3:0] ram_w4_l8192_id5_6_1_rdata;
  wire [3:0] ram_w4_l8192_id5_6_1_wdata;
  wire ram_w4_l8192_id5_6_1_wenable;
  wire [9:0] ram_w4_l8192_id5_7_0_addr;
  wire [3:0] ram_w4_l8192_id5_7_0_rdata;
  wire [3:0] ram_w4_l8192_id5_7_0_wdata;
  wire ram_w4_l8192_id5_7_0_wenable;
  wire [9:0] ram_w4_l8192_id5_7_1_addr;
  wire [3:0] ram_w4_l8192_id5_7_1_rdata;
  wire [3:0] ram_w4_l8192_id5_7_1_wdata;
  wire ram_w4_l8192_id5_7_1_wenable;
  wire [9:0] ram_w4_l8192_id6_0_0_addr;
  wire [3:0] ram_w4_l8192_id6_0_0_rdata;
  wire [3:0] ram_w4_l8192_id6_0_0_wdata;
  wire ram_w4_l8192_id6_0_0_wenable;
  wire [9:0] ram_w4_l8192_id6_0_1_addr;
  wire [3:0] ram_w4_l8192_id6_0_1_rdata;
  wire [3:0] ram_w4_l8192_id6_0_1_wdata;
  wire ram_w4_l8192_id6_0_1_wenable;
  wire [9:0] ram_w4_l8192_id6_1_0_addr;
  wire [3:0] ram_w4_l8192_id6_1_0_rdata;
  wire [3:0] ram_w4_l8192_id6_1_0_wdata;
  wire ram_w4_l8192_id6_1_0_wenable;
  wire [9:0] ram_w4_l8192_id6_1_1_addr;
  wire [3:0] ram_w4_l8192_id6_1_1_rdata;
  wire [3:0] ram_w4_l8192_id6_1_1_wdata;
  wire ram_w4_l8192_id6_1_1_wenable;
  wire [9:0] ram_w4_l8192_id6_2_0_addr;
  wire [3:0] ram_w4_l8192_id6_2_0_rdata;
  wire [3:0] ram_w4_l8192_id6_2_0_wdata;
  wire ram_w4_l8192_id6_2_0_wenable;
  wire [9:0] ram_w4_l8192_id6_2_1_addr;
  wire [3:0] ram_w4_l8192_id6_2_1_rdata;
  wire [3:0] ram_w4_l8192_id6_2_1_wdata;
  wire ram_w4_l8192_id6_2_1_wenable;
  wire [9:0] ram_w4_l8192_id6_3_0_addr;
  wire [3:0] ram_w4_l8192_id6_3_0_rdata;
  wire [3:0] ram_w4_l8192_id6_3_0_wdata;
  wire ram_w4_l8192_id6_3_0_wenable;
  wire [9:0] ram_w4_l8192_id6_3_1_addr;
  wire [3:0] ram_w4_l8192_id6_3_1_rdata;
  wire [3:0] ram_w4_l8192_id6_3_1_wdata;
  wire ram_w4_l8192_id6_3_1_wenable;
  wire [9:0] ram_w4_l8192_id6_4_0_addr;
  wire [3:0] ram_w4_l8192_id6_4_0_rdata;
  wire [3:0] ram_w4_l8192_id6_4_0_wdata;
  wire ram_w4_l8192_id6_4_0_wenable;
  wire [9:0] ram_w4_l8192_id6_4_1_addr;
  wire [3:0] ram_w4_l8192_id6_4_1_rdata;
  wire [3:0] ram_w4_l8192_id6_4_1_wdata;
  wire ram_w4_l8192_id6_4_1_wenable;
  wire [9:0] ram_w4_l8192_id6_5_0_addr;
  wire [3:0] ram_w4_l8192_id6_5_0_rdata;
  wire [3:0] ram_w4_l8192_id6_5_0_wdata;
  wire ram_w4_l8192_id6_5_0_wenable;
  wire [9:0] ram_w4_l8192_id6_5_1_addr;
  wire [3:0] ram_w4_l8192_id6_5_1_rdata;
  wire [3:0] ram_w4_l8192_id6_5_1_wdata;
  wire ram_w4_l8192_id6_5_1_wenable;
  wire [9:0] ram_w4_l8192_id6_6_0_addr;
  wire [3:0] ram_w4_l8192_id6_6_0_rdata;
  wire [3:0] ram_w4_l8192_id6_6_0_wdata;
  wire ram_w4_l8192_id6_6_0_wenable;
  wire [9:0] ram_w4_l8192_id6_6_1_addr;
  wire [3:0] ram_w4_l8192_id6_6_1_rdata;
  wire [3:0] ram_w4_l8192_id6_6_1_wdata;
  wire ram_w4_l8192_id6_6_1_wenable;
  wire [9:0] ram_w4_l8192_id6_7_0_addr;
  wire [3:0] ram_w4_l8192_id6_7_0_rdata;
  wire [3:0] ram_w4_l8192_id6_7_0_wdata;
  wire ram_w4_l8192_id6_7_0_wenable;
  wire [9:0] ram_w4_l8192_id6_7_1_addr;
  wire [3:0] ram_w4_l8192_id6_7_1_rdata;
  wire [3:0] ram_w4_l8192_id6_7_1_wdata;
  wire ram_w4_l8192_id6_7_1_wenable;
  wire [9:0] ram_w4_l8192_id7_0_0_addr;
  wire [3:0] ram_w4_l8192_id7_0_0_rdata;
  wire [3:0] ram_w4_l8192_id7_0_0_wdata;
  wire ram_w4_l8192_id7_0_0_wenable;
  wire [9:0] ram_w4_l8192_id7_0_1_addr;
  wire [3:0] ram_w4_l8192_id7_0_1_rdata;
  wire [3:0] ram_w4_l8192_id7_0_1_wdata;
  wire ram_w4_l8192_id7_0_1_wenable;
  wire [9:0] ram_w4_l8192_id7_1_0_addr;
  wire [3:0] ram_w4_l8192_id7_1_0_rdata;
  wire [3:0] ram_w4_l8192_id7_1_0_wdata;
  wire ram_w4_l8192_id7_1_0_wenable;
  wire [9:0] ram_w4_l8192_id7_1_1_addr;
  wire [3:0] ram_w4_l8192_id7_1_1_rdata;
  wire [3:0] ram_w4_l8192_id7_1_1_wdata;
  wire ram_w4_l8192_id7_1_1_wenable;
  wire [9:0] ram_w4_l8192_id7_2_0_addr;
  wire [3:0] ram_w4_l8192_id7_2_0_rdata;
  wire [3:0] ram_w4_l8192_id7_2_0_wdata;
  wire ram_w4_l8192_id7_2_0_wenable;
  wire [9:0] ram_w4_l8192_id7_2_1_addr;
  wire [3:0] ram_w4_l8192_id7_2_1_rdata;
  wire [3:0] ram_w4_l8192_id7_2_1_wdata;
  wire ram_w4_l8192_id7_2_1_wenable;
  wire [9:0] ram_w4_l8192_id7_3_0_addr;
  wire [3:0] ram_w4_l8192_id7_3_0_rdata;
  wire [3:0] ram_w4_l8192_id7_3_0_wdata;
  wire ram_w4_l8192_id7_3_0_wenable;
  wire [9:0] ram_w4_l8192_id7_3_1_addr;
  wire [3:0] ram_w4_l8192_id7_3_1_rdata;
  wire [3:0] ram_w4_l8192_id7_3_1_wdata;
  wire ram_w4_l8192_id7_3_1_wenable;
  wire [9:0] ram_w4_l8192_id7_4_0_addr;
  wire [3:0] ram_w4_l8192_id7_4_0_rdata;
  wire [3:0] ram_w4_l8192_id7_4_0_wdata;
  wire ram_w4_l8192_id7_4_0_wenable;
  wire [9:0] ram_w4_l8192_id7_4_1_addr;
  wire [3:0] ram_w4_l8192_id7_4_1_rdata;
  wire [3:0] ram_w4_l8192_id7_4_1_wdata;
  wire ram_w4_l8192_id7_4_1_wenable;
  wire [9:0] ram_w4_l8192_id7_5_0_addr;
  wire [3:0] ram_w4_l8192_id7_5_0_rdata;
  wire [3:0] ram_w4_l8192_id7_5_0_wdata;
  wire ram_w4_l8192_id7_5_0_wenable;
  wire [9:0] ram_w4_l8192_id7_5_1_addr;
  wire [3:0] ram_w4_l8192_id7_5_1_rdata;
  wire [3:0] ram_w4_l8192_id7_5_1_wdata;
  wire ram_w4_l8192_id7_5_1_wenable;
  wire [9:0] ram_w4_l8192_id7_6_0_addr;
  wire [3:0] ram_w4_l8192_id7_6_0_rdata;
  wire [3:0] ram_w4_l8192_id7_6_0_wdata;
  wire ram_w4_l8192_id7_6_0_wenable;
  wire [9:0] ram_w4_l8192_id7_6_1_addr;
  wire [3:0] ram_w4_l8192_id7_6_1_rdata;
  wire [3:0] ram_w4_l8192_id7_6_1_wdata;
  wire ram_w4_l8192_id7_6_1_wenable;
  wire [9:0] ram_w4_l8192_id7_7_0_addr;
  wire [3:0] ram_w4_l8192_id7_7_0_rdata;
  wire [3:0] ram_w4_l8192_id7_7_0_wdata;
  wire ram_w4_l8192_id7_7_0_wenable;
  wire [9:0] ram_w4_l8192_id7_7_1_addr;
  wire [3:0] ram_w4_l8192_id7_7_1_rdata;
  wire [3:0] ram_w4_l8192_id7_7_1_wdata;
  wire ram_w4_l8192_id7_7_1_wenable;
  wire [9:0] ram_w4_l8192_id8_0_0_addr;
  wire [3:0] ram_w4_l8192_id8_0_0_rdata;
  wire [3:0] ram_w4_l8192_id8_0_0_wdata;
  wire ram_w4_l8192_id8_0_0_wenable;
  wire [9:0] ram_w4_l8192_id8_0_1_addr;
  wire [3:0] ram_w4_l8192_id8_0_1_rdata;
  wire [3:0] ram_w4_l8192_id8_0_1_wdata;
  wire ram_w4_l8192_id8_0_1_wenable;
  wire [9:0] ram_w4_l8192_id8_1_0_addr;
  wire [3:0] ram_w4_l8192_id8_1_0_rdata;
  wire [3:0] ram_w4_l8192_id8_1_0_wdata;
  wire ram_w4_l8192_id8_1_0_wenable;
  wire [9:0] ram_w4_l8192_id8_1_1_addr;
  wire [3:0] ram_w4_l8192_id8_1_1_rdata;
  wire [3:0] ram_w4_l8192_id8_1_1_wdata;
  wire ram_w4_l8192_id8_1_1_wenable;
  wire [9:0] ram_w4_l8192_id8_2_0_addr;
  wire [3:0] ram_w4_l8192_id8_2_0_rdata;
  wire [3:0] ram_w4_l8192_id8_2_0_wdata;
  wire ram_w4_l8192_id8_2_0_wenable;
  wire [9:0] ram_w4_l8192_id8_2_1_addr;
  wire [3:0] ram_w4_l8192_id8_2_1_rdata;
  wire [3:0] ram_w4_l8192_id8_2_1_wdata;
  wire ram_w4_l8192_id8_2_1_wenable;
  wire [9:0] ram_w4_l8192_id8_3_0_addr;
  wire [3:0] ram_w4_l8192_id8_3_0_rdata;
  wire [3:0] ram_w4_l8192_id8_3_0_wdata;
  wire ram_w4_l8192_id8_3_0_wenable;
  wire [9:0] ram_w4_l8192_id8_3_1_addr;
  wire [3:0] ram_w4_l8192_id8_3_1_rdata;
  wire [3:0] ram_w4_l8192_id8_3_1_wdata;
  wire ram_w4_l8192_id8_3_1_wenable;
  wire [9:0] ram_w4_l8192_id8_4_0_addr;
  wire [3:0] ram_w4_l8192_id8_4_0_rdata;
  wire [3:0] ram_w4_l8192_id8_4_0_wdata;
  wire ram_w4_l8192_id8_4_0_wenable;
  wire [9:0] ram_w4_l8192_id8_4_1_addr;
  wire [3:0] ram_w4_l8192_id8_4_1_rdata;
  wire [3:0] ram_w4_l8192_id8_4_1_wdata;
  wire ram_w4_l8192_id8_4_1_wenable;
  wire [9:0] ram_w4_l8192_id8_5_0_addr;
  wire [3:0] ram_w4_l8192_id8_5_0_rdata;
  wire [3:0] ram_w4_l8192_id8_5_0_wdata;
  wire ram_w4_l8192_id8_5_0_wenable;
  wire [9:0] ram_w4_l8192_id8_5_1_addr;
  wire [3:0] ram_w4_l8192_id8_5_1_rdata;
  wire [3:0] ram_w4_l8192_id8_5_1_wdata;
  wire ram_w4_l8192_id8_5_1_wenable;
  wire [9:0] ram_w4_l8192_id8_6_0_addr;
  wire [3:0] ram_w4_l8192_id8_6_0_rdata;
  wire [3:0] ram_w4_l8192_id8_6_0_wdata;
  wire ram_w4_l8192_id8_6_0_wenable;
  wire [9:0] ram_w4_l8192_id8_6_1_addr;
  wire [3:0] ram_w4_l8192_id8_6_1_rdata;
  wire [3:0] ram_w4_l8192_id8_6_1_wdata;
  wire ram_w4_l8192_id8_6_1_wenable;
  wire [9:0] ram_w4_l8192_id8_7_0_addr;
  wire [3:0] ram_w4_l8192_id8_7_0_rdata;
  wire [3:0] ram_w4_l8192_id8_7_0_wdata;
  wire ram_w4_l8192_id8_7_0_wenable;
  wire [9:0] ram_w4_l8192_id8_7_1_addr;
  wire [3:0] ram_w4_l8192_id8_7_1_rdata;
  wire [3:0] ram_w4_l8192_id8_7_1_wdata;
  wire ram_w4_l8192_id8_7_1_wenable;
  wire [8:0] ram_w8_l2048_id0_0_0_addr;
  wire [7:0] ram_w8_l2048_id0_0_0_rdata;
  wire [7:0] ram_w8_l2048_id0_0_0_wdata;
  wire ram_w8_l2048_id0_0_0_wenable;
  wire [8:0] ram_w8_l2048_id0_0_1_addr;
  wire [7:0] ram_w8_l2048_id0_0_1_rdata;
  wire [7:0] ram_w8_l2048_id0_0_1_wdata;
  wire ram_w8_l2048_id0_0_1_wenable;
  wire [8:0] ram_w8_l2048_id0_1_0_addr;
  wire [7:0] ram_w8_l2048_id0_1_0_rdata;
  wire [7:0] ram_w8_l2048_id0_1_0_wdata;
  wire ram_w8_l2048_id0_1_0_wenable;
  wire [8:0] ram_w8_l2048_id0_1_1_addr;
  wire [7:0] ram_w8_l2048_id0_1_1_rdata;
  wire [7:0] ram_w8_l2048_id0_1_1_wdata;
  wire ram_w8_l2048_id0_1_1_wenable;
  wire [8:0] ram_w8_l2048_id0_2_0_addr;
  wire [7:0] ram_w8_l2048_id0_2_0_rdata;
  wire [7:0] ram_w8_l2048_id0_2_0_wdata;
  wire ram_w8_l2048_id0_2_0_wenable;
  wire [8:0] ram_w8_l2048_id0_2_1_addr;
  wire [7:0] ram_w8_l2048_id0_2_1_rdata;
  wire [7:0] ram_w8_l2048_id0_2_1_wdata;
  wire ram_w8_l2048_id0_2_1_wenable;
  wire [8:0] ram_w8_l2048_id0_3_0_addr;
  wire [7:0] ram_w8_l2048_id0_3_0_rdata;
  wire [7:0] ram_w8_l2048_id0_3_0_wdata;
  wire ram_w8_l2048_id0_3_0_wenable;
  wire [8:0] ram_w8_l2048_id0_3_1_addr;
  wire [7:0] ram_w8_l2048_id0_3_1_rdata;
  wire [7:0] ram_w8_l2048_id0_3_1_wdata;
  wire ram_w8_l2048_id0_3_1_wenable;
  wire [8:0] ram_w8_l2048_id10_0_0_addr;
  wire [7:0] ram_w8_l2048_id10_0_0_rdata;
  wire [7:0] ram_w8_l2048_id10_0_0_wdata;
  wire ram_w8_l2048_id10_0_0_wenable;
  wire [8:0] ram_w8_l2048_id10_0_1_addr;
  wire [7:0] ram_w8_l2048_id10_0_1_rdata;
  wire [7:0] ram_w8_l2048_id10_0_1_wdata;
  wire ram_w8_l2048_id10_0_1_wenable;
  wire [8:0] ram_w8_l2048_id10_1_0_addr;
  wire [7:0] ram_w8_l2048_id10_1_0_rdata;
  wire [7:0] ram_w8_l2048_id10_1_0_wdata;
  wire ram_w8_l2048_id10_1_0_wenable;
  wire [8:0] ram_w8_l2048_id10_1_1_addr;
  wire [7:0] ram_w8_l2048_id10_1_1_rdata;
  wire [7:0] ram_w8_l2048_id10_1_1_wdata;
  wire ram_w8_l2048_id10_1_1_wenable;
  wire [8:0] ram_w8_l2048_id10_2_0_addr;
  wire [7:0] ram_w8_l2048_id10_2_0_rdata;
  wire [7:0] ram_w8_l2048_id10_2_0_wdata;
  wire ram_w8_l2048_id10_2_0_wenable;
  wire [8:0] ram_w8_l2048_id10_2_1_addr;
  wire [7:0] ram_w8_l2048_id10_2_1_rdata;
  wire [7:0] ram_w8_l2048_id10_2_1_wdata;
  wire ram_w8_l2048_id10_2_1_wenable;
  wire [8:0] ram_w8_l2048_id10_3_0_addr;
  wire [7:0] ram_w8_l2048_id10_3_0_rdata;
  wire [7:0] ram_w8_l2048_id10_3_0_wdata;
  wire ram_w8_l2048_id10_3_0_wenable;
  wire [8:0] ram_w8_l2048_id10_3_1_addr;
  wire [7:0] ram_w8_l2048_id10_3_1_rdata;
  wire [7:0] ram_w8_l2048_id10_3_1_wdata;
  wire ram_w8_l2048_id10_3_1_wenable;
  wire [8:0] ram_w8_l2048_id11_0_0_addr;
  wire [7:0] ram_w8_l2048_id11_0_0_rdata;
  wire [7:0] ram_w8_l2048_id11_0_0_wdata;
  wire ram_w8_l2048_id11_0_0_wenable;
  wire [8:0] ram_w8_l2048_id11_0_1_addr;
  wire [7:0] ram_w8_l2048_id11_0_1_rdata;
  wire [7:0] ram_w8_l2048_id11_0_1_wdata;
  wire ram_w8_l2048_id11_0_1_wenable;
  wire [8:0] ram_w8_l2048_id11_1_0_addr;
  wire [7:0] ram_w8_l2048_id11_1_0_rdata;
  wire [7:0] ram_w8_l2048_id11_1_0_wdata;
  wire ram_w8_l2048_id11_1_0_wenable;
  wire [8:0] ram_w8_l2048_id11_1_1_addr;
  wire [7:0] ram_w8_l2048_id11_1_1_rdata;
  wire [7:0] ram_w8_l2048_id11_1_1_wdata;
  wire ram_w8_l2048_id11_1_1_wenable;
  wire [8:0] ram_w8_l2048_id11_2_0_addr;
  wire [7:0] ram_w8_l2048_id11_2_0_rdata;
  wire [7:0] ram_w8_l2048_id11_2_0_wdata;
  wire ram_w8_l2048_id11_2_0_wenable;
  wire [8:0] ram_w8_l2048_id11_2_1_addr;
  wire [7:0] ram_w8_l2048_id11_2_1_rdata;
  wire [7:0] ram_w8_l2048_id11_2_1_wdata;
  wire ram_w8_l2048_id11_2_1_wenable;
  wire [8:0] ram_w8_l2048_id11_3_0_addr;
  wire [7:0] ram_w8_l2048_id11_3_0_rdata;
  wire [7:0] ram_w8_l2048_id11_3_0_wdata;
  wire ram_w8_l2048_id11_3_0_wenable;
  wire [8:0] ram_w8_l2048_id11_3_1_addr;
  wire [7:0] ram_w8_l2048_id11_3_1_rdata;
  wire [7:0] ram_w8_l2048_id11_3_1_wdata;
  wire ram_w8_l2048_id11_3_1_wenable;
  wire [8:0] ram_w8_l2048_id1_0_0_addr;
  wire [7:0] ram_w8_l2048_id1_0_0_rdata;
  wire [7:0] ram_w8_l2048_id1_0_0_wdata;
  wire ram_w8_l2048_id1_0_0_wenable;
  wire [8:0] ram_w8_l2048_id1_0_1_addr;
  wire [7:0] ram_w8_l2048_id1_0_1_rdata;
  wire [7:0] ram_w8_l2048_id1_0_1_wdata;
  wire ram_w8_l2048_id1_0_1_wenable;
  wire [8:0] ram_w8_l2048_id1_1_0_addr;
  wire [7:0] ram_w8_l2048_id1_1_0_rdata;
  wire [7:0] ram_w8_l2048_id1_1_0_wdata;
  wire ram_w8_l2048_id1_1_0_wenable;
  wire [8:0] ram_w8_l2048_id1_1_1_addr;
  wire [7:0] ram_w8_l2048_id1_1_1_rdata;
  wire [7:0] ram_w8_l2048_id1_1_1_wdata;
  wire ram_w8_l2048_id1_1_1_wenable;
  wire [8:0] ram_w8_l2048_id1_2_0_addr;
  wire [7:0] ram_w8_l2048_id1_2_0_rdata;
  wire [7:0] ram_w8_l2048_id1_2_0_wdata;
  wire ram_w8_l2048_id1_2_0_wenable;
  wire [8:0] ram_w8_l2048_id1_2_1_addr;
  wire [7:0] ram_w8_l2048_id1_2_1_rdata;
  wire [7:0] ram_w8_l2048_id1_2_1_wdata;
  wire ram_w8_l2048_id1_2_1_wenable;
  wire [8:0] ram_w8_l2048_id1_3_0_addr;
  wire [7:0] ram_w8_l2048_id1_3_0_rdata;
  wire [7:0] ram_w8_l2048_id1_3_0_wdata;
  wire ram_w8_l2048_id1_3_0_wenable;
  wire [8:0] ram_w8_l2048_id1_3_1_addr;
  wire [7:0] ram_w8_l2048_id1_3_1_rdata;
  wire [7:0] ram_w8_l2048_id1_3_1_wdata;
  wire ram_w8_l2048_id1_3_1_wenable;
  wire [8:0] ram_w8_l2048_id2_0_0_addr;
  wire [7:0] ram_w8_l2048_id2_0_0_rdata;
  wire [7:0] ram_w8_l2048_id2_0_0_wdata;
  wire ram_w8_l2048_id2_0_0_wenable;
  wire [8:0] ram_w8_l2048_id2_0_1_addr;
  wire [7:0] ram_w8_l2048_id2_0_1_rdata;
  wire [7:0] ram_w8_l2048_id2_0_1_wdata;
  wire ram_w8_l2048_id2_0_1_wenable;
  wire [8:0] ram_w8_l2048_id2_1_0_addr;
  wire [7:0] ram_w8_l2048_id2_1_0_rdata;
  wire [7:0] ram_w8_l2048_id2_1_0_wdata;
  wire ram_w8_l2048_id2_1_0_wenable;
  wire [8:0] ram_w8_l2048_id2_1_1_addr;
  wire [7:0] ram_w8_l2048_id2_1_1_rdata;
  wire [7:0] ram_w8_l2048_id2_1_1_wdata;
  wire ram_w8_l2048_id2_1_1_wenable;
  wire [8:0] ram_w8_l2048_id2_2_0_addr;
  wire [7:0] ram_w8_l2048_id2_2_0_rdata;
  wire [7:0] ram_w8_l2048_id2_2_0_wdata;
  wire ram_w8_l2048_id2_2_0_wenable;
  wire [8:0] ram_w8_l2048_id2_2_1_addr;
  wire [7:0] ram_w8_l2048_id2_2_1_rdata;
  wire [7:0] ram_w8_l2048_id2_2_1_wdata;
  wire ram_w8_l2048_id2_2_1_wenable;
  wire [8:0] ram_w8_l2048_id2_3_0_addr;
  wire [7:0] ram_w8_l2048_id2_3_0_rdata;
  wire [7:0] ram_w8_l2048_id2_3_0_wdata;
  wire ram_w8_l2048_id2_3_0_wenable;
  wire [8:0] ram_w8_l2048_id2_3_1_addr;
  wire [7:0] ram_w8_l2048_id2_3_1_rdata;
  wire [7:0] ram_w8_l2048_id2_3_1_wdata;
  wire ram_w8_l2048_id2_3_1_wenable;
  wire [8:0] ram_w8_l2048_id3_0_0_addr;
  wire [7:0] ram_w8_l2048_id3_0_0_rdata;
  wire [7:0] ram_w8_l2048_id3_0_0_wdata;
  wire ram_w8_l2048_id3_0_0_wenable;
  wire [8:0] ram_w8_l2048_id3_0_1_addr;
  wire [7:0] ram_w8_l2048_id3_0_1_rdata;
  wire [7:0] ram_w8_l2048_id3_0_1_wdata;
  wire ram_w8_l2048_id3_0_1_wenable;
  wire [8:0] ram_w8_l2048_id3_1_0_addr;
  wire [7:0] ram_w8_l2048_id3_1_0_rdata;
  wire [7:0] ram_w8_l2048_id3_1_0_wdata;
  wire ram_w8_l2048_id3_1_0_wenable;
  wire [8:0] ram_w8_l2048_id3_1_1_addr;
  wire [7:0] ram_w8_l2048_id3_1_1_rdata;
  wire [7:0] ram_w8_l2048_id3_1_1_wdata;
  wire ram_w8_l2048_id3_1_1_wenable;
  wire [8:0] ram_w8_l2048_id3_2_0_addr;
  wire [7:0] ram_w8_l2048_id3_2_0_rdata;
  wire [7:0] ram_w8_l2048_id3_2_0_wdata;
  wire ram_w8_l2048_id3_2_0_wenable;
  wire [8:0] ram_w8_l2048_id3_2_1_addr;
  wire [7:0] ram_w8_l2048_id3_2_1_rdata;
  wire [7:0] ram_w8_l2048_id3_2_1_wdata;
  wire ram_w8_l2048_id3_2_1_wenable;
  wire [8:0] ram_w8_l2048_id3_3_0_addr;
  wire [7:0] ram_w8_l2048_id3_3_0_rdata;
  wire [7:0] ram_w8_l2048_id3_3_0_wdata;
  wire ram_w8_l2048_id3_3_0_wenable;
  wire [8:0] ram_w8_l2048_id3_3_1_addr;
  wire [7:0] ram_w8_l2048_id3_3_1_rdata;
  wire [7:0] ram_w8_l2048_id3_3_1_wdata;
  wire ram_w8_l2048_id3_3_1_wenable;
  wire [8:0] ram_w8_l2048_id4_0_0_addr;
  wire [7:0] ram_w8_l2048_id4_0_0_rdata;
  wire [7:0] ram_w8_l2048_id4_0_0_wdata;
  wire ram_w8_l2048_id4_0_0_wenable;
  wire [8:0] ram_w8_l2048_id4_0_1_addr;
  wire [7:0] ram_w8_l2048_id4_0_1_rdata;
  wire [7:0] ram_w8_l2048_id4_0_1_wdata;
  wire ram_w8_l2048_id4_0_1_wenable;
  wire [8:0] ram_w8_l2048_id4_1_0_addr;
  wire [7:0] ram_w8_l2048_id4_1_0_rdata;
  wire [7:0] ram_w8_l2048_id4_1_0_wdata;
  wire ram_w8_l2048_id4_1_0_wenable;
  wire [8:0] ram_w8_l2048_id4_1_1_addr;
  wire [7:0] ram_w8_l2048_id4_1_1_rdata;
  wire [7:0] ram_w8_l2048_id4_1_1_wdata;
  wire ram_w8_l2048_id4_1_1_wenable;
  wire [8:0] ram_w8_l2048_id4_2_0_addr;
  wire [7:0] ram_w8_l2048_id4_2_0_rdata;
  wire [7:0] ram_w8_l2048_id4_2_0_wdata;
  wire ram_w8_l2048_id4_2_0_wenable;
  wire [8:0] ram_w8_l2048_id4_2_1_addr;
  wire [7:0] ram_w8_l2048_id4_2_1_rdata;
  wire [7:0] ram_w8_l2048_id4_2_1_wdata;
  wire ram_w8_l2048_id4_2_1_wenable;
  wire [8:0] ram_w8_l2048_id4_3_0_addr;
  wire [7:0] ram_w8_l2048_id4_3_0_rdata;
  wire [7:0] ram_w8_l2048_id4_3_0_wdata;
  wire ram_w8_l2048_id4_3_0_wenable;
  wire [8:0] ram_w8_l2048_id4_3_1_addr;
  wire [7:0] ram_w8_l2048_id4_3_1_rdata;
  wire [7:0] ram_w8_l2048_id4_3_1_wdata;
  wire ram_w8_l2048_id4_3_1_wenable;
  wire [8:0] ram_w8_l2048_id5_0_0_addr;
  wire [7:0] ram_w8_l2048_id5_0_0_rdata;
  wire [7:0] ram_w8_l2048_id5_0_0_wdata;
  wire ram_w8_l2048_id5_0_0_wenable;
  wire [8:0] ram_w8_l2048_id5_0_1_addr;
  wire [7:0] ram_w8_l2048_id5_0_1_rdata;
  wire [7:0] ram_w8_l2048_id5_0_1_wdata;
  wire ram_w8_l2048_id5_0_1_wenable;
  wire [8:0] ram_w8_l2048_id5_1_0_addr;
  wire [7:0] ram_w8_l2048_id5_1_0_rdata;
  wire [7:0] ram_w8_l2048_id5_1_0_wdata;
  wire ram_w8_l2048_id5_1_0_wenable;
  wire [8:0] ram_w8_l2048_id5_1_1_addr;
  wire [7:0] ram_w8_l2048_id5_1_1_rdata;
  wire [7:0] ram_w8_l2048_id5_1_1_wdata;
  wire ram_w8_l2048_id5_1_1_wenable;
  wire [8:0] ram_w8_l2048_id5_2_0_addr;
  wire [7:0] ram_w8_l2048_id5_2_0_rdata;
  wire [7:0] ram_w8_l2048_id5_2_0_wdata;
  wire ram_w8_l2048_id5_2_0_wenable;
  wire [8:0] ram_w8_l2048_id5_2_1_addr;
  wire [7:0] ram_w8_l2048_id5_2_1_rdata;
  wire [7:0] ram_w8_l2048_id5_2_1_wdata;
  wire ram_w8_l2048_id5_2_1_wenable;
  wire [8:0] ram_w8_l2048_id5_3_0_addr;
  wire [7:0] ram_w8_l2048_id5_3_0_rdata;
  wire [7:0] ram_w8_l2048_id5_3_0_wdata;
  wire ram_w8_l2048_id5_3_0_wenable;
  wire [8:0] ram_w8_l2048_id5_3_1_addr;
  wire [7:0] ram_w8_l2048_id5_3_1_rdata;
  wire [7:0] ram_w8_l2048_id5_3_1_wdata;
  wire ram_w8_l2048_id5_3_1_wenable;
  wire [8:0] ram_w8_l2048_id6_0_0_addr;
  wire [7:0] ram_w8_l2048_id6_0_0_rdata;
  wire [7:0] ram_w8_l2048_id6_0_0_wdata;
  wire ram_w8_l2048_id6_0_0_wenable;
  wire [8:0] ram_w8_l2048_id6_0_1_addr;
  wire [7:0] ram_w8_l2048_id6_0_1_rdata;
  wire [7:0] ram_w8_l2048_id6_0_1_wdata;
  wire ram_w8_l2048_id6_0_1_wenable;
  wire [8:0] ram_w8_l2048_id6_1_0_addr;
  wire [7:0] ram_w8_l2048_id6_1_0_rdata;
  wire [7:0] ram_w8_l2048_id6_1_0_wdata;
  wire ram_w8_l2048_id6_1_0_wenable;
  wire [8:0] ram_w8_l2048_id6_1_1_addr;
  wire [7:0] ram_w8_l2048_id6_1_1_rdata;
  wire [7:0] ram_w8_l2048_id6_1_1_wdata;
  wire ram_w8_l2048_id6_1_1_wenable;
  wire [8:0] ram_w8_l2048_id6_2_0_addr;
  wire [7:0] ram_w8_l2048_id6_2_0_rdata;
  wire [7:0] ram_w8_l2048_id6_2_0_wdata;
  wire ram_w8_l2048_id6_2_0_wenable;
  wire [8:0] ram_w8_l2048_id6_2_1_addr;
  wire [7:0] ram_w8_l2048_id6_2_1_rdata;
  wire [7:0] ram_w8_l2048_id6_2_1_wdata;
  wire ram_w8_l2048_id6_2_1_wenable;
  wire [8:0] ram_w8_l2048_id6_3_0_addr;
  wire [7:0] ram_w8_l2048_id6_3_0_rdata;
  wire [7:0] ram_w8_l2048_id6_3_0_wdata;
  wire ram_w8_l2048_id6_3_0_wenable;
  wire [8:0] ram_w8_l2048_id6_3_1_addr;
  wire [7:0] ram_w8_l2048_id6_3_1_rdata;
  wire [7:0] ram_w8_l2048_id6_3_1_wdata;
  wire ram_w8_l2048_id6_3_1_wenable;
  wire [8:0] ram_w8_l2048_id7_0_0_addr;
  wire [7:0] ram_w8_l2048_id7_0_0_rdata;
  wire [7:0] ram_w8_l2048_id7_0_0_wdata;
  wire ram_w8_l2048_id7_0_0_wenable;
  wire [8:0] ram_w8_l2048_id7_0_1_addr;
  wire [7:0] ram_w8_l2048_id7_0_1_rdata;
  wire [7:0] ram_w8_l2048_id7_0_1_wdata;
  wire ram_w8_l2048_id7_0_1_wenable;
  wire [8:0] ram_w8_l2048_id7_1_0_addr;
  wire [7:0] ram_w8_l2048_id7_1_0_rdata;
  wire [7:0] ram_w8_l2048_id7_1_0_wdata;
  wire ram_w8_l2048_id7_1_0_wenable;
  wire [8:0] ram_w8_l2048_id7_1_1_addr;
  wire [7:0] ram_w8_l2048_id7_1_1_rdata;
  wire [7:0] ram_w8_l2048_id7_1_1_wdata;
  wire ram_w8_l2048_id7_1_1_wenable;
  wire [8:0] ram_w8_l2048_id7_2_0_addr;
  wire [7:0] ram_w8_l2048_id7_2_0_rdata;
  wire [7:0] ram_w8_l2048_id7_2_0_wdata;
  wire ram_w8_l2048_id7_2_0_wenable;
  wire [8:0] ram_w8_l2048_id7_2_1_addr;
  wire [7:0] ram_w8_l2048_id7_2_1_rdata;
  wire [7:0] ram_w8_l2048_id7_2_1_wdata;
  wire ram_w8_l2048_id7_2_1_wenable;
  wire [8:0] ram_w8_l2048_id7_3_0_addr;
  wire [7:0] ram_w8_l2048_id7_3_0_rdata;
  wire [7:0] ram_w8_l2048_id7_3_0_wdata;
  wire ram_w8_l2048_id7_3_0_wenable;
  wire [8:0] ram_w8_l2048_id7_3_1_addr;
  wire [7:0] ram_w8_l2048_id7_3_1_rdata;
  wire [7:0] ram_w8_l2048_id7_3_1_wdata;
  wire ram_w8_l2048_id7_3_1_wenable;
  wire [8:0] ram_w8_l2048_id8_0_0_addr;
  wire [7:0] ram_w8_l2048_id8_0_0_rdata;
  wire [7:0] ram_w8_l2048_id8_0_0_wdata;
  wire ram_w8_l2048_id8_0_0_wenable;
  wire [8:0] ram_w8_l2048_id8_0_1_addr;
  wire [7:0] ram_w8_l2048_id8_0_1_rdata;
  wire [7:0] ram_w8_l2048_id8_0_1_wdata;
  wire ram_w8_l2048_id8_0_1_wenable;
  wire [8:0] ram_w8_l2048_id8_1_0_addr;
  wire [7:0] ram_w8_l2048_id8_1_0_rdata;
  wire [7:0] ram_w8_l2048_id8_1_0_wdata;
  wire ram_w8_l2048_id8_1_0_wenable;
  wire [8:0] ram_w8_l2048_id8_1_1_addr;
  wire [7:0] ram_w8_l2048_id8_1_1_rdata;
  wire [7:0] ram_w8_l2048_id8_1_1_wdata;
  wire ram_w8_l2048_id8_1_1_wenable;
  wire [8:0] ram_w8_l2048_id8_2_0_addr;
  wire [7:0] ram_w8_l2048_id8_2_0_rdata;
  wire [7:0] ram_w8_l2048_id8_2_0_wdata;
  wire ram_w8_l2048_id8_2_0_wenable;
  wire [8:0] ram_w8_l2048_id8_2_1_addr;
  wire [7:0] ram_w8_l2048_id8_2_1_rdata;
  wire [7:0] ram_w8_l2048_id8_2_1_wdata;
  wire ram_w8_l2048_id8_2_1_wenable;
  wire [8:0] ram_w8_l2048_id8_3_0_addr;
  wire [7:0] ram_w8_l2048_id8_3_0_rdata;
  wire [7:0] ram_w8_l2048_id8_3_0_wdata;
  wire ram_w8_l2048_id8_3_0_wenable;
  wire [8:0] ram_w8_l2048_id8_3_1_addr;
  wire [7:0] ram_w8_l2048_id8_3_1_rdata;
  wire [7:0] ram_w8_l2048_id8_3_1_wdata;
  wire ram_w8_l2048_id8_3_1_wenable;
  wire [8:0] ram_w8_l2048_id9_0_0_addr;
  wire [7:0] ram_w8_l2048_id9_0_0_rdata;
  wire [7:0] ram_w8_l2048_id9_0_0_wdata;
  wire ram_w8_l2048_id9_0_0_wenable;
  wire [8:0] ram_w8_l2048_id9_0_1_addr;
  wire [7:0] ram_w8_l2048_id9_0_1_rdata;
  wire [7:0] ram_w8_l2048_id9_0_1_wdata;
  wire ram_w8_l2048_id9_0_1_wenable;
  wire [8:0] ram_w8_l2048_id9_1_0_addr;
  wire [7:0] ram_w8_l2048_id9_1_0_rdata;
  wire [7:0] ram_w8_l2048_id9_1_0_wdata;
  wire ram_w8_l2048_id9_1_0_wenable;
  wire [8:0] ram_w8_l2048_id9_1_1_addr;
  wire [7:0] ram_w8_l2048_id9_1_1_rdata;
  wire [7:0] ram_w8_l2048_id9_1_1_wdata;
  wire ram_w8_l2048_id9_1_1_wenable;
  wire [8:0] ram_w8_l2048_id9_2_0_addr;
  wire [7:0] ram_w8_l2048_id9_2_0_rdata;
  wire [7:0] ram_w8_l2048_id9_2_0_wdata;
  wire ram_w8_l2048_id9_2_0_wenable;
  wire [8:0] ram_w8_l2048_id9_2_1_addr;
  wire [7:0] ram_w8_l2048_id9_2_1_rdata;
  wire [7:0] ram_w8_l2048_id9_2_1_wdata;
  wire ram_w8_l2048_id9_2_1_wenable;
  wire [8:0] ram_w8_l2048_id9_3_0_addr;
  wire [7:0] ram_w8_l2048_id9_3_0_rdata;
  wire [7:0] ram_w8_l2048_id9_3_0_wdata;
  wire ram_w8_l2048_id9_3_0_wenable;
  wire [8:0] ram_w8_l2048_id9_3_1_addr;
  wire [7:0] ram_w8_l2048_id9_3_1_rdata;
  wire [7:0] ram_w8_l2048_id9_3_1_wdata;
  wire ram_w8_l2048_id9_3_1_wenable;
  wire [8:0] req_block_size_286;
  wire [9:0] req_block_size_33;
  wire [8:0] req_block_size_343;
  wire [8:0] req_block_size_400;
  wire rst_logic;
  wire set_req_287;
  wire set_req_34;
  wire set_req_344;
  wire set_req_401;
  wire [5:0] stream_conv2d_16_constant_0_data;
  wire stream_conv2d_16_constant_15_data;
  wire stream_conv2d_16_constant_16_data;
  wire [3:0] stream_conv2d_16_constant_17_data;
  wire [1:0] stream_conv2d_16_constant_1_data;
  wire [1:0] stream_conv2d_16_constant_2_data;
  wire [8:0] stream_conv2d_16_constant_3_data;
  wire [7:0] stream_conv2d_16_sink_37_data;
  wire stream_conv2d_16_sink_38_data;
  wire [7:0] stream_conv2d_16_source_10_data;
  wire [7:0] stream_conv2d_16_source_12_data;
  wire [7:0] stream_conv2d_16_source_14_data;
  wire [7:0] stream_conv2d_16_source_19_data;
  wire [7:0] stream_conv2d_16_source_20_data;
  wire [7:0] stream_conv2d_16_source_21_data;
  wire [7:0] stream_conv2d_16_source_22_data;
  wire [7:0] stream_conv2d_16_source_23_data;
  wire [7:0] stream_conv2d_16_source_24_data;
  wire [7:0] stream_conv2d_16_source_25_data;
  wire [7:0] stream_conv2d_16_source_26_data;
  wire [7:0] stream_conv2d_16_source_27_data;
  wire [3:0] stream_conv2d_16_source_28_data;
  wire [3:0] stream_conv2d_16_source_29_data;
  wire [3:0] stream_conv2d_16_source_30_data;
  wire [3:0] stream_conv2d_16_source_31_data;
  wire [3:0] stream_conv2d_16_source_32_data;
  wire [3:0] stream_conv2d_16_source_33_data;
  wire [3:0] stream_conv2d_16_source_34_data;
  wire [3:0] stream_conv2d_16_source_35_data;
  wire [3:0] stream_conv2d_16_source_36_data;
  wire [7:0] stream_conv2d_16_source_6_data;
  wire [7:0] stream_conv2d_16_source_8_data;
  wire [10:0] stream_matmul_29_constant_0_data;
  wire stream_matmul_29_constant_15_data;
  wire stream_matmul_29_constant_16_data;
  wire [3:0] stream_matmul_29_constant_17_data;
  wire [1:0] stream_matmul_29_constant_18_data;
  wire stream_matmul_29_constant_1_data;
  wire stream_matmul_29_constant_2_data;
  wire stream_matmul_29_constant_3_data;
  wire [7:0] stream_matmul_29_sink_21_data;
  wire stream_matmul_29_sink_22_data;
  wire [7:0] stream_matmul_29_source_10_data;
  wire [7:0] stream_matmul_29_source_12_data;
  wire [7:0] stream_matmul_29_source_14_data;
  wire [7:0] stream_matmul_29_source_19_data;
  wire [3:0] stream_matmul_29_source_20_data;
  wire [7:0] stream_matmul_29_source_6_data;
  wire [7:0] stream_matmul_29_source_8_data;
  wire [2:0] stream_max_pool_serial_18_constant_0_data;
  wire [3:0] stream_max_pool_serial_18_constant_2_data;
  wire [7:0] stream_max_pool_serial_18_sink_3_data;
  wire stream_max_pool_serial_18_sink_4_data;
  wire [7:0] stream_max_pool_serial_18_source_1_data;
  assign _24482_[9:0] = _tmp_50;
  assign _24483_[9:0] = _tmp_51;
  assign _24484_[9:0] = _tmp_52;
  assign _24485_[9:0] = _tmp_53;
  assign _24486_[9:0] = _tmp_54;
  assign _24487_[9:0] = _tmp_55;
  assign _24488_[9:0] = _tmp_56;
  assign _24489_[9:0] = _tmp_57;
  assign _24490_[9:0] = _tmp_58;
  assign _24491_[9:0] = _tmp_81;
  assign _24492_[9:0] = _tmp_82;
  assign _24493_[9:0] = _tmp_83;
  assign _24494_[9:0] = _tmp_84;
  assign _24495_[9:0] = _tmp_85;
  assign _24496_[9:0] = _tmp_86;
  assign _24497_[9:0] = _tmp_87;
  assign _24498_[9:0] = _tmp_88;
  assign _24499_[9:0] = _tmp_89;
  assign _24500_[9:0] = _tmp_112;
  assign _24501_[9:0] = _tmp_113;
  assign _24502_[9:0] = _tmp_114;
  assign _24503_[9:0] = _tmp_115;
  assign _24504_[9:0] = _tmp_116;
  assign _24505_[9:0] = _tmp_117;
  assign _24506_[9:0] = _tmp_118;
  assign _24507_[9:0] = _tmp_119;
  assign _24508_[9:0] = _tmp_120;
  assign _24509_[9:0] = _tmp_143;
  assign _24510_[9:0] = _tmp_144;
  assign _24511_[9:0] = _tmp_145;
  assign _24512_[9:0] = _tmp_146;
  assign _24513_[9:0] = _tmp_147;
  assign _24514_[9:0] = _tmp_148;
  assign _24515_[9:0] = _tmp_149;
  assign _24516_[9:0] = _tmp_150;
  assign _24517_[9:0] = _tmp_151;
  assign _24518_[9:0] = _tmp_174;
  assign _24519_[9:0] = _tmp_175;
  assign _24520_[9:0] = _tmp_176;
  assign _24521_[9:0] = _tmp_177;
  assign _24522_[9:0] = _tmp_178;
  assign _24523_[9:0] = _tmp_179;
  assign _24524_[9:0] = _tmp_180;
  assign _24525_[9:0] = _tmp_181;
  assign _24526_[9:0] = _tmp_182;
  assign _24527_[9:0] = _tmp_205;
  assign _24528_[9:0] = _tmp_206;
  assign _24529_[9:0] = _tmp_207;
  assign _24530_[9:0] = _tmp_208;
  assign _24531_[9:0] = _tmp_209;
  assign _24532_[9:0] = _tmp_210;
  assign _24533_[9:0] = _tmp_211;
  assign _24534_[9:0] = _tmp_212;
  assign _24535_[9:0] = _tmp_213;
  assign _24536_[9:0] = _tmp_236;
  assign _24537_[9:0] = _tmp_237;
  assign _24538_[9:0] = _tmp_238;
  assign _24539_[9:0] = _tmp_239;
  assign _24540_[9:0] = _tmp_240;
  assign _24541_[9:0] = _tmp_241;
  assign _24542_[9:0] = _tmp_242;
  assign _24543_[9:0] = _tmp_243;
  assign _24544_[9:0] = _tmp_244;
  assign _24545_[9:0] = _tmp_267;
  assign _24546_[9:0] = _tmp_268;
  assign _24547_[9:0] = _tmp_269;
  assign _24548_[9:0] = _tmp_270;
  assign _24549_[9:0] = _tmp_271;
  assign _24550_[9:0] = _tmp_272;
  assign _24551_[9:0] = _tmp_273;
  assign _24552_[9:0] = _tmp_274;
  assign _24553_[9:0] = _tmp_275;
  assign _24559_[8:0] = _tmp_297;
  assign _24560_[8:0] = _tmp_298;
  assign _24561_[8:0] = _tmp_299;
  assign _24562_[8:0] = _tmp_310;
  assign _24563_[8:0] = _tmp_311;
  assign _24564_[8:0] = _tmp_312;
  assign _24565_[8:0] = _tmp_323;
  assign _24566_[8:0] = _tmp_324;
  assign _24567_[8:0] = _tmp_325;
  assign _24568_[8:0] = _tmp_336;
  assign _24569_[8:0] = _tmp_337;
  assign _24570_[8:0] = _tmp_338;
  assign _24571_[8:0] = _tmp_354;
  assign _24572_[8:0] = _tmp_355;
  assign _24573_[8:0] = _tmp_356;
  assign _24574_[8:0] = _tmp_367;
  assign _24575_[8:0] = _tmp_368;
  assign _24576_[8:0] = _tmp_369;
  assign _24577_[8:0] = _tmp_380;
  assign _24578_[8:0] = _tmp_381;
  assign _24579_[8:0] = _tmp_382;
  assign _24580_[8:0] = _tmp_393;
  assign _24581_[8:0] = _tmp_394;
  assign _24582_[8:0] = _tmp_395;
  assign _24583_[8:0] = _tmp_411;
  assign _24584_[8:0] = _tmp_412;
  assign _24585_[8:0] = _tmp_413;
  assign _24586_[8:0] = _tmp_424;
  assign _24587_[8:0] = _tmp_425;
  assign _24588_[8:0] = _tmp_426;
  assign _24589_[8:0] = _tmp_437;
  assign _24590_[8:0] = _tmp_438;
  assign _24591_[8:0] = _tmp_439;
  assign _24592_[8:0] = _tmp_450;
  assign _24593_[8:0] = _tmp_451;
  assign _24594_[8:0] = _tmp_452;
  assign _28519_[32:31] = 2'h0;
  assign _28520_[32:31] = 2'h0;
  assign _28936_[32:2] = _28519_[30:0];
  assign _28940_[32:2] = _28520_[30:0];
  assign _28943_[15:0] = 16'h0000;
  assign _28944_[31:0] = 0;
  assign _28948_[49:0] = _28943_[65:16];
  assign _28949_[33:0] = _28944_[65:32];
  assign _28978_[30:23] = { _28978_[31], _28978_[31], _28978_[31], _28978_[31], _28978_[31], _28978_[31], _28978_[31], _28978_[31] };
  assign _28982_[31:8] = { _28978_[31], _28978_[22:0] };
  assign _28984_[38:31] = { _28984_[39], _28984_[39], _28984_[39], _28984_[39], _28984_[39], _28984_[39], _28984_[39], _28984_[39] };
  assign _28988_[39:8] = { _28984_[39], _28984_[30:0] };
  assign _28989_[10:3] = { _28989_[11], _28989_[11], _28989_[11], _28989_[11], _28989_[11], _28989_[11], _28989_[11], _28989_[11] };
  assign _28992_[11:8] = { _28989_[11], _28989_[2:0] };
  assign _28993_[10:3] = { _28993_[11], _28993_[11], _28993_[11], _28993_[11], _28993_[11], _28993_[11], _28993_[11], _28993_[11] };
  assign _28996_[11:8] = { _28993_[11], _28993_[2:0] };
  assign _28997_[10:3] = { _28997_[11], _28997_[11], _28997_[11], _28997_[11], _28997_[11], _28997_[11], _28997_[11], _28997_[11] };
  assign _29000_[11:8] = { _28997_[11], _28997_[2:0] };
  assign _29001_[10:3] = { _29001_[11], _29001_[11], _29001_[11], _29001_[11], _29001_[11], _29001_[11], _29001_[11], _29001_[11] };
  assign _29004_[11:8] = { _29001_[11], _29001_[2:0] };
  assign _29005_[10:3] = { _29005_[11], _29005_[11], _29005_[11], _29005_[11], _29005_[11], _29005_[11], _29005_[11], _29005_[11] };
  assign _29008_[11:8] = { _29005_[11], _29005_[2:0] };
  assign _29009_[10:3] = { _29009_[11], _29009_[11], _29009_[11], _29009_[11], _29009_[11], _29009_[11], _29009_[11], _29009_[11] };
  assign _29012_[11:8] = { _29009_[11], _29009_[2:0] };
  assign _29013_[10:3] = { _29013_[11], _29013_[11], _29013_[11], _29013_[11], _29013_[11], _29013_[11], _29013_[11], _29013_[11] };
  assign _29016_[11:8] = { _29013_[11], _29013_[2:0] };
  assign _29017_[10:3] = { _29017_[11], _29017_[11], _29017_[11], _29017_[11], _29017_[11], _29017_[11], _29017_[11], _29017_[11] };
  assign _29020_[11:8] = { _29017_[11], _29017_[2:0] };
  assign _29021_[10:3] = { _29021_[11], _29021_[11], _29021_[11], _29021_[11], _29021_[11], _29021_[11], _29021_[11], _29021_[11] };
  assign _29024_[11:8] = { _29021_[11], _29021_[2:0] };
  assign _29060_[0] = conv2d_16_mux_next_dma_flag_0;
  assign _29062_[0] = conv2d_16_mux_next_dma_flag_1;
  assign _29065_[0] = conv2d_16_mux_next_dma_flag_2;
  assign _29069_[7:0] = _tmp_1032;
  assign _29070_[7:0] = _stream_max_pool_serial_18_source_1_source_ram_rdata;
  assign _29071_[0] = _stream_max_pool_serial_18_start_flag;
  assign _29075_[7:0] = _tmp_1175;
  assign _29076_[7:0] = _stream_matmul_29_source_6_source_ram_rdata;
  assign _29080_[7:0] = _tmp_1186;
  assign _29081_[7:0] = _stream_matmul_29_source_8_source_ram_rdata;
  assign _29085_[7:0] = _tmp_1206;
  assign _29086_[7:0] = _stream_matmul_29_source_19_source_ram_rdata;
  assign _29094_[3:0] = _tmp_1220;
  assign _29095_[3:0] = _stream_matmul_29_source_20_source_ram_rdata;
  assign _29096_[0] = _stream_matmul_29_start_flag;
  assign _29099_[0] = _maxi_write_data_done;
  assign _29134_[0] = _tmp_7;
  assign _29234_[5:0] = cparam_conv2d_16_act_num_row;
  assign _29236_[6:0] = cparam_conv2d_16_bias_num;
  assign _29238_[3:0] = cparam_conv2d_16_cshamt_out_value;
  assign _29240_[4:0] = cparam_conv2d_16_max_col_count;
  assign _29242_[7:0] = cparam_conv2d_16_och_count_step;
  assign _29244_[5:0] = cparam_conv2d_16_inc_act_laddr_large;
  assign _29245_[6:0] = cparam_conv2d_16_act_read_step;
  assign _29247_[13:0] = cparam_conv2d_16_filter_base_step;
  assign _29249_[14:0] = cparam_conv2d_16_filter_read_size;
  assign _29250_[5:0] = cparam_conv2d_16_filter_read_block;
  assign _29252_[11:0] = cparam_conv2d_16_filter_read_step;
  assign _29253_[5:0] = cparam_conv2d_16_stream_reduce_size;
  assign _29255_[6:0] = cparam_conv2d_16_stream_act_local_large_offset;
  assign _29257_[5:0] = cparam_max_pool_serial_18_act_num_col;
  assign _29259_[4:0] = cparam_max_pool_serial_18_max_col_count;
  assign _29261_[6:0] = cparam_max_pool_serial_18_inc_out_laddr;
  assign _29263_[7:0] = cparam_max_pool_serial_18_inc_act_laddr;
  assign _29265_[8:0] = cparam_matmul_29_bias_num;
  assign _29267_[3:0] = cparam_matmul_29_cshamt_out_value;
  assign _29269_[0] = cparam_matmul_29_keep_filter;
  assign _29271_[7:0] = cparam_matmul_29_max_och_count;
  assign _29273_[5:0] = cparam_matmul_29_och_count_step;
  assign _29275_[10:0] = cparam_matmul_29_act_bat_step;
  assign _29277_[11:0] = cparam_matmul_29_filter_base_step;
  assign _29279_[12:0] = cparam_matmul_29_filter_read_size;
  assign _29283_[8:0] = cparam_matmul_29_out_bat_step;
  assign _29285_[4:0] = cparam_matmul_29_out_och_step;
  assign _29287_[4:0] = cparam_matmul_29_out_write_size;
  assign _29319_[7:0] = _tmp_469;
  assign _29320_[7:0] = _stream_conv2d_16_source_6_source_ram_rdata;
  assign _29324_[7:0] = _tmp_480;
  assign _29325_[7:0] = _stream_conv2d_16_source_8_source_ram_rdata;
  assign _29329_[7:0] = _tmp_500;
  assign _29330_[7:0] = _stream_conv2d_16_source_19_source_ram_rdata;
  assign _29334_[7:0] = _tmp_510;
  assign _29335_[7:0] = _stream_conv2d_16_source_20_source_ram_rdata;
  assign _29339_[7:0] = _tmp_520;
  assign _29340_[7:0] = _stream_conv2d_16_source_21_source_ram_rdata;
  assign _29344_[7:0] = _tmp_530;
  assign _29345_[7:0] = _stream_conv2d_16_source_22_source_ram_rdata;
  assign _29349_[7:0] = _tmp_540;
  assign _29350_[7:0] = _stream_conv2d_16_source_23_source_ram_rdata;
  assign _29354_[7:0] = _tmp_550;
  assign _29355_[7:0] = _stream_conv2d_16_source_24_source_ram_rdata;
  assign _29359_[7:0] = _tmp_560;
  assign _29360_[7:0] = _stream_conv2d_16_source_25_source_ram_rdata;
  assign _29364_[7:0] = _tmp_570;
  assign _29365_[7:0] = _stream_conv2d_16_source_26_source_ram_rdata;
  assign _29369_[7:0] = _tmp_580;
  assign _29370_[7:0] = _stream_conv2d_16_source_27_source_ram_rdata;
  assign _29378_[3:0] = _tmp_594;
  assign _29379_[3:0] = _stream_conv2d_16_source_28_source_ram_rdata;
  assign _29387_[3:0] = _tmp_608;
  assign _29388_[3:0] = _stream_conv2d_16_source_29_source_ram_rdata;
  assign _29396_[3:0] = _tmp_622;
  assign _29397_[3:0] = _stream_conv2d_16_source_30_source_ram_rdata;
  assign _29405_[3:0] = _tmp_636;
  assign _29406_[3:0] = _stream_conv2d_16_source_31_source_ram_rdata;
  assign _29414_[3:0] = _tmp_650;
  assign _29415_[3:0] = _stream_conv2d_16_source_32_source_ram_rdata;
  assign _29423_[3:0] = _tmp_664;
  assign _29424_[3:0] = _stream_conv2d_16_source_33_source_ram_rdata;
  assign _29432_[3:0] = _tmp_678;
  assign _29433_[3:0] = _stream_conv2d_16_source_34_source_ram_rdata;
  assign _29441_[3:0] = _tmp_692;
  assign _29442_[3:0] = _stream_conv2d_16_source_35_source_ram_rdata;
  assign _29450_[3:0] = _tmp_706;
  assign _29451_[3:0] = _stream_conv2d_16_source_36_source_ram_rdata;
  assign _29452_[0] = _stream_conv2d_16_start_flag;
  assign RESETN_inv_buf = _RESETN_inv_2;
  assign __delay_data_1007 = __delay_data_1262;
  assign __delay_data_1008 = __delay_data_1263;
  assign __delay_data_1009 = __delay_data_1264;
  assign __delay_data_1010 = __delay_data_1265;
  assign __delay_data_1011 = __delay_data_1266;
  assign __delay_data_1012 = __delay_data_1267;
  assign __delay_data_1013 = __delay_data_1021;
  assign __delay_data_1014 = __delay_data_1022;
  assign __delay_data_1015 = __delay_data_1023;
  assign __delay_data_1017 = __delay_data_1021;
  assign __delay_data_1018 = __delay_data_1022;
  assign __delay_data_1019 = __delay_data_1023;
  assign __delay_data_1025 = __delay_data_1234;
  assign __delay_data_1026 = __delay_data_1235;
  assign __delay_data_1027 = __delay_data_1236;
  assign __delay_data_1028 = __delay_data_1237;
  assign __delay_data_1029 = __delay_data_1238;
  assign __delay_data_1030 = __delay_data_1239;
  assign __delay_data_1031 = __delay_data_1240;
  assign __delay_data_1033 = __delay_data_1241;
  assign __delay_data_1034 = __delay_data_1242;
  assign __delay_data_1035 = __delay_data_1243;
  assign __delay_data_1036 = __delay_data_1244;
  assign __delay_data_1037 = __delay_data_1245;
  assign __delay_data_1055 = __delay_data_1262;
  assign __delay_data_1056 = __delay_data_1263;
  assign __delay_data_1057 = __delay_data_1264;
  assign __delay_data_1058 = __delay_data_1265;
  assign __delay_data_1059 = __delay_data_1266;
  assign __delay_data_1060 = __delay_data_1267;
  assign __delay_data_1061 = __delay_data_1234;
  assign __delay_data_1062 = __delay_data_1235;
  assign __delay_data_1063 = __delay_data_1236;
  assign __delay_data_1064 = __delay_data_1237;
  assign __delay_data_1065 = __delay_data_1238;
  assign __delay_data_1066 = __delay_data_1239;
  assign __delay_data_1067 = __delay_data_1240;
  assign __delay_data_1069 = __delay_data_1241;
  assign __delay_data_1070 = __delay_data_1242;
  assign __delay_data_1071 = __delay_data_1243;
  assign __delay_data_1072 = __delay_data_1244;
  assign __delay_data_1073 = __delay_data_1245;
  assign __delay_data_1090 = __delay_data_1262;
  assign __delay_data_1091 = __delay_data_1263;
  assign __delay_data_1092 = __delay_data_1264;
  assign __delay_data_1093 = __delay_data_1265;
  assign __delay_data_1094 = __delay_data_1266;
  assign __delay_data_1095 = __delay_data_1267;
  assign __delay_data_1096 = __delay_data_1234;
  assign __delay_data_1097 = __delay_data_1235;
  assign __delay_data_1098 = __delay_data_1236;
  assign __delay_data_1099 = __delay_data_1237;
  assign __delay_data_1100 = __delay_data_1238;
  assign __delay_data_1101 = __delay_data_1239;
  assign __delay_data_1102 = __delay_data_1240;
  assign __delay_data_1104 = __delay_data_1241;
  assign __delay_data_1105 = __delay_data_1242;
  assign __delay_data_1106 = __delay_data_1243;
  assign __delay_data_1107 = __delay_data_1244;
  assign __delay_data_1108 = __delay_data_1245;
  assign __delay_data_1125 = __delay_data_1262;
  assign __delay_data_1126 = __delay_data_1263;
  assign __delay_data_1127 = __delay_data_1264;
  assign __delay_data_1128 = __delay_data_1265;
  assign __delay_data_1129 = __delay_data_1266;
  assign __delay_data_1130 = __delay_data_1267;
  assign __delay_data_1131 = __delay_data_1234;
  assign __delay_data_1132 = __delay_data_1235;
  assign __delay_data_1133 = __delay_data_1236;
  assign __delay_data_1134 = __delay_data_1237;
  assign __delay_data_1135 = __delay_data_1238;
  assign __delay_data_1136 = __delay_data_1239;
  assign __delay_data_1137 = __delay_data_1240;
  assign __delay_data_1139 = __delay_data_1241;
  assign __delay_data_1140 = __delay_data_1242;
  assign __delay_data_1141 = __delay_data_1243;
  assign __delay_data_1142 = __delay_data_1244;
  assign __delay_data_1143 = __delay_data_1245;
  assign __delay_data_1160 = __delay_data_1262;
  assign __delay_data_1161 = __delay_data_1263;
  assign __delay_data_1162 = __delay_data_1264;
  assign __delay_data_1163 = __delay_data_1265;
  assign __delay_data_1164 = __delay_data_1266;
  assign __delay_data_1165 = __delay_data_1267;
  assign __delay_data_1166 = __delay_data_1234;
  assign __delay_data_1167 = __delay_data_1235;
  assign __delay_data_1168 = __delay_data_1236;
  assign __delay_data_1169 = __delay_data_1237;
  assign __delay_data_1170 = __delay_data_1238;
  assign __delay_data_1171 = __delay_data_1239;
  assign __delay_data_1172 = __delay_data_1240;
  assign __delay_data_1173 = __delay_data_1241;
  assign __delay_data_1174 = __delay_data_1242;
  assign __delay_data_1175 = __delay_data_1243;
  assign __delay_data_1176 = __delay_data_1244;
  assign __delay_data_1177 = __delay_data_1245;
  assign __delay_data_1194 = __delay_data_1262;
  assign __delay_data_1195 = __delay_data_1263;
  assign __delay_data_1196 = __delay_data_1264;
  assign __delay_data_1197 = __delay_data_1265;
  assign __delay_data_1198 = __delay_data_1266;
  assign __delay_data_1199 = __delay_data_1267;
  assign __delay_data_1200 = __delay_data_1234;
  assign __delay_data_1201 = __delay_data_1235;
  assign __delay_data_1202 = __delay_data_1236;
  assign __delay_data_1203 = __delay_data_1237;
  assign __delay_data_1204 = __delay_data_1238;
  assign __delay_data_1205 = __delay_data_1239;
  assign __delay_data_1206 = __delay_data_1240;
  assign __delay_data_1207 = __delay_data_1241;
  assign __delay_data_1208 = __delay_data_1242;
  assign __delay_data_1209 = __delay_data_1243;
  assign __delay_data_1210 = __delay_data_1244;
  assign __delay_data_1211 = __delay_data_1245;
  assign __delay_data_1228 = __delay_data_1262;
  assign __delay_data_1229 = __delay_data_1263;
  assign __delay_data_1230 = __delay_data_1264;
  assign __delay_data_1231 = __delay_data_1265;
  assign __delay_data_1232 = __delay_data_1266;
  assign __delay_data_1233 = __delay_data_1267;
  assign __delay_data_1397 = __delay_data_1528;
  assign __delay_data_1398 = __delay_data_1602;
  assign __delay_data_1399 = __delay_data_1603;
  assign __delay_data_1400 = __delay_data_1604;
  assign __delay_data_1401 = __delay_data_1605;
  assign __delay_data_1402 = __delay_data_1606;
  assign __delay_data_1403 = __delay_data_1607;
  assign __delay_data_1404 = __delay_data_1608;
  assign __delay_data_1405 = __delay_data_1609;
  assign __delay_data_1406 = __delay_data_1610;
  assign __delay_data_1407 = __delay_data_1611;
  assign __delay_data_1408 = __delay_data_1612;
  assign __delay_data_1409 = __delay_data_1613;
  assign __delay_data_1410 = __delay_data_1614;
  assign __delay_data_899 = __delay_data_1021;
  assign __delay_data_902 = __delay_data_1022;
  assign __delay_data_903 = __delay_data_1023;
  assign __delay_data_908 = __delay_data_1021;
  assign __delay_data_911 = __delay_data_1022;
  assign __delay_data_912 = __delay_data_1023;
  assign __delay_data_917 = __delay_data_1021;
  assign __delay_data_920 = __delay_data_1022;
  assign __delay_data_921 = __delay_data_1023;
  assign __delay_data_925 = __delay_data_1234;
  assign __delay_data_926 = __delay_data_1235;
  assign __delay_data_927 = __delay_data_1236;
  assign __delay_data_928 = __delay_data_1237;
  assign __delay_data_929 = __delay_data_1238;
  assign __delay_data_930 = __delay_data_1239;
  assign __delay_data_931 = __delay_data_1240;
  assign __delay_data_933 = __delay_data_1241;
  assign __delay_data_934 = __delay_data_1242;
  assign __delay_data_935 = __delay_data_1243;
  assign __delay_data_936 = __delay_data_1244;
  assign __delay_data_937 = __delay_data_1245;
  assign __delay_data_956 = __delay_data_1262;
  assign __delay_data_957 = __delay_data_1263;
  assign __delay_data_958 = __delay_data_1264;
  assign __delay_data_959 = __delay_data_1265;
  assign __delay_data_960 = __delay_data_1266;
  assign __delay_data_961 = __delay_data_1267;
  assign __delay_data_962 = __delay_data_1021;
  assign __delay_data_964 = __delay_data_1022;
  assign __delay_data_965 = __delay_data_1023;
  assign __delay_data_967 = __delay_data_1021;
  assign __delay_data_969 = __delay_data_1022;
  assign __delay_data_970 = __delay_data_1023;
  assign __delay_data_972 = __delay_data_1021;
  assign __delay_data_974 = __delay_data_1022;
  assign __delay_data_975 = __delay_data_1023;
  assign __delay_data_977 = __delay_data_1234;
  assign __delay_data_978 = __delay_data_1235;
  assign __delay_data_979 = __delay_data_1236;
  assign __delay_data_980 = __delay_data_1237;
  assign __delay_data_981 = __delay_data_1238;
  assign __delay_data_982 = __delay_data_1239;
  assign __delay_data_983 = __delay_data_1240;
  assign __delay_data_985 = __delay_data_1241;
  assign __delay_data_986 = __delay_data_1242;
  assign __delay_data_987 = __delay_data_1243;
  assign __delay_data_988 = __delay_data_1244;
  assign __delay_data_989 = __delay_data_1245;
  assign __muladd_data_103 = __muladd_madd_odata_reg_103;
  assign __muladd_data_120 = __muladd_madd_odata_reg_120;
  assign __muladd_data_137 = __muladd_madd_odata_reg_137;
  assign __muladd_data_154 = __muladd_madd_odata_reg_154;
  assign __muladd_data_171 = __muladd_madd_odata_reg_171;
  assign __muladd_data_188 = __muladd_madd_odata_reg_188;
  assign __muladd_data_205 = __muladd_madd_odata_reg_205;
  assign __muladd_data_69 = __muladd_madd_odata_reg_69;
  assign __muladd_data_86 = __muladd_madd_odata_reg_86;
  assign \__muladd_madd_103.CLK  = CLK;
  assign \__muladd_madd_103.a  = __delay_data_630;
  assign \__muladd_madd_103.b  = __delay_data_633;
  assign \__muladd_madd_103.c  = _cond_data_101;
  assign \__muladd_madd_103.d  = \__muladd_madd_103.madd._pipe_madd1 ;
  assign \__muladd_madd_103.madd.CLK  = CLK;
  assign \__muladd_madd_103.madd.a  = __delay_data_630;
  assign \__muladd_madd_103.madd.b  = __delay_data_633;
  assign \__muladd_madd_103.madd.c  = _cond_data_101;
  assign \__muladd_madd_103.madd.d  = \__muladd_madd_103.madd._pipe_madd1 ;
  assign \__muladd_madd_103.madd.update  = 1'h1;
  assign \__muladd_madd_103.update  = 1'h1;
  assign \__muladd_madd_120.CLK  = CLK;
  assign \__muladd_madd_120.a  = __delay_data_647;
  assign \__muladd_madd_120.b  = __delay_data_650;
  assign \__muladd_madd_120.c  = _cond_data_118;
  assign \__muladd_madd_120.d  = \__muladd_madd_120.madd._pipe_madd1 ;
  assign \__muladd_madd_120.madd.CLK  = CLK;
  assign \__muladd_madd_120.madd.a  = __delay_data_647;
  assign \__muladd_madd_120.madd.b  = __delay_data_650;
  assign \__muladd_madd_120.madd.c  = _cond_data_118;
  assign \__muladd_madd_120.madd.d  = \__muladd_madd_120.madd._pipe_madd1 ;
  assign \__muladd_madd_120.madd.update  = 1'h1;
  assign \__muladd_madd_120.update  = 1'h1;
  assign \__muladd_madd_137.CLK  = CLK;
  assign \__muladd_madd_137.a  = __delay_data_664;
  assign \__muladd_madd_137.b  = __delay_data_667;
  assign \__muladd_madd_137.c  = _cond_data_135;
  assign \__muladd_madd_137.d  = \__muladd_madd_137.madd._pipe_madd1 ;
  assign \__muladd_madd_137.madd.CLK  = CLK;
  assign \__muladd_madd_137.madd.a  = __delay_data_664;
  assign \__muladd_madd_137.madd.b  = __delay_data_667;
  assign \__muladd_madd_137.madd.c  = _cond_data_135;
  assign \__muladd_madd_137.madd.d  = \__muladd_madd_137.madd._pipe_madd1 ;
  assign \__muladd_madd_137.madd.update  = 1'h1;
  assign \__muladd_madd_137.update  = 1'h1;
  assign \__muladd_madd_154.CLK  = CLK;
  assign \__muladd_madd_154.a  = __delay_data_681;
  assign \__muladd_madd_154.b  = __delay_data_684;
  assign \__muladd_madd_154.c  = _cond_data_152;
  assign \__muladd_madd_154.d  = \__muladd_madd_154.madd._pipe_madd1 ;
  assign \__muladd_madd_154.madd.CLK  = CLK;
  assign \__muladd_madd_154.madd.a  = __delay_data_681;
  assign \__muladd_madd_154.madd.b  = __delay_data_684;
  assign \__muladd_madd_154.madd.c  = _cond_data_152;
  assign \__muladd_madd_154.madd.d  = \__muladd_madd_154.madd._pipe_madd1 ;
  assign \__muladd_madd_154.madd.update  = 1'h1;
  assign \__muladd_madd_154.update  = 1'h1;
  assign \__muladd_madd_171.CLK  = CLK;
  assign \__muladd_madd_171.a  = __delay_data_698;
  assign \__muladd_madd_171.b  = __delay_data_701;
  assign \__muladd_madd_171.c  = _cond_data_169;
  assign \__muladd_madd_171.d  = \__muladd_madd_171.madd._pipe_madd1 ;
  assign \__muladd_madd_171.madd.CLK  = CLK;
  assign \__muladd_madd_171.madd.a  = __delay_data_698;
  assign \__muladd_madd_171.madd.b  = __delay_data_701;
  assign \__muladd_madd_171.madd.c  = _cond_data_169;
  assign \__muladd_madd_171.madd.d  = \__muladd_madd_171.madd._pipe_madd1 ;
  assign \__muladd_madd_171.madd.update  = 1'h1;
  assign \__muladd_madd_171.update  = 1'h1;
  assign \__muladd_madd_188.CLK  = CLK;
  assign \__muladd_madd_188.a  = __delay_data_715;
  assign \__muladd_madd_188.b  = __delay_data_718;
  assign \__muladd_madd_188.c  = _cond_data_186;
  assign \__muladd_madd_188.d  = \__muladd_madd_188.madd._pipe_madd1 ;
  assign \__muladd_madd_188.madd.CLK  = CLK;
  assign \__muladd_madd_188.madd.a  = __delay_data_715;
  assign \__muladd_madd_188.madd.b  = __delay_data_718;
  assign \__muladd_madd_188.madd.c  = _cond_data_186;
  assign \__muladd_madd_188.madd.d  = \__muladd_madd_188.madd._pipe_madd1 ;
  assign \__muladd_madd_188.madd.update  = 1'h1;
  assign \__muladd_madd_188.update  = 1'h1;
  assign \__muladd_madd_205.CLK  = CLK;
  assign \__muladd_madd_205.a  = __delay_data_732;
  assign \__muladd_madd_205.b  = __delay_data_735;
  assign \__muladd_madd_205.c  = _cond_data_203;
  assign \__muladd_madd_205.d  = \__muladd_madd_205.madd._pipe_madd1 ;
  assign \__muladd_madd_205.madd.CLK  = CLK;
  assign \__muladd_madd_205.madd.a  = __delay_data_732;
  assign \__muladd_madd_205.madd.b  = __delay_data_735;
  assign \__muladd_madd_205.madd.c  = _cond_data_203;
  assign \__muladd_madd_205.madd.d  = \__muladd_madd_205.madd._pipe_madd1 ;
  assign \__muladd_madd_205.madd.update  = 1'h1;
  assign \__muladd_madd_205.update  = 1'h1;
  assign \__muladd_madd_69.CLK  = CLK;
  assign \__muladd_madd_69.a  = __delay_data_596;
  assign \__muladd_madd_69.b  = __delay_data_599;
  assign \__muladd_madd_69.c  = _cond_data_67;
  assign \__muladd_madd_69.d  = \__muladd_madd_69.madd._pipe_madd1 ;
  assign \__muladd_madd_69.madd.CLK  = CLK;
  assign \__muladd_madd_69.madd.a  = __delay_data_596;
  assign \__muladd_madd_69.madd.b  = __delay_data_599;
  assign \__muladd_madd_69.madd.c  = _cond_data_67;
  assign \__muladd_madd_69.madd.d  = \__muladd_madd_69.madd._pipe_madd1 ;
  assign \__muladd_madd_69.madd.update  = 1'h1;
  assign \__muladd_madd_69.update  = 1'h1;
  assign \__muladd_madd_86.CLK  = CLK;
  assign \__muladd_madd_86.a  = __delay_data_613;
  assign \__muladd_madd_86.b  = __delay_data_616;
  assign \__muladd_madd_86.c  = _cond_data_84;
  assign \__muladd_madd_86.d  = \__muladd_madd_86.madd._pipe_madd1 ;
  assign \__muladd_madd_86.madd.CLK  = CLK;
  assign \__muladd_madd_86.madd.a  = __delay_data_613;
  assign \__muladd_madd_86.madd.b  = __delay_data_616;
  assign \__muladd_madd_86.madd.c  = _cond_data_84;
  assign \__muladd_madd_86.madd.d  = \__muladd_madd_86.madd._pipe_madd1 ;
  assign \__muladd_madd_86.madd.update  = 1'h1;
  assign \__muladd_madd_86.update  = 1'h1;
  assign __muladd_madd_odata_103 = \__muladd_madd_103.madd._pipe_madd1 ;
  assign __muladd_madd_odata_120 = \__muladd_madd_120.madd._pipe_madd1 ;
  assign __muladd_madd_odata_137 = \__muladd_madd_137.madd._pipe_madd1 ;
  assign __muladd_madd_odata_154 = \__muladd_madd_154.madd._pipe_madd1 ;
  assign __muladd_madd_odata_171 = \__muladd_madd_171.madd._pipe_madd1 ;
  assign __muladd_madd_odata_188 = \__muladd_madd_188.madd._pipe_madd1 ;
  assign __muladd_madd_odata_205 = \__muladd_madd_205.madd._pipe_madd1 ;
  assign __muladd_madd_odata_69 = \__muladd_madd_69.madd._pipe_madd1 ;
  assign __muladd_madd_odata_86 = \__muladd_madd_86.madd._pipe_madd1 ;
  assign __muladd_madd_update_103 = 1'h1;
  assign __muladd_madd_update_120 = 1'h1;
  assign __muladd_madd_update_137 = 1'h1;
  assign __muladd_madd_update_154 = 1'h1;
  assign __muladd_madd_update_171 = 1'h1;
  assign __muladd_madd_update_188 = 1'h1;
  assign __muladd_madd_update_205 = 1'h1;
  assign __muladd_madd_update_69 = 1'h1;
  assign __muladd_madd_update_86 = 1'h1;
  assign __reduce_max_13_data_sink_wenable = 1'h0;
  assign __reduce_max_13_fsm = 0;
  assign __reduce_max_13_valid_sink_wenable = 1'h0;
  assign __reduce_max_13_x_idle = 1'h1;
  assign __reduce_max_13_x_source_ram_rvalid = 1'h0;
  assign __stream_seq_14_cond_2_1 = __set_flag_710_1;
  assign __stream_seq_14_cond_2_10 = __set_flag_710_10;
  assign __stream_seq_14_cond_2_11 = __set_flag_710_11;
  assign __stream_seq_14_cond_2_12 = __set_flag_710_12;
  assign __stream_seq_14_cond_2_13 = __set_flag_710_13;
  assign __stream_seq_14_cond_2_14 = __set_flag_710_14;
  assign __stream_seq_14_cond_2_15 = __set_flag_710_15;
  assign __stream_seq_14_cond_2_16 = __set_flag_710_16;
  assign __stream_seq_14_cond_2_17 = __set_flag_710_17;
  assign __stream_seq_14_cond_2_18 = __set_flag_710_18;
  assign __stream_seq_14_cond_2_19 = __set_flag_710_19;
  assign __stream_seq_14_cond_2_2 = __set_flag_710_2;
  assign __stream_seq_14_cond_2_20 = __set_flag_710_20;
  assign __stream_seq_14_cond_2_21 = __set_flag_710_21;
  assign __stream_seq_14_cond_2_22 = __set_flag_710_22;
  assign __stream_seq_14_cond_2_23 = __set_flag_710_23;
  assign __stream_seq_14_cond_2_24 = __set_flag_710_24;
  assign __stream_seq_14_cond_2_25 = __set_flag_710_25;
  assign __stream_seq_14_cond_2_26 = __set_flag_710_26;
  assign __stream_seq_14_cond_2_27 = __set_flag_710_27;
  assign __stream_seq_14_cond_2_28 = __set_flag_710_28;
  assign __stream_seq_14_cond_2_29 = __set_flag_710_29;
  assign __stream_seq_14_cond_2_3 = __set_flag_710_3;
  assign __stream_seq_14_cond_2_30 = __set_flag_710_30;
  assign __stream_seq_14_cond_2_31 = __set_flag_710_31;
  assign __stream_seq_14_cond_2_32 = __set_flag_710_32;
  assign __stream_seq_14_cond_2_33 = __set_flag_710_33;
  assign __stream_seq_14_cond_2_34 = __set_flag_710_34;
  assign __stream_seq_14_cond_2_35 = __set_flag_710_35;
  assign __stream_seq_14_cond_2_36 = __set_flag_710_36;
  assign __stream_seq_14_cond_2_37 = __set_flag_710_37;
  assign __stream_seq_14_cond_2_38 = __set_flag_710_38;
  assign __stream_seq_14_cond_2_39 = __set_flag_710_39;
  assign __stream_seq_14_cond_2_4 = __set_flag_710_4;
  assign __stream_seq_14_cond_2_40 = __set_flag_710_40;
  assign __stream_seq_14_cond_2_41 = __set_flag_710_41;
  assign __stream_seq_14_cond_2_42 = __set_flag_710_42;
  assign __stream_seq_14_cond_2_43 = __set_flag_710_43;
  assign __stream_seq_14_cond_2_44 = __set_flag_710_44;
  assign __stream_seq_14_cond_2_45 = __set_flag_710_45;
  assign __stream_seq_14_cond_2_5 = __set_flag_710_5;
  assign __stream_seq_14_cond_2_6 = __set_flag_710_6;
  assign __stream_seq_14_cond_2_7 = __set_flag_710_7;
  assign __stream_seq_14_cond_2_8 = __set_flag_710_8;
  assign __stream_seq_14_cond_2_9 = __set_flag_710_9;
  assign __stream_seq_15_cond_2_1 = __set_flag_1036_1;
  assign __stream_seq_15_cond_2_2 = __set_flag_1036_2;
  assign __stream_seq_15_cond_2_3 = __set_flag_1036_3;
  assign __stream_seq_15_cond_2_4 = __set_flag_1036_4;
  assign __stream_seq_15_cond_2_5 = __set_flag_1036_5;
  assign __stream_seq_15_cond_2_6 = __set_flag_1036_6;
  assign __stream_seq_15_cond_2_7 = __set_flag_1036_7;
  assign __stream_seq_15_cond_2_8 = __set_flag_1036_8;
  assign __stream_seq_15_cond_2_9 = __set_flag_1036_9;
  assign __stream_seq_16_cond_2_1 = __set_flag_1224_1;
  assign __stream_seq_16_cond_2_10 = __set_flag_1224_10;
  assign __stream_seq_16_cond_2_11 = __set_flag_1224_11;
  assign __stream_seq_16_cond_2_12 = __set_flag_1224_12;
  assign __stream_seq_16_cond_2_13 = __set_flag_1224_13;
  assign __stream_seq_16_cond_2_14 = __set_flag_1224_14;
  assign __stream_seq_16_cond_2_15 = __set_flag_1224_15;
  assign __stream_seq_16_cond_2_16 = __set_flag_1224_16;
  assign __stream_seq_16_cond_2_17 = __set_flag_1224_17;
  assign __stream_seq_16_cond_2_18 = __set_flag_1224_18;
  assign __stream_seq_16_cond_2_19 = __set_flag_1224_19;
  assign __stream_seq_16_cond_2_2 = __set_flag_1224_2;
  assign __stream_seq_16_cond_2_20 = __set_flag_1224_20;
  assign __stream_seq_16_cond_2_21 = __set_flag_1224_21;
  assign __stream_seq_16_cond_2_22 = __set_flag_1224_22;
  assign __stream_seq_16_cond_2_23 = __set_flag_1224_23;
  assign __stream_seq_16_cond_2_24 = __set_flag_1224_24;
  assign __stream_seq_16_cond_2_25 = __set_flag_1224_25;
  assign __stream_seq_16_cond_2_26 = __set_flag_1224_26;
  assign __stream_seq_16_cond_2_27 = __set_flag_1224_27;
  assign __stream_seq_16_cond_2_28 = __set_flag_1224_28;
  assign __stream_seq_16_cond_2_29 = __set_flag_1224_29;
  assign __stream_seq_16_cond_2_3 = __set_flag_1224_3;
  assign __stream_seq_16_cond_2_30 = __set_flag_1224_30;
  assign __stream_seq_16_cond_2_31 = __set_flag_1224_31;
  assign __stream_seq_16_cond_2_32 = __set_flag_1224_32;
  assign __stream_seq_16_cond_2_33 = __set_flag_1224_33;
  assign __stream_seq_16_cond_2_34 = __set_flag_1224_34;
  assign __stream_seq_16_cond_2_35 = __set_flag_1224_35;
  assign __stream_seq_16_cond_2_36 = __set_flag_1224_36;
  assign __stream_seq_16_cond_2_37 = __set_flag_1224_37;
  assign __stream_seq_16_cond_2_38 = __set_flag_1224_38;
  assign __stream_seq_16_cond_2_39 = __set_flag_1224_39;
  assign __stream_seq_16_cond_2_4 = __set_flag_1224_4;
  assign __stream_seq_16_cond_2_40 = __set_flag_1224_40;
  assign __stream_seq_16_cond_2_41 = __set_flag_1224_41;
  assign __stream_seq_16_cond_2_5 = __set_flag_1224_5;
  assign __stream_seq_16_cond_2_6 = __set_flag_1224_6;
  assign __stream_seq_16_cond_2_7 = __set_flag_1224_7;
  assign __stream_seq_16_cond_2_8 = __set_flag_1224_8;
  assign __stream_seq_16_cond_2_9 = __set_flag_1224_9;
  assign __substreamoutput_data_608 = __substreamoutput_data_876;
  assign __substreamoutput_data_760 = __substreamoutput_data_881;
  assign __substreamoutput_data_761 = __substreamoutput_data_882;
  assign __substreamoutput_data_771 = __substreamoutput_data_886;
  assign __tmp_1035_1 = _ram_w8_l2048_id1_0_cond_4_1;
  assign __tmp_1040_1 = __tmp_1046_1;
  assign __tmp_1040_2 = __tmp_1046_2;
  assign __tmp_1040_3 = __tmp_1046_3;
  assign __tmp_1040_4 = __tmp_1046_4;
  assign __tmp_1040_5 = __tmp_1046_5;
  assign __tmp_1042_1 = __tmp_1046_1;
  assign __tmp_1042_2 = __tmp_1046_2;
  assign __tmp_1042_3 = __tmp_1046_3;
  assign __tmp_1042_4 = __tmp_1046_4;
  assign __tmp_1042_5 = __tmp_1046_5;
  assign __tmp_1042_6 = __tmp_1046_6;
  assign __tmp_1042_7 = __tmp_1046_7;
  assign __tmp_1044_1 = __tmp_1046_1;
  assign __tmp_1044_2 = __tmp_1046_2;
  assign __tmp_1044_3 = __tmp_1046_3;
  assign __tmp_1044_4 = __tmp_1046_4;
  assign __tmp_1044_5 = __tmp_1046_5;
  assign __tmp_1044_6 = __tmp_1046_6;
  assign __tmp_1044_7 = __tmp_1046_7;
  assign __tmp_1048_1 = __tmp_1060_1;
  assign __tmp_1050_1 = __tmp_1060_1;
  assign __tmp_1050_2 = __tmp_1060_2;
  assign __tmp_1050_3 = __tmp_1060_3;
  assign __tmp_1050_4 = __tmp_1060_4;
  assign __tmp_1050_5 = __tmp_1060_5;
  assign __tmp_1052_1 = __tmp_1060_1;
  assign __tmp_1052_2 = __tmp_1060_2;
  assign __tmp_1052_3 = __tmp_1060_3;
  assign __tmp_1052_4 = __tmp_1060_4;
  assign __tmp_1054_1 = __tmp_1060_1;
  assign __tmp_1054_2 = __tmp_1060_2;
  assign __tmp_1054_3 = __tmp_1060_3;
  assign __tmp_1054_4 = __tmp_1060_4;
  assign __tmp_1056_1 = __tmp_1060_1;
  assign __tmp_1056_2 = __tmp_1060_2;
  assign __tmp_1056_3 = __tmp_1060_3;
  assign __tmp_1056_4 = __tmp_1060_4;
  assign __tmp_1056_5 = __tmp_1060_5;
  assign __tmp_1058_1 = __tmp_1060_1;
  assign __tmp_1058_2 = __tmp_1060_2;
  assign __tmp_1058_3 = __tmp_1060_3;
  assign __tmp_1058_4 = __tmp_1060_4;
  assign __tmp_1058_5 = __tmp_1060_5;
  assign __tmp_1062_1 = __tmp_1060_1;
  assign __tmp_1062_10 = __tmp_1068_10;
  assign __tmp_1062_2 = __tmp_1060_2;
  assign __tmp_1062_3 = __tmp_1060_3;
  assign __tmp_1062_4 = __tmp_1060_4;
  assign __tmp_1062_5 = __tmp_1060_5;
  assign __tmp_1062_6 = __tmp_1070_6;
  assign __tmp_1062_7 = __tmp_1068_7;
  assign __tmp_1062_8 = __tmp_1068_8;
  assign __tmp_1062_9 = __tmp_1068_9;
  assign __tmp_1064_1 = __tmp_1060_1;
  assign __tmp_1064_10 = __tmp_1068_10;
  assign __tmp_1064_2 = __tmp_1060_2;
  assign __tmp_1064_3 = __tmp_1060_3;
  assign __tmp_1064_4 = __tmp_1060_4;
  assign __tmp_1064_5 = __tmp_1060_5;
  assign __tmp_1064_6 = __tmp_1070_6;
  assign __tmp_1064_7 = __tmp_1068_7;
  assign __tmp_1064_8 = __tmp_1068_8;
  assign __tmp_1064_9 = __tmp_1068_9;
  assign __tmp_1066_1 = __tmp_1060_1;
  assign __tmp_1066_10 = __tmp_1068_10;
  assign __tmp_1066_2 = __tmp_1060_2;
  assign __tmp_1066_3 = __tmp_1060_3;
  assign __tmp_1066_4 = __tmp_1060_4;
  assign __tmp_1066_5 = __tmp_1060_5;
  assign __tmp_1066_6 = __tmp_1070_6;
  assign __tmp_1066_7 = __tmp_1068_7;
  assign __tmp_1066_8 = __tmp_1068_8;
  assign __tmp_1066_9 = __tmp_1068_9;
  assign __tmp_1068_1 = __tmp_1060_1;
  assign __tmp_1068_2 = __tmp_1060_2;
  assign __tmp_1068_3 = __tmp_1060_3;
  assign __tmp_1068_4 = __tmp_1060_4;
  assign __tmp_1068_5 = __tmp_1060_5;
  assign __tmp_1068_6 = __tmp_1070_6;
  assign __tmp_1070_1 = __tmp_1060_1;
  assign __tmp_1070_2 = __tmp_1060_2;
  assign __tmp_1070_3 = __tmp_1060_3;
  assign __tmp_1070_4 = __tmp_1060_4;
  assign __tmp_1070_5 = __tmp_1060_5;
  assign __tmp_1178_1 = _ram_w8_l2048_id2_0_cond_6_1;
  assign __tmp_1189_1 = _ram_w8_l2048_id0_3_cond_5_1;
  assign __tmp_1209_1 = _ram_w8_l2048_id3_0_cond_5_1;
  assign __tmp_1227_1 = __tmp_1249_1;
  assign __tmp_1227_2 = __tmp_1249_2;
  assign __tmp_1227_3 = __tmp_1249_3;
  assign __tmp_1227_4 = __tmp_1249_4;
  assign __tmp_1227_5 = __tmp_1249_5;
  assign __tmp_1229_1 = __tmp_1249_1;
  assign __tmp_1229_2 = __tmp_1249_2;
  assign __tmp_1229_3 = __tmp_1249_3;
  assign __tmp_1229_4 = __tmp_1249_4;
  assign __tmp_1229_5 = __tmp_1249_5;
  assign __tmp_1229_6 = __tmp_1249_6;
  assign __tmp_1229_7 = __tmp_1249_7;
  assign __tmp_1229_8 = __tmp_1249_8;
  assign __tmp_1231_1 = __tmp_1249_1;
  assign __tmp_1231_2 = __tmp_1249_2;
  assign __tmp_1231_3 = __tmp_1249_3;
  assign __tmp_1231_4 = __tmp_1249_4;
  assign __tmp_1231_5 = __tmp_1249_5;
  assign __tmp_1231_6 = __tmp_1249_6;
  assign __tmp_1231_7 = __tmp_1249_7;
  assign __tmp_1231_8 = __tmp_1249_8;
  assign __tmp_1233_1 = __tmp_1249_1;
  assign __tmp_1233_2 = __tmp_1249_2;
  assign __tmp_1233_3 = __tmp_1249_3;
  assign __tmp_1233_4 = __tmp_1249_4;
  assign __tmp_1233_5 = __tmp_1249_5;
  assign __tmp_1233_6 = __tmp_1249_6;
  assign __tmp_1233_7 = __tmp_1249_7;
  assign __tmp_1233_8 = __tmp_1249_8;
  assign __tmp_1235_1 = __tmp_1249_1;
  assign __tmp_1235_10 = __tmp_1249_10;
  assign __tmp_1235_11 = __tmp_1249_11;
  assign __tmp_1235_12 = __tmp_1249_12;
  assign __tmp_1235_13 = __tmp_1249_13;
  assign __tmp_1235_14 = __tmp_1249_14;
  assign __tmp_1235_15 = __tmp_1249_15;
  assign __tmp_1235_16 = __tmp_1249_16;
  assign __tmp_1235_17 = __tmp_1249_17;
  assign __tmp_1235_18 = __tmp_1249_18;
  assign __tmp_1235_2 = __tmp_1249_2;
  assign __tmp_1235_3 = __tmp_1249_3;
  assign __tmp_1235_4 = __tmp_1249_4;
  assign __tmp_1235_5 = __tmp_1249_5;
  assign __tmp_1235_6 = __tmp_1249_6;
  assign __tmp_1235_7 = __tmp_1249_7;
  assign __tmp_1235_8 = __tmp_1249_8;
  assign __tmp_1235_9 = __tmp_1249_9;
  assign __tmp_1237_1 = __tmp_1249_1;
  assign __tmp_1237_10 = __tmp_1249_10;
  assign __tmp_1237_11 = __tmp_1249_11;
  assign __tmp_1237_12 = __tmp_1249_12;
  assign __tmp_1237_13 = __tmp_1249_13;
  assign __tmp_1237_14 = __tmp_1249_14;
  assign __tmp_1237_15 = __tmp_1249_15;
  assign __tmp_1237_16 = __tmp_1249_16;
  assign __tmp_1237_17 = __tmp_1249_17;
  assign __tmp_1237_18 = __tmp_1249_18;
  assign __tmp_1237_19 = __tmp_1249_19;
  assign __tmp_1237_2 = __tmp_1249_2;
  assign __tmp_1237_20 = __tmp_1249_20;
  assign __tmp_1237_21 = __tmp_1249_21;
  assign __tmp_1237_22 = __tmp_1249_22;
  assign __tmp_1237_3 = __tmp_1249_3;
  assign __tmp_1237_4 = __tmp_1249_4;
  assign __tmp_1237_5 = __tmp_1249_5;
  assign __tmp_1237_6 = __tmp_1249_6;
  assign __tmp_1237_7 = __tmp_1249_7;
  assign __tmp_1237_8 = __tmp_1249_8;
  assign __tmp_1237_9 = __tmp_1249_9;
  assign __tmp_1239_1 = __tmp_1249_1;
  assign __tmp_1239_10 = __tmp_1249_10;
  assign __tmp_1239_11 = __tmp_1249_11;
  assign __tmp_1239_12 = __tmp_1249_12;
  assign __tmp_1239_13 = __tmp_1249_13;
  assign __tmp_1239_14 = __tmp_1249_14;
  assign __tmp_1239_15 = __tmp_1249_15;
  assign __tmp_1239_16 = __tmp_1249_16;
  assign __tmp_1239_17 = __tmp_1249_17;
  assign __tmp_1239_18 = __tmp_1249_18;
  assign __tmp_1239_19 = __tmp_1249_19;
  assign __tmp_1239_2 = __tmp_1249_2;
  assign __tmp_1239_20 = __tmp_1249_20;
  assign __tmp_1239_3 = __tmp_1249_3;
  assign __tmp_1239_4 = __tmp_1249_4;
  assign __tmp_1239_5 = __tmp_1249_5;
  assign __tmp_1239_6 = __tmp_1249_6;
  assign __tmp_1239_7 = __tmp_1249_7;
  assign __tmp_1239_8 = __tmp_1249_8;
  assign __tmp_1239_9 = __tmp_1249_9;
  assign __tmp_1241_1 = __tmp_1249_1;
  assign __tmp_1241_10 = __tmp_1249_10;
  assign __tmp_1241_11 = __tmp_1249_11;
  assign __tmp_1241_12 = __tmp_1249_12;
  assign __tmp_1241_13 = __tmp_1249_13;
  assign __tmp_1241_14 = __tmp_1249_14;
  assign __tmp_1241_15 = __tmp_1249_15;
  assign __tmp_1241_16 = __tmp_1249_16;
  assign __tmp_1241_17 = __tmp_1249_17;
  assign __tmp_1241_18 = __tmp_1249_18;
  assign __tmp_1241_19 = __tmp_1249_19;
  assign __tmp_1241_2 = __tmp_1249_2;
  assign __tmp_1241_20 = __tmp_1249_20;
  assign __tmp_1241_3 = __tmp_1249_3;
  assign __tmp_1241_4 = __tmp_1249_4;
  assign __tmp_1241_5 = __tmp_1249_5;
  assign __tmp_1241_6 = __tmp_1249_6;
  assign __tmp_1241_7 = __tmp_1249_7;
  assign __tmp_1241_8 = __tmp_1249_8;
  assign __tmp_1241_9 = __tmp_1249_9;
  assign __tmp_1243_1 = __tmp_1249_1;
  assign __tmp_1243_10 = __tmp_1249_10;
  assign __tmp_1243_11 = __tmp_1249_11;
  assign __tmp_1243_12 = __tmp_1249_12;
  assign __tmp_1243_13 = __tmp_1249_13;
  assign __tmp_1243_14 = __tmp_1249_14;
  assign __tmp_1243_15 = __tmp_1249_15;
  assign __tmp_1243_16 = __tmp_1249_16;
  assign __tmp_1243_17 = __tmp_1249_17;
  assign __tmp_1243_18 = __tmp_1249_18;
  assign __tmp_1243_19 = __tmp_1249_19;
  assign __tmp_1243_2 = __tmp_1249_2;
  assign __tmp_1243_20 = __tmp_1249_20;
  assign __tmp_1243_3 = __tmp_1249_3;
  assign __tmp_1243_4 = __tmp_1249_4;
  assign __tmp_1243_5 = __tmp_1249_5;
  assign __tmp_1243_6 = __tmp_1249_6;
  assign __tmp_1243_7 = __tmp_1249_7;
  assign __tmp_1243_8 = __tmp_1249_8;
  assign __tmp_1243_9 = __tmp_1249_9;
  assign __tmp_1245_1 = __tmp_1249_1;
  assign __tmp_1245_10 = __tmp_1249_10;
  assign __tmp_1245_11 = __tmp_1249_11;
  assign __tmp_1245_12 = __tmp_1249_12;
  assign __tmp_1245_13 = __tmp_1249_13;
  assign __tmp_1245_14 = __tmp_1249_14;
  assign __tmp_1245_15 = __tmp_1249_15;
  assign __tmp_1245_16 = __tmp_1249_16;
  assign __tmp_1245_17 = __tmp_1249_17;
  assign __tmp_1245_18 = __tmp_1249_18;
  assign __tmp_1245_19 = __tmp_1249_19;
  assign __tmp_1245_2 = __tmp_1249_2;
  assign __tmp_1245_20 = __tmp_1249_20;
  assign __tmp_1245_21 = __tmp_1249_21;
  assign __tmp_1245_22 = __tmp_1249_22;
  assign __tmp_1245_23 = __tmp_1249_23;
  assign __tmp_1245_24 = __tmp_1249_24;
  assign __tmp_1245_25 = __tmp_1249_25;
  assign __tmp_1245_26 = __tmp_1249_26;
  assign __tmp_1245_27 = __tmp_1249_27;
  assign __tmp_1245_28 = __tmp_1249_28;
  assign __tmp_1245_3 = __tmp_1249_3;
  assign __tmp_1245_4 = __tmp_1249_4;
  assign __tmp_1245_5 = __tmp_1249_5;
  assign __tmp_1245_6 = __tmp_1249_6;
  assign __tmp_1245_7 = __tmp_1249_7;
  assign __tmp_1245_8 = __tmp_1249_8;
  assign __tmp_1245_9 = __tmp_1249_9;
  assign __tmp_1247_1 = __tmp_1249_1;
  assign __tmp_1247_10 = __tmp_1249_10;
  assign __tmp_1247_11 = __tmp_1249_11;
  assign __tmp_1247_12 = __tmp_1249_12;
  assign __tmp_1247_13 = __tmp_1249_13;
  assign __tmp_1247_14 = __tmp_1249_14;
  assign __tmp_1247_15 = __tmp_1249_15;
  assign __tmp_1247_16 = __tmp_1249_16;
  assign __tmp_1247_17 = __tmp_1249_17;
  assign __tmp_1247_18 = __tmp_1249_18;
  assign __tmp_1247_19 = __tmp_1249_19;
  assign __tmp_1247_2 = __tmp_1249_2;
  assign __tmp_1247_20 = __tmp_1249_20;
  assign __tmp_1247_21 = __tmp_1249_21;
  assign __tmp_1247_22 = __tmp_1249_22;
  assign __tmp_1247_23 = __tmp_1249_23;
  assign __tmp_1247_24 = __tmp_1249_24;
  assign __tmp_1247_25 = __tmp_1249_25;
  assign __tmp_1247_26 = __tmp_1249_26;
  assign __tmp_1247_27 = __tmp_1249_27;
  assign __tmp_1247_28 = __tmp_1249_28;
  assign __tmp_1247_3 = __tmp_1249_3;
  assign __tmp_1247_4 = __tmp_1249_4;
  assign __tmp_1247_5 = __tmp_1249_5;
  assign __tmp_1247_6 = __tmp_1249_6;
  assign __tmp_1247_7 = __tmp_1249_7;
  assign __tmp_1247_8 = __tmp_1249_8;
  assign __tmp_1247_9 = __tmp_1249_9;
  assign __tmp_1251_1 = __tmp_1299_1;
  assign __tmp_1253_1 = __tmp_1299_1;
  assign __tmp_1253_2 = __tmp_1299_2;
  assign __tmp_1253_3 = __tmp_1299_3;
  assign __tmp_1253_4 = __tmp_1299_4;
  assign __tmp_1253_5 = __tmp_1299_5;
  assign __tmp_1255_1 = __tmp_1299_1;
  assign __tmp_1255_2 = __tmp_1299_2;
  assign __tmp_1255_3 = __tmp_1299_3;
  assign __tmp_1255_4 = __tmp_1299_4;
  assign __tmp_1255_5 = __tmp_1299_5;
  assign __tmp_1257_1 = __tmp_1299_1;
  assign __tmp_1257_2 = __tmp_1299_2;
  assign __tmp_1257_3 = __tmp_1299_3;
  assign __tmp_1257_4 = __tmp_1299_4;
  assign __tmp_1257_5 = __tmp_1299_5;
  assign __tmp_1259_1 = __tmp_1299_1;
  assign __tmp_1259_10 = __tmp_1299_10;
  assign __tmp_1259_11 = __tmp_1299_11;
  assign __tmp_1259_12 = __tmp_1299_12;
  assign __tmp_1259_2 = __tmp_1299_2;
  assign __tmp_1259_3 = __tmp_1299_3;
  assign __tmp_1259_4 = __tmp_1299_4;
  assign __tmp_1259_5 = __tmp_1299_5;
  assign __tmp_1259_6 = __tmp_1299_6;
  assign __tmp_1259_7 = __tmp_1299_7;
  assign __tmp_1259_8 = __tmp_1299_8;
  assign __tmp_1259_9 = __tmp_1299_9;
  assign __tmp_1261_1 = __tmp_1299_1;
  assign __tmp_1261_10 = __tmp_1299_10;
  assign __tmp_1261_11 = __tmp_1299_11;
  assign __tmp_1261_12 = __tmp_1299_12;
  assign __tmp_1261_2 = __tmp_1299_2;
  assign __tmp_1261_3 = __tmp_1299_3;
  assign __tmp_1261_4 = __tmp_1299_4;
  assign __tmp_1261_5 = __tmp_1299_5;
  assign __tmp_1261_6 = __tmp_1299_6;
  assign __tmp_1261_7 = __tmp_1299_7;
  assign __tmp_1261_8 = __tmp_1299_8;
  assign __tmp_1261_9 = __tmp_1299_9;
  assign __tmp_1263_1 = __tmp_1299_1;
  assign __tmp_1263_10 = __tmp_1299_10;
  assign __tmp_1263_11 = __tmp_1299_11;
  assign __tmp_1263_12 = __tmp_1299_12;
  assign __tmp_1263_2 = __tmp_1299_2;
  assign __tmp_1263_3 = __tmp_1299_3;
  assign __tmp_1263_4 = __tmp_1299_4;
  assign __tmp_1263_5 = __tmp_1299_5;
  assign __tmp_1263_6 = __tmp_1299_6;
  assign __tmp_1263_7 = __tmp_1299_7;
  assign __tmp_1263_8 = __tmp_1299_8;
  assign __tmp_1263_9 = __tmp_1299_9;
  assign __tmp_1265_1 = __tmp_1299_1;
  assign __tmp_1265_10 = __tmp_1299_10;
  assign __tmp_1265_11 = __tmp_1299_11;
  assign __tmp_1265_12 = __tmp_1299_12;
  assign __tmp_1265_13 = __tmp_1299_13;
  assign __tmp_1265_14 = __tmp_1299_14;
  assign __tmp_1265_15 = __tmp_1299_15;
  assign __tmp_1265_2 = __tmp_1299_2;
  assign __tmp_1265_3 = __tmp_1299_3;
  assign __tmp_1265_4 = __tmp_1299_4;
  assign __tmp_1265_5 = __tmp_1299_5;
  assign __tmp_1265_6 = __tmp_1299_6;
  assign __tmp_1265_7 = __tmp_1299_7;
  assign __tmp_1265_8 = __tmp_1299_8;
  assign __tmp_1265_9 = __tmp_1299_9;
  assign __tmp_1267_1 = __tmp_1299_1;
  assign __tmp_1267_2 = __tmp_1299_2;
  assign __tmp_1267_3 = __tmp_1299_3;
  assign __tmp_1267_4 = __tmp_1299_4;
  assign __tmp_1269_1 = __tmp_1299_1;
  assign __tmp_1269_2 = __tmp_1299_2;
  assign __tmp_1269_3 = __tmp_1299_3;
  assign __tmp_1269_4 = __tmp_1299_4;
  assign __tmp_1271_1 = __tmp_1299_1;
  assign __tmp_1271_2 = __tmp_1299_2;
  assign __tmp_1271_3 = __tmp_1299_3;
  assign __tmp_1271_4 = __tmp_1299_4;
  assign __tmp_1273_1 = __tmp_1299_1;
  assign __tmp_1273_10 = __tmp_1299_10;
  assign __tmp_1273_11 = __tmp_1299_11;
  assign __tmp_1273_12 = __tmp_1299_12;
  assign __tmp_1273_13 = __tmp_1299_13;
  assign __tmp_1273_14 = __tmp_1299_14;
  assign __tmp_1273_15 = __tmp_1299_15;
  assign __tmp_1273_16 = __tmp_1299_16;
  assign __tmp_1273_17 = __tmp_1299_17;
  assign __tmp_1273_18 = __tmp_1299_18;
  assign __tmp_1273_2 = __tmp_1299_2;
  assign __tmp_1273_3 = __tmp_1299_3;
  assign __tmp_1273_4 = __tmp_1299_4;
  assign __tmp_1273_5 = __tmp_1299_5;
  assign __tmp_1273_6 = __tmp_1299_6;
  assign __tmp_1273_7 = __tmp_1299_7;
  assign __tmp_1273_8 = __tmp_1299_8;
  assign __tmp_1273_9 = __tmp_1299_9;
  assign __tmp_1275_1 = __tmp_1299_1;
  assign __tmp_1275_10 = __tmp_1299_10;
  assign __tmp_1275_11 = __tmp_1299_11;
  assign __tmp_1275_12 = __tmp_1299_12;
  assign __tmp_1275_13 = __tmp_1299_13;
  assign __tmp_1275_14 = __tmp_1299_14;
  assign __tmp_1275_15 = __tmp_1299_15;
  assign __tmp_1275_16 = __tmp_1299_16;
  assign __tmp_1275_17 = __tmp_1299_17;
  assign __tmp_1275_2 = __tmp_1299_2;
  assign __tmp_1275_3 = __tmp_1299_3;
  assign __tmp_1275_4 = __tmp_1299_4;
  assign __tmp_1275_5 = __tmp_1299_5;
  assign __tmp_1275_6 = __tmp_1299_6;
  assign __tmp_1275_7 = __tmp_1299_7;
  assign __tmp_1275_8 = __tmp_1299_8;
  assign __tmp_1275_9 = __tmp_1299_9;
  assign __tmp_1277_1 = __tmp_1299_1;
  assign __tmp_1277_10 = __tmp_1299_10;
  assign __tmp_1277_11 = __tmp_1299_11;
  assign __tmp_1277_12 = __tmp_1299_12;
  assign __tmp_1277_13 = __tmp_1299_13;
  assign __tmp_1277_14 = __tmp_1299_14;
  assign __tmp_1277_15 = __tmp_1299_15;
  assign __tmp_1277_16 = __tmp_1299_16;
  assign __tmp_1277_17 = __tmp_1299_17;
  assign __tmp_1277_2 = __tmp_1299_2;
  assign __tmp_1277_3 = __tmp_1299_3;
  assign __tmp_1277_4 = __tmp_1299_4;
  assign __tmp_1277_5 = __tmp_1299_5;
  assign __tmp_1277_6 = __tmp_1299_6;
  assign __tmp_1277_7 = __tmp_1299_7;
  assign __tmp_1277_8 = __tmp_1299_8;
  assign __tmp_1277_9 = __tmp_1299_9;
  assign __tmp_1279_1 = __tmp_1299_1;
  assign __tmp_1279_10 = __tmp_1299_10;
  assign __tmp_1279_11 = __tmp_1299_11;
  assign __tmp_1279_12 = __tmp_1299_12;
  assign __tmp_1279_13 = __tmp_1299_13;
  assign __tmp_1279_14 = __tmp_1299_14;
  assign __tmp_1279_15 = __tmp_1299_15;
  assign __tmp_1279_16 = __tmp_1299_16;
  assign __tmp_1279_17 = __tmp_1299_17;
  assign __tmp_1279_2 = __tmp_1299_2;
  assign __tmp_1279_3 = __tmp_1299_3;
  assign __tmp_1279_4 = __tmp_1299_4;
  assign __tmp_1279_5 = __tmp_1299_5;
  assign __tmp_1279_6 = __tmp_1299_6;
  assign __tmp_1279_7 = __tmp_1299_7;
  assign __tmp_1279_8 = __tmp_1299_8;
  assign __tmp_1279_9 = __tmp_1299_9;
  assign __tmp_1281_1 = __tmp_1299_1;
  assign __tmp_1281_2 = __tmp_1299_2;
  assign __tmp_1281_3 = __tmp_1299_3;
  assign __tmp_1281_4 = __tmp_1299_4;
  assign __tmp_1281_5 = __tmp_1299_5;
  assign __tmp_1281_6 = __tmp_1299_6;
  assign __tmp_1281_7 = __tmp_1299_7;
  assign __tmp_1281_8 = __tmp_1299_8;
  assign __tmp_1281_9 = __tmp_1299_9;
  assign __tmp_1283_1 = __tmp_1299_1;
  assign __tmp_1283_2 = __tmp_1299_2;
  assign __tmp_1283_3 = __tmp_1299_3;
  assign __tmp_1283_4 = __tmp_1299_4;
  assign __tmp_1283_5 = __tmp_1299_5;
  assign __tmp_1283_6 = __tmp_1299_6;
  assign __tmp_1283_7 = __tmp_1299_7;
  assign __tmp_1283_8 = __tmp_1299_8;
  assign __tmp_1283_9 = __tmp_1299_9;
  assign __tmp_1285_1 = __tmp_1299_1;
  assign __tmp_1285_2 = __tmp_1299_2;
  assign __tmp_1285_3 = __tmp_1299_3;
  assign __tmp_1285_4 = __tmp_1299_4;
  assign __tmp_1285_5 = __tmp_1299_5;
  assign __tmp_1285_6 = __tmp_1299_6;
  assign __tmp_1285_7 = __tmp_1299_7;
  assign __tmp_1285_8 = __tmp_1299_8;
  assign __tmp_1285_9 = __tmp_1299_9;
  assign __tmp_1287_1 = __tmp_1299_1;
  assign __tmp_1287_10 = __tmp_1299_10;
  assign __tmp_1287_11 = __tmp_1299_11;
  assign __tmp_1287_12 = __tmp_1299_12;
  assign __tmp_1287_13 = __tmp_1299_13;
  assign __tmp_1287_14 = __tmp_1299_14;
  assign __tmp_1287_15 = __tmp_1299_15;
  assign __tmp_1287_16 = __tmp_1299_16;
  assign __tmp_1287_17 = __tmp_1299_17;
  assign __tmp_1287_18 = __tmp_1299_18;
  assign __tmp_1287_19 = __tmp_1299_19;
  assign __tmp_1287_2 = __tmp_1299_2;
  assign __tmp_1287_20 = __tmp_1291_20;
  assign __tmp_1287_21 = __tmp_1291_21;
  assign __tmp_1287_22 = __tmp_1291_22;
  assign __tmp_1287_23 = __tmp_1291_23;
  assign __tmp_1287_24 = __tmp_1291_24;
  assign __tmp_1287_25 = __tmp_1291_25;
  assign __tmp_1287_3 = __tmp_1299_3;
  assign __tmp_1287_4 = __tmp_1299_4;
  assign __tmp_1287_5 = __tmp_1299_5;
  assign __tmp_1287_6 = __tmp_1299_6;
  assign __tmp_1287_7 = __tmp_1299_7;
  assign __tmp_1287_8 = __tmp_1299_8;
  assign __tmp_1287_9 = __tmp_1299_9;
  assign __tmp_1289_1 = __tmp_1299_1;
  assign __tmp_1289_10 = __tmp_1299_10;
  assign __tmp_1289_11 = __tmp_1299_11;
  assign __tmp_1289_12 = __tmp_1299_12;
  assign __tmp_1289_13 = __tmp_1299_13;
  assign __tmp_1289_14 = __tmp_1299_14;
  assign __tmp_1289_15 = __tmp_1299_15;
  assign __tmp_1289_16 = __tmp_1299_16;
  assign __tmp_1289_17 = __tmp_1299_17;
  assign __tmp_1289_18 = __tmp_1299_18;
  assign __tmp_1289_19 = __tmp_1299_19;
  assign __tmp_1289_2 = __tmp_1299_2;
  assign __tmp_1289_20 = __tmp_1291_20;
  assign __tmp_1289_21 = __tmp_1291_21;
  assign __tmp_1289_22 = __tmp_1291_22;
  assign __tmp_1289_23 = __tmp_1291_23;
  assign __tmp_1289_24 = __tmp_1291_24;
  assign __tmp_1289_25 = __tmp_1291_25;
  assign __tmp_1289_3 = __tmp_1299_3;
  assign __tmp_1289_4 = __tmp_1299_4;
  assign __tmp_1289_5 = __tmp_1299_5;
  assign __tmp_1289_6 = __tmp_1299_6;
  assign __tmp_1289_7 = __tmp_1299_7;
  assign __tmp_1289_8 = __tmp_1299_8;
  assign __tmp_1289_9 = __tmp_1299_9;
  assign __tmp_1291_1 = __tmp_1299_1;
  assign __tmp_1291_10 = __tmp_1299_10;
  assign __tmp_1291_11 = __tmp_1299_11;
  assign __tmp_1291_12 = __tmp_1299_12;
  assign __tmp_1291_13 = __tmp_1299_13;
  assign __tmp_1291_14 = __tmp_1299_14;
  assign __tmp_1291_15 = __tmp_1299_15;
  assign __tmp_1291_16 = __tmp_1299_16;
  assign __tmp_1291_17 = __tmp_1299_17;
  assign __tmp_1291_18 = __tmp_1299_18;
  assign __tmp_1291_19 = __tmp_1299_19;
  assign __tmp_1291_2 = __tmp_1299_2;
  assign __tmp_1291_3 = __tmp_1299_3;
  assign __tmp_1291_4 = __tmp_1299_4;
  assign __tmp_1291_5 = __tmp_1299_5;
  assign __tmp_1291_6 = __tmp_1299_6;
  assign __tmp_1291_7 = __tmp_1299_7;
  assign __tmp_1291_8 = __tmp_1299_8;
  assign __tmp_1291_9 = __tmp_1299_9;
  assign __tmp_1293_1 = __tmp_1299_1;
  assign __tmp_1293_10 = __tmp_1299_10;
  assign __tmp_1293_11 = __tmp_1299_11;
  assign __tmp_1293_12 = __tmp_1299_12;
  assign __tmp_1293_2 = __tmp_1299_2;
  assign __tmp_1293_3 = __tmp_1299_3;
  assign __tmp_1293_4 = __tmp_1299_4;
  assign __tmp_1293_5 = __tmp_1299_5;
  assign __tmp_1293_6 = __tmp_1299_6;
  assign __tmp_1293_7 = __tmp_1299_7;
  assign __tmp_1293_8 = __tmp_1299_8;
  assign __tmp_1293_9 = __tmp_1299_9;
  assign __tmp_1295_1 = __tmp_1299_1;
  assign __tmp_1295_10 = __tmp_1299_10;
  assign __tmp_1295_11 = __tmp_1299_11;
  assign __tmp_1295_12 = __tmp_1299_12;
  assign __tmp_1295_2 = __tmp_1299_2;
  assign __tmp_1295_3 = __tmp_1299_3;
  assign __tmp_1295_4 = __tmp_1299_4;
  assign __tmp_1295_5 = __tmp_1299_5;
  assign __tmp_1295_6 = __tmp_1299_6;
  assign __tmp_1295_7 = __tmp_1299_7;
  assign __tmp_1295_8 = __tmp_1299_8;
  assign __tmp_1295_9 = __tmp_1299_9;
  assign __tmp_1297_1 = __tmp_1299_1;
  assign __tmp_1297_10 = __tmp_1299_10;
  assign __tmp_1297_11 = __tmp_1299_11;
  assign __tmp_1297_12 = __tmp_1299_12;
  assign __tmp_1297_2 = __tmp_1299_2;
  assign __tmp_1297_3 = __tmp_1299_3;
  assign __tmp_1297_4 = __tmp_1299_4;
  assign __tmp_1297_5 = __tmp_1299_5;
  assign __tmp_1297_6 = __tmp_1299_6;
  assign __tmp_1297_7 = __tmp_1299_7;
  assign __tmp_1297_8 = __tmp_1299_8;
  assign __tmp_1297_9 = __tmp_1299_9;
  assign __tmp_1299_20 = __tmp_1291_20;
  assign __tmp_1299_21 = __tmp_1291_21;
  assign __tmp_1299_22 = __tmp_1291_22;
  assign __tmp_1299_23 = __tmp_1291_23;
  assign __tmp_1299_24 = __tmp_1291_24;
  assign __tmp_1299_25 = __tmp_1291_25;
  assign __tmp_1299_26 = __tmp_1307_26;
  assign __tmp_1299_27 = __tmp_1307_27;
  assign __tmp_1299_28 = __tmp_1307_28;
  assign __tmp_1299_29 = __tmp_1307_29;
  assign __tmp_1299_30 = __tmp_1307_30;
  assign __tmp_1299_31 = __tmp_1307_31;
  assign __tmp_1299_32 = __tmp_1307_32;
  assign __tmp_1299_33 = __tmp_1307_33;
  assign __tmp_1299_34 = __tmp_1307_34;
  assign __tmp_1299_35 = __tmp_1307_35;
  assign __tmp_1299_36 = __tmp_1307_36;
  assign __tmp_1299_37 = __tmp_1307_37;
  assign __tmp_1299_38 = __tmp_1307_38;
  assign __tmp_1299_39 = __tmp_1305_39;
  assign __tmp_1299_40 = __tmp_1305_40;
  assign __tmp_1299_41 = __tmp_1305_41;
  assign __tmp_1299_42 = __tmp_1305_42;
  assign __tmp_1301_1 = __tmp_1299_1;
  assign __tmp_1301_10 = __tmp_1299_10;
  assign __tmp_1301_11 = __tmp_1299_11;
  assign __tmp_1301_12 = __tmp_1299_12;
  assign __tmp_1301_13 = __tmp_1299_13;
  assign __tmp_1301_14 = __tmp_1299_14;
  assign __tmp_1301_15 = __tmp_1299_15;
  assign __tmp_1301_16 = __tmp_1299_16;
  assign __tmp_1301_17 = __tmp_1299_17;
  assign __tmp_1301_18 = __tmp_1299_18;
  assign __tmp_1301_19 = __tmp_1299_19;
  assign __tmp_1301_2 = __tmp_1299_2;
  assign __tmp_1301_20 = __tmp_1291_20;
  assign __tmp_1301_21 = __tmp_1291_21;
  assign __tmp_1301_22 = __tmp_1291_22;
  assign __tmp_1301_23 = __tmp_1291_23;
  assign __tmp_1301_24 = __tmp_1291_24;
  assign __tmp_1301_25 = __tmp_1291_25;
  assign __tmp_1301_26 = __tmp_1307_26;
  assign __tmp_1301_27 = __tmp_1307_27;
  assign __tmp_1301_28 = __tmp_1307_28;
  assign __tmp_1301_29 = __tmp_1307_29;
  assign __tmp_1301_3 = __tmp_1299_3;
  assign __tmp_1301_30 = __tmp_1307_30;
  assign __tmp_1301_31 = __tmp_1307_31;
  assign __tmp_1301_32 = __tmp_1307_32;
  assign __tmp_1301_33 = __tmp_1307_33;
  assign __tmp_1301_34 = __tmp_1307_34;
  assign __tmp_1301_35 = __tmp_1307_35;
  assign __tmp_1301_36 = __tmp_1307_36;
  assign __tmp_1301_37 = __tmp_1307_37;
  assign __tmp_1301_38 = __tmp_1307_38;
  assign __tmp_1301_39 = __tmp_1305_39;
  assign __tmp_1301_4 = __tmp_1299_4;
  assign __tmp_1301_40 = __tmp_1305_40;
  assign __tmp_1301_41 = __tmp_1305_41;
  assign __tmp_1301_42 = __tmp_1305_42;
  assign __tmp_1301_5 = __tmp_1299_5;
  assign __tmp_1301_6 = __tmp_1299_6;
  assign __tmp_1301_7 = __tmp_1299_7;
  assign __tmp_1301_8 = __tmp_1299_8;
  assign __tmp_1301_9 = __tmp_1299_9;
  assign __tmp_1303_1 = __tmp_1299_1;
  assign __tmp_1303_10 = __tmp_1299_10;
  assign __tmp_1303_11 = __tmp_1299_11;
  assign __tmp_1303_12 = __tmp_1299_12;
  assign __tmp_1303_13 = __tmp_1299_13;
  assign __tmp_1303_14 = __tmp_1299_14;
  assign __tmp_1303_15 = __tmp_1299_15;
  assign __tmp_1303_16 = __tmp_1299_16;
  assign __tmp_1303_17 = __tmp_1299_17;
  assign __tmp_1303_18 = __tmp_1299_18;
  assign __tmp_1303_19 = __tmp_1299_19;
  assign __tmp_1303_2 = __tmp_1299_2;
  assign __tmp_1303_20 = __tmp_1291_20;
  assign __tmp_1303_21 = __tmp_1291_21;
  assign __tmp_1303_22 = __tmp_1291_22;
  assign __tmp_1303_23 = __tmp_1291_23;
  assign __tmp_1303_24 = __tmp_1291_24;
  assign __tmp_1303_25 = __tmp_1291_25;
  assign __tmp_1303_26 = __tmp_1307_26;
  assign __tmp_1303_27 = __tmp_1307_27;
  assign __tmp_1303_28 = __tmp_1307_28;
  assign __tmp_1303_29 = __tmp_1307_29;
  assign __tmp_1303_3 = __tmp_1299_3;
  assign __tmp_1303_30 = __tmp_1307_30;
  assign __tmp_1303_31 = __tmp_1307_31;
  assign __tmp_1303_32 = __tmp_1307_32;
  assign __tmp_1303_33 = __tmp_1307_33;
  assign __tmp_1303_34 = __tmp_1307_34;
  assign __tmp_1303_35 = __tmp_1307_35;
  assign __tmp_1303_36 = __tmp_1307_36;
  assign __tmp_1303_37 = __tmp_1307_37;
  assign __tmp_1303_38 = __tmp_1307_38;
  assign __tmp_1303_39 = __tmp_1305_39;
  assign __tmp_1303_4 = __tmp_1299_4;
  assign __tmp_1303_40 = __tmp_1305_40;
  assign __tmp_1303_41 = __tmp_1305_41;
  assign __tmp_1303_42 = __tmp_1305_42;
  assign __tmp_1303_5 = __tmp_1299_5;
  assign __tmp_1303_6 = __tmp_1299_6;
  assign __tmp_1303_7 = __tmp_1299_7;
  assign __tmp_1303_8 = __tmp_1299_8;
  assign __tmp_1303_9 = __tmp_1299_9;
  assign __tmp_1305_1 = __tmp_1299_1;
  assign __tmp_1305_10 = __tmp_1299_10;
  assign __tmp_1305_11 = __tmp_1299_11;
  assign __tmp_1305_12 = __tmp_1299_12;
  assign __tmp_1305_13 = __tmp_1299_13;
  assign __tmp_1305_14 = __tmp_1299_14;
  assign __tmp_1305_15 = __tmp_1299_15;
  assign __tmp_1305_16 = __tmp_1299_16;
  assign __tmp_1305_17 = __tmp_1299_17;
  assign __tmp_1305_18 = __tmp_1299_18;
  assign __tmp_1305_19 = __tmp_1299_19;
  assign __tmp_1305_2 = __tmp_1299_2;
  assign __tmp_1305_20 = __tmp_1291_20;
  assign __tmp_1305_21 = __tmp_1291_21;
  assign __tmp_1305_22 = __tmp_1291_22;
  assign __tmp_1305_23 = __tmp_1291_23;
  assign __tmp_1305_24 = __tmp_1291_24;
  assign __tmp_1305_25 = __tmp_1291_25;
  assign __tmp_1305_26 = __tmp_1307_26;
  assign __tmp_1305_27 = __tmp_1307_27;
  assign __tmp_1305_28 = __tmp_1307_28;
  assign __tmp_1305_29 = __tmp_1307_29;
  assign __tmp_1305_3 = __tmp_1299_3;
  assign __tmp_1305_30 = __tmp_1307_30;
  assign __tmp_1305_31 = __tmp_1307_31;
  assign __tmp_1305_32 = __tmp_1307_32;
  assign __tmp_1305_33 = __tmp_1307_33;
  assign __tmp_1305_34 = __tmp_1307_34;
  assign __tmp_1305_35 = __tmp_1307_35;
  assign __tmp_1305_36 = __tmp_1307_36;
  assign __tmp_1305_37 = __tmp_1307_37;
  assign __tmp_1305_38 = __tmp_1307_38;
  assign __tmp_1305_4 = __tmp_1299_4;
  assign __tmp_1305_5 = __tmp_1299_5;
  assign __tmp_1305_6 = __tmp_1299_6;
  assign __tmp_1305_7 = __tmp_1299_7;
  assign __tmp_1305_8 = __tmp_1299_8;
  assign __tmp_1305_9 = __tmp_1299_9;
  assign __tmp_1307_1 = __tmp_1299_1;
  assign __tmp_1307_10 = __tmp_1299_10;
  assign __tmp_1307_11 = __tmp_1299_11;
  assign __tmp_1307_12 = __tmp_1299_12;
  assign __tmp_1307_13 = __tmp_1299_13;
  assign __tmp_1307_14 = __tmp_1299_14;
  assign __tmp_1307_15 = __tmp_1299_15;
  assign __tmp_1307_16 = __tmp_1299_16;
  assign __tmp_1307_17 = __tmp_1299_17;
  assign __tmp_1307_18 = __tmp_1299_18;
  assign __tmp_1307_19 = __tmp_1299_19;
  assign __tmp_1307_2 = __tmp_1299_2;
  assign __tmp_1307_20 = __tmp_1291_20;
  assign __tmp_1307_21 = __tmp_1291_21;
  assign __tmp_1307_22 = __tmp_1291_22;
  assign __tmp_1307_23 = __tmp_1291_23;
  assign __tmp_1307_24 = __tmp_1291_24;
  assign __tmp_1307_25 = __tmp_1291_25;
  assign __tmp_1307_3 = __tmp_1299_3;
  assign __tmp_1307_4 = __tmp_1299_4;
  assign __tmp_1307_5 = __tmp_1299_5;
  assign __tmp_1307_6 = __tmp_1299_6;
  assign __tmp_1307_7 = __tmp_1299_7;
  assign __tmp_1307_8 = __tmp_1299_8;
  assign __tmp_1307_9 = __tmp_1299_9;
  assign __tmp_472_1 = _ram_w8_l2048_id1_0_cond_2_1;
  assign __tmp_483_1 = _ram_w8_l2048_id0_3_cond_2_1;
  assign __tmp_503_1 = _ram_w8_l2048_id2_0_cond_3_1;
  assign __tmp_513_1 = _ram_w8_l2048_id3_0_cond_2_1;
  assign __tmp_523_1 = _ram_w8_l2048_id4_0_cond_2_1;
  assign __tmp_533_1 = _ram_w8_l2048_id5_0_cond_3_1;
  assign __tmp_543_1 = _ram_w8_l2048_id6_0_cond_2_1;
  assign __tmp_553_1 = _ram_w8_l2048_id7_0_cond_2_1;
  assign __tmp_563_1 = _ram_w8_l2048_id8_0_cond_3_1;
  assign __tmp_573_1 = _ram_w8_l2048_id9_0_cond_2_1;
  assign __tmp_583_1 = _ram_w8_l2048_id10_0_cond_2_1;
  assign __tmp_597_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign __tmp_611_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign __tmp_625_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign __tmp_639_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign __tmp_653_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign __tmp_667_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign __tmp_681_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign __tmp_695_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign __tmp_709_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign __tmp_713_1 = __tmp_799_1;
  assign __tmp_713_2 = __tmp_799_2;
  assign __tmp_713_3 = __tmp_799_3;
  assign __tmp_713_4 = __tmp_799_4;
  assign __tmp_713_5 = __tmp_799_5;
  assign __tmp_715_1 = __tmp_799_1;
  assign __tmp_715_10 = __tmp_799_10;
  assign __tmp_715_11 = __tmp_799_11;
  assign __tmp_715_12 = __tmp_799_12;
  assign __tmp_715_2 = __tmp_799_2;
  assign __tmp_715_3 = __tmp_799_3;
  assign __tmp_715_4 = __tmp_799_4;
  assign __tmp_715_5 = __tmp_799_5;
  assign __tmp_715_6 = __tmp_799_6;
  assign __tmp_715_7 = __tmp_799_7;
  assign __tmp_715_8 = __tmp_799_8;
  assign __tmp_715_9 = __tmp_799_9;
  assign __tmp_717_1 = __tmp_799_1;
  assign __tmp_717_10 = __tmp_799_10;
  assign __tmp_717_11 = __tmp_799_11;
  assign __tmp_717_12 = __tmp_799_12;
  assign __tmp_717_2 = __tmp_799_2;
  assign __tmp_717_3 = __tmp_799_3;
  assign __tmp_717_4 = __tmp_799_4;
  assign __tmp_717_5 = __tmp_799_5;
  assign __tmp_717_6 = __tmp_799_6;
  assign __tmp_717_7 = __tmp_799_7;
  assign __tmp_717_8 = __tmp_799_8;
  assign __tmp_717_9 = __tmp_799_9;
  assign __tmp_719_1 = __tmp_799_1;
  assign __tmp_719_10 = __tmp_799_10;
  assign __tmp_719_11 = __tmp_799_11;
  assign __tmp_719_12 = __tmp_799_12;
  assign __tmp_719_2 = __tmp_799_2;
  assign __tmp_719_3 = __tmp_799_3;
  assign __tmp_719_4 = __tmp_799_4;
  assign __tmp_719_5 = __tmp_799_5;
  assign __tmp_719_6 = __tmp_799_6;
  assign __tmp_719_7 = __tmp_799_7;
  assign __tmp_719_8 = __tmp_799_8;
  assign __tmp_719_9 = __tmp_799_9;
  assign __tmp_721_1 = __tmp_799_1;
  assign __tmp_721_10 = __tmp_799_10;
  assign __tmp_721_11 = __tmp_799_11;
  assign __tmp_721_12 = __tmp_799_12;
  assign __tmp_721_2 = __tmp_799_2;
  assign __tmp_721_3 = __tmp_799_3;
  assign __tmp_721_4 = __tmp_799_4;
  assign __tmp_721_5 = __tmp_799_5;
  assign __tmp_721_6 = __tmp_799_6;
  assign __tmp_721_7 = __tmp_799_7;
  assign __tmp_721_8 = __tmp_799_8;
  assign __tmp_721_9 = __tmp_799_9;
  assign __tmp_723_1 = __tmp_799_1;
  assign __tmp_723_10 = __tmp_799_10;
  assign __tmp_723_11 = __tmp_799_11;
  assign __tmp_723_12 = __tmp_799_12;
  assign __tmp_723_2 = __tmp_799_2;
  assign __tmp_723_3 = __tmp_799_3;
  assign __tmp_723_4 = __tmp_799_4;
  assign __tmp_723_5 = __tmp_799_5;
  assign __tmp_723_6 = __tmp_799_6;
  assign __tmp_723_7 = __tmp_799_7;
  assign __tmp_723_8 = __tmp_799_8;
  assign __tmp_723_9 = __tmp_799_9;
  assign __tmp_725_1 = __tmp_799_1;
  assign __tmp_725_10 = __tmp_799_10;
  assign __tmp_725_11 = __tmp_799_11;
  assign __tmp_725_12 = __tmp_799_12;
  assign __tmp_725_2 = __tmp_799_2;
  assign __tmp_725_3 = __tmp_799_3;
  assign __tmp_725_4 = __tmp_799_4;
  assign __tmp_725_5 = __tmp_799_5;
  assign __tmp_725_6 = __tmp_799_6;
  assign __tmp_725_7 = __tmp_799_7;
  assign __tmp_725_8 = __tmp_799_8;
  assign __tmp_725_9 = __tmp_799_9;
  assign __tmp_727_1 = __tmp_799_1;
  assign __tmp_727_10 = __tmp_799_10;
  assign __tmp_727_11 = __tmp_799_11;
  assign __tmp_727_12 = __tmp_799_12;
  assign __tmp_727_2 = __tmp_799_2;
  assign __tmp_727_3 = __tmp_799_3;
  assign __tmp_727_4 = __tmp_799_4;
  assign __tmp_727_5 = __tmp_799_5;
  assign __tmp_727_6 = __tmp_799_6;
  assign __tmp_727_7 = __tmp_799_7;
  assign __tmp_727_8 = __tmp_799_8;
  assign __tmp_727_9 = __tmp_799_9;
  assign __tmp_729_1 = __tmp_799_1;
  assign __tmp_729_10 = __tmp_799_10;
  assign __tmp_729_11 = __tmp_799_11;
  assign __tmp_729_12 = __tmp_799_12;
  assign __tmp_729_2 = __tmp_799_2;
  assign __tmp_729_3 = __tmp_799_3;
  assign __tmp_729_4 = __tmp_799_4;
  assign __tmp_729_5 = __tmp_799_5;
  assign __tmp_729_6 = __tmp_799_6;
  assign __tmp_729_7 = __tmp_799_7;
  assign __tmp_729_8 = __tmp_799_8;
  assign __tmp_729_9 = __tmp_799_9;
  assign __tmp_731_1 = __tmp_799_1;
  assign __tmp_731_10 = __tmp_799_10;
  assign __tmp_731_11 = __tmp_799_11;
  assign __tmp_731_12 = __tmp_799_12;
  assign __tmp_731_2 = __tmp_799_2;
  assign __tmp_731_3 = __tmp_799_3;
  assign __tmp_731_4 = __tmp_799_4;
  assign __tmp_731_5 = __tmp_799_5;
  assign __tmp_731_6 = __tmp_799_6;
  assign __tmp_731_7 = __tmp_799_7;
  assign __tmp_731_8 = __tmp_799_8;
  assign __tmp_731_9 = __tmp_799_9;
  assign __tmp_733_1 = __tmp_799_1;
  assign __tmp_733_10 = __tmp_799_10;
  assign __tmp_733_11 = __tmp_799_11;
  assign __tmp_733_12 = __tmp_799_12;
  assign __tmp_733_2 = __tmp_799_2;
  assign __tmp_733_3 = __tmp_799_3;
  assign __tmp_733_4 = __tmp_799_4;
  assign __tmp_733_5 = __tmp_799_5;
  assign __tmp_733_6 = __tmp_799_6;
  assign __tmp_733_7 = __tmp_799_7;
  assign __tmp_733_8 = __tmp_799_8;
  assign __tmp_733_9 = __tmp_799_9;
  assign __tmp_735_1 = __tmp_799_1;
  assign __tmp_735_10 = __tmp_799_10;
  assign __tmp_735_11 = __tmp_799_11;
  assign __tmp_735_12 = __tmp_799_12;
  assign __tmp_735_2 = __tmp_799_2;
  assign __tmp_735_3 = __tmp_799_3;
  assign __tmp_735_4 = __tmp_799_4;
  assign __tmp_735_5 = __tmp_799_5;
  assign __tmp_735_6 = __tmp_799_6;
  assign __tmp_735_7 = __tmp_799_7;
  assign __tmp_735_8 = __tmp_799_8;
  assign __tmp_735_9 = __tmp_799_9;
  assign __tmp_737_1 = __tmp_799_1;
  assign __tmp_737_10 = __tmp_799_10;
  assign __tmp_737_11 = __tmp_799_11;
  assign __tmp_737_12 = __tmp_799_12;
  assign __tmp_737_2 = __tmp_799_2;
  assign __tmp_737_3 = __tmp_799_3;
  assign __tmp_737_4 = __tmp_799_4;
  assign __tmp_737_5 = __tmp_799_5;
  assign __tmp_737_6 = __tmp_799_6;
  assign __tmp_737_7 = __tmp_799_7;
  assign __tmp_737_8 = __tmp_799_8;
  assign __tmp_737_9 = __tmp_799_9;
  assign __tmp_739_1 = __tmp_799_1;
  assign __tmp_739_10 = __tmp_799_10;
  assign __tmp_739_11 = __tmp_799_11;
  assign __tmp_739_12 = __tmp_799_12;
  assign __tmp_739_2 = __tmp_799_2;
  assign __tmp_739_3 = __tmp_799_3;
  assign __tmp_739_4 = __tmp_799_4;
  assign __tmp_739_5 = __tmp_799_5;
  assign __tmp_739_6 = __tmp_799_6;
  assign __tmp_739_7 = __tmp_799_7;
  assign __tmp_739_8 = __tmp_799_8;
  assign __tmp_739_9 = __tmp_799_9;
  assign __tmp_741_1 = __tmp_799_1;
  assign __tmp_741_10 = __tmp_799_10;
  assign __tmp_741_11 = __tmp_799_11;
  assign __tmp_741_12 = __tmp_799_12;
  assign __tmp_741_2 = __tmp_799_2;
  assign __tmp_741_3 = __tmp_799_3;
  assign __tmp_741_4 = __tmp_799_4;
  assign __tmp_741_5 = __tmp_799_5;
  assign __tmp_741_6 = __tmp_799_6;
  assign __tmp_741_7 = __tmp_799_7;
  assign __tmp_741_8 = __tmp_799_8;
  assign __tmp_741_9 = __tmp_799_9;
  assign __tmp_743_1 = __tmp_799_1;
  assign __tmp_743_10 = __tmp_799_10;
  assign __tmp_743_11 = __tmp_799_11;
  assign __tmp_743_12 = __tmp_799_12;
  assign __tmp_743_2 = __tmp_799_2;
  assign __tmp_743_3 = __tmp_799_3;
  assign __tmp_743_4 = __tmp_799_4;
  assign __tmp_743_5 = __tmp_799_5;
  assign __tmp_743_6 = __tmp_799_6;
  assign __tmp_743_7 = __tmp_799_7;
  assign __tmp_743_8 = __tmp_799_8;
  assign __tmp_743_9 = __tmp_799_9;
  assign __tmp_745_1 = __tmp_799_1;
  assign __tmp_745_10 = __tmp_799_10;
  assign __tmp_745_11 = __tmp_799_11;
  assign __tmp_745_12 = __tmp_799_12;
  assign __tmp_745_2 = __tmp_799_2;
  assign __tmp_745_3 = __tmp_799_3;
  assign __tmp_745_4 = __tmp_799_4;
  assign __tmp_745_5 = __tmp_799_5;
  assign __tmp_745_6 = __tmp_799_6;
  assign __tmp_745_7 = __tmp_799_7;
  assign __tmp_745_8 = __tmp_799_8;
  assign __tmp_745_9 = __tmp_799_9;
  assign __tmp_747_1 = __tmp_799_1;
  assign __tmp_747_10 = __tmp_799_10;
  assign __tmp_747_11 = __tmp_799_11;
  assign __tmp_747_12 = __tmp_799_12;
  assign __tmp_747_2 = __tmp_799_2;
  assign __tmp_747_3 = __tmp_799_3;
  assign __tmp_747_4 = __tmp_799_4;
  assign __tmp_747_5 = __tmp_799_5;
  assign __tmp_747_6 = __tmp_799_6;
  assign __tmp_747_7 = __tmp_799_7;
  assign __tmp_747_8 = __tmp_799_8;
  assign __tmp_747_9 = __tmp_799_9;
  assign __tmp_749_1 = __tmp_799_1;
  assign __tmp_749_10 = __tmp_799_10;
  assign __tmp_749_11 = __tmp_799_11;
  assign __tmp_749_12 = __tmp_799_12;
  assign __tmp_749_2 = __tmp_799_2;
  assign __tmp_749_3 = __tmp_799_3;
  assign __tmp_749_4 = __tmp_799_4;
  assign __tmp_749_5 = __tmp_799_5;
  assign __tmp_749_6 = __tmp_799_6;
  assign __tmp_749_7 = __tmp_799_7;
  assign __tmp_749_8 = __tmp_799_8;
  assign __tmp_749_9 = __tmp_799_9;
  assign __tmp_751_1 = __tmp_799_1;
  assign __tmp_751_10 = __tmp_799_10;
  assign __tmp_751_11 = __tmp_799_11;
  assign __tmp_751_12 = __tmp_799_12;
  assign __tmp_751_2 = __tmp_799_2;
  assign __tmp_751_3 = __tmp_799_3;
  assign __tmp_751_4 = __tmp_799_4;
  assign __tmp_751_5 = __tmp_799_5;
  assign __tmp_751_6 = __tmp_799_6;
  assign __tmp_751_7 = __tmp_799_7;
  assign __tmp_751_8 = __tmp_799_8;
  assign __tmp_751_9 = __tmp_799_9;
  assign __tmp_753_1 = __tmp_799_1;
  assign __tmp_753_10 = __tmp_799_10;
  assign __tmp_753_11 = __tmp_799_11;
  assign __tmp_753_12 = __tmp_799_12;
  assign __tmp_753_2 = __tmp_799_2;
  assign __tmp_753_3 = __tmp_799_3;
  assign __tmp_753_4 = __tmp_799_4;
  assign __tmp_753_5 = __tmp_799_5;
  assign __tmp_753_6 = __tmp_799_6;
  assign __tmp_753_7 = __tmp_799_7;
  assign __tmp_753_8 = __tmp_799_8;
  assign __tmp_753_9 = __tmp_799_9;
  assign __tmp_755_1 = __tmp_799_1;
  assign __tmp_755_10 = __tmp_799_10;
  assign __tmp_755_11 = __tmp_799_11;
  assign __tmp_755_12 = __tmp_799_12;
  assign __tmp_755_2 = __tmp_799_2;
  assign __tmp_755_3 = __tmp_799_3;
  assign __tmp_755_4 = __tmp_799_4;
  assign __tmp_755_5 = __tmp_799_5;
  assign __tmp_755_6 = __tmp_799_6;
  assign __tmp_755_7 = __tmp_799_7;
  assign __tmp_755_8 = __tmp_799_8;
  assign __tmp_755_9 = __tmp_799_9;
  assign __tmp_757_1 = __tmp_799_1;
  assign __tmp_757_10 = __tmp_799_10;
  assign __tmp_757_11 = __tmp_799_11;
  assign __tmp_757_12 = __tmp_799_12;
  assign __tmp_757_2 = __tmp_799_2;
  assign __tmp_757_3 = __tmp_799_3;
  assign __tmp_757_4 = __tmp_799_4;
  assign __tmp_757_5 = __tmp_799_5;
  assign __tmp_757_6 = __tmp_799_6;
  assign __tmp_757_7 = __tmp_799_7;
  assign __tmp_757_8 = __tmp_799_8;
  assign __tmp_757_9 = __tmp_799_9;
  assign __tmp_759_1 = __tmp_799_1;
  assign __tmp_759_10 = __tmp_799_10;
  assign __tmp_759_11 = __tmp_799_11;
  assign __tmp_759_12 = __tmp_799_12;
  assign __tmp_759_2 = __tmp_799_2;
  assign __tmp_759_3 = __tmp_799_3;
  assign __tmp_759_4 = __tmp_799_4;
  assign __tmp_759_5 = __tmp_799_5;
  assign __tmp_759_6 = __tmp_799_6;
  assign __tmp_759_7 = __tmp_799_7;
  assign __tmp_759_8 = __tmp_799_8;
  assign __tmp_759_9 = __tmp_799_9;
  assign __tmp_761_1 = __tmp_799_1;
  assign __tmp_761_10 = __tmp_799_10;
  assign __tmp_761_11 = __tmp_799_11;
  assign __tmp_761_12 = __tmp_799_12;
  assign __tmp_761_2 = __tmp_799_2;
  assign __tmp_761_3 = __tmp_799_3;
  assign __tmp_761_4 = __tmp_799_4;
  assign __tmp_761_5 = __tmp_799_5;
  assign __tmp_761_6 = __tmp_799_6;
  assign __tmp_761_7 = __tmp_799_7;
  assign __tmp_761_8 = __tmp_799_8;
  assign __tmp_761_9 = __tmp_799_9;
  assign __tmp_763_1 = __tmp_799_1;
  assign __tmp_763_10 = __tmp_799_10;
  assign __tmp_763_11 = __tmp_799_11;
  assign __tmp_763_12 = __tmp_799_12;
  assign __tmp_763_2 = __tmp_799_2;
  assign __tmp_763_3 = __tmp_799_3;
  assign __tmp_763_4 = __tmp_799_4;
  assign __tmp_763_5 = __tmp_799_5;
  assign __tmp_763_6 = __tmp_799_6;
  assign __tmp_763_7 = __tmp_799_7;
  assign __tmp_763_8 = __tmp_799_8;
  assign __tmp_763_9 = __tmp_799_9;
  assign __tmp_765_1 = __tmp_799_1;
  assign __tmp_765_10 = __tmp_799_10;
  assign __tmp_765_11 = __tmp_799_11;
  assign __tmp_765_12 = __tmp_799_12;
  assign __tmp_765_2 = __tmp_799_2;
  assign __tmp_765_3 = __tmp_799_3;
  assign __tmp_765_4 = __tmp_799_4;
  assign __tmp_765_5 = __tmp_799_5;
  assign __tmp_765_6 = __tmp_799_6;
  assign __tmp_765_7 = __tmp_799_7;
  assign __tmp_765_8 = __tmp_799_8;
  assign __tmp_765_9 = __tmp_799_9;
  assign __tmp_767_1 = __tmp_799_1;
  assign __tmp_767_10 = __tmp_799_10;
  assign __tmp_767_11 = __tmp_799_11;
  assign __tmp_767_12 = __tmp_799_12;
  assign __tmp_767_2 = __tmp_799_2;
  assign __tmp_767_3 = __tmp_799_3;
  assign __tmp_767_4 = __tmp_799_4;
  assign __tmp_767_5 = __tmp_799_5;
  assign __tmp_767_6 = __tmp_799_6;
  assign __tmp_767_7 = __tmp_799_7;
  assign __tmp_767_8 = __tmp_799_8;
  assign __tmp_767_9 = __tmp_799_9;
  assign __tmp_769_1 = __tmp_799_1;
  assign __tmp_769_10 = __tmp_799_10;
  assign __tmp_769_11 = __tmp_799_11;
  assign __tmp_769_12 = __tmp_799_12;
  assign __tmp_769_13 = __tmp_799_13;
  assign __tmp_769_14 = __tmp_799_14;
  assign __tmp_769_15 = __tmp_799_15;
  assign __tmp_769_16 = __tmp_799_16;
  assign __tmp_769_17 = __tmp_799_17;
  assign __tmp_769_18 = __tmp_799_18;
  assign __tmp_769_19 = __tmp_799_19;
  assign __tmp_769_2 = __tmp_799_2;
  assign __tmp_769_20 = __tmp_799_20;
  assign __tmp_769_21 = __tmp_799_21;
  assign __tmp_769_22 = __tmp_799_22;
  assign __tmp_769_3 = __tmp_799_3;
  assign __tmp_769_4 = __tmp_799_4;
  assign __tmp_769_5 = __tmp_799_5;
  assign __tmp_769_6 = __tmp_799_6;
  assign __tmp_769_7 = __tmp_799_7;
  assign __tmp_769_8 = __tmp_799_8;
  assign __tmp_769_9 = __tmp_799_9;
  assign __tmp_771_1 = __tmp_799_1;
  assign __tmp_771_10 = __tmp_799_10;
  assign __tmp_771_11 = __tmp_799_11;
  assign __tmp_771_12 = __tmp_799_12;
  assign __tmp_771_13 = __tmp_799_13;
  assign __tmp_771_14 = __tmp_799_14;
  assign __tmp_771_15 = __tmp_799_15;
  assign __tmp_771_16 = __tmp_799_16;
  assign __tmp_771_17 = __tmp_799_17;
  assign __tmp_771_18 = __tmp_799_18;
  assign __tmp_771_19 = __tmp_799_19;
  assign __tmp_771_2 = __tmp_799_2;
  assign __tmp_771_20 = __tmp_799_20;
  assign __tmp_771_21 = __tmp_799_21;
  assign __tmp_771_22 = __tmp_799_22;
  assign __tmp_771_3 = __tmp_799_3;
  assign __tmp_771_4 = __tmp_799_4;
  assign __tmp_771_5 = __tmp_799_5;
  assign __tmp_771_6 = __tmp_799_6;
  assign __tmp_771_7 = __tmp_799_7;
  assign __tmp_771_8 = __tmp_799_8;
  assign __tmp_771_9 = __tmp_799_9;
  assign __tmp_773_1 = __tmp_799_1;
  assign __tmp_773_10 = __tmp_799_10;
  assign __tmp_773_11 = __tmp_799_11;
  assign __tmp_773_12 = __tmp_799_12;
  assign __tmp_773_13 = __tmp_799_13;
  assign __tmp_773_14 = __tmp_799_14;
  assign __tmp_773_15 = __tmp_799_15;
  assign __tmp_773_16 = __tmp_799_16;
  assign __tmp_773_17 = __tmp_799_17;
  assign __tmp_773_18 = __tmp_799_18;
  assign __tmp_773_19 = __tmp_799_19;
  assign __tmp_773_2 = __tmp_799_2;
  assign __tmp_773_20 = __tmp_799_20;
  assign __tmp_773_21 = __tmp_799_21;
  assign __tmp_773_22 = __tmp_799_22;
  assign __tmp_773_3 = __tmp_799_3;
  assign __tmp_773_4 = __tmp_799_4;
  assign __tmp_773_5 = __tmp_799_5;
  assign __tmp_773_6 = __tmp_799_6;
  assign __tmp_773_7 = __tmp_799_7;
  assign __tmp_773_8 = __tmp_799_8;
  assign __tmp_773_9 = __tmp_799_9;
  assign __tmp_775_1 = __tmp_799_1;
  assign __tmp_775_10 = __tmp_799_10;
  assign __tmp_775_11 = __tmp_799_11;
  assign __tmp_775_12 = __tmp_799_12;
  assign __tmp_775_13 = __tmp_799_13;
  assign __tmp_775_14 = __tmp_799_14;
  assign __tmp_775_15 = __tmp_799_15;
  assign __tmp_775_16 = __tmp_799_16;
  assign __tmp_775_17 = __tmp_799_17;
  assign __tmp_775_18 = __tmp_799_18;
  assign __tmp_775_19 = __tmp_799_19;
  assign __tmp_775_2 = __tmp_799_2;
  assign __tmp_775_20 = __tmp_799_20;
  assign __tmp_775_21 = __tmp_799_21;
  assign __tmp_775_22 = __tmp_799_22;
  assign __tmp_775_3 = __tmp_799_3;
  assign __tmp_775_4 = __tmp_799_4;
  assign __tmp_775_5 = __tmp_799_5;
  assign __tmp_775_6 = __tmp_799_6;
  assign __tmp_775_7 = __tmp_799_7;
  assign __tmp_775_8 = __tmp_799_8;
  assign __tmp_775_9 = __tmp_799_9;
  assign __tmp_777_1 = __tmp_799_1;
  assign __tmp_777_10 = __tmp_799_10;
  assign __tmp_777_11 = __tmp_799_11;
  assign __tmp_777_12 = __tmp_799_12;
  assign __tmp_777_13 = __tmp_799_13;
  assign __tmp_777_14 = __tmp_799_14;
  assign __tmp_777_15 = __tmp_799_15;
  assign __tmp_777_16 = __tmp_799_16;
  assign __tmp_777_17 = __tmp_799_17;
  assign __tmp_777_18 = __tmp_799_18;
  assign __tmp_777_19 = __tmp_799_19;
  assign __tmp_777_2 = __tmp_799_2;
  assign __tmp_777_20 = __tmp_799_20;
  assign __tmp_777_21 = __tmp_799_21;
  assign __tmp_777_22 = __tmp_799_22;
  assign __tmp_777_3 = __tmp_799_3;
  assign __tmp_777_4 = __tmp_799_4;
  assign __tmp_777_5 = __tmp_799_5;
  assign __tmp_777_6 = __tmp_799_6;
  assign __tmp_777_7 = __tmp_799_7;
  assign __tmp_777_8 = __tmp_799_8;
  assign __tmp_777_9 = __tmp_799_9;
  assign __tmp_779_1 = __tmp_799_1;
  assign __tmp_779_10 = __tmp_799_10;
  assign __tmp_779_11 = __tmp_799_11;
  assign __tmp_779_12 = __tmp_799_12;
  assign __tmp_779_13 = __tmp_799_13;
  assign __tmp_779_14 = __tmp_799_14;
  assign __tmp_779_15 = __tmp_799_15;
  assign __tmp_779_16 = __tmp_799_16;
  assign __tmp_779_17 = __tmp_799_17;
  assign __tmp_779_18 = __tmp_799_18;
  assign __tmp_779_19 = __tmp_799_19;
  assign __tmp_779_2 = __tmp_799_2;
  assign __tmp_779_20 = __tmp_799_20;
  assign __tmp_779_21 = __tmp_799_21;
  assign __tmp_779_22 = __tmp_799_22;
  assign __tmp_779_3 = __tmp_799_3;
  assign __tmp_779_4 = __tmp_799_4;
  assign __tmp_779_5 = __tmp_799_5;
  assign __tmp_779_6 = __tmp_799_6;
  assign __tmp_779_7 = __tmp_799_7;
  assign __tmp_779_8 = __tmp_799_8;
  assign __tmp_779_9 = __tmp_799_9;
  assign __tmp_781_1 = __tmp_799_1;
  assign __tmp_781_10 = __tmp_799_10;
  assign __tmp_781_11 = __tmp_799_11;
  assign __tmp_781_12 = __tmp_799_12;
  assign __tmp_781_13 = __tmp_799_13;
  assign __tmp_781_14 = __tmp_799_14;
  assign __tmp_781_15 = __tmp_799_15;
  assign __tmp_781_16 = __tmp_799_16;
  assign __tmp_781_17 = __tmp_799_17;
  assign __tmp_781_18 = __tmp_799_18;
  assign __tmp_781_19 = __tmp_799_19;
  assign __tmp_781_2 = __tmp_799_2;
  assign __tmp_781_20 = __tmp_799_20;
  assign __tmp_781_21 = __tmp_799_21;
  assign __tmp_781_22 = __tmp_799_22;
  assign __tmp_781_3 = __tmp_799_3;
  assign __tmp_781_4 = __tmp_799_4;
  assign __tmp_781_5 = __tmp_799_5;
  assign __tmp_781_6 = __tmp_799_6;
  assign __tmp_781_7 = __tmp_799_7;
  assign __tmp_781_8 = __tmp_799_8;
  assign __tmp_781_9 = __tmp_799_9;
  assign __tmp_783_1 = __tmp_799_1;
  assign __tmp_783_10 = __tmp_799_10;
  assign __tmp_783_11 = __tmp_799_11;
  assign __tmp_783_12 = __tmp_799_12;
  assign __tmp_783_13 = __tmp_799_13;
  assign __tmp_783_14 = __tmp_799_14;
  assign __tmp_783_15 = __tmp_799_15;
  assign __tmp_783_16 = __tmp_799_16;
  assign __tmp_783_17 = __tmp_799_17;
  assign __tmp_783_18 = __tmp_799_18;
  assign __tmp_783_19 = __tmp_799_19;
  assign __tmp_783_2 = __tmp_799_2;
  assign __tmp_783_20 = __tmp_799_20;
  assign __tmp_783_21 = __tmp_799_21;
  assign __tmp_783_22 = __tmp_799_22;
  assign __tmp_783_3 = __tmp_799_3;
  assign __tmp_783_4 = __tmp_799_4;
  assign __tmp_783_5 = __tmp_799_5;
  assign __tmp_783_6 = __tmp_799_6;
  assign __tmp_783_7 = __tmp_799_7;
  assign __tmp_783_8 = __tmp_799_8;
  assign __tmp_783_9 = __tmp_799_9;
  assign __tmp_785_1 = __tmp_799_1;
  assign __tmp_785_10 = __tmp_799_10;
  assign __tmp_785_11 = __tmp_799_11;
  assign __tmp_785_12 = __tmp_799_12;
  assign __tmp_785_13 = __tmp_799_13;
  assign __tmp_785_14 = __tmp_799_14;
  assign __tmp_785_15 = __tmp_799_15;
  assign __tmp_785_16 = __tmp_799_16;
  assign __tmp_785_17 = __tmp_799_17;
  assign __tmp_785_18 = __tmp_799_18;
  assign __tmp_785_19 = __tmp_799_19;
  assign __tmp_785_2 = __tmp_799_2;
  assign __tmp_785_20 = __tmp_799_20;
  assign __tmp_785_21 = __tmp_799_21;
  assign __tmp_785_22 = __tmp_799_22;
  assign __tmp_785_3 = __tmp_799_3;
  assign __tmp_785_4 = __tmp_799_4;
  assign __tmp_785_5 = __tmp_799_5;
  assign __tmp_785_6 = __tmp_799_6;
  assign __tmp_785_7 = __tmp_799_7;
  assign __tmp_785_8 = __tmp_799_8;
  assign __tmp_785_9 = __tmp_799_9;
  assign __tmp_787_1 = __tmp_799_1;
  assign __tmp_787_10 = __tmp_799_10;
  assign __tmp_787_11 = __tmp_799_11;
  assign __tmp_787_12 = __tmp_799_12;
  assign __tmp_787_13 = __tmp_799_13;
  assign __tmp_787_14 = __tmp_799_14;
  assign __tmp_787_15 = __tmp_799_15;
  assign __tmp_787_16 = __tmp_799_16;
  assign __tmp_787_17 = __tmp_799_17;
  assign __tmp_787_18 = __tmp_799_18;
  assign __tmp_787_19 = __tmp_799_19;
  assign __tmp_787_2 = __tmp_799_2;
  assign __tmp_787_20 = __tmp_799_20;
  assign __tmp_787_21 = __tmp_799_21;
  assign __tmp_787_22 = __tmp_799_22;
  assign __tmp_787_23 = __tmp_799_23;
  assign __tmp_787_24 = __tmp_799_24;
  assign __tmp_787_25 = __tmp_799_25;
  assign __tmp_787_26 = __tmp_799_26;
  assign __tmp_787_27 = __tmp_799_27;
  assign __tmp_787_28 = __tmp_799_28;
  assign __tmp_787_3 = __tmp_799_3;
  assign __tmp_787_4 = __tmp_799_4;
  assign __tmp_787_5 = __tmp_799_5;
  assign __tmp_787_6 = __tmp_799_6;
  assign __tmp_787_7 = __tmp_799_7;
  assign __tmp_787_8 = __tmp_799_8;
  assign __tmp_787_9 = __tmp_799_9;
  assign __tmp_789_1 = __tmp_799_1;
  assign __tmp_789_10 = __tmp_799_10;
  assign __tmp_789_11 = __tmp_799_11;
  assign __tmp_789_12 = __tmp_799_12;
  assign __tmp_789_13 = __tmp_799_13;
  assign __tmp_789_14 = __tmp_799_14;
  assign __tmp_789_15 = __tmp_799_15;
  assign __tmp_789_16 = __tmp_799_16;
  assign __tmp_789_17 = __tmp_799_17;
  assign __tmp_789_18 = __tmp_799_18;
  assign __tmp_789_19 = __tmp_799_19;
  assign __tmp_789_2 = __tmp_799_2;
  assign __tmp_789_20 = __tmp_799_20;
  assign __tmp_789_21 = __tmp_799_21;
  assign __tmp_789_22 = __tmp_799_22;
  assign __tmp_789_23 = __tmp_799_23;
  assign __tmp_789_24 = __tmp_799_24;
  assign __tmp_789_25 = __tmp_799_25;
  assign __tmp_789_26 = __tmp_799_26;
  assign __tmp_789_3 = __tmp_799_3;
  assign __tmp_789_4 = __tmp_799_4;
  assign __tmp_789_5 = __tmp_799_5;
  assign __tmp_789_6 = __tmp_799_6;
  assign __tmp_789_7 = __tmp_799_7;
  assign __tmp_789_8 = __tmp_799_8;
  assign __tmp_789_9 = __tmp_799_9;
  assign __tmp_791_1 = __tmp_799_1;
  assign __tmp_791_10 = __tmp_799_10;
  assign __tmp_791_11 = __tmp_799_11;
  assign __tmp_791_12 = __tmp_799_12;
  assign __tmp_791_13 = __tmp_799_13;
  assign __tmp_791_14 = __tmp_799_14;
  assign __tmp_791_15 = __tmp_799_15;
  assign __tmp_791_16 = __tmp_799_16;
  assign __tmp_791_17 = __tmp_799_17;
  assign __tmp_791_18 = __tmp_799_18;
  assign __tmp_791_19 = __tmp_799_19;
  assign __tmp_791_2 = __tmp_799_2;
  assign __tmp_791_20 = __tmp_799_20;
  assign __tmp_791_21 = __tmp_799_21;
  assign __tmp_791_22 = __tmp_799_22;
  assign __tmp_791_23 = __tmp_799_23;
  assign __tmp_791_24 = __tmp_799_24;
  assign __tmp_791_25 = __tmp_799_25;
  assign __tmp_791_26 = __tmp_799_26;
  assign __tmp_791_3 = __tmp_799_3;
  assign __tmp_791_4 = __tmp_799_4;
  assign __tmp_791_5 = __tmp_799_5;
  assign __tmp_791_6 = __tmp_799_6;
  assign __tmp_791_7 = __tmp_799_7;
  assign __tmp_791_8 = __tmp_799_8;
  assign __tmp_791_9 = __tmp_799_9;
  assign __tmp_793_1 = __tmp_799_1;
  assign __tmp_793_10 = __tmp_799_10;
  assign __tmp_793_11 = __tmp_799_11;
  assign __tmp_793_12 = __tmp_799_12;
  assign __tmp_793_13 = __tmp_799_13;
  assign __tmp_793_14 = __tmp_799_14;
  assign __tmp_793_15 = __tmp_799_15;
  assign __tmp_793_16 = __tmp_799_16;
  assign __tmp_793_17 = __tmp_799_17;
  assign __tmp_793_18 = __tmp_799_18;
  assign __tmp_793_19 = __tmp_799_19;
  assign __tmp_793_2 = __tmp_799_2;
  assign __tmp_793_20 = __tmp_799_20;
  assign __tmp_793_21 = __tmp_799_21;
  assign __tmp_793_22 = __tmp_799_22;
  assign __tmp_793_23 = __tmp_799_23;
  assign __tmp_793_24 = __tmp_799_24;
  assign __tmp_793_25 = __tmp_799_25;
  assign __tmp_793_26 = __tmp_799_26;
  assign __tmp_793_3 = __tmp_799_3;
  assign __tmp_793_4 = __tmp_799_4;
  assign __tmp_793_5 = __tmp_799_5;
  assign __tmp_793_6 = __tmp_799_6;
  assign __tmp_793_7 = __tmp_799_7;
  assign __tmp_793_8 = __tmp_799_8;
  assign __tmp_793_9 = __tmp_799_9;
  assign __tmp_795_1 = __tmp_799_1;
  assign __tmp_795_10 = __tmp_799_10;
  assign __tmp_795_11 = __tmp_799_11;
  assign __tmp_795_12 = __tmp_799_12;
  assign __tmp_795_13 = __tmp_799_13;
  assign __tmp_795_14 = __tmp_799_14;
  assign __tmp_795_15 = __tmp_799_15;
  assign __tmp_795_16 = __tmp_799_16;
  assign __tmp_795_17 = __tmp_799_17;
  assign __tmp_795_18 = __tmp_799_18;
  assign __tmp_795_19 = __tmp_799_19;
  assign __tmp_795_2 = __tmp_799_2;
  assign __tmp_795_20 = __tmp_799_20;
  assign __tmp_795_21 = __tmp_799_21;
  assign __tmp_795_22 = __tmp_799_22;
  assign __tmp_795_23 = __tmp_799_23;
  assign __tmp_795_24 = __tmp_799_24;
  assign __tmp_795_25 = __tmp_799_25;
  assign __tmp_795_26 = __tmp_799_26;
  assign __tmp_795_27 = __tmp_799_27;
  assign __tmp_795_28 = __tmp_799_28;
  assign __tmp_795_29 = __tmp_799_29;
  assign __tmp_795_3 = __tmp_799_3;
  assign __tmp_795_30 = __tmp_799_30;
  assign __tmp_795_31 = __tmp_799_31;
  assign __tmp_795_32 = __tmp_799_32;
  assign __tmp_795_33 = __tmp_799_33;
  assign __tmp_795_34 = __tmp_799_34;
  assign __tmp_795_4 = __tmp_799_4;
  assign __tmp_795_5 = __tmp_799_5;
  assign __tmp_795_6 = __tmp_799_6;
  assign __tmp_795_7 = __tmp_799_7;
  assign __tmp_795_8 = __tmp_799_8;
  assign __tmp_795_9 = __tmp_799_9;
  assign __tmp_797_1 = __tmp_799_1;
  assign __tmp_797_10 = __tmp_799_10;
  assign __tmp_797_11 = __tmp_799_11;
  assign __tmp_797_12 = __tmp_799_12;
  assign __tmp_797_13 = __tmp_799_13;
  assign __tmp_797_14 = __tmp_799_14;
  assign __tmp_797_15 = __tmp_799_15;
  assign __tmp_797_16 = __tmp_799_16;
  assign __tmp_797_17 = __tmp_799_17;
  assign __tmp_797_18 = __tmp_799_18;
  assign __tmp_797_19 = __tmp_799_19;
  assign __tmp_797_2 = __tmp_799_2;
  assign __tmp_797_20 = __tmp_799_20;
  assign __tmp_797_21 = __tmp_799_21;
  assign __tmp_797_22 = __tmp_799_22;
  assign __tmp_797_23 = __tmp_799_23;
  assign __tmp_797_24 = __tmp_799_24;
  assign __tmp_797_25 = __tmp_799_25;
  assign __tmp_797_26 = __tmp_799_26;
  assign __tmp_797_27 = __tmp_799_27;
  assign __tmp_797_28 = __tmp_799_28;
  assign __tmp_797_29 = __tmp_799_29;
  assign __tmp_797_3 = __tmp_799_3;
  assign __tmp_797_30 = __tmp_799_30;
  assign __tmp_797_31 = __tmp_799_31;
  assign __tmp_797_32 = __tmp_799_32;
  assign __tmp_797_33 = __tmp_799_33;
  assign __tmp_797_34 = __tmp_799_34;
  assign __tmp_797_4 = __tmp_799_4;
  assign __tmp_797_5 = __tmp_799_5;
  assign __tmp_797_6 = __tmp_799_6;
  assign __tmp_797_7 = __tmp_799_7;
  assign __tmp_797_8 = __tmp_799_8;
  assign __tmp_797_9 = __tmp_799_9;
  assign __tmp_801_1 = __tmp_947_1;
  assign __tmp_803_1 = __tmp_947_1;
  assign __tmp_803_2 = __tmp_947_2;
  assign __tmp_803_3 = __tmp_947_3;
  assign __tmp_803_4 = __tmp_947_4;
  assign __tmp_803_5 = __tmp_947_5;
  assign __tmp_803_6 = __tmp_947_6;
  assign __tmp_803_7 = __tmp_947_7;
  assign __tmp_803_8 = __tmp_947_8;
  assign __tmp_803_9 = __tmp_947_9;
  assign __tmp_805_1 = __tmp_947_1;
  assign __tmp_805_2 = __tmp_947_2;
  assign __tmp_805_3 = __tmp_947_3;
  assign __tmp_805_4 = __tmp_947_4;
  assign __tmp_805_5 = __tmp_947_5;
  assign __tmp_805_6 = __tmp_947_6;
  assign __tmp_805_7 = __tmp_947_7;
  assign __tmp_805_8 = __tmp_947_8;
  assign __tmp_805_9 = __tmp_947_9;
  assign __tmp_807_1 = __tmp_947_1;
  assign __tmp_807_2 = __tmp_947_2;
  assign __tmp_807_3 = __tmp_947_3;
  assign __tmp_807_4 = __tmp_947_4;
  assign __tmp_807_5 = __tmp_947_5;
  assign __tmp_807_6 = __tmp_947_6;
  assign __tmp_807_7 = __tmp_947_7;
  assign __tmp_807_8 = __tmp_947_8;
  assign __tmp_807_9 = __tmp_947_9;
  assign __tmp_809_1 = __tmp_947_1;
  assign __tmp_809_10 = __tmp_959_10;
  assign __tmp_809_11 = __tmp_959_11;
  assign __tmp_809_12 = __tmp_959_12;
  assign __tmp_809_2 = __tmp_947_2;
  assign __tmp_809_3 = __tmp_947_3;
  assign __tmp_809_4 = __tmp_947_4;
  assign __tmp_809_5 = __tmp_947_5;
  assign __tmp_809_6 = __tmp_947_6;
  assign __tmp_809_7 = __tmp_947_7;
  assign __tmp_809_8 = __tmp_947_8;
  assign __tmp_809_9 = __tmp_947_9;
  assign __tmp_811_1 = __tmp_947_1;
  assign __tmp_811_10 = __tmp_959_10;
  assign __tmp_811_11 = __tmp_959_11;
  assign __tmp_811_12 = __tmp_959_12;
  assign __tmp_811_2 = __tmp_947_2;
  assign __tmp_811_3 = __tmp_947_3;
  assign __tmp_811_4 = __tmp_947_4;
  assign __tmp_811_5 = __tmp_947_5;
  assign __tmp_811_6 = __tmp_947_6;
  assign __tmp_811_7 = __tmp_947_7;
  assign __tmp_811_8 = __tmp_947_8;
  assign __tmp_811_9 = __tmp_947_9;
  assign __tmp_813_1 = __tmp_947_1;
  assign __tmp_813_10 = __tmp_959_10;
  assign __tmp_813_11 = __tmp_959_11;
  assign __tmp_813_12 = __tmp_959_12;
  assign __tmp_813_2 = __tmp_947_2;
  assign __tmp_813_3 = __tmp_947_3;
  assign __tmp_813_4 = __tmp_947_4;
  assign __tmp_813_5 = __tmp_947_5;
  assign __tmp_813_6 = __tmp_947_6;
  assign __tmp_813_7 = __tmp_947_7;
  assign __tmp_813_8 = __tmp_947_8;
  assign __tmp_813_9 = __tmp_947_9;
  assign __tmp_815_1 = __tmp_947_1;
  assign __tmp_815_2 = __tmp_947_2;
  assign __tmp_815_3 = __tmp_947_3;
  assign __tmp_815_4 = __tmp_947_4;
  assign __tmp_815_5 = __tmp_947_5;
  assign __tmp_815_6 = __tmp_947_6;
  assign __tmp_815_7 = __tmp_947_7;
  assign __tmp_815_8 = __tmp_947_8;
  assign __tmp_815_9 = __tmp_947_9;
  assign __tmp_817_1 = __tmp_947_1;
  assign __tmp_817_2 = __tmp_947_2;
  assign __tmp_817_3 = __tmp_947_3;
  assign __tmp_817_4 = __tmp_947_4;
  assign __tmp_817_5 = __tmp_947_5;
  assign __tmp_817_6 = __tmp_947_6;
  assign __tmp_817_7 = __tmp_947_7;
  assign __tmp_817_8 = __tmp_947_8;
  assign __tmp_817_9 = __tmp_947_9;
  assign __tmp_819_1 = __tmp_947_1;
  assign __tmp_819_2 = __tmp_947_2;
  assign __tmp_819_3 = __tmp_947_3;
  assign __tmp_819_4 = __tmp_947_4;
  assign __tmp_819_5 = __tmp_947_5;
  assign __tmp_819_6 = __tmp_947_6;
  assign __tmp_819_7 = __tmp_947_7;
  assign __tmp_819_8 = __tmp_947_8;
  assign __tmp_819_9 = __tmp_947_9;
  assign __tmp_821_1 = __tmp_947_1;
  assign __tmp_821_10 = __tmp_959_10;
  assign __tmp_821_11 = __tmp_959_11;
  assign __tmp_821_12 = __tmp_959_12;
  assign __tmp_821_2 = __tmp_947_2;
  assign __tmp_821_3 = __tmp_947_3;
  assign __tmp_821_4 = __tmp_947_4;
  assign __tmp_821_5 = __tmp_947_5;
  assign __tmp_821_6 = __tmp_947_6;
  assign __tmp_821_7 = __tmp_947_7;
  assign __tmp_821_8 = __tmp_947_8;
  assign __tmp_821_9 = __tmp_947_9;
  assign __tmp_823_1 = __tmp_947_1;
  assign __tmp_823_10 = __tmp_959_10;
  assign __tmp_823_11 = __tmp_959_11;
  assign __tmp_823_12 = __tmp_959_12;
  assign __tmp_823_2 = __tmp_947_2;
  assign __tmp_823_3 = __tmp_947_3;
  assign __tmp_823_4 = __tmp_947_4;
  assign __tmp_823_5 = __tmp_947_5;
  assign __tmp_823_6 = __tmp_947_6;
  assign __tmp_823_7 = __tmp_947_7;
  assign __tmp_823_8 = __tmp_947_8;
  assign __tmp_823_9 = __tmp_947_9;
  assign __tmp_825_1 = __tmp_947_1;
  assign __tmp_825_10 = __tmp_959_10;
  assign __tmp_825_11 = __tmp_959_11;
  assign __tmp_825_12 = __tmp_959_12;
  assign __tmp_825_2 = __tmp_947_2;
  assign __tmp_825_3 = __tmp_947_3;
  assign __tmp_825_4 = __tmp_947_4;
  assign __tmp_825_5 = __tmp_947_5;
  assign __tmp_825_6 = __tmp_947_6;
  assign __tmp_825_7 = __tmp_947_7;
  assign __tmp_825_8 = __tmp_947_8;
  assign __tmp_825_9 = __tmp_947_9;
  assign __tmp_827_1 = __tmp_947_1;
  assign __tmp_827_2 = __tmp_947_2;
  assign __tmp_827_3 = __tmp_947_3;
  assign __tmp_827_4 = __tmp_947_4;
  assign __tmp_827_5 = __tmp_947_5;
  assign __tmp_827_6 = __tmp_947_6;
  assign __tmp_827_7 = __tmp_947_7;
  assign __tmp_827_8 = __tmp_947_8;
  assign __tmp_827_9 = __tmp_947_9;
  assign __tmp_829_1 = __tmp_947_1;
  assign __tmp_829_2 = __tmp_947_2;
  assign __tmp_829_3 = __tmp_947_3;
  assign __tmp_829_4 = __tmp_947_4;
  assign __tmp_829_5 = __tmp_947_5;
  assign __tmp_829_6 = __tmp_947_6;
  assign __tmp_829_7 = __tmp_947_7;
  assign __tmp_829_8 = __tmp_947_8;
  assign __tmp_829_9 = __tmp_947_9;
  assign __tmp_831_1 = __tmp_947_1;
  assign __tmp_831_2 = __tmp_947_2;
  assign __tmp_831_3 = __tmp_947_3;
  assign __tmp_831_4 = __tmp_947_4;
  assign __tmp_831_5 = __tmp_947_5;
  assign __tmp_831_6 = __tmp_947_6;
  assign __tmp_831_7 = __tmp_947_7;
  assign __tmp_831_8 = __tmp_947_8;
  assign __tmp_831_9 = __tmp_947_9;
  assign __tmp_833_1 = __tmp_947_1;
  assign __tmp_833_10 = __tmp_959_10;
  assign __tmp_833_11 = __tmp_959_11;
  assign __tmp_833_12 = __tmp_959_12;
  assign __tmp_833_2 = __tmp_947_2;
  assign __tmp_833_3 = __tmp_947_3;
  assign __tmp_833_4 = __tmp_947_4;
  assign __tmp_833_5 = __tmp_947_5;
  assign __tmp_833_6 = __tmp_947_6;
  assign __tmp_833_7 = __tmp_947_7;
  assign __tmp_833_8 = __tmp_947_8;
  assign __tmp_833_9 = __tmp_947_9;
  assign __tmp_835_1 = __tmp_947_1;
  assign __tmp_835_10 = __tmp_959_10;
  assign __tmp_835_11 = __tmp_959_11;
  assign __tmp_835_12 = __tmp_959_12;
  assign __tmp_835_2 = __tmp_947_2;
  assign __tmp_835_3 = __tmp_947_3;
  assign __tmp_835_4 = __tmp_947_4;
  assign __tmp_835_5 = __tmp_947_5;
  assign __tmp_835_6 = __tmp_947_6;
  assign __tmp_835_7 = __tmp_947_7;
  assign __tmp_835_8 = __tmp_947_8;
  assign __tmp_835_9 = __tmp_947_9;
  assign __tmp_837_1 = __tmp_947_1;
  assign __tmp_837_10 = __tmp_959_10;
  assign __tmp_837_11 = __tmp_959_11;
  assign __tmp_837_12 = __tmp_959_12;
  assign __tmp_837_2 = __tmp_947_2;
  assign __tmp_837_3 = __tmp_947_3;
  assign __tmp_837_4 = __tmp_947_4;
  assign __tmp_837_5 = __tmp_947_5;
  assign __tmp_837_6 = __tmp_947_6;
  assign __tmp_837_7 = __tmp_947_7;
  assign __tmp_837_8 = __tmp_947_8;
  assign __tmp_837_9 = __tmp_947_9;
  assign __tmp_839_1 = __tmp_947_1;
  assign __tmp_839_2 = __tmp_947_2;
  assign __tmp_839_3 = __tmp_947_3;
  assign __tmp_839_4 = __tmp_947_4;
  assign __tmp_839_5 = __tmp_947_5;
  assign __tmp_839_6 = __tmp_947_6;
  assign __tmp_839_7 = __tmp_947_7;
  assign __tmp_839_8 = __tmp_947_8;
  assign __tmp_839_9 = __tmp_947_9;
  assign __tmp_841_1 = __tmp_947_1;
  assign __tmp_841_2 = __tmp_947_2;
  assign __tmp_841_3 = __tmp_947_3;
  assign __tmp_841_4 = __tmp_947_4;
  assign __tmp_841_5 = __tmp_947_5;
  assign __tmp_841_6 = __tmp_947_6;
  assign __tmp_841_7 = __tmp_947_7;
  assign __tmp_841_8 = __tmp_947_8;
  assign __tmp_841_9 = __tmp_947_9;
  assign __tmp_843_1 = __tmp_947_1;
  assign __tmp_843_2 = __tmp_947_2;
  assign __tmp_843_3 = __tmp_947_3;
  assign __tmp_843_4 = __tmp_947_4;
  assign __tmp_843_5 = __tmp_947_5;
  assign __tmp_843_6 = __tmp_947_6;
  assign __tmp_843_7 = __tmp_947_7;
  assign __tmp_843_8 = __tmp_947_8;
  assign __tmp_843_9 = __tmp_947_9;
  assign __tmp_845_1 = __tmp_947_1;
  assign __tmp_845_10 = __tmp_959_10;
  assign __tmp_845_11 = __tmp_959_11;
  assign __tmp_845_12 = __tmp_959_12;
  assign __tmp_845_2 = __tmp_947_2;
  assign __tmp_845_3 = __tmp_947_3;
  assign __tmp_845_4 = __tmp_947_4;
  assign __tmp_845_5 = __tmp_947_5;
  assign __tmp_845_6 = __tmp_947_6;
  assign __tmp_845_7 = __tmp_947_7;
  assign __tmp_845_8 = __tmp_947_8;
  assign __tmp_845_9 = __tmp_947_9;
  assign __tmp_847_1 = __tmp_947_1;
  assign __tmp_847_10 = __tmp_959_10;
  assign __tmp_847_11 = __tmp_959_11;
  assign __tmp_847_12 = __tmp_959_12;
  assign __tmp_847_2 = __tmp_947_2;
  assign __tmp_847_3 = __tmp_947_3;
  assign __tmp_847_4 = __tmp_947_4;
  assign __tmp_847_5 = __tmp_947_5;
  assign __tmp_847_6 = __tmp_947_6;
  assign __tmp_847_7 = __tmp_947_7;
  assign __tmp_847_8 = __tmp_947_8;
  assign __tmp_847_9 = __tmp_947_9;
  assign __tmp_849_1 = __tmp_947_1;
  assign __tmp_849_10 = __tmp_959_10;
  assign __tmp_849_11 = __tmp_959_11;
  assign __tmp_849_12 = __tmp_959_12;
  assign __tmp_849_2 = __tmp_947_2;
  assign __tmp_849_3 = __tmp_947_3;
  assign __tmp_849_4 = __tmp_947_4;
  assign __tmp_849_5 = __tmp_947_5;
  assign __tmp_849_6 = __tmp_947_6;
  assign __tmp_849_7 = __tmp_947_7;
  assign __tmp_849_8 = __tmp_947_8;
  assign __tmp_849_9 = __tmp_947_9;
  assign __tmp_851_1 = __tmp_947_1;
  assign __tmp_851_2 = __tmp_947_2;
  assign __tmp_851_3 = __tmp_947_3;
  assign __tmp_851_4 = __tmp_947_4;
  assign __tmp_851_5 = __tmp_947_5;
  assign __tmp_851_6 = __tmp_947_6;
  assign __tmp_851_7 = __tmp_947_7;
  assign __tmp_851_8 = __tmp_947_8;
  assign __tmp_851_9 = __tmp_947_9;
  assign __tmp_853_1 = __tmp_947_1;
  assign __tmp_853_2 = __tmp_947_2;
  assign __tmp_853_3 = __tmp_947_3;
  assign __tmp_853_4 = __tmp_947_4;
  assign __tmp_853_5 = __tmp_947_5;
  assign __tmp_853_6 = __tmp_947_6;
  assign __tmp_853_7 = __tmp_947_7;
  assign __tmp_853_8 = __tmp_947_8;
  assign __tmp_853_9 = __tmp_947_9;
  assign __tmp_855_1 = __tmp_947_1;
  assign __tmp_855_2 = __tmp_947_2;
  assign __tmp_855_3 = __tmp_947_3;
  assign __tmp_855_4 = __tmp_947_4;
  assign __tmp_855_5 = __tmp_947_5;
  assign __tmp_855_6 = __tmp_947_6;
  assign __tmp_855_7 = __tmp_947_7;
  assign __tmp_855_8 = __tmp_947_8;
  assign __tmp_855_9 = __tmp_947_9;
  assign __tmp_857_1 = __tmp_947_1;
  assign __tmp_857_10 = __tmp_959_10;
  assign __tmp_857_11 = __tmp_959_11;
  assign __tmp_857_12 = __tmp_959_12;
  assign __tmp_857_2 = __tmp_947_2;
  assign __tmp_857_3 = __tmp_947_3;
  assign __tmp_857_4 = __tmp_947_4;
  assign __tmp_857_5 = __tmp_947_5;
  assign __tmp_857_6 = __tmp_947_6;
  assign __tmp_857_7 = __tmp_947_7;
  assign __tmp_857_8 = __tmp_947_8;
  assign __tmp_857_9 = __tmp_947_9;
  assign __tmp_859_1 = __tmp_947_1;
  assign __tmp_859_10 = __tmp_959_10;
  assign __tmp_859_11 = __tmp_959_11;
  assign __tmp_859_12 = __tmp_959_12;
  assign __tmp_859_2 = __tmp_947_2;
  assign __tmp_859_3 = __tmp_947_3;
  assign __tmp_859_4 = __tmp_947_4;
  assign __tmp_859_5 = __tmp_947_5;
  assign __tmp_859_6 = __tmp_947_6;
  assign __tmp_859_7 = __tmp_947_7;
  assign __tmp_859_8 = __tmp_947_8;
  assign __tmp_859_9 = __tmp_947_9;
  assign __tmp_861_1 = __tmp_947_1;
  assign __tmp_861_10 = __tmp_959_10;
  assign __tmp_861_11 = __tmp_959_11;
  assign __tmp_861_12 = __tmp_959_12;
  assign __tmp_861_2 = __tmp_947_2;
  assign __tmp_861_3 = __tmp_947_3;
  assign __tmp_861_4 = __tmp_947_4;
  assign __tmp_861_5 = __tmp_947_5;
  assign __tmp_861_6 = __tmp_947_6;
  assign __tmp_861_7 = __tmp_947_7;
  assign __tmp_861_8 = __tmp_947_8;
  assign __tmp_861_9 = __tmp_947_9;
  assign __tmp_863_1 = __tmp_947_1;
  assign __tmp_863_2 = __tmp_947_2;
  assign __tmp_863_3 = __tmp_947_3;
  assign __tmp_863_4 = __tmp_947_4;
  assign __tmp_863_5 = __tmp_947_5;
  assign __tmp_863_6 = __tmp_947_6;
  assign __tmp_863_7 = __tmp_947_7;
  assign __tmp_863_8 = __tmp_947_8;
  assign __tmp_863_9 = __tmp_947_9;
  assign __tmp_865_1 = __tmp_947_1;
  assign __tmp_865_2 = __tmp_947_2;
  assign __tmp_865_3 = __tmp_947_3;
  assign __tmp_865_4 = __tmp_947_4;
  assign __tmp_865_5 = __tmp_947_5;
  assign __tmp_865_6 = __tmp_947_6;
  assign __tmp_865_7 = __tmp_947_7;
  assign __tmp_865_8 = __tmp_947_8;
  assign __tmp_865_9 = __tmp_947_9;
  assign __tmp_867_1 = __tmp_947_1;
  assign __tmp_867_2 = __tmp_947_2;
  assign __tmp_867_3 = __tmp_947_3;
  assign __tmp_867_4 = __tmp_947_4;
  assign __tmp_867_5 = __tmp_947_5;
  assign __tmp_867_6 = __tmp_947_6;
  assign __tmp_867_7 = __tmp_947_7;
  assign __tmp_867_8 = __tmp_947_8;
  assign __tmp_867_9 = __tmp_947_9;
  assign __tmp_869_1 = __tmp_947_1;
  assign __tmp_869_10 = __tmp_959_10;
  assign __tmp_869_11 = __tmp_959_11;
  assign __tmp_869_12 = __tmp_959_12;
  assign __tmp_869_2 = __tmp_947_2;
  assign __tmp_869_3 = __tmp_947_3;
  assign __tmp_869_4 = __tmp_947_4;
  assign __tmp_869_5 = __tmp_947_5;
  assign __tmp_869_6 = __tmp_947_6;
  assign __tmp_869_7 = __tmp_947_7;
  assign __tmp_869_8 = __tmp_947_8;
  assign __tmp_869_9 = __tmp_947_9;
  assign __tmp_871_1 = __tmp_947_1;
  assign __tmp_871_10 = __tmp_959_10;
  assign __tmp_871_11 = __tmp_959_11;
  assign __tmp_871_12 = __tmp_959_12;
  assign __tmp_871_2 = __tmp_947_2;
  assign __tmp_871_3 = __tmp_947_3;
  assign __tmp_871_4 = __tmp_947_4;
  assign __tmp_871_5 = __tmp_947_5;
  assign __tmp_871_6 = __tmp_947_6;
  assign __tmp_871_7 = __tmp_947_7;
  assign __tmp_871_8 = __tmp_947_8;
  assign __tmp_871_9 = __tmp_947_9;
  assign __tmp_873_1 = __tmp_947_1;
  assign __tmp_873_10 = __tmp_959_10;
  assign __tmp_873_11 = __tmp_959_11;
  assign __tmp_873_12 = __tmp_959_12;
  assign __tmp_873_2 = __tmp_947_2;
  assign __tmp_873_3 = __tmp_947_3;
  assign __tmp_873_4 = __tmp_947_4;
  assign __tmp_873_5 = __tmp_947_5;
  assign __tmp_873_6 = __tmp_947_6;
  assign __tmp_873_7 = __tmp_947_7;
  assign __tmp_873_8 = __tmp_947_8;
  assign __tmp_873_9 = __tmp_947_9;
  assign __tmp_875_1 = __tmp_947_1;
  assign __tmp_875_2 = __tmp_947_2;
  assign __tmp_875_3 = __tmp_947_3;
  assign __tmp_875_4 = __tmp_947_4;
  assign __tmp_875_5 = __tmp_947_5;
  assign __tmp_875_6 = __tmp_947_6;
  assign __tmp_875_7 = __tmp_947_7;
  assign __tmp_875_8 = __tmp_947_8;
  assign __tmp_875_9 = __tmp_947_9;
  assign __tmp_877_1 = __tmp_947_1;
  assign __tmp_877_2 = __tmp_947_2;
  assign __tmp_877_3 = __tmp_947_3;
  assign __tmp_877_4 = __tmp_947_4;
  assign __tmp_877_5 = __tmp_947_5;
  assign __tmp_877_6 = __tmp_947_6;
  assign __tmp_877_7 = __tmp_947_7;
  assign __tmp_877_8 = __tmp_947_8;
  assign __tmp_877_9 = __tmp_947_9;
  assign __tmp_879_1 = __tmp_947_1;
  assign __tmp_879_2 = __tmp_947_2;
  assign __tmp_879_3 = __tmp_947_3;
  assign __tmp_879_4 = __tmp_947_4;
  assign __tmp_879_5 = __tmp_947_5;
  assign __tmp_879_6 = __tmp_947_6;
  assign __tmp_879_7 = __tmp_947_7;
  assign __tmp_879_8 = __tmp_947_8;
  assign __tmp_879_9 = __tmp_947_9;
  assign __tmp_881_1 = __tmp_947_1;
  assign __tmp_881_10 = __tmp_959_10;
  assign __tmp_881_11 = __tmp_959_11;
  assign __tmp_881_12 = __tmp_959_12;
  assign __tmp_881_2 = __tmp_947_2;
  assign __tmp_881_3 = __tmp_947_3;
  assign __tmp_881_4 = __tmp_947_4;
  assign __tmp_881_5 = __tmp_947_5;
  assign __tmp_881_6 = __tmp_947_6;
  assign __tmp_881_7 = __tmp_947_7;
  assign __tmp_881_8 = __tmp_947_8;
  assign __tmp_881_9 = __tmp_947_9;
  assign __tmp_883_1 = __tmp_947_1;
  assign __tmp_883_10 = __tmp_959_10;
  assign __tmp_883_11 = __tmp_959_11;
  assign __tmp_883_12 = __tmp_959_12;
  assign __tmp_883_2 = __tmp_947_2;
  assign __tmp_883_3 = __tmp_947_3;
  assign __tmp_883_4 = __tmp_947_4;
  assign __tmp_883_5 = __tmp_947_5;
  assign __tmp_883_6 = __tmp_947_6;
  assign __tmp_883_7 = __tmp_947_7;
  assign __tmp_883_8 = __tmp_947_8;
  assign __tmp_883_9 = __tmp_947_9;
  assign __tmp_885_1 = __tmp_947_1;
  assign __tmp_885_10 = __tmp_959_10;
  assign __tmp_885_11 = __tmp_959_11;
  assign __tmp_885_12 = __tmp_959_12;
  assign __tmp_885_2 = __tmp_947_2;
  assign __tmp_885_3 = __tmp_947_3;
  assign __tmp_885_4 = __tmp_947_4;
  assign __tmp_885_5 = __tmp_947_5;
  assign __tmp_885_6 = __tmp_947_6;
  assign __tmp_885_7 = __tmp_947_7;
  assign __tmp_885_8 = __tmp_947_8;
  assign __tmp_885_9 = __tmp_947_9;
  assign __tmp_887_1 = __tmp_947_1;
  assign __tmp_887_2 = __tmp_947_2;
  assign __tmp_887_3 = __tmp_947_3;
  assign __tmp_887_4 = __tmp_947_4;
  assign __tmp_887_5 = __tmp_947_5;
  assign __tmp_887_6 = __tmp_947_6;
  assign __tmp_887_7 = __tmp_947_7;
  assign __tmp_887_8 = __tmp_947_8;
  assign __tmp_887_9 = __tmp_947_9;
  assign __tmp_889_1 = __tmp_947_1;
  assign __tmp_889_2 = __tmp_947_2;
  assign __tmp_889_3 = __tmp_947_3;
  assign __tmp_889_4 = __tmp_947_4;
  assign __tmp_889_5 = __tmp_947_5;
  assign __tmp_889_6 = __tmp_947_6;
  assign __tmp_889_7 = __tmp_947_7;
  assign __tmp_889_8 = __tmp_947_8;
  assign __tmp_889_9 = __tmp_947_9;
  assign __tmp_891_1 = __tmp_947_1;
  assign __tmp_891_2 = __tmp_947_2;
  assign __tmp_891_3 = __tmp_947_3;
  assign __tmp_891_4 = __tmp_947_4;
  assign __tmp_891_5 = __tmp_947_5;
  assign __tmp_891_6 = __tmp_947_6;
  assign __tmp_891_7 = __tmp_947_7;
  assign __tmp_891_8 = __tmp_947_8;
  assign __tmp_891_9 = __tmp_947_9;
  assign __tmp_893_1 = __tmp_947_1;
  assign __tmp_893_10 = __tmp_959_10;
  assign __tmp_893_11 = __tmp_959_11;
  assign __tmp_893_12 = __tmp_959_12;
  assign __tmp_893_2 = __tmp_947_2;
  assign __tmp_893_3 = __tmp_947_3;
  assign __tmp_893_4 = __tmp_947_4;
  assign __tmp_893_5 = __tmp_947_5;
  assign __tmp_893_6 = __tmp_947_6;
  assign __tmp_893_7 = __tmp_947_7;
  assign __tmp_893_8 = __tmp_947_8;
  assign __tmp_893_9 = __tmp_947_9;
  assign __tmp_895_1 = __tmp_947_1;
  assign __tmp_895_10 = __tmp_959_10;
  assign __tmp_895_11 = __tmp_959_11;
  assign __tmp_895_12 = __tmp_959_12;
  assign __tmp_895_2 = __tmp_947_2;
  assign __tmp_895_3 = __tmp_947_3;
  assign __tmp_895_4 = __tmp_947_4;
  assign __tmp_895_5 = __tmp_947_5;
  assign __tmp_895_6 = __tmp_947_6;
  assign __tmp_895_7 = __tmp_947_7;
  assign __tmp_895_8 = __tmp_947_8;
  assign __tmp_895_9 = __tmp_947_9;
  assign __tmp_897_1 = __tmp_947_1;
  assign __tmp_897_10 = __tmp_959_10;
  assign __tmp_897_11 = __tmp_959_11;
  assign __tmp_897_12 = __tmp_959_12;
  assign __tmp_897_2 = __tmp_947_2;
  assign __tmp_897_3 = __tmp_947_3;
  assign __tmp_897_4 = __tmp_947_4;
  assign __tmp_897_5 = __tmp_947_5;
  assign __tmp_897_6 = __tmp_947_6;
  assign __tmp_897_7 = __tmp_947_7;
  assign __tmp_897_8 = __tmp_947_8;
  assign __tmp_897_9 = __tmp_947_9;
  assign __tmp_899_1 = __tmp_947_1;
  assign __tmp_899_2 = __tmp_947_2;
  assign __tmp_899_3 = __tmp_947_3;
  assign __tmp_899_4 = __tmp_947_4;
  assign __tmp_899_5 = __tmp_947_5;
  assign __tmp_899_6 = __tmp_947_6;
  assign __tmp_899_7 = __tmp_947_7;
  assign __tmp_899_8 = __tmp_947_8;
  assign __tmp_899_9 = __tmp_947_9;
  assign __tmp_901_1 = __tmp_947_1;
  assign __tmp_901_2 = __tmp_947_2;
  assign __tmp_901_3 = __tmp_947_3;
  assign __tmp_901_4 = __tmp_947_4;
  assign __tmp_901_5 = __tmp_947_5;
  assign __tmp_901_6 = __tmp_947_6;
  assign __tmp_901_7 = __tmp_947_7;
  assign __tmp_901_8 = __tmp_947_8;
  assign __tmp_901_9 = __tmp_947_9;
  assign __tmp_903_1 = __tmp_947_1;
  assign __tmp_903_2 = __tmp_947_2;
  assign __tmp_903_3 = __tmp_947_3;
  assign __tmp_903_4 = __tmp_947_4;
  assign __tmp_903_5 = __tmp_947_5;
  assign __tmp_903_6 = __tmp_947_6;
  assign __tmp_903_7 = __tmp_947_7;
  assign __tmp_903_8 = __tmp_947_8;
  assign __tmp_903_9 = __tmp_947_9;
  assign __tmp_905_1 = __tmp_947_1;
  assign __tmp_905_10 = __tmp_959_10;
  assign __tmp_905_11 = __tmp_959_11;
  assign __tmp_905_12 = __tmp_959_12;
  assign __tmp_905_2 = __tmp_947_2;
  assign __tmp_905_3 = __tmp_947_3;
  assign __tmp_905_4 = __tmp_947_4;
  assign __tmp_905_5 = __tmp_947_5;
  assign __tmp_905_6 = __tmp_947_6;
  assign __tmp_905_7 = __tmp_947_7;
  assign __tmp_905_8 = __tmp_947_8;
  assign __tmp_905_9 = __tmp_947_9;
  assign __tmp_907_1 = __tmp_947_1;
  assign __tmp_907_10 = __tmp_959_10;
  assign __tmp_907_11 = __tmp_959_11;
  assign __tmp_907_12 = __tmp_959_12;
  assign __tmp_907_2 = __tmp_947_2;
  assign __tmp_907_3 = __tmp_947_3;
  assign __tmp_907_4 = __tmp_947_4;
  assign __tmp_907_5 = __tmp_947_5;
  assign __tmp_907_6 = __tmp_947_6;
  assign __tmp_907_7 = __tmp_947_7;
  assign __tmp_907_8 = __tmp_947_8;
  assign __tmp_907_9 = __tmp_947_9;
  assign __tmp_909_1 = __tmp_947_1;
  assign __tmp_909_10 = __tmp_959_10;
  assign __tmp_909_11 = __tmp_959_11;
  assign __tmp_909_12 = __tmp_959_12;
  assign __tmp_909_2 = __tmp_947_2;
  assign __tmp_909_3 = __tmp_947_3;
  assign __tmp_909_4 = __tmp_947_4;
  assign __tmp_909_5 = __tmp_947_5;
  assign __tmp_909_6 = __tmp_947_6;
  assign __tmp_909_7 = __tmp_947_7;
  assign __tmp_909_8 = __tmp_947_8;
  assign __tmp_909_9 = __tmp_947_9;
  assign __tmp_911_1 = __tmp_947_1;
  assign __tmp_911_10 = __tmp_959_10;
  assign __tmp_911_11 = __tmp_959_11;
  assign __tmp_911_12 = __tmp_959_12;
  assign __tmp_911_13 = __tmp_969_13;
  assign __tmp_911_14 = __tmp_969_14;
  assign __tmp_911_15 = __tmp_969_15;
  assign __tmp_911_16 = __tmp_969_16;
  assign __tmp_911_17 = __tmp_969_17;
  assign __tmp_911_18 = __tmp_969_18;
  assign __tmp_911_19 = __tmp_969_19;
  assign __tmp_911_2 = __tmp_947_2;
  assign __tmp_911_3 = __tmp_947_3;
  assign __tmp_911_4 = __tmp_947_4;
  assign __tmp_911_5 = __tmp_947_5;
  assign __tmp_911_6 = __tmp_947_6;
  assign __tmp_911_7 = __tmp_947_7;
  assign __tmp_911_8 = __tmp_947_8;
  assign __tmp_911_9 = __tmp_947_9;
  assign __tmp_913_1 = __tmp_947_1;
  assign __tmp_913_10 = __tmp_959_10;
  assign __tmp_913_11 = __tmp_959_11;
  assign __tmp_913_12 = __tmp_959_12;
  assign __tmp_913_13 = __tmp_969_13;
  assign __tmp_913_14 = __tmp_969_14;
  assign __tmp_913_15 = __tmp_969_15;
  assign __tmp_913_16 = __tmp_969_16;
  assign __tmp_913_17 = __tmp_969_17;
  assign __tmp_913_18 = __tmp_969_18;
  assign __tmp_913_19 = __tmp_969_19;
  assign __tmp_913_2 = __tmp_947_2;
  assign __tmp_913_3 = __tmp_947_3;
  assign __tmp_913_4 = __tmp_947_4;
  assign __tmp_913_5 = __tmp_947_5;
  assign __tmp_913_6 = __tmp_947_6;
  assign __tmp_913_7 = __tmp_947_7;
  assign __tmp_913_8 = __tmp_947_8;
  assign __tmp_913_9 = __tmp_947_9;
  assign __tmp_915_1 = __tmp_947_1;
  assign __tmp_915_10 = __tmp_959_10;
  assign __tmp_915_11 = __tmp_959_11;
  assign __tmp_915_12 = __tmp_959_12;
  assign __tmp_915_13 = __tmp_969_13;
  assign __tmp_915_14 = __tmp_969_14;
  assign __tmp_915_15 = __tmp_969_15;
  assign __tmp_915_16 = __tmp_969_16;
  assign __tmp_915_17 = __tmp_969_17;
  assign __tmp_915_18 = __tmp_969_18;
  assign __tmp_915_19 = __tmp_969_19;
  assign __tmp_915_2 = __tmp_947_2;
  assign __tmp_915_3 = __tmp_947_3;
  assign __tmp_915_4 = __tmp_947_4;
  assign __tmp_915_5 = __tmp_947_5;
  assign __tmp_915_6 = __tmp_947_6;
  assign __tmp_915_7 = __tmp_947_7;
  assign __tmp_915_8 = __tmp_947_8;
  assign __tmp_915_9 = __tmp_947_9;
  assign __tmp_917_1 = __tmp_947_1;
  assign __tmp_917_10 = __tmp_959_10;
  assign __tmp_917_11 = __tmp_959_11;
  assign __tmp_917_12 = __tmp_959_12;
  assign __tmp_917_13 = __tmp_969_13;
  assign __tmp_917_14 = __tmp_969_14;
  assign __tmp_917_15 = __tmp_969_15;
  assign __tmp_917_16 = __tmp_969_16;
  assign __tmp_917_17 = __tmp_969_17;
  assign __tmp_917_18 = __tmp_969_18;
  assign __tmp_917_19 = __tmp_969_19;
  assign __tmp_917_2 = __tmp_947_2;
  assign __tmp_917_3 = __tmp_947_3;
  assign __tmp_917_4 = __tmp_947_4;
  assign __tmp_917_5 = __tmp_947_5;
  assign __tmp_917_6 = __tmp_947_6;
  assign __tmp_917_7 = __tmp_947_7;
  assign __tmp_917_8 = __tmp_947_8;
  assign __tmp_917_9 = __tmp_947_9;
  assign __tmp_919_1 = __tmp_947_1;
  assign __tmp_919_10 = __tmp_959_10;
  assign __tmp_919_11 = __tmp_959_11;
  assign __tmp_919_12 = __tmp_959_12;
  assign __tmp_919_13 = __tmp_969_13;
  assign __tmp_919_14 = __tmp_969_14;
  assign __tmp_919_15 = __tmp_969_15;
  assign __tmp_919_16 = __tmp_969_16;
  assign __tmp_919_17 = __tmp_969_17;
  assign __tmp_919_18 = __tmp_969_18;
  assign __tmp_919_19 = __tmp_969_19;
  assign __tmp_919_2 = __tmp_947_2;
  assign __tmp_919_3 = __tmp_947_3;
  assign __tmp_919_4 = __tmp_947_4;
  assign __tmp_919_5 = __tmp_947_5;
  assign __tmp_919_6 = __tmp_947_6;
  assign __tmp_919_7 = __tmp_947_7;
  assign __tmp_919_8 = __tmp_947_8;
  assign __tmp_919_9 = __tmp_947_9;
  assign __tmp_921_1 = __tmp_947_1;
  assign __tmp_921_10 = __tmp_959_10;
  assign __tmp_921_11 = __tmp_959_11;
  assign __tmp_921_12 = __tmp_959_12;
  assign __tmp_921_13 = __tmp_969_13;
  assign __tmp_921_14 = __tmp_969_14;
  assign __tmp_921_15 = __tmp_969_15;
  assign __tmp_921_16 = __tmp_969_16;
  assign __tmp_921_17 = __tmp_969_17;
  assign __tmp_921_18 = __tmp_969_18;
  assign __tmp_921_19 = __tmp_969_19;
  assign __tmp_921_2 = __tmp_947_2;
  assign __tmp_921_3 = __tmp_947_3;
  assign __tmp_921_4 = __tmp_947_4;
  assign __tmp_921_5 = __tmp_947_5;
  assign __tmp_921_6 = __tmp_947_6;
  assign __tmp_921_7 = __tmp_947_7;
  assign __tmp_921_8 = __tmp_947_8;
  assign __tmp_921_9 = __tmp_947_9;
  assign __tmp_923_1 = __tmp_947_1;
  assign __tmp_923_10 = __tmp_959_10;
  assign __tmp_923_11 = __tmp_959_11;
  assign __tmp_923_12 = __tmp_959_12;
  assign __tmp_923_13 = __tmp_969_13;
  assign __tmp_923_14 = __tmp_969_14;
  assign __tmp_923_15 = __tmp_969_15;
  assign __tmp_923_16 = __tmp_969_16;
  assign __tmp_923_17 = __tmp_969_17;
  assign __tmp_923_18 = __tmp_969_18;
  assign __tmp_923_19 = __tmp_969_19;
  assign __tmp_923_2 = __tmp_947_2;
  assign __tmp_923_3 = __tmp_947_3;
  assign __tmp_923_4 = __tmp_947_4;
  assign __tmp_923_5 = __tmp_947_5;
  assign __tmp_923_6 = __tmp_947_6;
  assign __tmp_923_7 = __tmp_947_7;
  assign __tmp_923_8 = __tmp_947_8;
  assign __tmp_923_9 = __tmp_947_9;
  assign __tmp_925_1 = __tmp_947_1;
  assign __tmp_925_10 = __tmp_959_10;
  assign __tmp_925_11 = __tmp_959_11;
  assign __tmp_925_12 = __tmp_959_12;
  assign __tmp_925_13 = __tmp_969_13;
  assign __tmp_925_14 = __tmp_969_14;
  assign __tmp_925_15 = __tmp_969_15;
  assign __tmp_925_16 = __tmp_969_16;
  assign __tmp_925_17 = __tmp_969_17;
  assign __tmp_925_18 = __tmp_969_18;
  assign __tmp_925_19 = __tmp_969_19;
  assign __tmp_925_2 = __tmp_947_2;
  assign __tmp_925_3 = __tmp_947_3;
  assign __tmp_925_4 = __tmp_947_4;
  assign __tmp_925_5 = __tmp_947_5;
  assign __tmp_925_6 = __tmp_947_6;
  assign __tmp_925_7 = __tmp_947_7;
  assign __tmp_925_8 = __tmp_947_8;
  assign __tmp_925_9 = __tmp_947_9;
  assign __tmp_927_1 = __tmp_947_1;
  assign __tmp_927_10 = __tmp_959_10;
  assign __tmp_927_11 = __tmp_959_11;
  assign __tmp_927_12 = __tmp_959_12;
  assign __tmp_927_13 = __tmp_969_13;
  assign __tmp_927_14 = __tmp_969_14;
  assign __tmp_927_15 = __tmp_969_15;
  assign __tmp_927_16 = __tmp_969_16;
  assign __tmp_927_17 = __tmp_969_17;
  assign __tmp_927_18 = __tmp_969_18;
  assign __tmp_927_19 = __tmp_969_19;
  assign __tmp_927_2 = __tmp_947_2;
  assign __tmp_927_3 = __tmp_947_3;
  assign __tmp_927_4 = __tmp_947_4;
  assign __tmp_927_5 = __tmp_947_5;
  assign __tmp_927_6 = __tmp_947_6;
  assign __tmp_927_7 = __tmp_947_7;
  assign __tmp_927_8 = __tmp_947_8;
  assign __tmp_927_9 = __tmp_947_9;
  assign __tmp_929_1 = __tmp_947_1;
  assign __tmp_929_2 = __tmp_947_2;
  assign __tmp_929_3 = __tmp_947_3;
  assign __tmp_929_4 = __tmp_947_4;
  assign __tmp_929_5 = __tmp_947_5;
  assign __tmp_929_6 = __tmp_947_6;
  assign __tmp_931_1 = __tmp_947_1;
  assign __tmp_931_2 = __tmp_947_2;
  assign __tmp_931_3 = __tmp_947_3;
  assign __tmp_931_4 = __tmp_947_4;
  assign __tmp_931_5 = __tmp_947_5;
  assign __tmp_931_6 = __tmp_947_6;
  assign __tmp_933_1 = __tmp_947_1;
  assign __tmp_933_2 = __tmp_947_2;
  assign __tmp_933_3 = __tmp_947_3;
  assign __tmp_933_4 = __tmp_947_4;
  assign __tmp_933_5 = __tmp_947_5;
  assign __tmp_933_6 = __tmp_947_6;
  assign __tmp_935_1 = __tmp_947_1;
  assign __tmp_935_10 = __tmp_959_10;
  assign __tmp_935_11 = __tmp_959_11;
  assign __tmp_935_12 = __tmp_959_12;
  assign __tmp_935_13 = __tmp_969_13;
  assign __tmp_935_14 = __tmp_969_14;
  assign __tmp_935_15 = __tmp_969_15;
  assign __tmp_935_16 = __tmp_969_16;
  assign __tmp_935_17 = __tmp_969_17;
  assign __tmp_935_18 = __tmp_969_18;
  assign __tmp_935_19 = __tmp_969_19;
  assign __tmp_935_2 = __tmp_947_2;
  assign __tmp_935_20 = __tmp_969_20;
  assign __tmp_935_21 = __tmp_969_21;
  assign __tmp_935_22 = __tmp_969_22;
  assign __tmp_935_23 = __tmp_969_23;
  assign __tmp_935_24 = __tmp_969_24;
  assign __tmp_935_3 = __tmp_947_3;
  assign __tmp_935_4 = __tmp_947_4;
  assign __tmp_935_5 = __tmp_947_5;
  assign __tmp_935_6 = __tmp_947_6;
  assign __tmp_935_7 = __tmp_947_7;
  assign __tmp_935_8 = __tmp_947_8;
  assign __tmp_935_9 = __tmp_947_9;
  assign __tmp_937_1 = __tmp_947_1;
  assign __tmp_937_10 = __tmp_959_10;
  assign __tmp_937_11 = __tmp_959_11;
  assign __tmp_937_12 = __tmp_959_12;
  assign __tmp_937_13 = __tmp_969_13;
  assign __tmp_937_14 = __tmp_969_14;
  assign __tmp_937_15 = __tmp_969_15;
  assign __tmp_937_16 = __tmp_969_16;
  assign __tmp_937_17 = __tmp_969_17;
  assign __tmp_937_18 = __tmp_969_18;
  assign __tmp_937_19 = __tmp_969_19;
  assign __tmp_937_2 = __tmp_947_2;
  assign __tmp_937_20 = __tmp_969_20;
  assign __tmp_937_21 = __tmp_969_21;
  assign __tmp_937_22 = __tmp_969_22;
  assign __tmp_937_23 = __tmp_969_23;
  assign __tmp_937_3 = __tmp_947_3;
  assign __tmp_937_4 = __tmp_947_4;
  assign __tmp_937_5 = __tmp_947_5;
  assign __tmp_937_6 = __tmp_947_6;
  assign __tmp_937_7 = __tmp_947_7;
  assign __tmp_937_8 = __tmp_947_8;
  assign __tmp_937_9 = __tmp_947_9;
  assign __tmp_939_1 = __tmp_947_1;
  assign __tmp_939_10 = __tmp_959_10;
  assign __tmp_939_11 = __tmp_959_11;
  assign __tmp_939_12 = __tmp_959_12;
  assign __tmp_939_13 = __tmp_969_13;
  assign __tmp_939_14 = __tmp_969_14;
  assign __tmp_939_15 = __tmp_969_15;
  assign __tmp_939_16 = __tmp_969_16;
  assign __tmp_939_17 = __tmp_969_17;
  assign __tmp_939_18 = __tmp_969_18;
  assign __tmp_939_19 = __tmp_969_19;
  assign __tmp_939_2 = __tmp_947_2;
  assign __tmp_939_20 = __tmp_969_20;
  assign __tmp_939_21 = __tmp_969_21;
  assign __tmp_939_22 = __tmp_969_22;
  assign __tmp_939_23 = __tmp_969_23;
  assign __tmp_939_3 = __tmp_947_3;
  assign __tmp_939_4 = __tmp_947_4;
  assign __tmp_939_5 = __tmp_947_5;
  assign __tmp_939_6 = __tmp_947_6;
  assign __tmp_939_7 = __tmp_947_7;
  assign __tmp_939_8 = __tmp_947_8;
  assign __tmp_939_9 = __tmp_947_9;
  assign __tmp_941_1 = __tmp_947_1;
  assign __tmp_941_10 = __tmp_959_10;
  assign __tmp_941_11 = __tmp_959_11;
  assign __tmp_941_12 = __tmp_959_12;
  assign __tmp_941_13 = __tmp_969_13;
  assign __tmp_941_14 = __tmp_969_14;
  assign __tmp_941_15 = __tmp_969_15;
  assign __tmp_941_16 = __tmp_969_16;
  assign __tmp_941_17 = __tmp_969_17;
  assign __tmp_941_18 = __tmp_969_18;
  assign __tmp_941_19 = __tmp_969_19;
  assign __tmp_941_2 = __tmp_947_2;
  assign __tmp_941_20 = __tmp_969_20;
  assign __tmp_941_21 = __tmp_969_21;
  assign __tmp_941_22 = __tmp_969_22;
  assign __tmp_941_23 = __tmp_969_23;
  assign __tmp_941_3 = __tmp_947_3;
  assign __tmp_941_4 = __tmp_947_4;
  assign __tmp_941_5 = __tmp_947_5;
  assign __tmp_941_6 = __tmp_947_6;
  assign __tmp_941_7 = __tmp_947_7;
  assign __tmp_941_8 = __tmp_947_8;
  assign __tmp_941_9 = __tmp_947_9;
  assign __tmp_943_1 = __tmp_947_1;
  assign __tmp_943_2 = __tmp_947_2;
  assign __tmp_943_3 = __tmp_947_3;
  assign __tmp_943_4 = __tmp_947_4;
  assign __tmp_943_5 = __tmp_947_5;
  assign __tmp_943_6 = __tmp_947_6;
  assign __tmp_943_7 = __tmp_947_7;
  assign __tmp_943_8 = __tmp_947_8;
  assign __tmp_943_9 = __tmp_947_9;
  assign __tmp_945_1 = __tmp_947_1;
  assign __tmp_945_2 = __tmp_947_2;
  assign __tmp_945_3 = __tmp_947_3;
  assign __tmp_945_4 = __tmp_947_4;
  assign __tmp_945_5 = __tmp_947_5;
  assign __tmp_945_6 = __tmp_947_6;
  assign __tmp_945_7 = __tmp_947_7;
  assign __tmp_945_8 = __tmp_947_8;
  assign __tmp_945_9 = __tmp_947_9;
  assign __tmp_949_1 = __tmp_947_1;
  assign __tmp_949_10 = __tmp_959_10;
  assign __tmp_949_11 = __tmp_959_11;
  assign __tmp_949_12 = __tmp_959_12;
  assign __tmp_949_13 = __tmp_969_13;
  assign __tmp_949_14 = __tmp_969_14;
  assign __tmp_949_15 = __tmp_969_15;
  assign __tmp_949_16 = __tmp_969_16;
  assign __tmp_949_17 = __tmp_969_17;
  assign __tmp_949_18 = __tmp_969_18;
  assign __tmp_949_19 = __tmp_969_19;
  assign __tmp_949_2 = __tmp_947_2;
  assign __tmp_949_20 = __tmp_969_20;
  assign __tmp_949_21 = __tmp_969_21;
  assign __tmp_949_22 = __tmp_969_22;
  assign __tmp_949_23 = __tmp_969_23;
  assign __tmp_949_24 = __tmp_969_24;
  assign __tmp_949_25 = __tmp_969_25;
  assign __tmp_949_26 = __tmp_969_26;
  assign __tmp_949_27 = __tmp_969_27;
  assign __tmp_949_28 = __tmp_969_28;
  assign __tmp_949_29 = __tmp_969_29;
  assign __tmp_949_3 = __tmp_947_3;
  assign __tmp_949_30 = __tmp_969_30;
  assign __tmp_949_31 = __tmp_969_31;
  assign __tmp_949_4 = __tmp_947_4;
  assign __tmp_949_5 = __tmp_947_5;
  assign __tmp_949_6 = __tmp_947_6;
  assign __tmp_949_7 = __tmp_947_7;
  assign __tmp_949_8 = __tmp_947_8;
  assign __tmp_949_9 = __tmp_947_9;
  assign __tmp_951_1 = __tmp_947_1;
  assign __tmp_951_10 = __tmp_959_10;
  assign __tmp_951_11 = __tmp_959_11;
  assign __tmp_951_12 = __tmp_959_12;
  assign __tmp_951_13 = __tmp_969_13;
  assign __tmp_951_14 = __tmp_969_14;
  assign __tmp_951_15 = __tmp_969_15;
  assign __tmp_951_16 = __tmp_969_16;
  assign __tmp_951_17 = __tmp_969_17;
  assign __tmp_951_18 = __tmp_969_18;
  assign __tmp_951_19 = __tmp_969_19;
  assign __tmp_951_2 = __tmp_947_2;
  assign __tmp_951_20 = __tmp_969_20;
  assign __tmp_951_21 = __tmp_969_21;
  assign __tmp_951_22 = __tmp_969_22;
  assign __tmp_951_23 = __tmp_969_23;
  assign __tmp_951_24 = __tmp_969_24;
  assign __tmp_951_25 = __tmp_969_25;
  assign __tmp_951_26 = __tmp_969_26;
  assign __tmp_951_27 = __tmp_969_27;
  assign __tmp_951_28 = __tmp_969_28;
  assign __tmp_951_29 = __tmp_969_29;
  assign __tmp_951_3 = __tmp_947_3;
  assign __tmp_951_30 = __tmp_969_30;
  assign __tmp_951_31 = __tmp_969_31;
  assign __tmp_951_4 = __tmp_947_4;
  assign __tmp_951_5 = __tmp_947_5;
  assign __tmp_951_6 = __tmp_947_6;
  assign __tmp_951_7 = __tmp_947_7;
  assign __tmp_951_8 = __tmp_947_8;
  assign __tmp_951_9 = __tmp_947_9;
  assign __tmp_953_1 = __tmp_947_1;
  assign __tmp_953_10 = __tmp_959_10;
  assign __tmp_953_11 = __tmp_959_11;
  assign __tmp_953_12 = __tmp_959_12;
  assign __tmp_953_13 = __tmp_969_13;
  assign __tmp_953_14 = __tmp_969_14;
  assign __tmp_953_15 = __tmp_969_15;
  assign __tmp_953_16 = __tmp_969_16;
  assign __tmp_953_17 = __tmp_969_17;
  assign __tmp_953_18 = __tmp_969_18;
  assign __tmp_953_19 = __tmp_969_19;
  assign __tmp_953_2 = __tmp_947_2;
  assign __tmp_953_20 = __tmp_969_20;
  assign __tmp_953_21 = __tmp_969_21;
  assign __tmp_953_22 = __tmp_969_22;
  assign __tmp_953_23 = __tmp_969_23;
  assign __tmp_953_24 = __tmp_969_24;
  assign __tmp_953_25 = __tmp_969_25;
  assign __tmp_953_26 = __tmp_969_26;
  assign __tmp_953_27 = __tmp_969_27;
  assign __tmp_953_28 = __tmp_969_28;
  assign __tmp_953_29 = __tmp_969_29;
  assign __tmp_953_3 = __tmp_947_3;
  assign __tmp_953_30 = __tmp_969_30;
  assign __tmp_953_31 = __tmp_969_31;
  assign __tmp_953_4 = __tmp_947_4;
  assign __tmp_953_5 = __tmp_947_5;
  assign __tmp_953_6 = __tmp_947_6;
  assign __tmp_953_7 = __tmp_947_7;
  assign __tmp_953_8 = __tmp_947_8;
  assign __tmp_953_9 = __tmp_947_9;
  assign __tmp_955_1 = __tmp_947_1;
  assign __tmp_955_10 = __tmp_959_10;
  assign __tmp_955_11 = __tmp_959_11;
  assign __tmp_955_12 = __tmp_959_12;
  assign __tmp_955_2 = __tmp_947_2;
  assign __tmp_955_3 = __tmp_947_3;
  assign __tmp_955_4 = __tmp_947_4;
  assign __tmp_955_5 = __tmp_947_5;
  assign __tmp_955_6 = __tmp_947_6;
  assign __tmp_955_7 = __tmp_947_7;
  assign __tmp_955_8 = __tmp_947_8;
  assign __tmp_955_9 = __tmp_947_9;
  assign __tmp_957_1 = __tmp_947_1;
  assign __tmp_957_10 = __tmp_959_10;
  assign __tmp_957_11 = __tmp_959_11;
  assign __tmp_957_12 = __tmp_959_12;
  assign __tmp_957_2 = __tmp_947_2;
  assign __tmp_957_3 = __tmp_947_3;
  assign __tmp_957_4 = __tmp_947_4;
  assign __tmp_957_5 = __tmp_947_5;
  assign __tmp_957_6 = __tmp_947_6;
  assign __tmp_957_7 = __tmp_947_7;
  assign __tmp_957_8 = __tmp_947_8;
  assign __tmp_957_9 = __tmp_947_9;
  assign __tmp_959_1 = __tmp_947_1;
  assign __tmp_959_2 = __tmp_947_2;
  assign __tmp_959_3 = __tmp_947_3;
  assign __tmp_959_4 = __tmp_947_4;
  assign __tmp_959_5 = __tmp_947_5;
  assign __tmp_959_6 = __tmp_947_6;
  assign __tmp_959_7 = __tmp_947_7;
  assign __tmp_959_8 = __tmp_947_8;
  assign __tmp_959_9 = __tmp_947_9;
  assign __tmp_961_1 = __tmp_947_1;
  assign __tmp_961_10 = __tmp_959_10;
  assign __tmp_961_11 = __tmp_959_11;
  assign __tmp_961_12 = __tmp_959_12;
  assign __tmp_961_13 = __tmp_969_13;
  assign __tmp_961_14 = __tmp_969_14;
  assign __tmp_961_15 = __tmp_969_15;
  assign __tmp_961_16 = __tmp_969_16;
  assign __tmp_961_17 = __tmp_969_17;
  assign __tmp_961_18 = __tmp_969_18;
  assign __tmp_961_19 = __tmp_969_19;
  assign __tmp_961_2 = __tmp_947_2;
  assign __tmp_961_20 = __tmp_969_20;
  assign __tmp_961_21 = __tmp_969_21;
  assign __tmp_961_22 = __tmp_969_22;
  assign __tmp_961_23 = __tmp_969_23;
  assign __tmp_961_24 = __tmp_969_24;
  assign __tmp_961_25 = __tmp_969_25;
  assign __tmp_961_26 = __tmp_969_26;
  assign __tmp_961_27 = __tmp_969_27;
  assign __tmp_961_28 = __tmp_969_28;
  assign __tmp_961_29 = __tmp_969_29;
  assign __tmp_961_3 = __tmp_947_3;
  assign __tmp_961_30 = __tmp_969_30;
  assign __tmp_961_31 = __tmp_969_31;
  assign __tmp_961_32 = __tmp_969_32;
  assign __tmp_961_33 = __tmp_969_33;
  assign __tmp_961_34 = __tmp_969_34;
  assign __tmp_961_35 = __tmp_969_35;
  assign __tmp_961_36 = __tmp_969_36;
  assign __tmp_961_37 = __tmp_969_37;
  assign __tmp_961_38 = __tmp_969_38;
  assign __tmp_961_39 = __tmp_969_39;
  assign __tmp_961_4 = __tmp_947_4;
  assign __tmp_961_40 = __tmp_969_40;
  assign __tmp_961_41 = __tmp_969_41;
  assign __tmp_961_42 = __tmp_969_42;
  assign __tmp_961_43 = __tmp_967_43;
  assign __tmp_961_44 = __tmp_967_44;
  assign __tmp_961_45 = __tmp_967_45;
  assign __tmp_961_46 = __tmp_967_46;
  assign __tmp_961_5 = __tmp_947_5;
  assign __tmp_961_6 = __tmp_947_6;
  assign __tmp_961_7 = __tmp_947_7;
  assign __tmp_961_8 = __tmp_947_8;
  assign __tmp_961_9 = __tmp_947_9;
  assign __tmp_963_1 = __tmp_947_1;
  assign __tmp_963_10 = __tmp_959_10;
  assign __tmp_963_11 = __tmp_959_11;
  assign __tmp_963_12 = __tmp_959_12;
  assign __tmp_963_13 = __tmp_969_13;
  assign __tmp_963_14 = __tmp_969_14;
  assign __tmp_963_15 = __tmp_969_15;
  assign __tmp_963_16 = __tmp_969_16;
  assign __tmp_963_17 = __tmp_969_17;
  assign __tmp_963_18 = __tmp_969_18;
  assign __tmp_963_19 = __tmp_969_19;
  assign __tmp_963_2 = __tmp_947_2;
  assign __tmp_963_20 = __tmp_969_20;
  assign __tmp_963_21 = __tmp_969_21;
  assign __tmp_963_22 = __tmp_969_22;
  assign __tmp_963_23 = __tmp_969_23;
  assign __tmp_963_24 = __tmp_969_24;
  assign __tmp_963_25 = __tmp_969_25;
  assign __tmp_963_26 = __tmp_969_26;
  assign __tmp_963_27 = __tmp_969_27;
  assign __tmp_963_28 = __tmp_969_28;
  assign __tmp_963_29 = __tmp_969_29;
  assign __tmp_963_3 = __tmp_947_3;
  assign __tmp_963_30 = __tmp_969_30;
  assign __tmp_963_31 = __tmp_969_31;
  assign __tmp_963_32 = __tmp_969_32;
  assign __tmp_963_33 = __tmp_969_33;
  assign __tmp_963_34 = __tmp_969_34;
  assign __tmp_963_35 = __tmp_969_35;
  assign __tmp_963_36 = __tmp_969_36;
  assign __tmp_963_37 = __tmp_969_37;
  assign __tmp_963_38 = __tmp_969_38;
  assign __tmp_963_39 = __tmp_969_39;
  assign __tmp_963_4 = __tmp_947_4;
  assign __tmp_963_40 = __tmp_969_40;
  assign __tmp_963_41 = __tmp_969_41;
  assign __tmp_963_42 = __tmp_969_42;
  assign __tmp_963_43 = __tmp_967_43;
  assign __tmp_963_44 = __tmp_967_44;
  assign __tmp_963_45 = __tmp_967_45;
  assign __tmp_963_46 = __tmp_967_46;
  assign __tmp_963_5 = __tmp_947_5;
  assign __tmp_963_6 = __tmp_947_6;
  assign __tmp_963_7 = __tmp_947_7;
  assign __tmp_963_8 = __tmp_947_8;
  assign __tmp_963_9 = __tmp_947_9;
  assign __tmp_965_1 = __tmp_947_1;
  assign __tmp_965_10 = __tmp_959_10;
  assign __tmp_965_11 = __tmp_959_11;
  assign __tmp_965_12 = __tmp_959_12;
  assign __tmp_965_13 = __tmp_969_13;
  assign __tmp_965_14 = __tmp_969_14;
  assign __tmp_965_15 = __tmp_969_15;
  assign __tmp_965_16 = __tmp_969_16;
  assign __tmp_965_17 = __tmp_969_17;
  assign __tmp_965_18 = __tmp_969_18;
  assign __tmp_965_19 = __tmp_969_19;
  assign __tmp_965_2 = __tmp_947_2;
  assign __tmp_965_20 = __tmp_969_20;
  assign __tmp_965_21 = __tmp_969_21;
  assign __tmp_965_22 = __tmp_969_22;
  assign __tmp_965_23 = __tmp_969_23;
  assign __tmp_965_24 = __tmp_969_24;
  assign __tmp_965_25 = __tmp_969_25;
  assign __tmp_965_26 = __tmp_969_26;
  assign __tmp_965_27 = __tmp_969_27;
  assign __tmp_965_28 = __tmp_969_28;
  assign __tmp_965_29 = __tmp_969_29;
  assign __tmp_965_3 = __tmp_947_3;
  assign __tmp_965_30 = __tmp_969_30;
  assign __tmp_965_31 = __tmp_969_31;
  assign __tmp_965_32 = __tmp_969_32;
  assign __tmp_965_33 = __tmp_969_33;
  assign __tmp_965_34 = __tmp_969_34;
  assign __tmp_965_35 = __tmp_969_35;
  assign __tmp_965_36 = __tmp_969_36;
  assign __tmp_965_37 = __tmp_969_37;
  assign __tmp_965_38 = __tmp_969_38;
  assign __tmp_965_39 = __tmp_969_39;
  assign __tmp_965_4 = __tmp_947_4;
  assign __tmp_965_40 = __tmp_969_40;
  assign __tmp_965_41 = __tmp_969_41;
  assign __tmp_965_42 = __tmp_969_42;
  assign __tmp_965_43 = __tmp_967_43;
  assign __tmp_965_44 = __tmp_967_44;
  assign __tmp_965_45 = __tmp_967_45;
  assign __tmp_965_46 = __tmp_967_46;
  assign __tmp_965_5 = __tmp_947_5;
  assign __tmp_965_6 = __tmp_947_6;
  assign __tmp_965_7 = __tmp_947_7;
  assign __tmp_965_8 = __tmp_947_8;
  assign __tmp_965_9 = __tmp_947_9;
  assign __tmp_967_1 = __tmp_947_1;
  assign __tmp_967_10 = __tmp_959_10;
  assign __tmp_967_11 = __tmp_959_11;
  assign __tmp_967_12 = __tmp_959_12;
  assign __tmp_967_13 = __tmp_969_13;
  assign __tmp_967_14 = __tmp_969_14;
  assign __tmp_967_15 = __tmp_969_15;
  assign __tmp_967_16 = __tmp_969_16;
  assign __tmp_967_17 = __tmp_969_17;
  assign __tmp_967_18 = __tmp_969_18;
  assign __tmp_967_19 = __tmp_969_19;
  assign __tmp_967_2 = __tmp_947_2;
  assign __tmp_967_20 = __tmp_969_20;
  assign __tmp_967_21 = __tmp_969_21;
  assign __tmp_967_22 = __tmp_969_22;
  assign __tmp_967_23 = __tmp_969_23;
  assign __tmp_967_24 = __tmp_969_24;
  assign __tmp_967_25 = __tmp_969_25;
  assign __tmp_967_26 = __tmp_969_26;
  assign __tmp_967_27 = __tmp_969_27;
  assign __tmp_967_28 = __tmp_969_28;
  assign __tmp_967_29 = __tmp_969_29;
  assign __tmp_967_3 = __tmp_947_3;
  assign __tmp_967_30 = __tmp_969_30;
  assign __tmp_967_31 = __tmp_969_31;
  assign __tmp_967_32 = __tmp_969_32;
  assign __tmp_967_33 = __tmp_969_33;
  assign __tmp_967_34 = __tmp_969_34;
  assign __tmp_967_35 = __tmp_969_35;
  assign __tmp_967_36 = __tmp_969_36;
  assign __tmp_967_37 = __tmp_969_37;
  assign __tmp_967_38 = __tmp_969_38;
  assign __tmp_967_39 = __tmp_969_39;
  assign __tmp_967_4 = __tmp_947_4;
  assign __tmp_967_40 = __tmp_969_40;
  assign __tmp_967_41 = __tmp_969_41;
  assign __tmp_967_42 = __tmp_969_42;
  assign __tmp_967_5 = __tmp_947_5;
  assign __tmp_967_6 = __tmp_947_6;
  assign __tmp_967_7 = __tmp_947_7;
  assign __tmp_967_8 = __tmp_947_8;
  assign __tmp_967_9 = __tmp_947_9;
  assign __tmp_969_1 = __tmp_947_1;
  assign __tmp_969_10 = __tmp_959_10;
  assign __tmp_969_11 = __tmp_959_11;
  assign __tmp_969_12 = __tmp_959_12;
  assign __tmp_969_2 = __tmp_947_2;
  assign __tmp_969_3 = __tmp_947_3;
  assign __tmp_969_4 = __tmp_947_4;
  assign __tmp_969_5 = __tmp_947_5;
  assign __tmp_969_6 = __tmp_947_6;
  assign __tmp_969_7 = __tmp_947_7;
  assign __tmp_969_8 = __tmp_947_8;
  assign __tmp_969_9 = __tmp_947_9;
  assign _acc_0_fsm = 0;
  assign _acc_0_rshift_idle = 1'h1;
  assign _acc_0_rshift_source_ram_rvalid = 1'h0;
  assign _acc_0_sum_sink_wenable = 1'h0;
  assign _acc_0_valid_sink_wenable = 1'h0;
  assign _acc_0_x_idle = 1'h1;
  assign _acc_0_x_source_ram_rvalid = 1'h0;
  assign _add_tree_1_fsm = 0;
  assign _add_tree_1_sum_sink_wenable = 1'h0;
  assign _add_tree_1_var0_idle = 1'h1;
  assign _add_tree_1_var0_source_ram_rvalid = 1'h0;
  assign _add_tree_2_fsm = 0;
  assign _add_tree_2_sum_sink_wenable = 1'h0;
  assign _add_tree_2_var0_idle = 1'h1;
  assign _add_tree_2_var0_source_ram_rvalid = 1'h0;
  assign _add_tree_2_var1_idle = 1'h1;
  assign _add_tree_2_var1_source_ram_rvalid = 1'h0;
  assign _add_tree_2_var2_idle = 1'h1;
  assign _add_tree_2_var2_source_ram_rvalid = 1'h0;
  assign _add_tree_2_var3_idle = 1'h1;
  assign _add_tree_2_var3_source_ram_rvalid = 1'h0;
  assign _add_tree_2_var4_idle = 1'h1;
  assign _add_tree_2_var4_source_ram_rvalid = 1'h0;
  assign _add_tree_2_var5_idle = 1'h1;
  assign _add_tree_2_var5_source_ram_rvalid = 1'h0;
  assign _add_tree_2_var6_idle = 1'h1;
  assign _add_tree_2_var6_source_ram_rvalid = 1'h0;
  assign _add_tree_2_var7_idle = 1'h1;
  assign _add_tree_2_var7_source_ram_rvalid = 1'h0;
  assign _add_tree_2_var8_idle = 1'h1;
  assign _add_tree_2_var8_source_ram_rvalid = 1'h0;
  assign _cast_data_23 = __variable_wdata_22;
  assign _cast_src_23 = __variable_wdata_22;
  assign _cond_data_775 = _cond_data_890;
  assign _dataflow_cat_odata_107 = _dataflow_cat_data_107;
  assign _dataflow_cat_odata_167 = _dataflow_cat_data_167;
  assign _dataflow_cat_odata_98 = _dataflow_cat_data_98;
  assign _dataflow_cat_ovalid_107 = _dataflow_cat_valid_107;
  assign _dataflow_cat_ovalid_167 = _dataflow_cat_valid_167;
  assign _dataflow_cat_ovalid_98 = _dataflow_cat_valid_98;
  assign _dataflow_slice_odata_111 = _dataflow_slice_data_111;
  assign _dataflow_slice_odata_114 = _dataflow_slice_data_114;
  assign _dataflow_slice_odata_117 = _dataflow_slice_data_117;
  assign _dataflow_slice_odata_12 = _dataflow_slice_data_12;
  assign _dataflow_slice_odata_120 = _dataflow_slice_data_120;
  assign _dataflow_slice_odata_124 = _dataflow_slice_data_124;
  assign _dataflow_slice_odata_127 = _dataflow_slice_data_127;
  assign _dataflow_slice_odata_130 = _dataflow_slice_data_130;
  assign _dataflow_slice_odata_133 = _dataflow_slice_data_133;
  assign _dataflow_slice_odata_136 = _dataflow_slice_data_136;
  assign _dataflow_slice_odata_139 = _dataflow_slice_data_139;
  assign _dataflow_slice_odata_142 = _dataflow_slice_data_142;
  assign _dataflow_slice_odata_145 = _dataflow_slice_data_145;
  assign _dataflow_slice_odata_149 = _dataflow_slice_data_149;
  assign _dataflow_slice_odata_152 = _dataflow_slice_data_152;
  assign _dataflow_slice_odata_155 = _dataflow_slice_data_155;
  assign _dataflow_slice_odata_158 = _dataflow_slice_data_158;
  assign _dataflow_slice_odata_16 = _dataflow_slice_data_16;
  assign _dataflow_slice_odata_19 = _dataflow_slice_data_19;
  assign _dataflow_slice_odata_22 = _dataflow_slice_data_22;
  assign _dataflow_slice_odata_25 = _dataflow_slice_data_25;
  assign _dataflow_slice_odata_29 = _dataflow_slice_data_29;
  assign _dataflow_slice_odata_3 = _dataflow_slice_data_3;
  assign _dataflow_slice_odata_32 = _dataflow_slice_data_32;
  assign _dataflow_slice_odata_35 = _dataflow_slice_data_35;
  assign _dataflow_slice_odata_38 = _dataflow_slice_data_38;
  assign _dataflow_slice_odata_41 = _dataflow_slice_data_41;
  assign _dataflow_slice_odata_44 = _dataflow_slice_data_44;
  assign _dataflow_slice_odata_47 = _dataflow_slice_data_47;
  assign _dataflow_slice_odata_50 = _dataflow_slice_data_50;
  assign _dataflow_slice_odata_54 = _dataflow_slice_data_54;
  assign _dataflow_slice_odata_57 = _dataflow_slice_data_57;
  assign _dataflow_slice_odata_6 = _dataflow_slice_data_6;
  assign _dataflow_slice_odata_60 = _dataflow_slice_data_60;
  assign _dataflow_slice_odata_63 = _dataflow_slice_data_63;
  assign _dataflow_slice_odata_67 = _dataflow_slice_data_67;
  assign _dataflow_slice_odata_70 = _dataflow_slice_data_70;
  assign _dataflow_slice_odata_73 = _dataflow_slice_data_73;
  assign _dataflow_slice_odata_76 = _dataflow_slice_data_76;
  assign _dataflow_slice_odata_80 = _dataflow_slice_data_80;
  assign _dataflow_slice_odata_83 = _dataflow_slice_data_83;
  assign _dataflow_slice_odata_86 = _dataflow_slice_data_86;
  assign _dataflow_slice_odata_89 = _dataflow_slice_data_89;
  assign _dataflow_slice_odata_9 = _dataflow_slice_data_9;
  assign _dataflow_slice_ovalid_111 = _dataflow_slice_valid_111;
  assign _dataflow_slice_ovalid_114 = _dataflow_slice_valid_114;
  assign _dataflow_slice_ovalid_117 = _dataflow_slice_valid_117;
  assign _dataflow_slice_ovalid_12 = _dataflow_slice_valid_12;
  assign _dataflow_slice_ovalid_120 = _dataflow_slice_valid_120;
  assign _dataflow_slice_ovalid_124 = _dataflow_slice_valid_124;
  assign _dataflow_slice_ovalid_127 = _dataflow_slice_valid_127;
  assign _dataflow_slice_ovalid_130 = _dataflow_slice_valid_130;
  assign _dataflow_slice_ovalid_133 = _dataflow_slice_valid_133;
  assign _dataflow_slice_ovalid_136 = _dataflow_slice_valid_136;
  assign _dataflow_slice_ovalid_139 = _dataflow_slice_valid_139;
  assign _dataflow_slice_ovalid_142 = _dataflow_slice_valid_142;
  assign _dataflow_slice_ovalid_145 = _dataflow_slice_valid_145;
  assign _dataflow_slice_ovalid_149 = _dataflow_slice_valid_149;
  assign _dataflow_slice_ovalid_152 = _dataflow_slice_valid_152;
  assign _dataflow_slice_ovalid_155 = _dataflow_slice_valid_155;
  assign _dataflow_slice_ovalid_158 = _dataflow_slice_valid_158;
  assign _dataflow_slice_ovalid_16 = _dataflow_slice_valid_16;
  assign _dataflow_slice_ovalid_19 = _dataflow_slice_valid_19;
  assign _dataflow_slice_ovalid_22 = _dataflow_slice_valid_22;
  assign _dataflow_slice_ovalid_25 = _dataflow_slice_valid_25;
  assign _dataflow_slice_ovalid_29 = _dataflow_slice_valid_29;
  assign _dataflow_slice_ovalid_3 = _dataflow_slice_valid_3;
  assign _dataflow_slice_ovalid_32 = _dataflow_slice_valid_32;
  assign _dataflow_slice_ovalid_35 = _dataflow_slice_valid_35;
  assign _dataflow_slice_ovalid_38 = _dataflow_slice_valid_38;
  assign _dataflow_slice_ovalid_41 = _dataflow_slice_valid_41;
  assign _dataflow_slice_ovalid_44 = _dataflow_slice_valid_44;
  assign _dataflow_slice_ovalid_47 = _dataflow_slice_valid_47;
  assign _dataflow_slice_ovalid_50 = _dataflow_slice_valid_50;
  assign _dataflow_slice_ovalid_54 = _dataflow_slice_valid_54;
  assign _dataflow_slice_ovalid_57 = _dataflow_slice_valid_57;
  assign _dataflow_slice_ovalid_6 = _dataflow_slice_valid_6;
  assign _dataflow_slice_ovalid_60 = _dataflow_slice_valid_60;
  assign _dataflow_slice_ovalid_63 = _dataflow_slice_valid_63;
  assign _dataflow_slice_ovalid_67 = _dataflow_slice_valid_67;
  assign _dataflow_slice_ovalid_70 = _dataflow_slice_valid_70;
  assign _dataflow_slice_ovalid_73 = _dataflow_slice_valid_73;
  assign _dataflow_slice_ovalid_76 = _dataflow_slice_valid_76;
  assign _dataflow_slice_ovalid_80 = _dataflow_slice_valid_80;
  assign _dataflow_slice_ovalid_83 = _dataflow_slice_valid_83;
  assign _dataflow_slice_ovalid_86 = _dataflow_slice_valid_86;
  assign _dataflow_slice_ovalid_89 = _dataflow_slice_valid_89;
  assign _dataflow_slice_ovalid_9 = _dataflow_slice_valid_9;
  assign _eq_data_277 = _eq_data_357;
  assign _eq_data_281 = _eq_data_361;
  assign _eq_data_284 = _eq_data_364;
  assign _eq_data_287 = _eq_data_357;
  assign _eq_data_291 = _eq_data_361;
  assign _eq_data_294 = _eq_data_364;
  assign _eq_data_297 = _eq_data_357;
  assign _eq_data_301 = _eq_data_361;
  assign _eq_data_304 = _eq_data_364;
  assign _eq_data_307 = _eq_data_357;
  assign _eq_data_311 = _eq_data_361;
  assign _eq_data_314 = _eq_data_364;
  assign _eq_data_317 = _eq_data_357;
  assign _eq_data_321 = _eq_data_361;
  assign _eq_data_324 = _eq_data_364;
  assign _eq_data_327 = _eq_data_357;
  assign _eq_data_331 = _eq_data_361;
  assign _eq_data_334 = _eq_data_364;
  assign _eq_data_337 = _eq_data_357;
  assign _eq_data_341 = _eq_data_361;
  assign _eq_data_344 = _eq_data_364;
  assign _eq_data_347 = _eq_data_357;
  assign _eq_data_351 = _eq_data_361;
  assign _eq_data_354 = _eq_data_364;
  assign _eq_data_367 = _eq_data_447;
  assign _eq_data_371 = _eq_data_451;
  assign _eq_data_374 = _eq_data_454;
  assign _eq_data_377 = _eq_data_447;
  assign _eq_data_381 = _eq_data_451;
  assign _eq_data_384 = _eq_data_454;
  assign _eq_data_387 = _eq_data_447;
  assign _eq_data_391 = _eq_data_451;
  assign _eq_data_394 = _eq_data_454;
  assign _eq_data_397 = _eq_data_447;
  assign _eq_data_401 = _eq_data_451;
  assign _eq_data_404 = _eq_data_454;
  assign _eq_data_407 = _eq_data_447;
  assign _eq_data_411 = _eq_data_451;
  assign _eq_data_414 = _eq_data_454;
  assign _eq_data_417 = _eq_data_447;
  assign _eq_data_421 = _eq_data_451;
  assign _eq_data_424 = _eq_data_454;
  assign _eq_data_427 = _eq_data_447;
  assign _eq_data_431 = _eq_data_451;
  assign _eq_data_434 = _eq_data_454;
  assign _eq_data_437 = _eq_data_447;
  assign _eq_data_441 = _eq_data_451;
  assign _eq_data_444 = _eq_data_454;
  assign _greaterthan_data_773 = _greaterthan_data_888;
  assign _maxi_cond_0_1 = _saxi_cond_0_1;
  assign _maxi_cond_1_1 = _saxi_cond_0_1;
  assign _maxi_cond_2_1 = _saxi_cond_0_1;
  assign _maxi_cond_3_1 = _saxi_cond_0_1;
  assign _maxi_cond_4_1 = _saxi_cond_0_1;
  assign _mul_10_fsm = 0;
  assign _mul_10_rshift_idle = 1'h1;
  assign _mul_10_rshift_source_ram_rvalid = 1'h0;
  assign _mul_10_x_idle = 1'h1;
  assign _mul_10_x_source_ram_rvalid = 1'h0;
  assign _mul_10_y_idle = 1'h1;
  assign _mul_10_y_source_ram_rvalid = 1'h0;
  assign _mul_10_z_sink_wenable = 1'h0;
  assign _mul_11_fsm = 0;
  assign _mul_11_rshift_idle = 1'h1;
  assign _mul_11_rshift_source_ram_rvalid = 1'h0;
  assign _mul_11_x_idle = 1'h1;
  assign _mul_11_x_source_ram_rvalid = 1'h0;
  assign _mul_11_y_idle = 1'h1;
  assign _mul_11_y_source_ram_rvalid = 1'h0;
  assign _mul_11_z_sink_wenable = 1'h0;
  assign _mul_12_fsm = 0;
  assign _mul_12_rshift_idle = 1'h1;
  assign _mul_12_rshift_source_ram_rvalid = 1'h0;
  assign _mul_12_x_idle = 1'h1;
  assign _mul_12_x_source_ram_rvalid = 1'h0;
  assign _mul_12_y_idle = 1'h1;
  assign _mul_12_y_source_ram_rvalid = 1'h0;
  assign _mul_12_z_sink_wenable = 1'h0;
  assign _mul_4_fsm = 0;
  assign _mul_4_rshift_idle = 1'h1;
  assign _mul_4_rshift_source_ram_rvalid = 1'h0;
  assign _mul_4_x_idle = 1'h1;
  assign _mul_4_x_source_ram_rvalid = 1'h0;
  assign _mul_4_y_idle = 1'h1;
  assign _mul_4_y_source_ram_rvalid = 1'h0;
  assign _mul_4_z_sink_wenable = 1'h0;
  assign _mul_5_fsm = 0;
  assign _mul_5_rshift_idle = 1'h1;
  assign _mul_5_rshift_source_ram_rvalid = 1'h0;
  assign _mul_5_x_idle = 1'h1;
  assign _mul_5_x_source_ram_rvalid = 1'h0;
  assign _mul_5_y_idle = 1'h1;
  assign _mul_5_y_source_ram_rvalid = 1'h0;
  assign _mul_5_z_sink_wenable = 1'h0;
  assign _mul_6_fsm = 0;
  assign _mul_6_rshift_idle = 1'h1;
  assign _mul_6_rshift_source_ram_rvalid = 1'h0;
  assign _mul_6_x_idle = 1'h1;
  assign _mul_6_x_source_ram_rvalid = 1'h0;
  assign _mul_6_y_idle = 1'h1;
  assign _mul_6_y_source_ram_rvalid = 1'h0;
  assign _mul_6_z_sink_wenable = 1'h0;
  assign _mul_7_fsm = 0;
  assign _mul_7_rshift_idle = 1'h1;
  assign _mul_7_rshift_source_ram_rvalid = 1'h0;
  assign _mul_7_x_idle = 1'h1;
  assign _mul_7_x_source_ram_rvalid = 1'h0;
  assign _mul_7_y_idle = 1'h1;
  assign _mul_7_y_source_ram_rvalid = 1'h0;
  assign _mul_7_z_sink_wenable = 1'h0;
  assign _mul_8_fsm = 0;
  assign _mul_8_rshift_idle = 1'h1;
  assign _mul_8_rshift_source_ram_rvalid = 1'h0;
  assign _mul_8_x_idle = 1'h1;
  assign _mul_8_x_source_ram_rvalid = 1'h0;
  assign _mul_8_y_idle = 1'h1;
  assign _mul_8_y_source_ram_rvalid = 1'h0;
  assign _mul_8_z_sink_wenable = 1'h0;
  assign _mul_9_fsm = 0;
  assign _mul_9_rshift_idle = 1'h1;
  assign _mul_9_rshift_source_ram_rvalid = 1'h0;
  assign _mul_9_x_idle = 1'h1;
  assign _mul_9_x_source_ram_rvalid = 1'h0;
  assign _mul_9_y_idle = 1'h1;
  assign _mul_9_y_source_ram_rvalid = 1'h0;
  assign _mul_9_z_sink_wenable = 1'h0;
  assign _mul_rshift_clip_3_fsm = 0;
  assign _mul_rshift_clip_3_rshift_idle = 1'h1;
  assign _mul_rshift_clip_3_rshift_source_ram_rvalid = 1'h0;
  assign _mul_rshift_clip_3_x_idle = 1'h1;
  assign _mul_rshift_clip_3_x_source_ram_rvalid = 1'h0;
  assign _mul_rshift_clip_3_y_idle = 1'h1;
  assign _mul_rshift_clip_3_y_source_ram_rvalid = 1'h0;
  assign _mul_rshift_clip_3_z_sink_wenable = 1'h0;
  assign _plus_data_607 = _plus_data_743;
  assign _plus_data_624 = _plus_data_743;
  assign _plus_data_641 = _plus_data_743;
  assign _plus_data_658 = _plus_data_743;
  assign _plus_data_675 = _plus_data_743;
  assign _plus_data_692 = _plus_data_743;
  assign _plus_data_709 = _plus_data_743;
  assign _plus_data_726 = _plus_data_743;
  assign _pointer_data_556 = __variable_wdata_217[0];
  assign _pointer_data_558 = __variable_wdata_217[1];
  assign _pointer_data_560 = __variable_wdata_217[2];
  assign _pointer_data_562 = __variable_wdata_217[3];
  assign _pointer_data_564 = __variable_wdata_217[4];
  assign _pointer_data_566 = __variable_wdata_217[5];
  assign _pointer_data_568 = __variable_wdata_217[6];
  assign _pointer_data_570 = __variable_wdata_217[7];
  assign _pointer_data_572 = __variable_wdata_217[8];
  assign _pointer_data_870 = __variable_wdata_799;
  assign _ram_w4_l8192_id0_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_0_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_0_cond_2_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_0_cond_3_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_0_cond_4_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_0_cond_5_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_0_cond_6_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_1_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_1_cond_2_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_1_cond_3_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_1_cond_4_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_1_cond_5_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_1_cond_6_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_2_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_2_cond_2_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_2_cond_3_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_2_cond_4_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_2_cond_5_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_2_cond_6_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_3_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_3_cond_2_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_3_cond_3_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_3_cond_4_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_3_cond_5_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_3_cond_6_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_4_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_4_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_4_cond_2_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_4_cond_3_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_4_cond_4_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_4_cond_5_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_4_cond_6_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_5_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_5_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_5_cond_2_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_5_cond_3_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_5_cond_4_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_5_cond_5_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_5_cond_6_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_6_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_6_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_6_cond_2_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_6_cond_3_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_6_cond_4_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_6_cond_5_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_6_cond_6_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_7_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_7_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_7_cond_3_1 = _ram_w4_l8192_id0_7_cond_2_1;
  assign _ram_w4_l8192_id0_7_cond_4_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id0_7_cond_5_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id0_7_cond_6_1 = __tmp_1223_1;
  assign _ram_w4_l8192_id1_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id1_0_cond_1_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_0_cond_2_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id1_1_cond_1_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_1_cond_2_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id1_2_cond_1_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_2_cond_2_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id1_3_cond_1_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_3_cond_2_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_4_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id1_4_cond_1_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_4_cond_2_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_5_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id1_5_cond_1_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_5_cond_2_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_6_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id1_6_cond_1_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_6_cond_2_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id1_7_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id1_7_cond_2_1 = _ram_w4_l8192_id1_7_cond_1_1;
  assign _ram_w4_l8192_id2_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id2_0_cond_1_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_0_cond_2_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id2_1_cond_1_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_1_cond_2_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id2_2_cond_1_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_2_cond_2_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id2_3_cond_1_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_3_cond_2_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_4_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id2_4_cond_1_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_4_cond_2_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_5_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id2_5_cond_1_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_5_cond_2_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_6_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id2_6_cond_1_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_6_cond_2_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id2_7_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id2_7_cond_2_1 = _ram_w4_l8192_id2_7_cond_1_1;
  assign _ram_w4_l8192_id3_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id3_0_cond_1_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_0_cond_2_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id3_1_cond_1_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_1_cond_2_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id3_2_cond_1_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_2_cond_2_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id3_3_cond_1_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_3_cond_2_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_4_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id3_4_cond_1_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_4_cond_2_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_5_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id3_5_cond_1_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_5_cond_2_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_6_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id3_6_cond_1_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_6_cond_2_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id3_7_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id3_7_cond_2_1 = _ram_w4_l8192_id3_7_cond_1_1;
  assign _ram_w4_l8192_id4_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id4_0_cond_1_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_0_cond_2_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id4_1_cond_1_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_1_cond_2_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id4_2_cond_1_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_2_cond_2_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id4_3_cond_1_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_3_cond_2_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_4_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id4_4_cond_1_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_4_cond_2_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_5_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id4_5_cond_1_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_5_cond_2_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_6_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id4_6_cond_1_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_6_cond_2_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id4_7_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id4_7_cond_2_1 = _ram_w4_l8192_id4_7_cond_1_1;
  assign _ram_w4_l8192_id5_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id5_0_cond_1_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_0_cond_2_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id5_1_cond_1_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_1_cond_2_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id5_2_cond_1_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_2_cond_2_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id5_3_cond_1_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_3_cond_2_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_4_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id5_4_cond_1_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_4_cond_2_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_5_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id5_5_cond_1_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_5_cond_2_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_6_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id5_6_cond_1_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_6_cond_2_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id5_7_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id5_7_cond_1_1 = _ram_w4_l8192_id5_7_cond_2_1;
  assign _ram_w4_l8192_id6_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id6_0_cond_1_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_0_cond_2_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id6_1_cond_1_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_1_cond_2_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id6_2_cond_2_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id6_3_cond_1_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_3_cond_2_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_4_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id6_4_cond_1_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_4_cond_2_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_5_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id6_5_cond_1_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_5_cond_2_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_6_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id6_6_cond_1_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_6_cond_2_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_7_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id6_7_cond_1_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id6_7_cond_2_1 = _ram_w4_l8192_id6_2_cond_1_1;
  assign _ram_w4_l8192_id7_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id7_0_cond_1_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_0_cond_2_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id7_1_cond_1_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_1_cond_2_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id7_2_cond_1_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_2_cond_2_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id7_3_cond_1_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_3_cond_2_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_4_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id7_4_cond_1_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_4_cond_2_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_5_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id7_5_cond_1_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_5_cond_2_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_6_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id7_6_cond_1_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_6_cond_2_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id7_7_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id7_7_cond_2_1 = _ram_w4_l8192_id7_7_cond_1_1;
  assign _ram_w4_l8192_id8_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id8_0_cond_2_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id8_1_cond_1_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_1_cond_2_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id8_2_cond_1_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_2_cond_2_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id8_3_cond_1_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_3_cond_2_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_4_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id8_4_cond_1_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_4_cond_2_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_5_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id8_5_cond_1_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_5_cond_2_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_6_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id8_6_cond_1_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_6_cond_2_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_7_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w4_l8192_id8_7_cond_1_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w4_l8192_id8_7_cond_2_1 = _ram_w4_l8192_id8_0_cond_1_1;
  assign _ram_w8_l2048_id0_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id0_0_cond_1_1 = _ram_w8_l2048_id0_3_cond_2_1;
  assign _ram_w8_l2048_id0_0_cond_2_1 = _ram_w8_l2048_id0_3_cond_2_1;
  assign _ram_w8_l2048_id0_0_cond_4_1 = _ram_w8_l2048_id0_3_cond_5_1;
  assign _ram_w8_l2048_id0_0_cond_5_1 = _ram_w8_l2048_id0_3_cond_5_1;
  assign _ram_w8_l2048_id0_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id0_1_cond_1_1 = _ram_w8_l2048_id0_3_cond_2_1;
  assign _ram_w8_l2048_id0_1_cond_2_1 = _ram_w8_l2048_id0_3_cond_2_1;
  assign _ram_w8_l2048_id0_1_cond_4_1 = _ram_w8_l2048_id0_3_cond_5_1;
  assign _ram_w8_l2048_id0_1_cond_5_1 = _ram_w8_l2048_id0_3_cond_5_1;
  assign _ram_w8_l2048_id0_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id0_2_cond_1_1 = _ram_w8_l2048_id0_3_cond_2_1;
  assign _ram_w8_l2048_id0_2_cond_2_1 = _ram_w8_l2048_id0_3_cond_2_1;
  assign _ram_w8_l2048_id0_2_cond_4_1 = _ram_w8_l2048_id0_3_cond_5_1;
  assign _ram_w8_l2048_id0_2_cond_5_1 = _ram_w8_l2048_id0_3_cond_5_1;
  assign _ram_w8_l2048_id0_3_cond_1_1 = _ram_w8_l2048_id0_3_cond_2_1;
  assign _ram_w8_l2048_id0_3_cond_4_1 = _ram_w8_l2048_id0_3_cond_5_1;
  assign _ram_w8_l2048_id10_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id10_0_cond_1_1 = _ram_w8_l2048_id10_0_cond_2_1;
  assign _ram_w8_l2048_id10_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id10_1_cond_1_1 = _ram_w8_l2048_id10_0_cond_2_1;
  assign _ram_w8_l2048_id10_1_cond_2_1 = _ram_w8_l2048_id10_0_cond_2_1;
  assign _ram_w8_l2048_id10_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id10_2_cond_1_1 = _ram_w8_l2048_id10_0_cond_2_1;
  assign _ram_w8_l2048_id10_2_cond_2_1 = _ram_w8_l2048_id10_0_cond_2_1;
  assign _ram_w8_l2048_id10_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id10_3_cond_1_1 = _ram_w8_l2048_id10_0_cond_2_1;
  assign _ram_w8_l2048_id10_3_cond_2_1 = _ram_w8_l2048_id10_0_cond_2_1;
  assign _ram_w8_l2048_id1_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id1_0_cond_1_1 = _ram_w8_l2048_id1_0_cond_2_1;
  assign _ram_w8_l2048_id1_0_cond_3_1 = _ram_w8_l2048_id1_0_cond_4_1;
  assign _ram_w8_l2048_id1_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id1_1_cond_1_1 = _ram_w8_l2048_id1_0_cond_2_1;
  assign _ram_w8_l2048_id1_1_cond_2_1 = _ram_w8_l2048_id1_0_cond_2_1;
  assign _ram_w8_l2048_id1_1_cond_3_1 = _ram_w8_l2048_id1_0_cond_4_1;
  assign _ram_w8_l2048_id1_1_cond_4_1 = _ram_w8_l2048_id1_0_cond_4_1;
  assign _ram_w8_l2048_id1_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id1_2_cond_1_1 = _ram_w8_l2048_id1_0_cond_2_1;
  assign _ram_w8_l2048_id1_2_cond_2_1 = _ram_w8_l2048_id1_0_cond_2_1;
  assign _ram_w8_l2048_id1_2_cond_3_1 = _ram_w8_l2048_id1_0_cond_4_1;
  assign _ram_w8_l2048_id1_2_cond_4_1 = _ram_w8_l2048_id1_0_cond_4_1;
  assign _ram_w8_l2048_id1_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id1_3_cond_1_1 = _ram_w8_l2048_id1_0_cond_2_1;
  assign _ram_w8_l2048_id1_3_cond_2_1 = _ram_w8_l2048_id1_0_cond_2_1;
  assign _ram_w8_l2048_id1_3_cond_3_1 = _ram_w8_l2048_id1_0_cond_4_1;
  assign _ram_w8_l2048_id1_3_cond_4_1 = _ram_w8_l2048_id1_0_cond_4_1;
  assign _ram_w8_l2048_id2_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id2_0_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id2_0_cond_2_1 = _ram_w8_l2048_id2_0_cond_3_1;
  assign _ram_w8_l2048_id2_0_cond_4_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id2_0_cond_5_1 = _ram_w8_l2048_id2_0_cond_6_1;
  assign _ram_w8_l2048_id2_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id2_1_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id2_1_cond_2_1 = _ram_w8_l2048_id2_0_cond_3_1;
  assign _ram_w8_l2048_id2_1_cond_3_1 = _ram_w8_l2048_id2_0_cond_3_1;
  assign _ram_w8_l2048_id2_1_cond_4_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id2_1_cond_5_1 = _ram_w8_l2048_id2_0_cond_6_1;
  assign _ram_w8_l2048_id2_1_cond_6_1 = _ram_w8_l2048_id2_0_cond_6_1;
  assign _ram_w8_l2048_id2_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id2_2_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id2_2_cond_2_1 = _ram_w8_l2048_id2_0_cond_3_1;
  assign _ram_w8_l2048_id2_2_cond_3_1 = _ram_w8_l2048_id2_0_cond_3_1;
  assign _ram_w8_l2048_id2_2_cond_4_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id2_2_cond_5_1 = _ram_w8_l2048_id2_0_cond_6_1;
  assign _ram_w8_l2048_id2_2_cond_6_1 = _ram_w8_l2048_id2_0_cond_6_1;
  assign _ram_w8_l2048_id2_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id2_3_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id2_3_cond_2_1 = _ram_w8_l2048_id2_0_cond_3_1;
  assign _ram_w8_l2048_id2_3_cond_3_1 = _ram_w8_l2048_id2_0_cond_3_1;
  assign _ram_w8_l2048_id2_3_cond_4_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id2_3_cond_5_1 = _ram_w8_l2048_id2_0_cond_6_1;
  assign _ram_w8_l2048_id2_3_cond_6_1 = _ram_w8_l2048_id2_0_cond_6_1;
  assign _ram_w8_l2048_id3_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id3_0_cond_1_1 = _ram_w8_l2048_id3_0_cond_2_1;
  assign _ram_w8_l2048_id3_0_cond_3_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id3_0_cond_4_1 = _ram_w8_l2048_id3_0_cond_5_1;
  assign _ram_w8_l2048_id3_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id3_1_cond_1_1 = _ram_w8_l2048_id3_0_cond_2_1;
  assign _ram_w8_l2048_id3_1_cond_2_1 = _ram_w8_l2048_id3_0_cond_2_1;
  assign _ram_w8_l2048_id3_1_cond_3_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id3_1_cond_4_1 = _ram_w8_l2048_id3_0_cond_5_1;
  assign _ram_w8_l2048_id3_1_cond_5_1 = _ram_w8_l2048_id3_0_cond_5_1;
  assign _ram_w8_l2048_id3_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id3_2_cond_1_1 = _ram_w8_l2048_id3_0_cond_2_1;
  assign _ram_w8_l2048_id3_2_cond_2_1 = _ram_w8_l2048_id3_0_cond_2_1;
  assign _ram_w8_l2048_id3_2_cond_3_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id3_2_cond_4_1 = _ram_w8_l2048_id3_0_cond_5_1;
  assign _ram_w8_l2048_id3_2_cond_5_1 = _ram_w8_l2048_id3_0_cond_5_1;
  assign _ram_w8_l2048_id3_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id3_3_cond_1_1 = _ram_w8_l2048_id3_0_cond_2_1;
  assign _ram_w8_l2048_id3_3_cond_2_1 = _ram_w8_l2048_id3_0_cond_2_1;
  assign _ram_w8_l2048_id3_3_cond_3_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id3_3_cond_4_1 = _ram_w8_l2048_id3_0_cond_5_1;
  assign _ram_w8_l2048_id3_3_cond_5_1 = _ram_w8_l2048_id3_0_cond_5_1;
  assign _ram_w8_l2048_id4_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id4_0_cond_1_1 = _ram_w8_l2048_id4_0_cond_2_1;
  assign _ram_w8_l2048_id4_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id4_1_cond_1_1 = _ram_w8_l2048_id4_0_cond_2_1;
  assign _ram_w8_l2048_id4_1_cond_2_1 = _ram_w8_l2048_id4_0_cond_2_1;
  assign _ram_w8_l2048_id4_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id4_2_cond_1_1 = _ram_w8_l2048_id4_0_cond_2_1;
  assign _ram_w8_l2048_id4_2_cond_2_1 = _ram_w8_l2048_id4_0_cond_2_1;
  assign _ram_w8_l2048_id4_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id4_3_cond_1_1 = _ram_w8_l2048_id4_0_cond_2_1;
  assign _ram_w8_l2048_id4_3_cond_2_1 = _ram_w8_l2048_id4_0_cond_2_1;
  assign _ram_w8_l2048_id5_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id5_0_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id5_0_cond_2_1 = _ram_w8_l2048_id5_0_cond_3_1;
  assign _ram_w8_l2048_id5_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id5_1_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id5_1_cond_2_1 = _ram_w8_l2048_id5_0_cond_3_1;
  assign _ram_w8_l2048_id5_1_cond_3_1 = _ram_w8_l2048_id5_0_cond_3_1;
  assign _ram_w8_l2048_id5_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id5_2_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id5_2_cond_2_1 = _ram_w8_l2048_id5_0_cond_3_1;
  assign _ram_w8_l2048_id5_2_cond_3_1 = _ram_w8_l2048_id5_0_cond_3_1;
  assign _ram_w8_l2048_id5_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id5_3_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id5_3_cond_2_1 = _ram_w8_l2048_id5_0_cond_3_1;
  assign _ram_w8_l2048_id5_3_cond_3_1 = _ram_w8_l2048_id5_0_cond_3_1;
  assign _ram_w8_l2048_id6_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id6_0_cond_1_1 = _ram_w8_l2048_id6_0_cond_2_1;
  assign _ram_w8_l2048_id6_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id6_1_cond_1_1 = _ram_w8_l2048_id6_0_cond_2_1;
  assign _ram_w8_l2048_id6_1_cond_2_1 = _ram_w8_l2048_id6_0_cond_2_1;
  assign _ram_w8_l2048_id6_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id6_2_cond_1_1 = _ram_w8_l2048_id6_0_cond_2_1;
  assign _ram_w8_l2048_id6_2_cond_2_1 = _ram_w8_l2048_id6_0_cond_2_1;
  assign _ram_w8_l2048_id6_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id6_3_cond_1_1 = _ram_w8_l2048_id6_0_cond_2_1;
  assign _ram_w8_l2048_id6_3_cond_2_1 = _ram_w8_l2048_id6_0_cond_2_1;
  assign _ram_w8_l2048_id7_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id7_0_cond_1_1 = _ram_w8_l2048_id7_0_cond_2_1;
  assign _ram_w8_l2048_id7_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id7_1_cond_1_1 = _ram_w8_l2048_id7_0_cond_2_1;
  assign _ram_w8_l2048_id7_1_cond_2_1 = _ram_w8_l2048_id7_0_cond_2_1;
  assign _ram_w8_l2048_id7_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id7_2_cond_1_1 = _ram_w8_l2048_id7_0_cond_2_1;
  assign _ram_w8_l2048_id7_2_cond_2_1 = _ram_w8_l2048_id7_0_cond_2_1;
  assign _ram_w8_l2048_id7_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id7_3_cond_1_1 = _ram_w8_l2048_id7_0_cond_2_1;
  assign _ram_w8_l2048_id7_3_cond_2_1 = _ram_w8_l2048_id7_0_cond_2_1;
  assign _ram_w8_l2048_id8_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id8_0_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id8_0_cond_2_1 = _ram_w8_l2048_id8_0_cond_3_1;
  assign _ram_w8_l2048_id8_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id8_1_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id8_1_cond_2_1 = _ram_w8_l2048_id8_0_cond_3_1;
  assign _ram_w8_l2048_id8_1_cond_3_1 = _ram_w8_l2048_id8_0_cond_3_1;
  assign _ram_w8_l2048_id8_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id8_2_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id8_2_cond_2_1 = _ram_w8_l2048_id8_0_cond_3_1;
  assign _ram_w8_l2048_id8_2_cond_3_1 = _ram_w8_l2048_id8_0_cond_3_1;
  assign _ram_w8_l2048_id8_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id8_3_cond_1_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id8_3_cond_2_1 = _ram_w8_l2048_id8_0_cond_3_1;
  assign _ram_w8_l2048_id8_3_cond_3_1 = _ram_w8_l2048_id8_0_cond_3_1;
  assign _ram_w8_l2048_id9_0_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id9_0_cond_1_1 = _ram_w8_l2048_id9_0_cond_2_1;
  assign _ram_w8_l2048_id9_1_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id9_1_cond_1_1 = _ram_w8_l2048_id9_0_cond_2_1;
  assign _ram_w8_l2048_id9_1_cond_2_1 = _ram_w8_l2048_id9_0_cond_2_1;
  assign _ram_w8_l2048_id9_2_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id9_2_cond_1_1 = _ram_w8_l2048_id9_0_cond_2_1;
  assign _ram_w8_l2048_id9_2_cond_2_1 = _ram_w8_l2048_id9_0_cond_2_1;
  assign _ram_w8_l2048_id9_3_cond_0_1 = _ram_w8_l2048_id0_3_cond_0_1;
  assign _ram_w8_l2048_id9_3_cond_1_1 = _ram_w8_l2048_id9_0_cond_2_1;
  assign _ram_w8_l2048_id9_3_cond_2_1 = _ram_w8_l2048_id9_0_cond_2_1;
  assign _reduce_max_13_data_data = _reducemax_data_211;
  assign _reduce_max_13_size_data = __variable_wdata_208;
  assign _reduce_max_13_valid_data = _pulse_data_213;
  assign _reduce_max_13_x_data = __variable_wdata_207;
  assign _reinterpretcast_data_234 = __variable_wdata_230;
  assign _reinterpretcast_data_241 = __variable_wdata_237;
  assign _reinterpretcast_data_248 = __variable_wdata_244;
  assign _reinterpretcast_data_255 = __variable_wdata_251;
  assign _reinterpretcast_data_262 = __variable_wdata_258;
  assign _reinterpretcast_data_493 = _cond_data_376;
  assign _reinterpretcast_data_494 = _cond_data_406;
  assign _reinterpretcast_data_495 = _cond_data_436;
  assign _reinterpretcast_data_496 = _cond_data_386;
  assign _reinterpretcast_data_497 = _cond_data_416;
  assign _reinterpretcast_data_498 = _cond_data_446;
  assign _reinterpretcast_data_499 = _cond_data_396;
  assign _reinterpretcast_data_500 = _cond_data_426;
  assign _reinterpretcast_data_501 = _cond_data_456;
  assign _reinterpretcast_data_547 = __variable_wdata_502;
  assign _reinterpretcast_data_548 = __variable_wdata_503;
  assign _reinterpretcast_data_549 = __variable_wdata_504;
  assign _reinterpretcast_data_550 = __variable_wdata_505;
  assign _reinterpretcast_data_551 = __variable_wdata_506;
  assign _reinterpretcast_data_552 = __variable_wdata_507;
  assign _reinterpretcast_data_553 = __variable_wdata_508;
  assign _reinterpretcast_data_554 = __variable_wdata_509;
  assign _reinterpretcast_data_555 = __variable_wdata_510;
  assign _reinterpretcast_data_776 = _cond_data_890;
  assign _reinterpretcast_data_789 = __variable_wdata_778;
  assign _reinterpretcast_data_795 = __substreamoutput_data_793;
  assign _reinterpretcast_data_816 = __variable_wdata_812;
  assign _reinterpretcast_data_823 = __variable_wdata_819;
  assign _reinterpretcast_data_830 = __variable_wdata_826;
  assign _reinterpretcast_data_837 = __variable_wdata_833;
  assign _reinterpretcast_data_844 = __variable_wdata_840;
  assign _reinterpretcast_data_863 = _cond_data_857;
  assign _reinterpretcast_data_869 = __variable_wdata_864;
  assign _reinterpretcast_data_897 = _cond_data_896;
  assign _reinterpretcast_src_234 = __variable_wdata_230;
  assign _reinterpretcast_src_241 = __variable_wdata_237;
  assign _reinterpretcast_src_248 = __variable_wdata_244;
  assign _reinterpretcast_src_255 = __variable_wdata_251;
  assign _reinterpretcast_src_262 = __variable_wdata_258;
  assign _reinterpretcast_src_493 = _cond_data_376;
  assign _reinterpretcast_src_494 = _cond_data_406;
  assign _reinterpretcast_src_495 = _cond_data_436;
  assign _reinterpretcast_src_496 = _cond_data_386;
  assign _reinterpretcast_src_497 = _cond_data_416;
  assign _reinterpretcast_src_498 = _cond_data_446;
  assign _reinterpretcast_src_499 = _cond_data_396;
  assign _reinterpretcast_src_500 = _cond_data_426;
  assign _reinterpretcast_src_501 = _cond_data_456;
  assign _reinterpretcast_src_547 = __variable_wdata_502;
  assign _reinterpretcast_src_548 = __variable_wdata_503;
  assign _reinterpretcast_src_549 = __variable_wdata_504;
  assign _reinterpretcast_src_550 = __variable_wdata_505;
  assign _reinterpretcast_src_551 = __variable_wdata_506;
  assign _reinterpretcast_src_552 = __variable_wdata_507;
  assign _reinterpretcast_src_553 = __variable_wdata_508;
  assign _reinterpretcast_src_554 = __variable_wdata_509;
  assign _reinterpretcast_src_555 = __variable_wdata_510;
  assign _reinterpretcast_src_776 = _cond_data_890;
  assign _reinterpretcast_src_789 = __variable_wdata_778;
  assign _reinterpretcast_src_795 = __substreamoutput_data_793;
  assign _reinterpretcast_src_816 = __variable_wdata_812;
  assign _reinterpretcast_src_823 = __variable_wdata_819;
  assign _reinterpretcast_src_830 = __variable_wdata_826;
  assign _reinterpretcast_src_837 = __variable_wdata_833;
  assign _reinterpretcast_src_844 = __variable_wdata_840;
  assign _reinterpretcast_src_863 = _cond_data_857;
  assign _reinterpretcast_src_869 = __variable_wdata_864;
  assign _reinterpretcast_src_897 = _cond_data_896;
  assign _set_flag_1024 = _set_flag_1036;
  assign _set_flag_1025 = _set_flag_1036;
  assign _set_flag_1026 = _set_flag_1036;
  assign _set_flag_1163 = _set_flag_1224;
  assign _set_flag_1164 = _set_flag_1224;
  assign _set_flag_1165 = _set_flag_1224;
  assign _set_flag_1166 = _set_flag_1224;
  assign _set_flag_1167 = _set_flag_1224;
  assign _set_flag_1168 = _set_flag_1224;
  assign _set_flag_1169 = _set_flag_1224;
  assign _set_flag_1179 = _set_flag_1224;
  assign _set_flag_1180 = _set_flag_1224;
  assign _set_flag_1190 = _set_flag_1224;
  assign _set_flag_1191 = _set_flag_1224;
  assign _set_flag_1192 = _set_flag_1224;
  assign _set_flag_1193 = _set_flag_1224;
  assign _set_flag_1194 = _set_flag_1224;
  assign _set_flag_1195 = _set_flag_1224;
  assign _set_flag_1196 = _set_flag_1224;
  assign _set_flag_1197 = _set_flag_1224;
  assign _set_flag_1198 = _set_flag_1224;
  assign _set_flag_1199 = _set_flag_1224;
  assign _set_flag_1200 = _set_flag_1224;
  assign _set_flag_1210 = _set_flag_1224;
  assign _set_flag_457 = _set_flag_710;
  assign _set_flag_458 = _set_flag_710;
  assign _set_flag_459 = _set_flag_710;
  assign _set_flag_460 = _set_flag_710;
  assign _set_flag_461 = _set_flag_710;
  assign _set_flag_462 = _set_flag_710;
  assign _set_flag_463 = _set_flag_710;
  assign _set_flag_473 = _set_flag_710;
  assign _set_flag_474 = _set_flag_710;
  assign _set_flag_484 = _set_flag_710;
  assign _set_flag_485 = _set_flag_710;
  assign _set_flag_486 = _set_flag_710;
  assign _set_flag_487 = _set_flag_710;
  assign _set_flag_488 = _set_flag_710;
  assign _set_flag_489 = _set_flag_710;
  assign _set_flag_490 = _set_flag_710;
  assign _set_flag_491 = _set_flag_710;
  assign _set_flag_492 = _set_flag_710;
  assign _set_flag_493 = _set_flag_710;
  assign _set_flag_494 = _set_flag_710;
  assign _set_flag_504 = _set_flag_710;
  assign _set_flag_514 = _set_flag_710;
  assign _set_flag_524 = _set_flag_710;
  assign _set_flag_534 = _set_flag_710;
  assign _set_flag_544 = _set_flag_710;
  assign _set_flag_554 = _set_flag_710;
  assign _set_flag_564 = _set_flag_710;
  assign _set_flag_574 = _set_flag_710;
  assign _set_flag_584 = _set_flag_710;
  assign _set_flag_598 = _set_flag_710;
  assign _set_flag_612 = _set_flag_710;
  assign _set_flag_626 = _set_flag_710;
  assign _set_flag_640 = _set_flag_710;
  assign _set_flag_654 = _set_flag_710;
  assign _set_flag_668 = _set_flag_710;
  assign _set_flag_682 = _set_flag_710;
  assign _set_flag_696 = _set_flag_710;
  assign _slice_data_233 = __variable_wdata_230;
  assign _slice_data_240 = __variable_wdata_237;
  assign _slice_data_247 = __variable_wdata_244;
  assign _slice_data_254 = __variable_wdata_251;
  assign _slice_data_261 = __variable_wdata_258;
  assign _slice_data_815 = __variable_wdata_812;
  assign _slice_data_822 = __variable_wdata_819;
  assign _slice_data_829 = __variable_wdata_826;
  assign _slice_data_836 = __variable_wdata_833;
  assign _slice_data_843 = __variable_wdata_840;
  assign _stream_conv2d_16_sink_38_sink_wenable = 1'h0;
  assign _stream_conv2d_16_source_10_source_ram_rvalid = 1'h0;
  assign _stream_conv2d_16_source_12_source_ram_rvalid = 1'h0;
  assign _stream_conv2d_16_source_14_source_ram_rvalid = 1'h0;
  assign _stream_matmul_29_sink_22_sink_wenable = 1'h0;
  assign _stream_matmul_29_source_10_source_ram_rvalid = 1'h0;
  assign _stream_matmul_29_source_12_source_ram_rvalid = 1'h0;
  assign _stream_matmul_29_source_14_source_ram_rvalid = 1'h0;
  assign _stream_max_pool_serial_18_done = _stream_max_pool_serial_18_source_1_idle;
  assign _stream_max_pool_serial_18_sink_4_sink_wenable = 1'h0;
  assign _times_data_41 = _times_mul_odata_reg_41;
  assign \_times_mul_41.CLK  = CLK;
  assign \_times_mul_41.a  = __variable_wdata_38;
  assign \_times_mul_41.b  = __variable_wdata_39;
  assign \_times_mul_41.c  = \_times_mul_41.mult._pipe_mul1 ;
  assign \_times_mul_41.mult.CLK  = CLK;
  assign \_times_mul_41.mult.a  = __variable_wdata_38;
  assign \_times_mul_41.mult.b  = __variable_wdata_39;
  assign \_times_mul_41.mult.c  = \_times_mul_41.mult._pipe_mul1 ;
  assign \_times_mul_41.mult.update  = 1'h1;
  assign \_times_mul_41.update  = 1'h1;
  assign _times_mul_odata_41 = \_times_mul_41.mult._pipe_mul1 ;
  assign _times_mul_update_41 = 1'h1;
  assign _tmp_1010 = 1'h1;
  assign _tmp_1027 = _stream_max_pool_serial_18_source_1_source_ram_raddr[1:0];
  assign _tmp_1037 = _stream_max_pool_serial_18_sink_3_sink_waddr[1:0];
  assign _tmp_1042 = _tmp_1040;
  assign _tmp_1044 = _tmp_1040;
  assign _tmp_1046 = _tmp_1040;
  assign _tmp_1048 = _tmp_1056;
  assign _tmp_1050 = _tmp_1056;
  assign _tmp_1052 = _tmp_1056;
  assign _tmp_1054 = _tmp_1056;
  assign _tmp_1058 = _tmp_1056;
  assign _tmp_1060 = _tmp_1056;
  assign _tmp_1062 = _tmp_1056;
  assign _tmp_1064 = _tmp_1056;
  assign _tmp_1066 = _tmp_1056;
  assign _tmp_1068 = _tmp_1056;
  assign _tmp_1070 = _tmp_1056;
  assign _tmp_1075 = 1'h1;
  assign _tmp_1087 = 1'h1;
  assign _tmp_1099 = 1'h1;
  assign _tmp_1111 = 1'h1;
  assign _tmp_1170 = _stream_matmul_29_source_6_source_ram_raddr[1:0];
  assign _tmp_1181 = _stream_matmul_29_source_8_source_ram_raddr[1:0];
  assign _tmp_1201 = _stream_matmul_29_source_19_source_ram_raddr[1:0];
  assign _tmp_121 = _tmp_112;
  assign _tmp_1211 = _stream_matmul_29_source_20_source_ram_raddr[2:0];
  assign _tmp_122 = _tmp_113;
  assign _tmp_1225 = _stream_matmul_29_sink_21_sink_waddr[1:0];
  assign _tmp_1229 = _tmp_1227;
  assign _tmp_123 = _tmp_114;
  assign _tmp_1231 = _tmp_1227;
  assign _tmp_1233 = _tmp_1227;
  assign _tmp_1235 = _tmp_1227;
  assign _tmp_1237 = _tmp_1227;
  assign _tmp_1239 = _tmp_1227;
  assign _tmp_124 = _tmp_115;
  assign _tmp_1241 = _tmp_1227;
  assign _tmp_1243 = _tmp_1227;
  assign _tmp_1245 = _tmp_1227;
  assign _tmp_1247 = _tmp_1227;
  assign _tmp_1249 = _tmp_1227;
  assign _tmp_125 = _tmp_116;
  assign _tmp_1251 = _tmp_1281;
  assign _tmp_1253 = _tmp_1281;
  assign _tmp_1255 = _tmp_1281;
  assign _tmp_1257 = _tmp_1281;
  assign _tmp_1259 = _tmp_1281;
  assign _tmp_126 = _tmp_117;
  assign _tmp_1261 = _tmp_1281;
  assign _tmp_1263 = _tmp_1281;
  assign _tmp_1265 = _tmp_1281;
  assign _tmp_1267 = _tmp_1281;
  assign _tmp_1269 = _tmp_1281;
  assign _tmp_127 = _tmp_118;
  assign _tmp_1271 = _tmp_1281;
  assign _tmp_1273 = _tmp_1281;
  assign _tmp_1275 = _tmp_1281;
  assign _tmp_1277 = _tmp_1281;
  assign _tmp_1279 = _tmp_1281;
  assign _tmp_128 = _tmp_119;
  assign _tmp_1283 = _tmp_1281;
  assign _tmp_1285 = _tmp_1281;
  assign _tmp_1287 = _tmp_1281;
  assign _tmp_1289 = _tmp_1281;
  assign _tmp_129 = _tmp_120;
  assign _tmp_1291 = _tmp_1281;
  assign _tmp_1293 = _tmp_1281;
  assign _tmp_1295 = _tmp_1281;
  assign _tmp_1297 = _tmp_1281;
  assign _tmp_1299 = _tmp_1281;
  assign _tmp_1301 = _tmp_1281;
  assign _tmp_1303 = _tmp_1281;
  assign _tmp_1305 = _tmp_1281;
  assign _tmp_1307 = _tmp_1281;
  assign _tmp_1312 = 1'h1;
  assign _tmp_1324 = 1'h1;
  assign _tmp_1336 = 1'h1;
  assign _tmp_1348 = 1'h1;
  assign _tmp_152 = _tmp_143;
  assign _tmp_153 = _tmp_144;
  assign _tmp_154 = _tmp_145;
  assign _tmp_155 = _tmp_146;
  assign _tmp_156 = _tmp_147;
  assign _tmp_157 = _tmp_148;
  assign _tmp_158 = _tmp_149;
  assign _tmp_159 = _tmp_150;
  assign _tmp_160 = _tmp_151;
  assign _tmp_183 = _tmp_174;
  assign _tmp_184 = _tmp_175;
  assign _tmp_185 = _tmp_176;
  assign _tmp_186 = _tmp_177;
  assign _tmp_187 = _tmp_178;
  assign _tmp_188 = _tmp_179;
  assign _tmp_189 = _tmp_180;
  assign _tmp_190 = _tmp_181;
  assign _tmp_191 = _tmp_182;
  assign _tmp_214 = _tmp_205;
  assign _tmp_215 = _tmp_206;
  assign _tmp_216 = _tmp_207;
  assign _tmp_217 = _tmp_208;
  assign _tmp_218 = _tmp_209;
  assign _tmp_219 = _tmp_210;
  assign _tmp_220 = _tmp_211;
  assign _tmp_221 = _tmp_212;
  assign _tmp_222 = _tmp_213;
  assign _tmp_245 = _tmp_236;
  assign _tmp_246 = _tmp_237;
  assign _tmp_247 = _tmp_238;
  assign _tmp_248 = _tmp_239;
  assign _tmp_249 = _tmp_240;
  assign _tmp_250 = _tmp_241;
  assign _tmp_251 = _tmp_242;
  assign _tmp_252 = _tmp_243;
  assign _tmp_253 = _tmp_244;
  assign _tmp_276 = _tmp_267;
  assign _tmp_277 = _tmp_268;
  assign _tmp_278 = _tmp_269;
  assign _tmp_279 = _tmp_270;
  assign _tmp_280 = _tmp_271;
  assign _tmp_281 = _tmp_272;
  assign _tmp_282 = _tmp_273;
  assign _tmp_283 = _tmp_274;
  assign _tmp_284 = _tmp_275;
  assign _tmp_300 = _tmp_297;
  assign _tmp_301 = _tmp_298;
  assign _tmp_302 = _tmp_299;
  assign _tmp_313 = _tmp_310;
  assign _tmp_314 = _tmp_311;
  assign _tmp_315 = _tmp_312;
  assign _tmp_326 = _tmp_323;
  assign _tmp_327 = _tmp_324;
  assign _tmp_328 = _tmp_325;
  assign _tmp_339 = _tmp_336;
  assign _tmp_340 = _tmp_337;
  assign _tmp_341 = _tmp_338;
  assign _tmp_357 = _tmp_354;
  assign _tmp_358 = _tmp_355;
  assign _tmp_359 = _tmp_356;
  assign _tmp_370 = _tmp_367;
  assign _tmp_371 = _tmp_368;
  assign _tmp_372 = _tmp_369;
  assign _tmp_383 = _tmp_380;
  assign _tmp_384 = _tmp_381;
  assign _tmp_385 = _tmp_382;
  assign _tmp_396 = _tmp_393;
  assign _tmp_397 = _tmp_394;
  assign _tmp_398 = _tmp_395;
  assign _tmp_414 = _tmp_411;
  assign _tmp_415 = _tmp_412;
  assign _tmp_416 = _tmp_413;
  assign _tmp_427 = _tmp_424;
  assign _tmp_428 = _tmp_425;
  assign _tmp_429 = _tmp_426;
  assign _tmp_440 = _tmp_437;
  assign _tmp_441 = _tmp_438;
  assign _tmp_442 = _tmp_439;
  assign _tmp_453 = _tmp_450;
  assign _tmp_454 = _tmp_451;
  assign _tmp_455 = _tmp_452;
  assign _tmp_464 = _stream_conv2d_16_source_6_source_ram_raddr[1:0];
  assign _tmp_475 = _stream_conv2d_16_source_8_source_ram_raddr[1:0];
  assign _tmp_495 = _stream_conv2d_16_source_19_source_ram_raddr[1:0];
  assign _tmp_505 = _stream_conv2d_16_source_20_source_ram_raddr[1:0];
  assign _tmp_515 = _stream_conv2d_16_source_21_source_ram_raddr[1:0];
  assign _tmp_525 = _stream_conv2d_16_source_22_source_ram_raddr[1:0];
  assign _tmp_535 = _stream_conv2d_16_source_23_source_ram_raddr[1:0];
  assign _tmp_545 = _stream_conv2d_16_source_24_source_ram_raddr[1:0];
  assign _tmp_555 = _stream_conv2d_16_source_25_source_ram_raddr[1:0];
  assign _tmp_565 = _stream_conv2d_16_source_26_source_ram_raddr[1:0];
  assign _tmp_575 = _stream_conv2d_16_source_27_source_ram_raddr[1:0];
  assign _tmp_585 = _stream_conv2d_16_source_28_source_ram_raddr[2:0];
  assign _tmp_59 = _tmp_50;
  assign _tmp_599 = _stream_conv2d_16_source_29_source_ram_raddr[2:0];
  assign _tmp_60 = _tmp_51;
  assign _tmp_61 = _tmp_52;
  assign _tmp_613 = _stream_conv2d_16_source_30_source_ram_raddr[2:0];
  assign _tmp_62 = _tmp_53;
  assign _tmp_627 = _stream_conv2d_16_source_31_source_ram_raddr[2:0];
  assign _tmp_63 = _tmp_54;
  assign _tmp_64 = _tmp_55;
  assign _tmp_641 = _stream_conv2d_16_source_32_source_ram_raddr[2:0];
  assign _tmp_65 = _tmp_56;
  assign _tmp_655 = _stream_conv2d_16_source_33_source_ram_raddr[2:0];
  assign _tmp_66 = _tmp_57;
  assign _tmp_669 = _stream_conv2d_16_source_34_source_ram_raddr[2:0];
  assign _tmp_67 = _tmp_58;
  assign _tmp_683 = _stream_conv2d_16_source_35_source_ram_raddr[2:0];
  assign _tmp_697 = _stream_conv2d_16_source_36_source_ram_raddr[2:0];
  assign _tmp_711 = _stream_conv2d_16_sink_37_sink_waddr[1:0];
  assign _tmp_715 = _tmp_713;
  assign _tmp_717 = _tmp_713;
  assign _tmp_719 = _tmp_713;
  assign _tmp_721 = _tmp_713;
  assign _tmp_723 = _tmp_713;
  assign _tmp_725 = _tmp_713;
  assign _tmp_727 = _tmp_713;
  assign _tmp_729 = _tmp_713;
  assign _tmp_731 = _tmp_713;
  assign _tmp_733 = _tmp_713;
  assign _tmp_735 = _tmp_713;
  assign _tmp_737 = _tmp_713;
  assign _tmp_739 = _tmp_713;
  assign _tmp_741 = _tmp_713;
  assign _tmp_743 = _tmp_713;
  assign _tmp_745 = _tmp_713;
  assign _tmp_747 = _tmp_713;
  assign _tmp_749 = _tmp_713;
  assign _tmp_751 = _tmp_713;
  assign _tmp_753 = _tmp_713;
  assign _tmp_755 = _tmp_713;
  assign _tmp_757 = _tmp_713;
  assign _tmp_759 = _tmp_713;
  assign _tmp_761 = _tmp_713;
  assign _tmp_763 = _tmp_713;
  assign _tmp_765 = _tmp_713;
  assign _tmp_767 = _tmp_713;
  assign _tmp_769 = _tmp_713;
  assign _tmp_771 = _tmp_713;
  assign _tmp_773 = _tmp_713;
  assign _tmp_775 = _tmp_713;
  assign _tmp_777 = _tmp_713;
  assign _tmp_779 = _tmp_713;
  assign _tmp_781 = _tmp_713;
  assign _tmp_783 = _tmp_713;
  assign _tmp_785 = _tmp_713;
  assign _tmp_787 = _tmp_713;
  assign _tmp_789 = _tmp_713;
  assign _tmp_791 = _tmp_713;
  assign _tmp_793 = _tmp_713;
  assign _tmp_795 = _tmp_713;
  assign _tmp_797 = _tmp_713;
  assign _tmp_799 = _tmp_713;
  assign _tmp_801 = _tmp_943;
  assign _tmp_803 = _tmp_943;
  assign _tmp_805 = _tmp_943;
  assign _tmp_807 = _tmp_943;
  assign _tmp_809 = _tmp_943;
  assign _tmp_811 = _tmp_943;
  assign _tmp_813 = _tmp_943;
  assign _tmp_815 = _tmp_943;
  assign _tmp_817 = _tmp_943;
  assign _tmp_819 = _tmp_943;
  assign _tmp_821 = _tmp_943;
  assign _tmp_823 = _tmp_943;
  assign _tmp_825 = _tmp_943;
  assign _tmp_827 = _tmp_943;
  assign _tmp_829 = _tmp_943;
  assign _tmp_831 = _tmp_943;
  assign _tmp_833 = _tmp_943;
  assign _tmp_835 = _tmp_943;
  assign _tmp_837 = _tmp_943;
  assign _tmp_839 = _tmp_943;
  assign _tmp_841 = _tmp_943;
  assign _tmp_843 = _tmp_943;
  assign _tmp_845 = _tmp_943;
  assign _tmp_847 = _tmp_943;
  assign _tmp_849 = _tmp_943;
  assign _tmp_851 = _tmp_943;
  assign _tmp_853 = _tmp_943;
  assign _tmp_855 = _tmp_943;
  assign _tmp_857 = _tmp_943;
  assign _tmp_859 = _tmp_943;
  assign _tmp_861 = _tmp_943;
  assign _tmp_863 = _tmp_943;
  assign _tmp_865 = _tmp_943;
  assign _tmp_867 = _tmp_943;
  assign _tmp_869 = _tmp_943;
  assign _tmp_871 = _tmp_943;
  assign _tmp_873 = _tmp_943;
  assign _tmp_875 = _tmp_943;
  assign _tmp_877 = _tmp_943;
  assign _tmp_879 = _tmp_943;
  assign _tmp_881 = _tmp_943;
  assign _tmp_883 = _tmp_943;
  assign _tmp_885 = _tmp_943;
  assign _tmp_887 = _tmp_943;
  assign _tmp_889 = _tmp_943;
  assign _tmp_891 = _tmp_943;
  assign _tmp_893 = _tmp_943;
  assign _tmp_895 = _tmp_943;
  assign _tmp_897 = _tmp_943;
  assign _tmp_899 = _tmp_943;
  assign _tmp_90 = _tmp_81;
  assign _tmp_901 = _tmp_943;
  assign _tmp_903 = _tmp_943;
  assign _tmp_905 = _tmp_943;
  assign _tmp_907 = _tmp_943;
  assign _tmp_909 = _tmp_943;
  assign _tmp_91 = _tmp_82;
  assign _tmp_911 = _tmp_943;
  assign _tmp_913 = _tmp_943;
  assign _tmp_915 = _tmp_943;
  assign _tmp_917 = _tmp_943;
  assign _tmp_919 = _tmp_943;
  assign _tmp_92 = _tmp_83;
  assign _tmp_921 = _tmp_943;
  assign _tmp_923 = _tmp_943;
  assign _tmp_925 = _tmp_943;
  assign _tmp_927 = _tmp_943;
  assign _tmp_929 = _tmp_943;
  assign _tmp_93 = _tmp_84;
  assign _tmp_931 = _tmp_943;
  assign _tmp_933 = _tmp_943;
  assign _tmp_935 = _tmp_943;
  assign _tmp_937 = _tmp_943;
  assign _tmp_939 = _tmp_943;
  assign _tmp_94 = _tmp_85;
  assign _tmp_941 = _tmp_943;
  assign _tmp_945 = _tmp_943;
  assign _tmp_947 = _tmp_943;
  assign _tmp_949 = _tmp_943;
  assign _tmp_95 = _tmp_86;
  assign _tmp_951 = _tmp_943;
  assign _tmp_953 = _tmp_943;
  assign _tmp_955 = _tmp_943;
  assign _tmp_957 = _tmp_943;
  assign _tmp_959 = _tmp_943;
  assign _tmp_96 = _tmp_87;
  assign _tmp_961 = _tmp_943;
  assign _tmp_963 = _tmp_943;
  assign _tmp_965 = _tmp_943;
  assign _tmp_967 = _tmp_943;
  assign _tmp_969 = _tmp_943;
  assign _tmp_97 = _tmp_88;
  assign _tmp_974 = 1'h1;
  assign _tmp_98 = _tmp_89;
  assign _tmp_986 = 1'h1;
  assign _tmp_998 = 1'h1;
  assign acc_0_rshift_data = __variable_wdata_1;
  assign acc_0_size_data = __variable_wdata_2;
  assign acc_0_sum_data = _sra_data_21;
  assign acc_0_valid_data = __delay_data_758;
  assign acc_0_x_data = __variable_wdata_0;
  assign add_tree_1_sum_data = __variable_wdata_22;
  assign add_tree_1_var0_data = __variable_wdata_22;
  assign add_tree_2_sum_data = __plusn_data_37;
  assign add_tree_2_var0_data = __variable_wdata_24;
  assign add_tree_2_var1_data = __variable_wdata_25;
  assign add_tree_2_var2_data = __variable_wdata_26;
  assign add_tree_2_var3_data = __variable_wdata_27;
  assign add_tree_2_var4_data = __variable_wdata_28;
  assign add_tree_2_var5_data = __variable_wdata_29;
  assign add_tree_2_var6_data = __variable_wdata_30;
  assign add_tree_2_var7_data = __variable_wdata_31;
  assign add_tree_2_var8_data = __variable_wdata_32;
  assign conv2d_16_stream_out_local = conv2d_16_stream_out_local_col;
  assign conv2d_16_stream_out_local_val = 0;
  assign conv2d_16_update_act = 1'h1;
  assign cparam_conv2d_16_act_func_index = 1'h0;
  assign cparam_conv2d_16_act_num_col = cparam_conv2d_16_act_num_row;
  assign cparam_conv2d_16_act_offset_values_1 = 0;
  assign cparam_conv2d_16_act_read_block = cparam_conv2d_16_inc_act_laddr_large;
  assign cparam_conv2d_16_act_read_size = cparam_conv2d_16_act_offset_values_2[8:0];
  assign cparam_conv2d_16_act_row_step = cparam_conv2d_16_act_offset_values_2[8:0];
  assign cparam_conv2d_16_bias_scala = 1'h0;
  assign cparam_conv2d_16_col_select_initval = 2'h2;
  assign cparam_conv2d_16_cshamt_mul_value = 1'h0;
  assign cparam_conv2d_16_cshamt_sum_value = 1'h0;
  assign cparam_conv2d_16_data_stationary = 1'h0;
  assign cparam_conv2d_16_dma_flag_conds_0 = 1'h1;
  assign cparam_conv2d_16_dma_flag_conds_1 = 1'h0;
  assign cparam_conv2d_16_dma_flag_conds_2 = 1'h0;
  assign cparam_conv2d_16_filter_num_col_minus_stride_col_mod = 2'h2;
  assign cparam_conv2d_16_inc_act_laddr_conds_0 = 1'h1;
  assign cparam_conv2d_16_inc_act_laddr_conds_1 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_10 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_11 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_12 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_13 = 1'h1;
  assign cparam_conv2d_16_inc_act_laddr_conds_14 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_15 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_16 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_17 = 1'h1;
  assign cparam_conv2d_16_inc_act_laddr_conds_18 = 1'h1;
  assign cparam_conv2d_16_inc_act_laddr_conds_19 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_2 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_20 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_21 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_22 = 1'h1;
  assign cparam_conv2d_16_inc_act_laddr_conds_23 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_24 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_25 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_26 = 1'h1;
  assign cparam_conv2d_16_inc_act_laddr_conds_3 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_4 = 1'h1;
  assign cparam_conv2d_16_inc_act_laddr_conds_5 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_6 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_7 = 1'h0;
  assign cparam_conv2d_16_inc_act_laddr_conds_8 = 1'h1;
  assign cparam_conv2d_16_inc_act_laddr_conds_9 = 1'h1;
  assign cparam_conv2d_16_inc_act_laddr_small = 1'h0;
  assign cparam_conv2d_16_inc_out_laddr_col = cparam_conv2d_16_bias_num;
  assign cparam_conv2d_16_inc_sync_out = cparam_conv2d_16_act_num_row;
  assign cparam_conv2d_16_inc_sync_out_res = 1'h0;
  assign cparam_conv2d_16_keep_filter = 1'h1;
  assign cparam_conv2d_16_keep_input = 1'h1;
  assign cparam_conv2d_16_max_bat_count = 1'h0;
  assign cparam_conv2d_16_max_och_count = 1'h0;
  assign cparam_conv2d_16_max_row_count = cparam_conv2d_16_max_col_count;
  assign cparam_conv2d_16_out_col_step = cparam_conv2d_16_bias_num;
  assign cparam_conv2d_16_out_num_col = cparam_conv2d_16_act_num_row;
  assign cparam_conv2d_16_out_num_row = cparam_conv2d_16_act_num_row;
  assign cparam_conv2d_16_out_och_step = cparam_conv2d_16_bias_num;
  assign cparam_conv2d_16_out_offset_values_0 = 1'h0;
  assign cparam_conv2d_16_out_row_step = 10'h200;
  assign cparam_conv2d_16_out_write_size = 10'h200;
  assign cparam_conv2d_16_out_write_size_res = 10'h200;
  assign cparam_conv2d_16_pad_col_left = 1'h1;
  assign cparam_conv2d_16_pad_row_top = 1'h1;
  assign cparam_conv2d_16_scale_num = 1'h1;
  assign cparam_conv2d_16_scale_scala = 1'h1;
  assign cparam_conv2d_16_stream_act_local_large_flags_0 = 1'h0;
  assign cparam_conv2d_16_stream_act_local_large_flags_1 = 1'h0;
  assign cparam_conv2d_16_stream_act_local_large_flags_2 = 1'h1;
  assign cparam_conv2d_16_stream_act_local_small_flags_0 = 1'h0;
  assign cparam_conv2d_16_stream_act_local_small_flags_1 = 1'h0;
  assign cparam_conv2d_16_stream_act_local_small_flags_2 = 1'h1;
  assign cparam_conv2d_16_stream_act_local_small_offset = 1'h0;
  assign cparam_conv2d_16_stream_aligned_reduce_size = cparam_conv2d_16_filter_read_block;
  assign cparam_conv2d_16_stream_num_ops = cparam_conv2d_16_bias_num;
  assign cparam_conv2d_16_stream_num_ops_res = cparam_conv2d_16_bias_num;
  assign cparam_conv2d_16_stream_omit_mask = 1'h0;
  assign cparam_conv2d_16_stride_col_mod_filter_num = 1'h1;
  assign cparam_conv2d_16_stride_col_par_col = 1'h1;
  assign cparam_conv2d_16_stride_row_par_row = 1'h1;
  assign cparam_conv2d_16_vshamt_mul_num = 1'h0;
  assign cparam_conv2d_16_vshamt_mul_scala = 1'h0;
  assign cparam_conv2d_16_vshamt_out_num = 1'h0;
  assign cparam_conv2d_16_vshamt_out_scala = 1'h0;
  assign cparam_conv2d_16_vshamt_sum_num = 1'h0;
  assign cparam_conv2d_16_vshamt_sum_scala = 1'h0;
  assign cparam_matmul_29_act_func_index = cparam_matmul_29_keep_filter;
  assign cparam_matmul_29_act_num_col = 1'h1;
  assign cparam_matmul_29_act_num_row = 1'h1;
  assign cparam_matmul_29_act_offset_values_0 = 0;
  assign cparam_matmul_29_act_read_size = cparam_matmul_29_act_bat_step;
  assign cparam_matmul_29_act_read_step = cparam_matmul_29_act_bat_step;
  assign cparam_matmul_29_act_row_step = cparam_matmul_29_act_bat_step;
  assign cparam_matmul_29_bias_scala = 1'h0;
  assign cparam_matmul_29_col_select_initval = 1'h0;
  assign cparam_matmul_29_cshamt_mul_value = 1'h0;
  assign cparam_matmul_29_cshamt_sum_value = 1'h0;
  assign cparam_matmul_29_data_stationary = 1'h0;
  assign cparam_matmul_29_dma_flag_conds_0 = 1'h1;
  assign cparam_matmul_29_filter_num_col_minus_stride_col_mod = 1'h1;
  assign cparam_matmul_29_filter_read_step = cparam_matmul_29_filter_read_size;
  assign cparam_matmul_29_inc_act_laddr_conds_0 = 1'h0;
  assign cparam_matmul_29_inc_act_laddr_large = cparam_matmul_29_act_bat_step;
  assign cparam_matmul_29_inc_act_laddr_small = cparam_matmul_29_act_bat_step;
  assign cparam_matmul_29_inc_out_laddr_col = cparam_matmul_29_bias_num;
  assign cparam_matmul_29_inc_sync_out = 1'h1;
  assign cparam_matmul_29_inc_sync_out_res = 1'h0;
  assign cparam_matmul_29_keep_input = 1'h1;
  assign cparam_matmul_29_max_bat_count = 1'h0;
  assign cparam_matmul_29_max_col_count = 1'h0;
  assign cparam_matmul_29_max_row_count = 1'h0;
  assign cparam_matmul_29_out_col_step = cparam_matmul_29_out_bat_step;
  assign cparam_matmul_29_out_num_col = 1'h1;
  assign cparam_matmul_29_out_num_row = 1'h1;
  assign cparam_matmul_29_out_offset_values_0 = 1'h0;
  assign cparam_matmul_29_out_row_step = cparam_matmul_29_out_bat_step;
  assign cparam_matmul_29_out_write_size_res = cparam_matmul_29_out_write_size;
  assign cparam_matmul_29_pad_col_left = 1'h0;
  assign cparam_matmul_29_pad_row_top = 1'h0;
  assign cparam_matmul_29_scale_num = 1'h1;
  assign cparam_matmul_29_scale_scala = 1'h1;
  assign cparam_matmul_29_stream_act_local_large_flags_0 = 1'h0;
  assign cparam_matmul_29_stream_act_local_large_offset = 1'h0;
  assign cparam_matmul_29_stream_act_local_small_flags_0 = 1'h0;
  assign cparam_matmul_29_stream_act_local_small_offset = 1'h0;
  assign cparam_matmul_29_stream_aligned_reduce_size = cparam_matmul_29_act_bat_step;
  assign cparam_matmul_29_stream_num_ops = cparam_matmul_29_out_write_size;
  assign cparam_matmul_29_stream_num_ops_res = cparam_matmul_29_out_write_size;
  assign cparam_matmul_29_stream_omit_mask = 1'h0;
  assign cparam_matmul_29_stream_reduce_size = cparam_matmul_29_act_bat_step;
  assign cparam_matmul_29_stride_col_mod_filter_num = 1'h0;
  assign cparam_matmul_29_stride_col_par_col = 1'h1;
  assign cparam_matmul_29_stride_row_par_row = 1'h1;
  assign cparam_matmul_29_vshamt_mul_num = 1'h0;
  assign cparam_matmul_29_vshamt_mul_scala = 1'h0;
  assign cparam_matmul_29_vshamt_out_num = 1'h0;
  assign cparam_matmul_29_vshamt_out_scala = 1'h0;
  assign cparam_matmul_29_vshamt_sum_num = 1'h0;
  assign cparam_matmul_29_vshamt_sum_scala = 1'h0;
  assign cparam_max_pool_serial_18_act_num_row = cparam_max_pool_serial_18_act_num_col;
  assign cparam_max_pool_serial_18_act_offset_values_0 = 0;
  assign cparam_max_pool_serial_18_act_offset_values_1 = 512;
  assign cparam_max_pool_serial_18_act_read_block = cparam_max_pool_serial_18_inc_out_laddr;
  assign cparam_max_pool_serial_18_act_read_size = 10'h200;
  assign cparam_max_pool_serial_18_act_row_step = 11'h400;
  assign cparam_max_pool_serial_18_col_select_initval = 1'h0;
  assign cparam_max_pool_serial_18_ksize_col_minus_stride_col_mod = 2'h2;
  assign cparam_max_pool_serial_18_local_pad_offset = 1'h0;
  assign cparam_max_pool_serial_18_max_bat_count = 1'h0;
  assign cparam_max_pool_serial_18_max_row_count = cparam_max_pool_serial_18_max_col_count;
  assign cparam_max_pool_serial_18_out_row_step = 9'h100;
  assign cparam_max_pool_serial_18_out_write_size = 9'h100;
  assign cparam_max_pool_serial_18_pad_col_left = 1'h0;
  assign cparam_max_pool_serial_18_pad_row_top = 1'h0;
  assign cparam_max_pool_serial_18_stream_size = cparam_max_pool_serial_18_inc_out_laddr;
  assign cparam_max_pool_serial_18_stride_col = 2'h2;
  assign cparam_max_pool_serial_18_stride_col_mod_ksize = 1'h0;
  assign cparam_max_pool_serial_18_stride_row = 2'h2;
  assign matmul_29_stream_out_local = matmul_29_stream_out_local_col;
  assign matmul_29_stream_out_local_val = 0;
  assign matmul_29_update_act = 1'h1;
  assign matmul_29_update_filter = 1'h1;
  assign maxi_arburst = 2'h1;
  assign maxi_arcache = 4'h3;
  assign maxi_arlock = 1'h0;
  assign maxi_arprot = 3'h0;
  assign maxi_arqos = 4'h0;
  assign maxi_arsize = 3'h2;
  assign maxi_aruser = 2'h0;
  assign maxi_awburst = 2'h1;
  assign maxi_awcache = 4'h3;
  assign maxi_awlock = 1'h0;
  assign maxi_awprot = 3'h0;
  assign maxi_awqos = 4'h0;
  assign maxi_awsize = 3'h2;
  assign maxi_awuser = 2'h0;
  assign maxi_bready = 1'h1;
  assign mul_10_rshift_data = __variable_wdata_158;
  assign mul_10_x_data = __variable_wdata_156;
  assign mul_10_y_data = __variable_wdata_157;
  assign mul_10_z_data = _sra_data_172;
  assign mul_11_rshift_data = __variable_wdata_175;
  assign mul_11_x_data = __variable_wdata_173;
  assign mul_11_y_data = __variable_wdata_174;
  assign mul_11_z_data = _sra_data_189;
  assign mul_12_rshift_data = __variable_wdata_192;
  assign mul_12_x_data = __variable_wdata_190;
  assign mul_12_y_data = __variable_wdata_191;
  assign mul_12_z_data = _sra_data_206;
  assign mul_4_rshift_data = __variable_wdata_56;
  assign mul_4_x_data = __variable_wdata_54;
  assign mul_4_y_data = __variable_wdata_55;
  assign mul_4_z_data = _sra_data_70;
  assign mul_5_rshift_data = __variable_wdata_73;
  assign mul_5_x_data = __variable_wdata_71;
  assign mul_5_y_data = __variable_wdata_72;
  assign mul_5_z_data = _sra_data_87;
  assign mul_6_rshift_data = __variable_wdata_90;
  assign mul_6_x_data = __variable_wdata_88;
  assign mul_6_y_data = __variable_wdata_89;
  assign mul_6_z_data = _sra_data_104;
  assign mul_7_rshift_data = __variable_wdata_107;
  assign mul_7_x_data = __variable_wdata_105;
  assign mul_7_y_data = __variable_wdata_106;
  assign mul_7_z_data = _sra_data_121;
  assign mul_8_rshift_data = __variable_wdata_124;
  assign mul_8_x_data = __variable_wdata_122;
  assign mul_8_y_data = __variable_wdata_123;
  assign mul_8_z_data = _sra_data_138;
  assign mul_9_rshift_data = __variable_wdata_141;
  assign mul_9_x_data = __variable_wdata_139;
  assign mul_9_y_data = __variable_wdata_140;
  assign mul_9_z_data = _sra_data_155;
  assign mul_rshift_clip_3_rshift_data = __variable_wdata_40;
  assign mul_rshift_clip_3_x_data = __variable_wdata_38;
  assign mul_rshift_clip_3_y_data = __variable_wdata_39;
  assign mul_rshift_clip_3_z_data = _cond_data_53;
  assign ram_w4_l8192_id0_0_0_wdata = 4'h0;
  assign ram_w4_l8192_id0_0_0_wenable = 1'h0;
  assign ram_w4_l8192_id0_1_0_wdata = 4'h0;
  assign ram_w4_l8192_id0_1_0_wenable = 1'h0;
  assign ram_w4_l8192_id0_2_0_wdata = 4'h0;
  assign ram_w4_l8192_id0_2_0_wenable = 1'h0;
  assign ram_w4_l8192_id0_3_0_wdata = 4'h0;
  assign ram_w4_l8192_id0_3_0_wenable = 1'h0;
  assign ram_w4_l8192_id0_4_0_wdata = 4'h0;
  assign ram_w4_l8192_id0_4_0_wenable = 1'h0;
  assign ram_w4_l8192_id0_5_0_wdata = 4'h0;
  assign ram_w4_l8192_id0_5_0_wenable = 1'h0;
  assign ram_w4_l8192_id0_6_0_wdata = 4'h0;
  assign ram_w4_l8192_id0_6_0_wenable = 1'h0;
  assign ram_w4_l8192_id0_7_0_wdata = 4'h0;
  assign ram_w4_l8192_id0_7_0_wenable = 1'h0;
  assign ram_w4_l8192_id1_0_0_wdata = 4'h0;
  assign ram_w4_l8192_id1_0_0_wenable = 1'h0;
  assign ram_w4_l8192_id1_1_0_wdata = 4'h0;
  assign ram_w4_l8192_id1_1_0_wenable = 1'h0;
  assign ram_w4_l8192_id1_2_0_wdata = 4'h0;
  assign ram_w4_l8192_id1_2_0_wenable = 1'h0;
  assign ram_w4_l8192_id1_3_0_wdata = 4'h0;
  assign ram_w4_l8192_id1_3_0_wenable = 1'h0;
  assign ram_w4_l8192_id1_4_0_wdata = 4'h0;
  assign ram_w4_l8192_id1_4_0_wenable = 1'h0;
  assign ram_w4_l8192_id1_5_0_wdata = 4'h0;
  assign ram_w4_l8192_id1_5_0_wenable = 1'h0;
  assign ram_w4_l8192_id1_6_0_wdata = 4'h0;
  assign ram_w4_l8192_id1_6_0_wenable = 1'h0;
  assign ram_w4_l8192_id1_7_0_wdata = 4'h0;
  assign ram_w4_l8192_id1_7_0_wenable = 1'h0;
  assign ram_w4_l8192_id2_0_0_wdata = 4'h0;
  assign ram_w4_l8192_id2_0_0_wenable = 1'h0;
  assign ram_w4_l8192_id2_1_0_wdata = 4'h0;
  assign ram_w4_l8192_id2_1_0_wenable = 1'h0;
  assign ram_w4_l8192_id2_2_0_wdata = 4'h0;
  assign ram_w4_l8192_id2_2_0_wenable = 1'h0;
  assign ram_w4_l8192_id2_3_0_wdata = 4'h0;
  assign ram_w4_l8192_id2_3_0_wenable = 1'h0;
  assign ram_w4_l8192_id2_4_0_wdata = 4'h0;
  assign ram_w4_l8192_id2_4_0_wenable = 1'h0;
  assign ram_w4_l8192_id2_5_0_wdata = 4'h0;
  assign ram_w4_l8192_id2_5_0_wenable = 1'h0;
  assign ram_w4_l8192_id2_6_0_wdata = 4'h0;
  assign ram_w4_l8192_id2_6_0_wenable = 1'h0;
  assign ram_w4_l8192_id2_7_0_wdata = 4'h0;
  assign ram_w4_l8192_id2_7_0_wenable = 1'h0;
  assign ram_w4_l8192_id3_0_0_wdata = 4'h0;
  assign ram_w4_l8192_id3_0_0_wenable = 1'h0;
  assign ram_w4_l8192_id3_1_0_wdata = 4'h0;
  assign ram_w4_l8192_id3_1_0_wenable = 1'h0;
  assign ram_w4_l8192_id3_2_0_wdata = 4'h0;
  assign ram_w4_l8192_id3_2_0_wenable = 1'h0;
  assign ram_w4_l8192_id3_3_0_wdata = 4'h0;
  assign ram_w4_l8192_id3_3_0_wenable = 1'h0;
  assign ram_w4_l8192_id3_4_0_wdata = 4'h0;
  assign ram_w4_l8192_id3_4_0_wenable = 1'h0;
  assign ram_w4_l8192_id3_5_0_wdata = 4'h0;
  assign ram_w4_l8192_id3_5_0_wenable = 1'h0;
  assign ram_w4_l8192_id3_6_0_wdata = 4'h0;
  assign ram_w4_l8192_id3_6_0_wenable = 1'h0;
  assign ram_w4_l8192_id3_7_0_wdata = 4'h0;
  assign ram_w4_l8192_id3_7_0_wenable = 1'h0;
  assign ram_w4_l8192_id4_0_0_wdata = 4'h0;
  assign ram_w4_l8192_id4_0_0_wenable = 1'h0;
  assign ram_w4_l8192_id4_1_0_wdata = 4'h0;
  assign ram_w4_l8192_id4_1_0_wenable = 1'h0;
  assign ram_w4_l8192_id4_2_0_wdata = 4'h0;
  assign ram_w4_l8192_id4_2_0_wenable = 1'h0;
  assign ram_w4_l8192_id4_3_0_wdata = 4'h0;
  assign ram_w4_l8192_id4_3_0_wenable = 1'h0;
  assign ram_w4_l8192_id4_4_0_wdata = 4'h0;
  assign ram_w4_l8192_id4_4_0_wenable = 1'h0;
  assign ram_w4_l8192_id4_5_0_wdata = 4'h0;
  assign ram_w4_l8192_id4_5_0_wenable = 1'h0;
  assign ram_w4_l8192_id4_6_0_wdata = 4'h0;
  assign ram_w4_l8192_id4_6_0_wenable = 1'h0;
  assign ram_w4_l8192_id4_7_0_wdata = 4'h0;
  assign ram_w4_l8192_id4_7_0_wenable = 1'h0;
  assign ram_w4_l8192_id5_0_0_wdata = 4'h0;
  assign ram_w4_l8192_id5_0_0_wenable = 1'h0;
  assign ram_w4_l8192_id5_1_0_wdata = 4'h0;
  assign ram_w4_l8192_id5_1_0_wenable = 1'h0;
  assign ram_w4_l8192_id5_2_0_wdata = 4'h0;
  assign ram_w4_l8192_id5_2_0_wenable = 1'h0;
  assign ram_w4_l8192_id5_3_0_wdata = 4'h0;
  assign ram_w4_l8192_id5_3_0_wenable = 1'h0;
  assign ram_w4_l8192_id5_4_0_wdata = 4'h0;
  assign ram_w4_l8192_id5_4_0_wenable = 1'h0;
  assign ram_w4_l8192_id5_5_0_wdata = 4'h0;
  assign ram_w4_l8192_id5_5_0_wenable = 1'h0;
  assign ram_w4_l8192_id5_6_0_wdata = 4'h0;
  assign ram_w4_l8192_id5_6_0_wenable = 1'h0;
  assign ram_w4_l8192_id5_7_0_wdata = 4'h0;
  assign ram_w4_l8192_id5_7_0_wenable = 1'h0;
  assign ram_w4_l8192_id6_0_0_wdata = 4'h0;
  assign ram_w4_l8192_id6_0_0_wenable = 1'h0;
  assign ram_w4_l8192_id6_1_0_wdata = 4'h0;
  assign ram_w4_l8192_id6_1_0_wenable = 1'h0;
  assign ram_w4_l8192_id6_2_0_wdata = 4'h0;
  assign ram_w4_l8192_id6_2_0_wenable = 1'h0;
  assign ram_w4_l8192_id6_3_0_wdata = 4'h0;
  assign ram_w4_l8192_id6_3_0_wenable = 1'h0;
  assign ram_w4_l8192_id6_4_0_wdata = 4'h0;
  assign ram_w4_l8192_id6_4_0_wenable = 1'h0;
  assign ram_w4_l8192_id6_5_0_wdata = 4'h0;
  assign ram_w4_l8192_id6_5_0_wenable = 1'h0;
  assign ram_w4_l8192_id6_6_0_wdata = 4'h0;
  assign ram_w4_l8192_id6_6_0_wenable = 1'h0;
  assign ram_w4_l8192_id6_7_0_wdata = 4'h0;
  assign ram_w4_l8192_id6_7_0_wenable = 1'h0;
  assign ram_w4_l8192_id7_0_0_wdata = 4'h0;
  assign ram_w4_l8192_id7_0_0_wenable = 1'h0;
  assign ram_w4_l8192_id7_1_0_wdata = 4'h0;
  assign ram_w4_l8192_id7_1_0_wenable = 1'h0;
  assign ram_w4_l8192_id7_2_0_wdata = 4'h0;
  assign ram_w4_l8192_id7_2_0_wenable = 1'h0;
  assign ram_w4_l8192_id7_3_0_wdata = 4'h0;
  assign ram_w4_l8192_id7_3_0_wenable = 1'h0;
  assign ram_w4_l8192_id7_4_0_wdata = 4'h0;
  assign ram_w4_l8192_id7_4_0_wenable = 1'h0;
  assign ram_w4_l8192_id7_5_0_wdata = 4'h0;
  assign ram_w4_l8192_id7_5_0_wenable = 1'h0;
  assign ram_w4_l8192_id7_6_0_wdata = 4'h0;
  assign ram_w4_l8192_id7_6_0_wenable = 1'h0;
  assign ram_w4_l8192_id7_7_0_wdata = 4'h0;
  assign ram_w4_l8192_id7_7_0_wenable = 1'h0;
  assign ram_w4_l8192_id8_0_0_wdata = 4'h0;
  assign ram_w4_l8192_id8_0_0_wenable = 1'h0;
  assign ram_w4_l8192_id8_1_0_wdata = 4'h0;
  assign ram_w4_l8192_id8_1_0_wenable = 1'h0;
  assign ram_w4_l8192_id8_2_0_wdata = 4'h0;
  assign ram_w4_l8192_id8_2_0_wenable = 1'h0;
  assign ram_w4_l8192_id8_3_0_wdata = 4'h0;
  assign ram_w4_l8192_id8_3_0_wenable = 1'h0;
  assign ram_w4_l8192_id8_4_0_wdata = 4'h0;
  assign ram_w4_l8192_id8_4_0_wenable = 1'h0;
  assign ram_w4_l8192_id8_5_0_wdata = 4'h0;
  assign ram_w4_l8192_id8_5_0_wenable = 1'h0;
  assign ram_w4_l8192_id8_6_0_wdata = 4'h0;
  assign ram_w4_l8192_id8_6_0_wenable = 1'h0;
  assign ram_w4_l8192_id8_7_0_wdata = 4'h0;
  assign ram_w4_l8192_id8_7_0_wenable = 1'h0;
  assign ram_w8_l2048_id10_0_0_wdata = 8'h00;
  assign ram_w8_l2048_id10_0_0_wenable = 1'h0;
  assign ram_w8_l2048_id10_1_0_wdata = 8'h00;
  assign ram_w8_l2048_id10_1_0_wenable = 1'h0;
  assign ram_w8_l2048_id10_2_0_wdata = 8'h00;
  assign ram_w8_l2048_id10_2_0_wenable = 1'h0;
  assign ram_w8_l2048_id10_3_0_wdata = 8'h00;
  assign ram_w8_l2048_id10_3_0_wenable = 1'h0;
  assign ram_w8_l2048_id11_0_1_wdata = 8'h00;
  assign ram_w8_l2048_id11_0_1_wenable = 1'h0;
  assign ram_w8_l2048_id11_1_1_wdata = 8'h00;
  assign ram_w8_l2048_id11_1_1_wenable = 1'h0;
  assign ram_w8_l2048_id11_2_1_wdata = 8'h00;
  assign ram_w8_l2048_id11_2_1_wenable = 1'h0;
  assign ram_w8_l2048_id11_3_1_wdata = 8'h00;
  assign ram_w8_l2048_id11_3_1_wenable = 1'h0;
  assign ram_w8_l2048_id2_0_0_wdata = 8'h00;
  assign ram_w8_l2048_id2_0_0_wenable = 1'h0;
  assign ram_w8_l2048_id2_1_0_wdata = 8'h00;
  assign ram_w8_l2048_id2_1_0_wenable = 1'h0;
  assign ram_w8_l2048_id2_2_0_wdata = 8'h00;
  assign ram_w8_l2048_id2_2_0_wenable = 1'h0;
  assign ram_w8_l2048_id2_3_0_wdata = 8'h00;
  assign ram_w8_l2048_id2_3_0_wenable = 1'h0;
  assign ram_w8_l2048_id3_0_0_wdata = 8'h00;
  assign ram_w8_l2048_id3_0_0_wenable = 1'h0;
  assign ram_w8_l2048_id3_1_0_wdata = 8'h00;
  assign ram_w8_l2048_id3_1_0_wenable = 1'h0;
  assign ram_w8_l2048_id3_2_0_wdata = 8'h00;
  assign ram_w8_l2048_id3_2_0_wenable = 1'h0;
  assign ram_w8_l2048_id3_3_0_wdata = 8'h00;
  assign ram_w8_l2048_id3_3_0_wenable = 1'h0;
  assign ram_w8_l2048_id4_0_0_wdata = 8'h00;
  assign ram_w8_l2048_id4_0_0_wenable = 1'h0;
  assign ram_w8_l2048_id4_1_0_wdata = 8'h00;
  assign ram_w8_l2048_id4_1_0_wenable = 1'h0;
  assign ram_w8_l2048_id4_2_0_wdata = 8'h00;
  assign ram_w8_l2048_id4_2_0_wenable = 1'h0;
  assign ram_w8_l2048_id4_3_0_wdata = 8'h00;
  assign ram_w8_l2048_id4_3_0_wenable = 1'h0;
  assign ram_w8_l2048_id5_0_0_wdata = 8'h00;
  assign ram_w8_l2048_id5_0_0_wenable = 1'h0;
  assign ram_w8_l2048_id5_1_0_wdata = 8'h00;
  assign ram_w8_l2048_id5_1_0_wenable = 1'h0;
  assign ram_w8_l2048_id5_2_0_wdata = 8'h00;
  assign ram_w8_l2048_id5_2_0_wenable = 1'h0;
  assign ram_w8_l2048_id5_3_0_wdata = 8'h00;
  assign ram_w8_l2048_id5_3_0_wenable = 1'h0;
  assign ram_w8_l2048_id6_0_0_wdata = 8'h00;
  assign ram_w8_l2048_id6_0_0_wenable = 1'h0;
  assign ram_w8_l2048_id6_1_0_wdata = 8'h00;
  assign ram_w8_l2048_id6_1_0_wenable = 1'h0;
  assign ram_w8_l2048_id6_2_0_wdata = 8'h00;
  assign ram_w8_l2048_id6_2_0_wenable = 1'h0;
  assign ram_w8_l2048_id6_3_0_wdata = 8'h00;
  assign ram_w8_l2048_id6_3_0_wenable = 1'h0;
  assign ram_w8_l2048_id7_0_0_wdata = 8'h00;
  assign ram_w8_l2048_id7_0_0_wenable = 1'h0;
  assign ram_w8_l2048_id7_1_0_wdata = 8'h00;
  assign ram_w8_l2048_id7_1_0_wenable = 1'h0;
  assign ram_w8_l2048_id7_2_0_wdata = 8'h00;
  assign ram_w8_l2048_id7_2_0_wenable = 1'h0;
  assign ram_w8_l2048_id7_3_0_wdata = 8'h00;
  assign ram_w8_l2048_id7_3_0_wenable = 1'h0;
  assign ram_w8_l2048_id8_0_0_wdata = 8'h00;
  assign ram_w8_l2048_id8_0_0_wenable = 1'h0;
  assign ram_w8_l2048_id8_1_0_wdata = 8'h00;
  assign ram_w8_l2048_id8_1_0_wenable = 1'h0;
  assign ram_w8_l2048_id8_2_0_wdata = 8'h00;
  assign ram_w8_l2048_id8_2_0_wenable = 1'h0;
  assign ram_w8_l2048_id8_3_0_wdata = 8'h00;
  assign ram_w8_l2048_id8_3_0_wenable = 1'h0;
  assign ram_w8_l2048_id9_0_0_wdata = 8'h00;
  assign ram_w8_l2048_id9_0_0_wenable = 1'h0;
  assign ram_w8_l2048_id9_1_0_wdata = 8'h00;
  assign ram_w8_l2048_id9_1_0_wenable = 1'h0;
  assign ram_w8_l2048_id9_2_0_wdata = 8'h00;
  assign ram_w8_l2048_id9_2_0_wenable = 1'h0;
  assign ram_w8_l2048_id9_3_0_wdata = 8'h00;
  assign ram_w8_l2048_id9_3_0_wenable = 1'h0;
  assign saxi_bresp = 2'h0;
  assign saxi_rresp = 2'h0;
  assign stream_conv2d_16_constant_0_data = __variable_wdata_214;
  assign stream_conv2d_16_constant_15_data = __variable_wdata_264;
  assign stream_conv2d_16_constant_16_data = __variable_wdata_265;
  assign stream_conv2d_16_constant_17_data = __variable_wdata_266;
  assign stream_conv2d_16_constant_1_data = __variable_wdata_215;
  assign stream_conv2d_16_constant_2_data = __variable_wdata_216;
  assign stream_conv2d_16_constant_3_data = __variable_wdata_217;
  assign stream_conv2d_16_sink_37_data = _cond_data_890;
  assign stream_conv2d_16_sink_38_data = __delay_data_1614;
  assign stream_conv2d_16_source_10_data = __variable_wdata_244;
  assign stream_conv2d_16_source_12_data = __variable_wdata_251;
  assign stream_conv2d_16_source_14_data = __variable_wdata_258;
  assign stream_conv2d_16_source_19_data = __variable_wdata_268;
  assign stream_conv2d_16_source_20_data = __variable_wdata_269;
  assign stream_conv2d_16_source_21_data = __variable_wdata_270;
  assign stream_conv2d_16_source_22_data = __variable_wdata_271;
  assign stream_conv2d_16_source_23_data = __variable_wdata_272;
  assign stream_conv2d_16_source_24_data = __variable_wdata_273;
  assign stream_conv2d_16_source_25_data = __variable_wdata_274;
  assign stream_conv2d_16_source_26_data = __variable_wdata_275;
  assign stream_conv2d_16_source_27_data = __variable_wdata_276;
  assign stream_conv2d_16_source_28_data = __variable_wdata_502;
  assign stream_conv2d_16_source_29_data = __variable_wdata_503;
  assign stream_conv2d_16_source_30_data = __variable_wdata_504;
  assign stream_conv2d_16_source_31_data = __variable_wdata_505;
  assign stream_conv2d_16_source_32_data = __variable_wdata_506;
  assign stream_conv2d_16_source_33_data = __variable_wdata_507;
  assign stream_conv2d_16_source_34_data = __variable_wdata_508;
  assign stream_conv2d_16_source_35_data = __variable_wdata_509;
  assign stream_conv2d_16_source_36_data = __variable_wdata_510;
  assign stream_conv2d_16_source_6_data = __variable_wdata_230;
  assign stream_conv2d_16_source_8_data = __variable_wdata_237;
  assign stream_matmul_29_constant_0_data = __variable_wdata_796;
  assign stream_matmul_29_constant_15_data = __variable_wdata_846;
  assign stream_matmul_29_constant_16_data = __variable_wdata_847;
  assign stream_matmul_29_constant_17_data = __variable_wdata_848;
  assign stream_matmul_29_constant_18_data = __variable_wdata_849;
  assign stream_matmul_29_constant_1_data = __variable_wdata_797;
  assign stream_matmul_29_constant_2_data = __variable_wdata_798;
  assign stream_matmul_29_constant_3_data = __variable_wdata_799;
  assign stream_matmul_29_sink_21_data = _cond_data_896;
  assign stream_matmul_29_sink_22_data = __delay_data_1616;
  assign stream_matmul_29_source_10_data = __variable_wdata_826;
  assign stream_matmul_29_source_12_data = __variable_wdata_833;
  assign stream_matmul_29_source_14_data = __variable_wdata_840;
  assign stream_matmul_29_source_19_data = __variable_wdata_850;
  assign stream_matmul_29_source_20_data = __variable_wdata_864;
  assign stream_matmul_29_source_6_data = __variable_wdata_812;
  assign stream_matmul_29_source_8_data = __variable_wdata_819;
  assign stream_max_pool_serial_18_constant_0_data = __variable_wdata_777;
  assign stream_max_pool_serial_18_constant_2_data = __variable_wdata_779;
  assign stream_max_pool_serial_18_sink_3_data = __substreamoutput_data_793;
  assign stream_max_pool_serial_18_sink_4_data = __substreamoutput_data_794;
  assign stream_max_pool_serial_18_source_1_data = __variable_wdata_778;
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29453_ ( .A({ _06896_, _06886_ }), .Y(_05728_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29454_ ( .A({ _06887_, _06891_, main_fsm[4] }), .Y(_06886_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _29455_ ( .A({ _06888_, _06890_, _06889_, main_fsm[5] }), .Y(_06887_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29456_ ( .A(main_fsm[15:12]), .Y(_06888_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29457_ ( .A(main_fsm[11:8]), .Y(_06889_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29458_ ( .A({ main_fsm[6], main_fsm[7] }), .Y(_06890_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29459_ ( .A({ _06895_, _06894_, _06893_, _06892_ }), .Y(_06891_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29460_ ( .A(main_fsm[23:20]), .Y(_06892_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29461_ ( .A(main_fsm[19:16]), .Y(_06893_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29462_ ( .A(main_fsm[31:28]), .Y(_06894_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29463_ ( .A(main_fsm[27:24]), .Y(_06895_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _29464_ ( .A({ main_fsm[0], main_fsm[1], main_fsm[2], main_fsm[3] }), .Y(_06896_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29465_ ( .A({ _06897_, _06886_ }), .Y(_05729_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29466_ ( .A({ main_fsm[0], main_fsm[2:1], main_fsm[3] }), .Y(_06897_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _29467_ ( .A({ main_fsm[4], _06900_, _06898_, _06891_ }), .Y(_05730_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29468_ ( .A({ main_fsm[5], _06899_, _06889_, _06888_ }), .Y(_06898_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _29469_ ( .A({ main_fsm[6], main_fsm[7] }), .Y(_06899_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _29470_ ( .A({ main_fsm[0], main_fsm[2:1], main_fsm[3] }), .Y(_06900_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29471_ ( .A({ _06902_, _06901_ }), .Y(_05731_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29472_ ( .A({ main_fsm[4], _06898_, _06891_ }), .Y(_06901_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29473_ ( .A({ main_fsm[2], main_fsm[0], main_fsm[1], main_fsm[3] }), .Y(_06902_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _29474_ ( .A({ main_fsm[4], _06897_, _06898_, _06891_ }), .Y(_05732_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29475_ ( .A({ _06904_, _06903_ }), .Y(_05733_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29476_ ( .A({ _06891_, _06898_, main_fsm[4] }), .Y(_06903_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _29477_ ( .A({ main_fsm[0], main_fsm[2], main_fsm[3], main_fsm[1] }), .Y(_06904_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29478_ ( .A({ _06891_, _06905_, _06898_, main_fsm[4] }), .Y(_05734_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _29479_ ( .A({ main_fsm[1], main_fsm[2], main_fsm[0], main_fsm[3] }), .Y(_06905_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29480_ ( .A({ _06896_, _06903_ }), .Y(_05735_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _29481_ ( .A({ main_fsm[4], _06907_, _06906_, _06891_ }), .Y(_05736_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _29482_ ( .A({ _06888_, _06899_, _06889_, main_fsm[5] }), .Y(_06906_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29483_ ( .A({ main_fsm[0], main_fsm[2:1], main_fsm[3] }), .Y(_06907_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29484_ ( .A({ _06909_, _06908_ }), .Y(_05737_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29485_ ( .A({ main_fsm[4], _06906_, _06891_ }), .Y(_06908_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _29486_ ( .A({ main_fsm[3:2], main_fsm[0], main_fsm[1] }), .Y(_06909_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29487_ ( .A({ _06910_, _06908_ }), .Y(_05738_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _29488_ ( .A({ main_fsm[0], main_fsm[2:1], main_fsm[3] }), .Y(_06910_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _29489_ ( .A({ main_fsm[4], _06911_, _06906_, _06891_ }), .Y(_05739_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29490_ ( .A({ main_fsm[1:0], main_fsm[2], main_fsm[3] }), .Y(_06911_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _29491_ ( .A({ _06914_, _06912_, _06891_ }), .Y(_05740_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29492_ ( .A({ _06913_, _06899_, _06889_, _06888_ }), .Y(_06912_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _29493_ ( .A(main_fsm[5:4]), .Y(_06913_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _29494_ ( .A(main_fsm[3:0]), .Y(_06914_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29495_ ( .A({ _06916_, _06915_ }), .Y(_05741_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29496_ ( .A({ _06912_, _06891_ }), .Y(_06915_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _29497_ ( .A({ main_fsm[0], main_fsm[3], main_fsm[1], main_fsm[2] }), .Y(_06916_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _29498_ ( .A({ _06911_, _06912_, _06891_ }), .Y(_05742_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _29499_ ( .A({ _06917_, _06915_ }), .Y(_05743_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29500_ ( .A({ main_fsm[0], main_fsm[2:1], main_fsm[3] }), .Y(_06917_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29501_ ( .A({ _06021_, _06930_ }), .Y(_05514_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _29502_ ( .A({ _06928_, _06923_, _06920_, _06918_ }), .Y(_06021_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29503_ ( .A({ control_conv2d_16[1], _06919_, control_conv2d_16[0] }), .Y(_06918_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _29504_ ( .A(control_conv2d_16[3:2]), .Y(_06919_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29505_ ( .A({ _06922_, _06921_ }), .Y(_06920_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29506_ ( .A(control_conv2d_16[15:12]), .Y(_06921_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29507_ ( .A(control_conv2d_16[11:8]), .Y(_06922_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29508_ ( .A({ _06927_, _06926_, _06925_, _06924_ }), .Y(_06923_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29509_ ( .A(control_conv2d_16[23:20]), .Y(_06924_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29510_ ( .A(control_conv2d_16[19:16]), .Y(_06925_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29511_ ( .A(control_conv2d_16[31:28]), .Y(_06926_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29512_ ( .A(control_conv2d_16[27:24]), .Y(_06927_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29513_ ( .A({ _06929_, control_conv2d_16[4] }), .Y(_06928_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _29514_ ( .A(control_conv2d_16[7:5]), .Y(_06929_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29515_ ( .A({ _06933_, _06931_, _06923_, _06920_ }), .Y(_06930_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29516_ ( .A({ control_conv2d_16[4], _06932_ }), .Y(_06931_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29517_ ( .A({ control_conv2d_16[5], control_conv2d_16[7:6] }), .Y(_06932_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _29518_ ( .A({ control_conv2d_16[2], control_conv2d_16[0], control_conv2d_16[1], control_conv2d_16[3] }), .Y(_06933_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29519_ ( .A({ _05959_, _06934_ }), .Y(_24054_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29520_ ( .A({ _06935_, _06940_, _stream_conv2d_16_source_32_source_pat_fsm_15[0] }), .Y(_06934_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29521_ ( .A({ _06939_, _06938_, _06936_ }), .Y(_06935_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29522_ ( .A({ _06937_, _stream_conv2d_16_source_32_source_pat_fsm_15[3:2] }), .Y(_06936_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29523_ ( .A(_stream_conv2d_16_source_32_source_pat_fsm_15[7:4]), .Y(_06937_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29524_ ( .A(_stream_conv2d_16_source_32_source_pat_fsm_15[15:12]), .Y(_06938_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29525_ ( .A(_stream_conv2d_16_source_32_source_pat_fsm_15[11:8]), .Y(_06939_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29526_ ( .A({ _06944_, _06943_, _06942_, _06941_ }), .Y(_06940_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29527_ ( .A(_stream_conv2d_16_source_32_source_pat_fsm_15[23:20]), .Y(_06941_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29528_ ( .A(_stream_conv2d_16_source_32_source_pat_fsm_15[19:16]), .Y(_06942_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29529_ ( .A(_stream_conv2d_16_source_32_source_pat_fsm_15[31:28]), .Y(_06943_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29530_ ( .A(_stream_conv2d_16_source_32_source_pat_fsm_15[27:24]), .Y(_06944_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29531_ ( .A({ _06935_, _stream_conv2d_16_source_32_source_pat_fsm_15[0], _06940_, _stream_conv2d_16_source_32_source_pat_fsm_15[1] }), .Y(_05959_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29532_ ( .A({ _17775_, _06945_, _17743_, _05959_ }), .Y(_17711_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29533_ ( .A({ _06934_, _stream_conv2d_16_source_32_source_pat_fsm_15[1] }), .Y(_06945_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29534_ ( .A({ _17786_, _06945_, _17754_, _05959_ }), .Y(_17722_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29535_ ( .A({ _17797_, _06945_, _17765_, _05959_ }), .Y(_17733_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29536_ ( .A({ _17800_, _06945_, _17768_, _05959_ }), .Y(_17736_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29537_ ( .A({ _17801_, _06945_, _17769_, _05959_ }), .Y(_17737_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29538_ ( .A({ _17802_, _06945_, _17770_, _05959_ }), .Y(_17738_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29539_ ( .A({ _17803_, _06945_, _17771_, _05959_ }), .Y(_17739_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29540_ ( .A({ _17804_, _06945_, _17772_, _05959_ }), .Y(_17740_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29541_ ( .A({ _17805_, _06945_, _17773_, _05959_ }), .Y(_17741_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29542_ ( .A({ _17806_, _06945_, _17774_, _05959_ }), .Y(_17742_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29543_ ( .A({ _17776_, _06945_, _17744_, _05959_ }), .Y(_17712_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29544_ ( .A({ _17777_, _06945_, _17745_, _05959_ }), .Y(_17713_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29545_ ( .A({ _17778_, _06945_, _17746_, _05959_ }), .Y(_17714_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29546_ ( .A({ _17779_, _06945_, _17747_, _05959_ }), .Y(_17715_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29547_ ( .A({ _17780_, _06945_, _17748_, _05959_ }), .Y(_17716_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29548_ ( .A({ _17781_, _06945_, _17749_, _05959_ }), .Y(_17717_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29549_ ( .A({ _17782_, _06945_, _17750_, _05959_ }), .Y(_17718_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29550_ ( .A({ _17783_, _06945_, _17751_, _05959_ }), .Y(_17719_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29551_ ( .A({ _17784_, _06945_, _17752_, _05959_ }), .Y(_17720_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29552_ ( .A({ _17785_, _06945_, _17753_, _05959_ }), .Y(_17721_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29553_ ( .A({ _17787_, _06945_, _17755_, _05959_ }), .Y(_17723_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29554_ ( .A({ _17788_, _06945_, _17756_, _05959_ }), .Y(_17724_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29555_ ( .A({ _17789_, _06945_, _17757_, _05959_ }), .Y(_17725_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29556_ ( .A({ _17790_, _06945_, _17758_, _05959_ }), .Y(_17726_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29557_ ( .A({ _17791_, _06945_, _17759_, _05959_ }), .Y(_17727_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29558_ ( .A({ _17792_, _06945_, _17760_, _05959_ }), .Y(_17728_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29559_ ( .A({ _17793_, _06945_, _17761_, _05959_ }), .Y(_17729_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29560_ ( .A({ _17794_, _06945_, _17762_, _05959_ }), .Y(_17730_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29561_ ( .A({ _17795_, _06945_, _17763_, _05959_ }), .Y(_17731_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29562_ ( .A({ _17796_, _06945_, _17764_, _05959_ }), .Y(_17732_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29563_ ( .A({ _17798_, _06945_, _17766_, _05959_ }), .Y(_17734_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29564_ ( .A({ _17799_, _06945_, _17767_, _05959_ }), .Y(_17735_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29565_ ( .A({ _05956_, _06946_ }), .Y(_24053_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29566_ ( .A({ _06947_, _06952_, _stream_conv2d_16_source_33_source_pat_fsm_16[0] }), .Y(_06946_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29567_ ( .A({ _06951_, _06950_, _06948_ }), .Y(_06947_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29568_ ( .A({ _06949_, _stream_conv2d_16_source_33_source_pat_fsm_16[3:2] }), .Y(_06948_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29569_ ( .A(_stream_conv2d_16_source_33_source_pat_fsm_16[7:4]), .Y(_06949_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29570_ ( .A(_stream_conv2d_16_source_33_source_pat_fsm_16[15:12]), .Y(_06950_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29571_ ( .A(_stream_conv2d_16_source_33_source_pat_fsm_16[11:8]), .Y(_06951_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29572_ ( .A({ _06956_, _06955_, _06954_, _06953_ }), .Y(_06952_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29573_ ( .A(_stream_conv2d_16_source_33_source_pat_fsm_16[23:20]), .Y(_06953_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29574_ ( .A(_stream_conv2d_16_source_33_source_pat_fsm_16[19:16]), .Y(_06954_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29575_ ( .A(_stream_conv2d_16_source_33_source_pat_fsm_16[31:28]), .Y(_06955_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29576_ ( .A(_stream_conv2d_16_source_33_source_pat_fsm_16[27:24]), .Y(_06956_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29577_ ( .A({ _06947_, _stream_conv2d_16_source_33_source_pat_fsm_16[0], _06952_, _stream_conv2d_16_source_33_source_pat_fsm_16[1] }), .Y(_05956_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29578_ ( .A({ _17679_, _06957_, _17647_, _05956_ }), .Y(_17615_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29579_ ( .A({ _06946_, _stream_conv2d_16_source_33_source_pat_fsm_16[1] }), .Y(_06957_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29580_ ( .A({ _17690_, _06957_, _17658_, _05956_ }), .Y(_17626_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29581_ ( .A({ _17701_, _06957_, _17669_, _05956_ }), .Y(_17637_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29582_ ( .A({ _17704_, _06957_, _17672_, _05956_ }), .Y(_17640_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29583_ ( .A({ _17705_, _06957_, _17673_, _05956_ }), .Y(_17641_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29584_ ( .A({ _17706_, _06957_, _17674_, _05956_ }), .Y(_17642_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29585_ ( .A({ _17707_, _06957_, _17675_, _05956_ }), .Y(_17643_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29586_ ( .A({ _17708_, _06957_, _17676_, _05956_ }), .Y(_17644_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29587_ ( .A({ _17709_, _06957_, _17677_, _05956_ }), .Y(_17645_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29588_ ( .A({ _17710_, _06957_, _17678_, _05956_ }), .Y(_17646_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29589_ ( .A({ _17680_, _06957_, _17648_, _05956_ }), .Y(_17616_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29590_ ( .A({ _17681_, _06957_, _17649_, _05956_ }), .Y(_17617_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29591_ ( .A({ _17682_, _06957_, _17650_, _05956_ }), .Y(_17618_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29592_ ( .A({ _17683_, _06957_, _17651_, _05956_ }), .Y(_17619_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29593_ ( .A({ _17684_, _06957_, _17652_, _05956_ }), .Y(_17620_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29594_ ( .A({ _17685_, _06957_, _17653_, _05956_ }), .Y(_17621_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29595_ ( .A({ _17686_, _06957_, _17654_, _05956_ }), .Y(_17622_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29596_ ( .A({ _17687_, _06957_, _17655_, _05956_ }), .Y(_17623_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29597_ ( .A({ _17688_, _06957_, _17656_, _05956_ }), .Y(_17624_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29598_ ( .A({ _17689_, _06957_, _17657_, _05956_ }), .Y(_17625_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29599_ ( .A({ _17691_, _06957_, _17659_, _05956_ }), .Y(_17627_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29600_ ( .A({ _17692_, _06957_, _17660_, _05956_ }), .Y(_17628_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29601_ ( .A({ _17693_, _06957_, _17661_, _05956_ }), .Y(_17629_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29602_ ( .A({ _17694_, _06957_, _17662_, _05956_ }), .Y(_17630_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29603_ ( .A({ _17695_, _06957_, _17663_, _05956_ }), .Y(_17631_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29604_ ( .A({ _17696_, _06957_, _17664_, _05956_ }), .Y(_17632_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29605_ ( .A({ _17697_, _06957_, _17665_, _05956_ }), .Y(_17633_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29606_ ( .A({ _17698_, _06957_, _17666_, _05956_ }), .Y(_17634_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29607_ ( .A({ _17699_, _06957_, _17667_, _05956_ }), .Y(_17635_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29608_ ( .A({ _17700_, _06957_, _17668_, _05956_ }), .Y(_17636_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29609_ ( .A({ _17702_, _06957_, _17670_, _05956_ }), .Y(_17638_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29610_ ( .A({ _17703_, _06957_, _17671_, _05956_ }), .Y(_17639_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29611_ ( .A({ _05954_, _06958_ }), .Y(_24052_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29612_ ( .A({ _06959_, _06964_, _stream_conv2d_16_source_34_source_pat_fsm_17[0] }), .Y(_06958_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29613_ ( .A({ _06963_, _06962_, _06960_ }), .Y(_06959_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29614_ ( .A({ _06961_, _stream_conv2d_16_source_34_source_pat_fsm_17[3:2] }), .Y(_06960_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29615_ ( .A(_stream_conv2d_16_source_34_source_pat_fsm_17[7:4]), .Y(_06961_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29616_ ( .A(_stream_conv2d_16_source_34_source_pat_fsm_17[15:12]), .Y(_06962_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29617_ ( .A(_stream_conv2d_16_source_34_source_pat_fsm_17[11:8]), .Y(_06963_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29618_ ( .A({ _06968_, _06967_, _06966_, _06965_ }), .Y(_06964_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29619_ ( .A(_stream_conv2d_16_source_34_source_pat_fsm_17[23:20]), .Y(_06965_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29620_ ( .A(_stream_conv2d_16_source_34_source_pat_fsm_17[19:16]), .Y(_06966_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29621_ ( .A(_stream_conv2d_16_source_34_source_pat_fsm_17[31:28]), .Y(_06967_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29622_ ( .A(_stream_conv2d_16_source_34_source_pat_fsm_17[27:24]), .Y(_06968_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29623_ ( .A({ _06959_, _stream_conv2d_16_source_34_source_pat_fsm_17[0], _06964_, _stream_conv2d_16_source_34_source_pat_fsm_17[1] }), .Y(_05954_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29624_ ( .A({ _17583_, _06969_, _17551_, _05954_ }), .Y(_17519_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29625_ ( .A({ _06958_, _stream_conv2d_16_source_34_source_pat_fsm_17[1] }), .Y(_06969_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29626_ ( .A({ _17594_, _06969_, _17562_, _05954_ }), .Y(_17530_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29627_ ( .A({ _17605_, _06969_, _17573_, _05954_ }), .Y(_17541_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29628_ ( .A({ _17608_, _06969_, _17576_, _05954_ }), .Y(_17544_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29629_ ( .A({ _17609_, _06969_, _17577_, _05954_ }), .Y(_17545_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29630_ ( .A({ _17610_, _06969_, _17578_, _05954_ }), .Y(_17546_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29631_ ( .A({ _17611_, _06969_, _17579_, _05954_ }), .Y(_17547_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29632_ ( .A({ _17612_, _06969_, _17580_, _05954_ }), .Y(_17548_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29633_ ( .A({ _17613_, _06969_, _17581_, _05954_ }), .Y(_17549_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29634_ ( .A({ _17614_, _06969_, _17582_, _05954_ }), .Y(_17550_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29635_ ( .A({ _17584_, _06969_, _17552_, _05954_ }), .Y(_17520_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29636_ ( .A({ _17585_, _06969_, _17553_, _05954_ }), .Y(_17521_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29637_ ( .A({ _17586_, _06969_, _17554_, _05954_ }), .Y(_17522_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29638_ ( .A({ _17587_, _06969_, _17555_, _05954_ }), .Y(_17523_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29639_ ( .A({ _17588_, _06969_, _17556_, _05954_ }), .Y(_17524_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29640_ ( .A({ _17589_, _06969_, _17557_, _05954_ }), .Y(_17525_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29641_ ( .A({ _17590_, _06969_, _17558_, _05954_ }), .Y(_17526_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29642_ ( .A({ _17591_, _06969_, _17559_, _05954_ }), .Y(_17527_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29643_ ( .A({ _17592_, _06969_, _17560_, _05954_ }), .Y(_17528_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29644_ ( .A({ _17593_, _06969_, _17561_, _05954_ }), .Y(_17529_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29645_ ( .A({ _17595_, _06969_, _17563_, _05954_ }), .Y(_17531_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29646_ ( .A({ _17596_, _06969_, _17564_, _05954_ }), .Y(_17532_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29647_ ( .A({ _17597_, _06969_, _17565_, _05954_ }), .Y(_17533_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29648_ ( .A({ _17598_, _06969_, _17566_, _05954_ }), .Y(_17534_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29649_ ( .A({ _17599_, _06969_, _17567_, _05954_ }), .Y(_17535_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29650_ ( .A({ _17600_, _06969_, _17568_, _05954_ }), .Y(_17536_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29651_ ( .A({ _17601_, _06969_, _17569_, _05954_ }), .Y(_17537_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29652_ ( .A({ _17602_, _06969_, _17570_, _05954_ }), .Y(_17538_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29653_ ( .A({ _17603_, _06969_, _17571_, _05954_ }), .Y(_17539_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29654_ ( .A({ _17604_, _06969_, _17572_, _05954_ }), .Y(_17540_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29655_ ( .A({ _17606_, _06969_, _17574_, _05954_ }), .Y(_17542_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29656_ ( .A({ _17607_, _06969_, _17575_, _05954_ }), .Y(_17543_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29657_ ( .A({ _05949_, _06970_ }), .Y(_24050_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29658_ ( .A({ _06979_, _06976_, _06971_ }), .Y(_06970_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29659_ ( .A({ _06975_, _06974_, _06973_, _06972_ }), .Y(_06971_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29660_ ( .A(_stream_conv2d_16_source_36_source_pat_fsm_19[23:20]), .Y(_06972_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29661_ ( .A(_stream_conv2d_16_source_36_source_pat_fsm_19[19:16]), .Y(_06973_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29662_ ( .A(_stream_conv2d_16_source_36_source_pat_fsm_19[31:28]), .Y(_06974_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29663_ ( .A(_stream_conv2d_16_source_36_source_pat_fsm_19[27:24]), .Y(_06975_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29664_ ( .A({ _06978_, _06977_ }), .Y(_06976_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29665_ ( .A(_stream_conv2d_16_source_36_source_pat_fsm_19[15:12]), .Y(_06977_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29666_ ( .A(_stream_conv2d_16_source_36_source_pat_fsm_19[11:8]), .Y(_06978_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29667_ ( .A({ _06980_, _stream_conv2d_16_source_36_source_pat_fsm_19[3:2], _stream_conv2d_16_source_36_source_pat_fsm_19[0] }), .Y(_06979_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29668_ ( .A(_stream_conv2d_16_source_36_source_pat_fsm_19[7:4]), .Y(_06980_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _29669_ ( .A({ _06981_, _06980_, _06976_, _06971_ }), .Y(_05949_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29670_ ( .A({ _stream_conv2d_16_source_36_source_pat_fsm_19[0], _stream_conv2d_16_source_36_source_pat_fsm_19[3:1] }), .Y(_06981_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29671_ ( .A({ _17391_, _06982_, _17359_, _05949_ }), .Y(_17327_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29672_ ( .A({ _06970_, _stream_conv2d_16_source_36_source_pat_fsm_19[1] }), .Y(_06982_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29673_ ( .A({ _17402_, _06982_, _17370_, _05949_ }), .Y(_17338_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29674_ ( .A({ _17413_, _06982_, _17381_, _05949_ }), .Y(_17349_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29675_ ( .A({ _17416_, _06982_, _17384_, _05949_ }), .Y(_17352_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29676_ ( .A({ _17417_, _06982_, _17385_, _05949_ }), .Y(_17353_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29677_ ( .A({ _17418_, _06982_, _17386_, _05949_ }), .Y(_17354_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29678_ ( .A({ _17419_, _06982_, _17387_, _05949_ }), .Y(_17355_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29679_ ( .A({ _17420_, _06982_, _17388_, _05949_ }), .Y(_17356_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29680_ ( .A({ _17421_, _06982_, _17389_, _05949_ }), .Y(_17357_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29681_ ( .A({ _17422_, _06982_, _17390_, _05949_ }), .Y(_17358_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29682_ ( .A({ _17392_, _06982_, _17360_, _05949_ }), .Y(_17328_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29683_ ( .A({ _17393_, _06982_, _17361_, _05949_ }), .Y(_17329_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29684_ ( .A({ _17394_, _06982_, _17362_, _05949_ }), .Y(_17330_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29685_ ( .A({ _17395_, _06982_, _17363_, _05949_ }), .Y(_17331_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29686_ ( .A({ _17396_, _06982_, _17364_, _05949_ }), .Y(_17332_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29687_ ( .A({ _17397_, _06982_, _17365_, _05949_ }), .Y(_17333_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29688_ ( .A({ _17398_, _06982_, _17366_, _05949_ }), .Y(_17334_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29689_ ( .A({ _17399_, _06982_, _17367_, _05949_ }), .Y(_17335_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29690_ ( .A({ _17400_, _06982_, _17368_, _05949_ }), .Y(_17336_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29691_ ( .A({ _17401_, _06982_, _17369_, _05949_ }), .Y(_17337_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29692_ ( .A({ _17403_, _06982_, _17371_, _05949_ }), .Y(_17339_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29693_ ( .A({ _17404_, _06982_, _17372_, _05949_ }), .Y(_17340_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29694_ ( .A({ _17405_, _06982_, _17373_, _05949_ }), .Y(_17341_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29695_ ( .A({ _17406_, _06982_, _17374_, _05949_ }), .Y(_17342_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29696_ ( .A({ _17407_, _06982_, _17375_, _05949_ }), .Y(_17343_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29697_ ( .A({ _17408_, _06982_, _17376_, _05949_ }), .Y(_17344_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29698_ ( .A({ _17409_, _06982_, _17377_, _05949_ }), .Y(_17345_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29699_ ( .A({ _17410_, _06982_, _17378_, _05949_ }), .Y(_17346_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29700_ ( .A({ _17411_, _06982_, _17379_, _05949_ }), .Y(_17347_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29701_ ( .A({ _17412_, _06982_, _17380_, _05949_ }), .Y(_17348_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29702_ ( .A({ _17414_, _06982_, _17382_, _05949_ }), .Y(_17350_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29703_ ( .A({ _17415_, _06982_, _17383_, _05949_ }), .Y(_17351_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29704_ ( .A({ _05952_, _06983_ }), .Y(_24051_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29705_ ( .A({ _06984_, _06989_, _stream_conv2d_16_source_35_source_pat_fsm_18[0] }), .Y(_06983_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29706_ ( .A({ _06988_, _06987_, _06985_ }), .Y(_06984_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29707_ ( .A({ _06986_, _stream_conv2d_16_source_35_source_pat_fsm_18[3:2] }), .Y(_06985_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29708_ ( .A(_stream_conv2d_16_source_35_source_pat_fsm_18[7:4]), .Y(_06986_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29709_ ( .A(_stream_conv2d_16_source_35_source_pat_fsm_18[15:12]), .Y(_06987_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29710_ ( .A(_stream_conv2d_16_source_35_source_pat_fsm_18[11:8]), .Y(_06988_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29711_ ( .A({ _06993_, _06992_, _06991_, _06990_ }), .Y(_06989_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29712_ ( .A(_stream_conv2d_16_source_35_source_pat_fsm_18[23:20]), .Y(_06990_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29713_ ( .A(_stream_conv2d_16_source_35_source_pat_fsm_18[19:16]), .Y(_06991_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29714_ ( .A(_stream_conv2d_16_source_35_source_pat_fsm_18[31:28]), .Y(_06992_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29715_ ( .A(_stream_conv2d_16_source_35_source_pat_fsm_18[27:24]), .Y(_06993_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29716_ ( .A({ _06984_, _stream_conv2d_16_source_35_source_pat_fsm_18[0], _06989_, _stream_conv2d_16_source_35_source_pat_fsm_18[1] }), .Y(_05952_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29717_ ( .A({ _17487_, _06994_, _17455_, _05952_ }), .Y(_17423_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _29718_ ( .A({ _06983_, _stream_conv2d_16_source_35_source_pat_fsm_18[1] }), .Y(_06994_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29719_ ( .A({ _17498_, _06994_, _17466_, _05952_ }), .Y(_17434_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29720_ ( .A({ _17509_, _06994_, _17477_, _05952_ }), .Y(_17445_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29721_ ( .A({ _17512_, _06994_, _17480_, _05952_ }), .Y(_17448_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29722_ ( .A({ _17513_, _06994_, _17481_, _05952_ }), .Y(_17449_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29723_ ( .A({ _17514_, _06994_, _17482_, _05952_ }), .Y(_17450_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29724_ ( .A({ _17515_, _06994_, _17483_, _05952_ }), .Y(_17451_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29725_ ( .A({ _17516_, _06994_, _17484_, _05952_ }), .Y(_17452_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29726_ ( .A({ _17517_, _06994_, _17485_, _05952_ }), .Y(_17453_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29727_ ( .A({ _17518_, _06994_, _17486_, _05952_ }), .Y(_17454_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29728_ ( .A({ _17488_, _06994_, _17456_, _05952_ }), .Y(_17424_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29729_ ( .A({ _17489_, _06994_, _17457_, _05952_ }), .Y(_17425_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29730_ ( .A({ _17490_, _06994_, _17458_, _05952_ }), .Y(_17426_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29731_ ( .A({ _17491_, _06994_, _17459_, _05952_ }), .Y(_17427_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29732_ ( .A({ _17492_, _06994_, _17460_, _05952_ }), .Y(_17428_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29733_ ( .A({ _17493_, _06994_, _17461_, _05952_ }), .Y(_17429_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29734_ ( .A({ _17494_, _06994_, _17462_, _05952_ }), .Y(_17430_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29735_ ( .A({ _17495_, _06994_, _17463_, _05952_ }), .Y(_17431_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29736_ ( .A({ _17496_, _06994_, _17464_, _05952_ }), .Y(_17432_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29737_ ( .A({ _17497_, _06994_, _17465_, _05952_ }), .Y(_17433_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29738_ ( .A({ _17499_, _06994_, _17467_, _05952_ }), .Y(_17435_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29739_ ( .A({ _17500_, _06994_, _17468_, _05952_ }), .Y(_17436_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29740_ ( .A({ _17501_, _06994_, _17469_, _05952_ }), .Y(_17437_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29741_ ( .A({ _17502_, _06994_, _17470_, _05952_ }), .Y(_17438_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29742_ ( .A({ _17503_, _06994_, _17471_, _05952_ }), .Y(_17439_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29743_ ( .A({ _17504_, _06994_, _17472_, _05952_ }), .Y(_17440_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29744_ ( .A({ _17505_, _06994_, _17473_, _05952_ }), .Y(_17441_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29745_ ( .A({ _17506_, _06994_, _17474_, _05952_ }), .Y(_17442_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29746_ ( .A({ _17507_, _06994_, _17475_, _05952_ }), .Y(_17443_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29747_ ( .A({ _17508_, _06994_, _17476_, _05952_ }), .Y(_17444_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29748_ ( .A({ _17510_, _06994_, _17478_, _05952_ }), .Y(_17446_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29749_ ( .A({ _17511_, _06994_, _17479_, _05952_ }), .Y(_17447_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29750_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18247_, _18279_ }), .Y(_18215_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29751_ ( .A({ _06996_, _07004_, _stream_conv2d_16_source_27_source_pat_fsm_10[1] }), .Y(_06995_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29752_ ( .A({ _07003_, _07002_, _06997_ }), .Y(_06996_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29753_ ( .A({ _07001_, _07000_, _06999_, _06998_ }), .Y(_06997_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29754_ ( .A(_stream_conv2d_16_source_27_source_pat_fsm_10[23:20]), .Y(_06998_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29755_ ( .A(_stream_conv2d_16_source_27_source_pat_fsm_10[19:16]), .Y(_06999_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29756_ ( .A(_stream_conv2d_16_source_27_source_pat_fsm_10[31:28]), .Y(_07000_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29757_ ( .A(_stream_conv2d_16_source_27_source_pat_fsm_10[27:24]), .Y(_07001_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29758_ ( .A(_stream_conv2d_16_source_27_source_pat_fsm_10[15:12]), .Y(_07002_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29759_ ( .A(_stream_conv2d_16_source_27_source_pat_fsm_10[11:8]), .Y(_07003_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29760_ ( .A({ _07005_, _stream_conv2d_16_source_27_source_pat_fsm_10[3:2] }), .Y(_07004_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29761_ ( .A(_stream_conv2d_16_source_27_source_pat_fsm_10[7:4]), .Y(_07005_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29762_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18246_, _18278_ }), .Y(_18214_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29763_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18244_, _18276_ }), .Y(_18212_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29764_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18243_, _18275_ }), .Y(_18211_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29765_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18242_, _18274_ }), .Y(_18210_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29766_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18241_, _18273_ }), .Y(_18209_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29767_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18240_, _18272_ }), .Y(_18208_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29768_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18239_, _18271_ }), .Y(_18207_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29769_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18238_, _18270_ }), .Y(_18206_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29770_ ( .A({ _07014_, _07006_ }), .Y(_24049_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29771_ ( .A({ _07013_, _07012_, _07009_, _07007_ }), .Y(_07006_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29772_ ( .A({ _07008_, _stream_conv2d_16_sink_37_sink_fsm_20[31:29] }), .Y(_07007_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29773_ ( .A({ _stream_conv2d_16_sink_37_sink_fsm_20[27:26], _stream_conv2d_16_sink_37_sink_fsm_20[24], _stream_conv2d_16_sink_37_sink_fsm_20[21] }), .Y(_07008_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _29774_ ( .A({ _07011_, _07010_, _stream_conv2d_16_sink_37_sink_fsm_20[11:10] }), .Y(_07009_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29775_ ( .A({ _stream_conv2d_16_sink_37_sink_fsm_20[28], _stream_conv2d_16_sink_37_sink_fsm_20[25], _stream_conv2d_16_sink_37_sink_fsm_20[23:22] }), .Y(_07010_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29776_ ( .A({ _stream_conv2d_16_sink_37_sink_fsm_20[19:18], _stream_conv2d_16_sink_37_sink_fsm_20[16], _stream_conv2d_16_sink_37_sink_fsm_20[13] }), .Y(_07011_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29777_ ( .A({ _stream_conv2d_16_sink_37_sink_fsm_20[12], _stream_conv2d_16_sink_37_sink_fsm_20[9:8], _stream_conv2d_16_sink_37_sink_fsm_20[1] }), .Y(_07012_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29778_ ( .A({ _stream_conv2d_16_sink_37_sink_fsm_20[20], _stream_conv2d_16_sink_37_sink_fsm_20[17], _stream_conv2d_16_sink_37_sink_fsm_20[15:14] }), .Y(_07013_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29779_ ( .A({ _07015_, _stream_conv2d_16_sink_37_sink_fsm_20[6:5] }), .Y(_07014_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29780_ ( .A({ _stream_conv2d_16_sink_37_sink_fsm_20[7], _stream_conv2d_16_sink_37_sink_fsm_20[4:2] }), .Y(_07015_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29781_ ( .A({ _17231_, _07016_, _17295_, _07017_ }), .Y(_17263_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29782_ ( .A({ _stream_conv2d_16_sink_37_sink_fsm_20[0], _24049_ }), .Y(_07016_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29783_ ( .A({ _07006_, _07014_, _stream_conv2d_16_sink_37_sink_fsm_20[0] }), .Y(_07017_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29784_ ( .A({ _17242_, _07016_, _17306_, _07017_ }), .Y(_17274_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29785_ ( .A({ _17253_, _07016_, _17317_, _07017_ }), .Y(_17285_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29786_ ( .A({ _17256_, _07016_, _17320_, _07017_ }), .Y(_17288_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29787_ ( .A({ _17257_, _07016_, _17321_, _07017_ }), .Y(_17289_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29788_ ( .A({ _17258_, _07016_, _17322_, _07017_ }), .Y(_17290_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29789_ ( .A({ _17259_, _07016_, _17323_, _07017_ }), .Y(_17291_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29790_ ( .A({ _17260_, _07016_, _17324_, _07017_ }), .Y(_17292_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29791_ ( .A({ _17261_, _07016_, _17325_, _07017_ }), .Y(_17293_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29792_ ( .A({ _17262_, _07016_, _17326_, _07017_ }), .Y(_17294_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29793_ ( .A({ _17232_, _07016_, _17296_, _07017_ }), .Y(_17264_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29794_ ( .A({ _17233_, _07016_, _17297_, _07017_ }), .Y(_17265_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29795_ ( .A({ _17234_, _07016_, _17298_, _07017_ }), .Y(_17266_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29796_ ( .A({ _17235_, _07016_, _17299_, _07017_ }), .Y(_17267_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29797_ ( .A({ _17236_, _07016_, _17300_, _07017_ }), .Y(_17268_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29798_ ( .A({ _17237_, _07016_, _17301_, _07017_ }), .Y(_17269_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29799_ ( .A({ _17238_, _07016_, _17302_, _07017_ }), .Y(_17270_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29800_ ( .A({ _17239_, _07016_, _17303_, _07017_ }), .Y(_17271_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29801_ ( .A({ _17240_, _07016_, _17304_, _07017_ }), .Y(_17272_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29802_ ( .A({ _17241_, _07016_, _17305_, _07017_ }), .Y(_17273_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29803_ ( .A({ _17243_, _07016_, _17307_, _07017_ }), .Y(_17275_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29804_ ( .A({ _17244_, _07016_, _17308_, _07017_ }), .Y(_17276_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29805_ ( .A({ _17245_, _07016_, _17309_, _07017_ }), .Y(_17277_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29806_ ( .A({ _17246_, _07016_, _17310_, _07017_ }), .Y(_17278_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29807_ ( .A({ _17247_, _07016_, _17311_, _07017_ }), .Y(_17279_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29808_ ( .A({ _17248_, _07016_, _17312_, _07017_ }), .Y(_17280_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29809_ ( .A({ _17249_, _07016_, _17313_, _07017_ }), .Y(_17281_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29810_ ( .A({ _17250_, _07016_, _17314_, _07017_ }), .Y(_17282_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29811_ ( .A({ _17251_, _07016_, _17315_, _07017_ }), .Y(_17283_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29812_ ( .A({ _17252_, _07016_, _17316_, _07017_ }), .Y(_17284_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29813_ ( .A({ _17254_, _07016_, _17318_, _07017_ }), .Y(_17286_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29814_ ( .A({ _17255_, _07016_, _17319_, _07017_ }), .Y(_17287_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29815_ ( .A({ _05948_, _07018_ }), .Y(_05516_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _29816_ ( .A({ _07027_, _07019_, _maxi_write_fsm[0], _maxi_write_fsm[1] }), .Y(_07018_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _29817_ ( .A({ _07026_, _07025_, _07020_ }), .Y(_07019_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29818_ ( .A({ _07024_, _07023_, _07022_, _07021_ }), .Y(_07020_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29819_ ( .A(_maxi_write_fsm[23:20]), .Y(_07021_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29820_ ( .A(_maxi_write_fsm[19:16]), .Y(_07022_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29821_ ( .A(_maxi_write_fsm[31:28]), .Y(_07023_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29822_ ( .A(_maxi_write_fsm[27:24]), .Y(_07024_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29823_ ( .A(_maxi_write_fsm[15:12]), .Y(_07025_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29824_ ( .A(_maxi_write_fsm[11:8]), .Y(_07026_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _29825_ ( .A({ _07028_, _maxi_write_fsm[2], _maxi_write_fsm[3] }), .Y(_07027_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _29826_ ( .A(_maxi_write_fsm[7:4]), .Y(_07028_) );
  \$lut  #( .LUT(16'hefff), .WIDTH(4) ) _29827_ ( .A({ _07029_, _07019_, _maxi_write_fsm[2], _maxi_write_fsm[3] }), .Y(_05948_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29828_ ( .A({ _maxi_write_fsm[0], _07028_, _maxi_write_fsm[1] }), .Y(_07029_) );
  \$lut  #( .LUT(16'hfeff), .WIDTH(4) ) _29829_ ( .A({ _05947_, _07033_, _07031_, _24047_ }), .Y(_24048_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _29830_ ( .A({ _07030_, _07018_ }), .Y(_24047_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29831_ ( .A({ _maxi_write_fsm[0], _maxi_write_fsm[1], _07027_, _07019_ }), .Y(_07030_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29832_ ( .A({ _07019_, _07029_, _maxi_write_fsm[3] }), .Y(_07031_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _29833_ ( .A({ _07032_, _07028_, _07019_ }), .Y(_05947_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29834_ ( .A({ _maxi_write_fsm[2], _maxi_write_fsm[0], _maxi_write_fsm[1], _maxi_write_fsm[3] }), .Y(_07032_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _29835_ ( .A({ _07019_, _maxi_write_fsm[1], _07027_, _maxi_write_fsm[0] }), .Y(_07033_) );
  \$lut  #( .LUT(16'h8fff), .WIDTH(4) ) _29836_ ( .A({ _07034_, _05947_, _07018_, _17199_ }), .Y(_17103_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29837_ ( .A({ _17135_, _07030_, _17167_, _07033_ }), .Y(_07034_) );
  \$lut  #( .LUT(16'h8fff), .WIDTH(4) ) _29838_ ( .A({ _05948_, _07035_, _07030_, _17146_ }), .Y(_17114_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29839_ ( .A({ _17210_, _07018_, _07033_, _17178_ }), .Y(_07035_) );
  \$lut  #( .LUT(16'h8fff), .WIDTH(4) ) _29840_ ( .A({ _07036_, _05947_, _07018_, _17221_ }), .Y(_17125_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29841_ ( .A({ _17157_, _07030_, _17189_, _07033_ }), .Y(_07036_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29842_ ( .A({ _07037_, _17160_, _07030_ }), .Y(_17128_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29843_ ( .A({ _17224_, _07018_, _07033_, _17192_ }), .Y(_07037_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29844_ ( .A({ _07038_, _17161_, _07030_ }), .Y(_17129_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29845_ ( .A({ _17225_, _07018_, _07033_, _17193_ }), .Y(_07038_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29846_ ( .A({ _07039_, _17162_, _07030_ }), .Y(_17130_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29847_ ( .A({ _17226_, _07018_, _07033_, _17194_ }), .Y(_07039_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29848_ ( .A({ _07040_, _17163_, _07030_ }), .Y(_17131_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29849_ ( .A({ _17227_, _07018_, _07033_, _17195_ }), .Y(_07040_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29850_ ( .A({ _07041_, _17164_, _07030_ }), .Y(_17132_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29851_ ( .A({ _17228_, _07018_, _07033_, _17196_ }), .Y(_07041_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29852_ ( .A({ _07042_, _17197_, _07033_ }), .Y(_17133_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29853_ ( .A({ _17229_, _07018_, _07030_, _17165_ }), .Y(_07042_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29854_ ( .A({ _07043_, _17198_, _07033_ }), .Y(_17134_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29855_ ( .A({ _17230_, _07018_, _07030_, _17166_ }), .Y(_07043_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29856_ ( .A({ _07044_, _17136_, _07030_ }), .Y(_17104_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29857_ ( .A({ _17200_, _07018_, _07033_, _17168_ }), .Y(_07044_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29858_ ( .A({ _07045_, _17169_, _07033_ }), .Y(_17105_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29859_ ( .A({ _17201_, _07018_, _07030_, _17137_ }), .Y(_07045_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29860_ ( .A({ _07046_, _17170_, _07033_ }), .Y(_17106_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29861_ ( .A({ _17202_, _07018_, _07030_, _17138_ }), .Y(_07046_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29862_ ( .A({ _07047_, _17139_, _07030_ }), .Y(_17107_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29863_ ( .A({ _17203_, _07018_, _07033_, _17171_ }), .Y(_07047_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29864_ ( .A({ _07048_, _17172_, _07033_ }), .Y(_17108_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29865_ ( .A({ _17204_, _07018_, _07030_, _17140_ }), .Y(_07048_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29866_ ( .A({ _07049_, _17173_, _07033_ }), .Y(_17109_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29867_ ( .A({ _17205_, _07018_, _07030_, _17141_ }), .Y(_07049_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29868_ ( .A({ _07050_, _17142_, _07030_ }), .Y(_17110_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29869_ ( .A({ _17206_, _07018_, _07033_, _17174_ }), .Y(_07050_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29870_ ( .A({ _07051_, _17175_, _07033_ }), .Y(_17111_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29871_ ( .A({ _17207_, _07018_, _07030_, _17143_ }), .Y(_07051_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29872_ ( .A({ _07052_, _17144_, _07030_ }), .Y(_17112_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29873_ ( .A({ _17208_, _07018_, _07033_, _17176_ }), .Y(_07052_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29874_ ( .A({ _07053_, _17145_, _07030_ }), .Y(_17113_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29875_ ( .A({ _17209_, _07018_, _07033_, _17177_ }), .Y(_07053_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29876_ ( .A({ _07054_, _17147_, _07030_ }), .Y(_17115_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29877_ ( .A({ _17211_, _07018_, _07033_, _17179_ }), .Y(_07054_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29878_ ( .A({ _07055_, _17148_, _07030_ }), .Y(_17116_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29879_ ( .A({ _17212_, _07018_, _07033_, _17180_ }), .Y(_07055_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29880_ ( .A({ _07056_, _17149_, _07030_ }), .Y(_17117_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29881_ ( .A({ _17213_, _07018_, _07033_, _17181_ }), .Y(_07056_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29882_ ( .A({ _07057_, _17150_, _07030_ }), .Y(_17118_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29883_ ( .A({ _17214_, _07018_, _07033_, _17182_ }), .Y(_07057_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29884_ ( .A({ _07058_, _17151_, _07030_ }), .Y(_17119_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29885_ ( .A({ _17215_, _07018_, _07033_, _17183_ }), .Y(_07058_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29886_ ( .A({ _07059_, _17152_, _07030_ }), .Y(_17120_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29887_ ( .A({ _17216_, _07018_, _07033_, _17184_ }), .Y(_07059_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29888_ ( .A({ _07060_, _17153_, _07030_ }), .Y(_17121_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29889_ ( .A({ _17217_, _07018_, _07033_, _17185_ }), .Y(_07060_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29890_ ( .A({ _07061_, _17186_, _07033_ }), .Y(_17122_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29891_ ( .A({ _17218_, _07018_, _07030_, _17154_ }), .Y(_07061_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29892_ ( .A({ _07062_, _17187_, _07033_ }), .Y(_17123_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29893_ ( .A({ _17219_, _07018_, _07030_, _17155_ }), .Y(_07062_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29894_ ( .A({ _07063_, _17156_, _07030_ }), .Y(_17124_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29895_ ( .A({ _17220_, _07018_, _07033_, _17188_ }), .Y(_07063_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29896_ ( .A({ _07064_, _17190_, _07033_ }), .Y(_17126_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29897_ ( .A({ _17222_, _07018_, _07030_, _17158_ }), .Y(_07064_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29898_ ( .A({ _07065_, _17191_, _07033_ }), .Y(_17127_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _29899_ ( .A({ _17223_, _07018_, _07030_, _17159_ }), .Y(_07065_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29900_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18237_, _18269_ }), .Y(_18205_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29901_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18236_, _18268_ }), .Y(_18204_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29902_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18235_, _18267_ }), .Y(_18203_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29903_ ( .A({ _17071_, _07018_, _07030_, _17007_ }), .Y(_17039_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29904_ ( .A({ _17082_, _07018_, _07030_, _17018_ }), .Y(_17050_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29905_ ( .A({ _17093_, _07018_, _07030_, _17029_ }), .Y(_17061_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29906_ ( .A({ _17096_, _07018_, _07030_, _17032_ }), .Y(_17064_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29907_ ( .A({ _17097_, _07018_, _07030_, _17033_ }), .Y(_17065_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29908_ ( .A({ _17098_, _07018_, _07030_, _17034_ }), .Y(_17066_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29909_ ( .A({ _17099_, _07018_, _07030_, _17035_ }), .Y(_17067_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29910_ ( .A({ _17100_, _07018_, _07030_, _17036_ }), .Y(_17068_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29911_ ( .A({ _17101_, _07018_, _07030_, _17037_ }), .Y(_17069_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29912_ ( .A({ _17102_, _07018_, _07030_, _17038_ }), .Y(_17070_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29913_ ( .A({ _17072_, _07018_, _07030_, _17008_ }), .Y(_17040_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29914_ ( .A({ _17073_, _07018_, _07030_, _17009_ }), .Y(_17041_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29915_ ( .A({ _17074_, _07018_, _07030_, _17010_ }), .Y(_17042_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29916_ ( .A({ _17075_, _07018_, _07030_, _17011_ }), .Y(_17043_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29917_ ( .A({ _17076_, _07018_, _07030_, _17012_ }), .Y(_17044_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29918_ ( .A({ _17077_, _07018_, _07030_, _17013_ }), .Y(_17045_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29919_ ( .A({ _17078_, _07018_, _07030_, _17014_ }), .Y(_17046_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29920_ ( .A({ _17079_, _07018_, _07030_, _17015_ }), .Y(_17047_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29921_ ( .A({ _17080_, _07018_, _07030_, _17016_ }), .Y(_17048_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29922_ ( .A({ _17081_, _07018_, _07030_, _17017_ }), .Y(_17049_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29923_ ( .A({ _17083_, _07018_, _07030_, _17019_ }), .Y(_17051_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29924_ ( .A({ _17084_, _07018_, _07030_, _17020_ }), .Y(_17052_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29925_ ( .A({ _17085_, _07018_, _07030_, _17021_ }), .Y(_17053_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29926_ ( .A({ _17086_, _07018_, _07030_, _17022_ }), .Y(_17054_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29927_ ( .A({ _17087_, _07018_, _07030_, _17023_ }), .Y(_17055_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29928_ ( .A({ _17088_, _07018_, _07030_, _17024_ }), .Y(_17056_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29929_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18233_, _18265_ }), .Y(_18201_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29930_ ( .A({ _17089_, _07018_, _07030_, _17025_ }), .Y(_17057_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29931_ ( .A({ _17090_, _07018_, _07030_, _17026_ }), .Y(_17058_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29932_ ( .A({ _17091_, _07018_, _07030_, _17027_ }), .Y(_17059_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29933_ ( .A({ _17092_, _07018_, _07030_, _17028_ }), .Y(_17060_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29934_ ( .A({ _17094_, _07018_, _07030_, _17030_ }), .Y(_17062_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29935_ ( .A({ _17095_, _07018_, _07030_, _17031_ }), .Y(_17063_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29936_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18232_, _18264_ }), .Y(_18200_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29937_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18231_, _18263_ }), .Y(_18199_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29938_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18230_, _18262_ }), .Y(_18198_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29939_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18229_, _18261_ }), .Y(_18197_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29940_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18226_, _18258_ }), .Y(_18194_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29941_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18228_, _18260_ }), .Y(_18196_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29942_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18227_, _18259_ }), .Y(_18195_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29943_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18225_, _18257_ }), .Y(_18193_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29944_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18224_, _18256_ }), .Y(_18192_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29945_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18252_, _18284_ }), .Y(_18220_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29946_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18254_, _18286_ }), .Y(_18222_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29947_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18253_, _18285_ }), .Y(_18221_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29948_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18251_, _18283_ }), .Y(_18219_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29949_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18250_, _18282_ }), .Y(_18218_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29950_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18245_, _18277_ }), .Y(_18213_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29951_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18249_, _18281_ }), .Y(_18217_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29952_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18248_, _18280_ }), .Y(_18216_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29953_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18234_, _18266_ }), .Y(_18202_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _29954_ ( .A({ _06995_, _stream_conv2d_16_source_27_source_pat_fsm_10[0], _18223_, _18255_ }), .Y(_18191_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29955_ ( .A({ _05967_, _06995_ }), .Y(_24059_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _29956_ ( .A({ _stream_conv2d_16_source_27_source_pat_fsm_10[1], _06996_, _07004_, _stream_conv2d_16_source_27_source_pat_fsm_10[0] }), .Y(_05967_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29957_ ( .A({ _16974_, _07018_, _16908_, _05948_ }), .Y(_16941_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29958_ ( .A({ _16985_, _07018_, _16919_, _05948_ }), .Y(_16952_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29959_ ( .A({ _16996_, _07018_, _16930_, _05948_ }), .Y(_16963_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29960_ ( .A({ _17000_, _07018_, _16934_, _05948_ }), .Y(_16967_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29961_ ( .A({ _17001_, _07018_, _16935_, _05948_ }), .Y(_16968_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29962_ ( .A({ _17002_, _07018_, _16936_, _05948_ }), .Y(_16969_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29963_ ( .A({ _17003_, _07018_, _16937_, _05948_ }), .Y(_16970_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29964_ ( .A({ _17004_, _07018_, _16938_, _05948_ }), .Y(_16971_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29965_ ( .A({ _17005_, _07018_, _16939_, _05948_ }), .Y(_16972_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29966_ ( .A({ _17006_, _07018_, _16940_, _05948_ }), .Y(_16973_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29967_ ( .A({ _16975_, _07018_, _16909_, _05948_ }), .Y(_16942_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29968_ ( .A({ _16976_, _07018_, _16910_, _05948_ }), .Y(_16943_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29969_ ( .A({ _16977_, _07018_, _16911_, _05948_ }), .Y(_16944_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29970_ ( .A({ _16978_, _07018_, _16912_, _05948_ }), .Y(_16945_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29971_ ( .A({ _16979_, _07018_, _16913_, _05948_ }), .Y(_16946_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29972_ ( .A({ _16980_, _07018_, _16914_, _05948_ }), .Y(_16947_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29973_ ( .A({ _16981_, _07018_, _16915_, _05948_ }), .Y(_16948_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29974_ ( .A({ _16982_, _07018_, _16916_, _05948_ }), .Y(_16949_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29975_ ( .A({ _16983_, _07018_, _16917_, _05948_ }), .Y(_16950_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29976_ ( .A({ _16984_, _07018_, _16918_, _05948_ }), .Y(_16951_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29977_ ( .A({ _16986_, _07018_, _16920_, _05948_ }), .Y(_16953_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29978_ ( .A({ _16987_, _07018_, _16921_, _05948_ }), .Y(_16954_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29979_ ( .A({ _16988_, _07018_, _16922_, _05948_ }), .Y(_16955_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29980_ ( .A({ _16989_, _07018_, _16923_, _05948_ }), .Y(_16956_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29981_ ( .A({ _16990_, _07018_, _16924_, _05948_ }), .Y(_16957_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29982_ ( .A({ _16991_, _07018_, _16925_, _05948_ }), .Y(_16958_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29983_ ( .A({ _16992_, _07018_, _16926_, _05948_ }), .Y(_16959_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29984_ ( .A({ _16993_, _07018_, _16927_, _05948_ }), .Y(_16960_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29985_ ( .A({ _16994_, _07018_, _16928_, _05948_ }), .Y(_16961_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29986_ ( .A({ _16995_, _07018_, _16929_, _05948_ }), .Y(_16962_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29987_ ( .A({ _16997_, _07018_, _16931_, _05948_ }), .Y(_16964_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29988_ ( .A({ _16998_, _07018_, _16932_, _05948_ }), .Y(_16965_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _29989_ ( .A({ _16999_, _07018_, _16933_, _05948_ }), .Y(_16966_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _29990_ ( .A({ _06021_, _07066_ }), .Y(_24075_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _29991_ ( .A({ _07067_, _06931_, _06923_, _06920_ }), .Y(_07066_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _29992_ ( .A({ control_conv2d_16[2:0], control_conv2d_16[3] }), .Y(_07067_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _29993_ ( .A({ _06021_, _21579_, _06930_ }), .Y(_21580_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _29994_ ( .A({ _21247_, _06930_, _07066_, _21279_ }), .Y(_05517_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _29995_ ( .A({ _07099_, _07093_, _07068_ }), .Y(_24046_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _29996_ ( .A({ _07087_, _07069_, _05945_, _07085_ }), .Y(_07068_) );
  \$lut  #( .LUT(16'hebff), .WIDTH(4) ) _29997_ ( .A({ _07070_, control_max_pool_serial_18[2], _07080_, control_max_pool_serial_18[3] }), .Y(_07069_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _29998_ ( .A({ control_max_pool_serial_18[4], _07071_, control_max_pool_serial_18[5] }), .Y(_07070_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _29999_ ( .A({ _07077_, _07072_ }), .Y(_07071_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30000_ ( .A({ _07076_, _07075_, _07074_, _07073_ }), .Y(_07072_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30001_ ( .A(control_max_pool_serial_18[31:28]), .Y(_07073_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30002_ ( .A({ control_max_pool_serial_18[26:25], control_max_pool_serial_18[23], control_max_pool_serial_18[20] }), .Y(_07074_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30003_ ( .A({ control_max_pool_serial_18[11], control_max_pool_serial_18[8:6] }), .Y(_07075_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30004_ ( .A({ control_max_pool_serial_18[19], control_max_pool_serial_18[16], control_max_pool_serial_18[14:13] }), .Y(_07076_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30005_ ( .A({ _07079_, _07078_, control_max_pool_serial_18[10:9] }), .Y(_07077_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30006_ ( .A({ control_max_pool_serial_18[27], control_max_pool_serial_18[24], control_max_pool_serial_18[22:21] }), .Y(_07078_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30007_ ( .A({ control_max_pool_serial_18[18:17], control_max_pool_serial_18[15], control_max_pool_serial_18[12] }), .Y(_07079_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30008_ ( .A({ control_max_pool_serial_18[0], control_max_pool_serial_18[1] }), .Y(_07080_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30009_ ( .A({ _07084_, _07081_ }), .Y(_05945_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30010_ ( .A({ _07083_, _07082_, _07071_ }), .Y(_07081_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _30011_ ( .A(control_max_pool_serial_18[3:2]), .Y(_07082_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _30012_ ( .A({ control_max_pool_serial_18[4], control_max_pool_serial_18[5] }), .Y(_07083_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30013_ ( .A(control_max_pool_serial_18[1:0]), .Y(_07084_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30014_ ( .A({ _07086_, _07080_, _07070_ }), .Y(_07085_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30015_ ( .A({ control_max_pool_serial_18[2], control_max_pool_serial_18[3] }), .Y(_07086_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30016_ ( .A({ _05942_, _07092_, _07088_ }), .Y(_07087_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30017_ ( .A({ control_max_pool_serial_18[3:2], _07083_, _07071_ }), .Y(_07088_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _30018_ ( .A({ control_max_pool_serial_18[4], _07071_, _07089_, control_max_pool_serial_18[5] }), .Y(_05942_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30019_ ( .A({ _07091_, _07090_ }), .Y(_07089_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30020_ ( .A(control_max_pool_serial_18[3:2]), .Y(_07090_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30021_ ( .A({ control_max_pool_serial_18[0], control_max_pool_serial_18[1] }), .Y(_07091_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30022_ ( .A({ _07083_, _07086_, _07071_ }), .Y(_07092_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _30023_ ( .A({ _07097_, _07094_, _07081_ }), .Y(_07093_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30024_ ( .A({ _07096_, _07095_ }), .Y(_07094_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30025_ ( .A({ _07090_, _07083_, _07071_ }), .Y(_07095_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _30026_ ( .A({ control_max_pool_serial_18[0], control_max_pool_serial_18[1] }), .Y(_07096_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30027_ ( .A({ _07082_, _07098_ }), .Y(_07097_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30028_ ( .A({ control_max_pool_serial_18[4], _07071_, _07096_, control_max_pool_serial_18[5] }), .Y(_07098_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30029_ ( .A({ _07095_, _07102_, _07101_, _07100_ }), .Y(_07099_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30030_ ( .A({ _07084_, _07082_, _07070_ }), .Y(_07100_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30031_ ( .A({ _07090_, _07098_ }), .Y(_07101_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30032_ ( .A({ _07091_, _07082_, _07070_ }), .Y(_07102_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30033_ ( .A({ _21246_, _06930_, _07066_, _21278_ }), .Y(_05518_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30034_ ( .A({ _21244_, _06930_, _07066_, _21276_ }), .Y(_05519_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30035_ ( .A({ _21243_, _06930_, _07066_, _21275_ }), .Y(_05520_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30036_ ( .A({ _21242_, _06930_, _07066_, _21274_ }), .Y(_05521_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30037_ ( .A({ _07083_, _07089_, _07071_ }), .Y(_07103_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30038_ ( .A({ _16614_, _07084_, _07082_, _07070_ }), .Y(_07104_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30039_ ( .A({ _16902_, _07106_ }), .Y(_07105_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30040_ ( .A({ _07096_, _07083_, _07082_, _07071_ }), .Y(_07106_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30041_ ( .A({ _16582_, _07086_, _07070_ }), .Y(_07107_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30042_ ( .A({ _16710_, _07084_, _07088_ }), .Y(_07108_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30043_ ( .A({ _16838_, _07096_, _07092_ }), .Y(_07109_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30044_ ( .A({ _16646_, _07091_, _07082_, _07070_ }), .Y(_07110_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30045_ ( .A({ _21241_, _06930_, _07066_, _21273_ }), .Y(_05522_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30046_ ( .A({ _16588_, _07084_, _07082_, _07070_ }), .Y(_07111_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30047_ ( .A({ _16556_, _07086_, _07080_, _07070_ }), .Y(_07112_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _30048_ ( .A({ _24044_, _07115_, _07114_, _16812_ }), .Y(_07113_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30049_ ( .A({ _07096_, _07092_ }), .Y(_07114_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _30050_ ( .A({ _07084_, _07081_, _07086_, _07070_ }), .Y(_24044_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30051_ ( .A({ _16620_, _07091_, _07082_, _07070_ }), .Y(_07115_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _30052_ ( .A({ _07117_, _07118_, _07097_, _16652_ }), .Y(_07116_) );
  \$lut  #( .LUT(16'hf4ff), .WIDTH(4) ) _30053_ ( .A({ _07088_, control_max_pool_serial_18[0], control_max_pool_serial_18[1], _16684_ }), .Y(_07117_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30054_ ( .A({ _16876_, _07106_ }), .Y(_07118_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30055_ ( .A({ _07127_, _07122_, _07120_, _07119_ }), .Y(_16522_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30056_ ( .A({ _16618_, _07100_, _16842_, _07114_ }), .Y(_07119_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30057_ ( .A({ _16554_, _07101_, _16746_, _07121_ }), .Y(_07120_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30058_ ( .A({ _07084_, _07095_ }), .Y(_07121_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30059_ ( .A({ _07126_, _07125_, _07124_, _07123_ }), .Y(_07122_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30060_ ( .A({ _16586_, _07086_, _07080_, _07070_ }), .Y(_07123_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30061_ ( .A({ _16874_, _07080_, _07081_ }), .Y(_07124_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30062_ ( .A({ _16906_, _07106_ }), .Y(_07125_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30063_ ( .A({ _16682_, _07082_, _07098_ }), .Y(_07126_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30064_ ( .A({ _07129_, _07131_, _07130_, _07128_ }), .Y(_07127_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30065_ ( .A({ _16650_, _07091_, _07082_, _07070_ }), .Y(_07128_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30066_ ( .A({ _16490_, _05942_, _16778_, _07103_ }), .Y(_07129_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30067_ ( .A({ _16810_, _07096_, _07095_ }), .Y(_07130_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30068_ ( .A({ _16714_, _07084_, _07088_ }), .Y(_07131_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30069_ ( .A({ _16855_, _07080_, _07081_ }), .Y(_07132_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _30070_ ( .A({ _07091_, _07081_, _07086_, _07070_ }), .Y(_07133_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30071_ ( .A({ _16471_, _05942_, _16759_, _07103_ }), .Y(_07134_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _30072_ ( .A({ _07092_, _07091_, _07084_ }), .Y(_07135_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30073_ ( .A({ _16567_, _07086_, _07080_, _07070_ }), .Y(_07136_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30074_ ( .A({ _16887_, _07106_ }), .Y(_07137_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30075_ ( .A({ _16535_, _07090_, _07098_ }), .Y(_07138_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30076_ ( .A({ _16866_, _07080_, _07081_ }), .Y(_07139_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30077_ ( .A({ _16578_, _07086_, _07070_ }), .Y(_07140_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30078_ ( .A({ _07069_, _07142_, _07135_, _07143_ }), .Y(_07141_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30079_ ( .A({ _16482_, _05942_, _16770_, _07103_ }), .Y(_07142_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30080_ ( .A({ _16898_, _07106_ }), .Y(_07143_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30081_ ( .A({ _07084_, _07088_ }), .Y(_07144_) );
  \$lut  #( .LUT(16'h770f), .WIDTH(4) ) _30082_ ( .A({ control_max_pool_serial_18[1], _07088_, control_max_pool_serial_18[0], _07095_ }), .Y(_07145_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30083_ ( .A({ _16738_, _07084_, _07095_ }), .Y(_07146_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30084_ ( .A({ _16642_, _07091_, _07082_, _07070_ }), .Y(_07147_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30085_ ( .A({ _16610_, _07084_, _07082_, _07070_ }), .Y(_07148_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30086_ ( .A({ _16645_, _07091_, _07082_, _07070_ }), .Y(_07149_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30087_ ( .A({ _16613_, _07084_, _07082_, _07070_ }), .Y(_07150_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30088_ ( .A({ _16869_, _07080_, _07081_ }), .Y(_07151_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30089_ ( .A({ _16709_, _07084_, _07088_ }), .Y(_07152_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30090_ ( .A({ _16581_, _07086_, _07080_, _07070_ }), .Y(_07153_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30091_ ( .A({ _16901_, _07106_ }), .Y(_07154_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30092_ ( .A({ _21240_, _06930_, _07066_, _21272_ }), .Y(_05523_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30093_ ( .A({ _16839_, _07096_, _07092_ }), .Y(_07155_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30094_ ( .A({ _16647_, _07091_, _07082_, _07070_ }), .Y(_07156_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30095_ ( .A({ _16711_, _07144_, _16903_, _07106_ }), .Y(_07157_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30096_ ( .A({ _16807_, _07094_, _16871_, _07159_ }), .Y(_07158_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30097_ ( .A({ _07080_, _07081_ }), .Y(_07159_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30098_ ( .A({ _07162_, _07164_, _07163_, _07161_ }), .Y(_07160_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30099_ ( .A({ _16615_, _07084_, _07082_, _07070_ }), .Y(_07161_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30100_ ( .A({ _16487_, _05942_, _16775_, _07103_ }), .Y(_07162_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30101_ ( .A({ _16583_, _07086_, _07080_, _07070_ }), .Y(_07163_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30102_ ( .A({ _16743_, _07084_, _07095_ }), .Y(_07164_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30103_ ( .A({ _07172_, _07171_, _07170_, _07165_ }), .Y(_16520_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30104_ ( .A({ _07169_, _07168_, _07167_, _07166_ }), .Y(_07165_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30105_ ( .A({ _16616_, _07084_, _07082_, _07070_ }), .Y(_07166_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30106_ ( .A({ _16552_, _07090_, _07098_ }), .Y(_07167_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30107_ ( .A({ _16904_, _07106_ }), .Y(_07168_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30108_ ( .A({ _16648_, _07091_, _07082_, _07070_ }), .Y(_07169_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30109_ ( .A({ _16584_, _07085_, _16744_, _07121_ }), .Y(_07170_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30110_ ( .A({ _16680_, _07097_, _16840_, _07114_ }), .Y(_07171_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30111_ ( .A({ _07174_, _07176_, _07175_, _07173_ }), .Y(_07172_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30112_ ( .A({ _16808_, _07096_, _07095_ }), .Y(_07173_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30113_ ( .A({ _16488_, _05942_, _16776_, _07103_ }), .Y(_07174_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30114_ ( .A({ _16712_, _07084_, _07088_ }), .Y(_07175_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30115_ ( .A({ _16872_, _07080_, _07081_ }), .Y(_07176_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30116_ ( .A({ _16841_, _07096_, _07092_ }), .Y(_07177_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30117_ ( .A({ _16713_, _07144_, _16905_, _07106_ }), .Y(_07178_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30118_ ( .A({ _16585_, _07085_, _16873_, _07159_ }), .Y(_07179_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30119_ ( .A({ _16553_, _07090_, _07098_ }), .Y(_07180_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30120_ ( .A({ _16489_, _05942_, _16777_, _07103_ }), .Y(_07181_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30121_ ( .A({ _16782_, _07096_, _07095_ }), .Y(_07182_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30122_ ( .A({ _16878_, _07106_ }), .Y(_07183_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30123_ ( .A({ _16558_, _07085_, _07144_, _16686_ }), .Y(_07184_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30124_ ( .A({ _16718_, _07121_, _16814_, _07114_ }), .Y(_07185_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30125_ ( .A({ _07188_, _07190_, _07189_, _07187_ }), .Y(_07186_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30126_ ( .A({ _16590_, _07084_, _07082_, _07070_ }), .Y(_07187_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30127_ ( .A({ _16462_, _05942_, _16750_, _07103_ }), .Y(_07188_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30128_ ( .A({ _16622_, _07091_, _07082_, _07070_ }), .Y(_07189_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30129_ ( .A({ _16846_, _07080_, _07081_ }), .Y(_07190_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30130_ ( .A({ _16619_, _07084_, _07082_, _07070_ }), .Y(_07191_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30131_ ( .A({ _16907_, _07106_ }), .Y(_07192_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30132_ ( .A({ _16651_, _07091_, _07082_, _07070_ }), .Y(_07193_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30133_ ( .A({ _16587_, _07085_, _16683_, _07097_ }), .Y(_07194_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30134_ ( .A({ _16555_, _07101_, _16843_, _07114_ }), .Y(_07195_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30135_ ( .A({ _16491_, _05942_, _16779_, _07103_ }), .Y(_07196_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30136_ ( .A({ _16715_, _07084_, _07088_ }), .Y(_07197_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30137_ ( .A({ _16875_, _07080_, _07081_ }), .Y(_07198_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30138_ ( .A({ _16621_, _07102_, _16813_, _07114_ }), .Y(_07199_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30139_ ( .A({ _16557_, _07085_, _16589_, _07100_ }), .Y(_07200_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30140_ ( .A({ _16877_, _07106_ }), .Y(_07201_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30141_ ( .A({ _16845_, _07080_, _07081_ }), .Y(_07202_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30142_ ( .A({ _16461_, _05942_, _16749_, _07103_ }), .Y(_07203_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30143_ ( .A({ _16781_, _07096_, _07095_ }), .Y(_07204_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30144_ ( .A({ _21239_, _06930_, _07066_, _21271_ }), .Y(_05524_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30145_ ( .A({ _16594_, _07084_, _07082_, _07070_ }), .Y(_07205_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30146_ ( .A({ _16882_, _07106_ }), .Y(_07206_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30147_ ( .A({ _16626_, _07091_, _07082_, _07070_ }), .Y(_07207_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30148_ ( .A({ _16658_, _07097_, _16850_, _07159_ }), .Y(_07208_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30149_ ( .A({ _16530_, _07101_, _16818_, _07114_ }), .Y(_07209_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30150_ ( .A({ _16466_, _05942_, _16754_, _07103_ }), .Y(_07210_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30151_ ( .A({ _16690_, _07084_, _07088_ }), .Y(_07211_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30152_ ( .A({ _16562_, _07086_, _07080_, _07070_ }), .Y(_07212_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30153_ ( .A({ _16815_, _07096_, _07092_ }), .Y(_07213_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30154_ ( .A({ _16783_, _07094_, _07144_, _16687_ }), .Y(_07214_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30155_ ( .A({ _16559_, _07085_, _16879_, _07106_ }), .Y(_07215_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30156_ ( .A({ _07218_, _07220_, _07219_, _07217_ }), .Y(_07216_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30157_ ( .A({ _16719_, _07084_, _07095_ }), .Y(_07217_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30158_ ( .A({ _16463_, _05942_, _16751_, _07103_ }), .Y(_07218_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30159_ ( .A({ _16847_, _07080_, _07081_ }), .Y(_07219_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30160_ ( .A({ _16527_, _07090_, _07098_ }), .Y(_07220_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30161_ ( .A({ _16816_, _07096_, _07092_ }), .Y(_07221_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30162_ ( .A({ _16784_, _07094_, _07144_, _16688_ }), .Y(_07222_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30163_ ( .A({ _16848_, _07159_, _16880_, _07106_ }), .Y(_07223_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30164_ ( .A({ _07226_, _07228_, _07227_, _07225_ }), .Y(_07224_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30165_ ( .A({ _16720_, _07084_, _07095_ }), .Y(_07225_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30166_ ( .A({ _16464_, _05942_, _16752_, _07103_ }), .Y(_07226_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30167_ ( .A({ _16560_, _07086_, _07080_, _07070_ }), .Y(_07227_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30168_ ( .A({ _16528_, _07090_, _07098_ }), .Y(_07228_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30169_ ( .A({ _16785_, _07096_, _07095_ }), .Y(_07229_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30170_ ( .A({ _16881_, _07106_ }), .Y(_07230_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30171_ ( .A({ _16561_, _07085_, _07144_, _16689_ }), .Y(_07231_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30172_ ( .A({ _16721_, _07121_, _16817_, _07114_ }), .Y(_07232_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30173_ ( .A({ _07235_, _07237_, _07236_, _07234_ }), .Y(_07233_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30174_ ( .A({ _16593_, _07084_, _07082_, _07070_ }), .Y(_07234_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30175_ ( .A({ _16465_, _05942_, _16753_, _07103_ }), .Y(_07235_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30176_ ( .A({ _16625_, _07091_, _07082_, _07070_ }), .Y(_07236_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30177_ ( .A({ _16849_, _07080_, _07081_ }), .Y(_07237_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30178_ ( .A({ _07242_, _07241_, _07240_, _07239_ }), .Y(_07238_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30179_ ( .A({ _16883_, _07106_ }), .Y(_07239_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30180_ ( .A({ _16563_, _07086_, _07080_, _07070_ }), .Y(_07240_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30181_ ( .A({ _16659_, _07082_, _07098_ }), .Y(_07241_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30182_ ( .A({ _16595_, _07084_, _07082_, _07070_ }), .Y(_07242_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30183_ ( .A({ _16531_, _07101_, _16819_, _07114_ }), .Y(_07243_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30184_ ( .A({ _16627_, _07102_, _07144_, _16691_ }), .Y(_07244_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30185_ ( .A({ _16467_, _05942_, _16755_, _07103_ }), .Y(_07245_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30186_ ( .A({ _16851_, _07080_, _07081_ }), .Y(_07246_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30187_ ( .A({ _07254_, _07249_, _07248_, _07247_ }), .Y(_16506_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30188_ ( .A({ _16666_, _07097_, _16730_, _07121_ }), .Y(_07247_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30189_ ( .A({ _16794_, _07094_, _07144_, _16698_ }), .Y(_07248_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30190_ ( .A({ _07253_, _07252_, _07251_, _07250_ }), .Y(_07249_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30191_ ( .A({ _16890_, _07106_ }), .Y(_07250_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30192_ ( .A({ _16826_, _07096_, _07092_ }), .Y(_07251_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30193_ ( .A({ _16602_, _07084_, _07082_, _07070_ }), .Y(_07252_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30194_ ( .A({ _16538_, _07090_, _07098_ }), .Y(_07253_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30195_ ( .A({ _07256_, _07258_, _07257_, _07255_ }), .Y(_07254_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30196_ ( .A({ _16570_, _07086_, _07080_, _07070_ }), .Y(_07255_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30197_ ( .A({ _16474_, _05942_, _16762_, _07103_ }), .Y(_07256_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30198_ ( .A({ _16634_, _07091_, _07082_, _07070_ }), .Y(_07257_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30199_ ( .A({ _16858_, _07080_, _07081_ }), .Y(_07258_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30200_ ( .A({ _16596_, _07100_, _07101_, _16532_ }), .Y(_07259_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30201_ ( .A({ _16628_, _07102_, _16852_, _07159_ }), .Y(_07260_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30202_ ( .A({ _16884_, _07106_ }), .Y(_07261_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30203_ ( .A({ _16660_, _07082_, _07098_ }), .Y(_07262_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30204_ ( .A({ _16820_, _07096_, _07092_ }), .Y(_07263_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30205_ ( .A({ _16468_, _05942_, _16756_, _07103_ }), .Y(_07264_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30206_ ( .A({ _16692_, _07084_, _07088_ }), .Y(_07265_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30207_ ( .A({ _16564_, _07086_, _07080_, _07070_ }), .Y(_07266_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30208_ ( .A({ _16597_, _07084_, _07082_, _07070_ }), .Y(_07267_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30209_ ( .A({ _16661_, _07082_, _07098_ }), .Y(_07268_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30210_ ( .A({ _16533_, _07101_, _16853_, _07159_ }), .Y(_07269_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30211_ ( .A({ _16693_, _07144_, _16821_, _07114_ }), .Y(_07270_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30212_ ( .A({ _07273_, _07275_, _07274_, _07272_ }), .Y(_07271_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30213_ ( .A({ _16565_, _07086_, _07080_, _07070_ }), .Y(_07272_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30214_ ( .A({ _16469_, _05942_, _16757_, _07103_ }), .Y(_07273_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30215_ ( .A({ _16885_, _07106_ }), .Y(_07274_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30216_ ( .A({ _16629_, _07091_, _07082_, _07070_ }), .Y(_07275_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30217_ ( .A({ _16822_, _07096_, _07092_ }), .Y(_07276_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30218_ ( .A({ _16694_, _07144_, _16886_, _07106_ }), .Y(_07277_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30219_ ( .A({ _16566_, _07085_, _16854_, _07159_ }), .Y(_07278_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30220_ ( .A({ _16534_, _07090_, _07098_ }), .Y(_07279_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30221_ ( .A({ _16470_, _05942_, _16758_, _07103_ }), .Y(_07280_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30222_ ( .A({ _16600_, _07100_, _07101_, _16536_ }), .Y(_07281_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30223_ ( .A({ _16664_, _07097_, _07102_, _16632_ }), .Y(_07282_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30224_ ( .A({ _16888_, _07106_ }), .Y(_07283_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30225_ ( .A({ _16568_, _07086_, _07080_, _07070_ }), .Y(_07284_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30226_ ( .A({ _16472_, _05942_, _16760_, _07103_ }), .Y(_07285_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30227_ ( .A({ _16856_, _07080_, _07081_ }), .Y(_07286_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30228_ ( .A({ _16825_, _07096_, _07092_ }), .Y(_07287_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30229_ ( .A({ _16697_, _07144_, _16889_, _07106_ }), .Y(_07288_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30230_ ( .A({ _16569_, _07085_, _16857_, _07159_ }), .Y(_07289_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30231_ ( .A({ _16537_, _07090_, _07098_ }), .Y(_07290_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30232_ ( .A({ _16473_, _05942_, _16761_, _07103_ }), .Y(_07291_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30233_ ( .A({ _16893_, _07106_ }), .Y(_07292_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30234_ ( .A({ _16669_, _07082_, _07098_ }), .Y(_07293_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30235_ ( .A({ _16573_, _07086_, _07080_, _07070_ }), .Y(_07294_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30236_ ( .A({ _16701_, _07144_, _16829_, _07114_ }), .Y(_07295_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30237_ ( .A({ _16605_, _07100_, _07101_, _16541_ }), .Y(_07296_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30238_ ( .A({ _16477_, _05942_, _16765_, _07103_ }), .Y(_07297_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30239_ ( .A({ _16637_, _07091_, _07082_, _07070_ }), .Y(_07298_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30240_ ( .A({ _16861_, _07080_, _07081_ }), .Y(_07299_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30241_ ( .A({ _16635_, _07091_, _07082_, _07070_ }), .Y(_07300_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30242_ ( .A({ _16827_, _07096_, _07092_ }), .Y(_07301_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30243_ ( .A({ _16731_, _07084_, _07095_ }), .Y(_07302_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30244_ ( .A({ _16795_, _07094_, _07144_, _16699_ }), .Y(_07303_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30245_ ( .A({ _16859_, _07159_, _16891_, _07106_ }), .Y(_07304_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30246_ ( .A({ _16603_, _07084_, _07082_, _07070_ }), .Y(_07305_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30247_ ( .A({ _16475_, _05942_, _16763_, _07103_ }), .Y(_07306_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30248_ ( .A({ _16571_, _07086_, _07080_, _07070_ }), .Y(_07307_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30249_ ( .A({ _07315_, _07310_, _07309_, _07308_ }), .Y(_16508_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30250_ ( .A({ _16668_, _07097_, _16828_, _07114_ }), .Y(_07308_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30251_ ( .A({ _16604_, _07100_, _16732_, _07121_ }), .Y(_07309_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30252_ ( .A({ _07314_, _07313_, _07312_, _07311_ }), .Y(_07310_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30253_ ( .A({ _16860_, _07080_, _07081_ }), .Y(_07311_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30254_ ( .A({ _16892_, _07106_ }), .Y(_07312_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30255_ ( .A({ _16572_, _07086_, _07080_, _07070_ }), .Y(_07313_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30256_ ( .A({ _16540_, _07090_, _07098_ }), .Y(_07314_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30257_ ( .A({ _07317_, _07319_, _07318_, _07316_ }), .Y(_07315_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30258_ ( .A({ _16636_, _07091_, _07082_, _07070_ }), .Y(_07316_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30259_ ( .A({ _16476_, _05942_, _16764_, _07103_ }), .Y(_07317_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30260_ ( .A({ _16796_, _07096_, _07095_ }), .Y(_07318_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30261_ ( .A({ _16700_, _07084_, _07088_ }), .Y(_07319_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30262_ ( .A({ _21238_, _06930_, _07066_, _21270_ }), .Y(_05525_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30263_ ( .A({ _07323_, _07322_, _07321_, _13037_ }), .Y(_16510_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30264_ ( .A({ _16542_, _07090_, _07098_ }), .Y(_07320_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30265_ ( .A({ _16798_, _07094_, _16862_, _07159_ }), .Y(_07321_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30266_ ( .A({ _16670_, _07097_, _16734_, _07121_ }), .Y(_07322_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30267_ ( .A({ _07325_, _07327_, _07326_, _07324_ }), .Y(_07323_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30268_ ( .A({ _16830_, _07096_, _07092_ }), .Y(_07324_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30269_ ( .A({ _16478_, _05942_, _16766_, _07103_ }), .Y(_07325_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30270_ ( .A({ _16894_, _07106_ }), .Y(_07326_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30271_ ( .A({ _16702_, _07084_, _07088_ }), .Y(_07327_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30272_ ( .A({ _07335_, _07334_, _07333_, _07328_ }), .Y(_16512_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30273_ ( .A({ _07332_, _07331_, _07330_, _07329_ }), .Y(_07328_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30274_ ( .A({ _16608_, _07084_, _07082_, _07070_ }), .Y(_07329_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30275_ ( .A({ _16544_, _07090_, _07098_ }), .Y(_07330_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30276_ ( .A({ _16896_, _07106_ }), .Y(_07331_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30277_ ( .A({ _16640_, _07091_, _07082_, _07070_ }), .Y(_07332_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30278_ ( .A({ _16576_, _07085_, _16736_, _07121_ }), .Y(_07333_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30279_ ( .A({ _16672_, _07097_, _16832_, _07114_ }), .Y(_07334_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30280_ ( .A({ _07337_, _07339_, _07338_, _07336_ }), .Y(_07335_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30281_ ( .A({ _16800_, _07096_, _07095_ }), .Y(_07336_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30282_ ( .A({ _16480_, _05942_, _16768_, _07103_ }), .Y(_07337_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30283_ ( .A({ _16704_, _07084_, _07088_ }), .Y(_07338_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30284_ ( .A({ _16864_, _07080_, _07081_ }), .Y(_07339_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30285_ ( .A({ _16831_, _07096_, _07092_ }), .Y(_07340_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30286_ ( .A({ _16703_, _07144_, _16895_, _07106_ }), .Y(_07341_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30287_ ( .A({ _16575_, _07085_, _16863_, _07159_ }), .Y(_07342_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30288_ ( .A({ _16543_, _07090_, _07098_ }), .Y(_07343_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30289_ ( .A({ _16479_, _05942_, _16767_, _07103_ }), .Y(_07344_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30290_ ( .A({ _16609_, _07100_, _07101_, _16545_ }), .Y(_07345_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30291_ ( .A({ _16673_, _07097_, _16737_, _07121_ }), .Y(_07346_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30292_ ( .A({ _16865_, _07080_, _07081_ }), .Y(_07347_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30293_ ( .A({ _16897_, _07106_ }), .Y(_07348_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30294_ ( .A({ _07351_, _07353_, _07352_, _07350_ }), .Y(_07349_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30295_ ( .A({ _16641_, _07091_, _07082_, _07070_ }), .Y(_07350_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30296_ ( .A({ _16481_, _05942_, _16769_, _07103_ }), .Y(_07351_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30297_ ( .A({ _16577_, _07086_, _07080_, _07070_ }), .Y(_07352_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30298_ ( .A({ _16705_, _07084_, _07088_ }), .Y(_07353_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30299_ ( .A({ _07361_, _07356_, _07355_, _07354_ }), .Y(_16515_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30300_ ( .A({ _16611_, _07100_, _16835_, _07114_ }), .Y(_07354_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30301_ ( .A({ _16547_, _07101_, _16739_, _07121_ }), .Y(_07355_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30302_ ( .A({ _07360_, _07359_, _07358_, _07357_ }), .Y(_07356_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30303_ ( .A({ _16579_, _07086_, _07080_, _07070_ }), .Y(_07357_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30304_ ( .A({ _16867_, _07080_, _07081_ }), .Y(_07358_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30305_ ( .A({ _16899_, _07106_ }), .Y(_07359_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30306_ ( .A({ _16675_, _07082_, _07098_ }), .Y(_07360_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30307_ ( .A({ _07363_, _07365_, _07364_, _07362_ }), .Y(_07361_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30308_ ( .A({ _16643_, _07091_, _07082_, _07070_ }), .Y(_07362_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30309_ ( .A({ _16483_, _05942_, _16771_, _07103_ }), .Y(_07363_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30310_ ( .A({ _16803_, _07096_, _07095_ }), .Y(_07364_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30311_ ( .A({ _16707_, _07084_, _07088_ }), .Y(_07365_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30312_ ( .A({ _16612_, _07100_, _16836_, _07114_ }), .Y(_07366_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30313_ ( .A({ _16644_, _07102_, _16868_, _07159_ }), .Y(_07367_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30314_ ( .A({ _16900_, _07106_ }), .Y(_07368_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30315_ ( .A({ _16484_, _05942_, _16772_, _07103_ }), .Y(_07369_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30316_ ( .A({ _16708_, _07084_, _07088_ }), .Y(_07370_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30317_ ( .A({ _16580_, _07086_, _07080_, _07070_ }), .Y(_07371_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30318_ ( .A({ _21237_, _06930_, _07066_, _21269_ }), .Y(_05526_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30319_ ( .A({ _21236_, _06930_, _07066_, _21268_ }), .Y(_05527_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30320_ ( .A({ _21235_, _06930_, _07066_, _21267_ }), .Y(_05528_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30321_ ( .A({ _21233_, _06930_, _07066_, _21265_ }), .Y(_05529_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30322_ ( .A({ _21232_, _06930_, _07066_, _21264_ }), .Y(_05530_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30323_ ( .A({ _21231_, _06930_, _07066_, _21263_ }), .Y(_05531_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30324_ ( .A({ _21230_, _06930_, _07066_, _21262_ }), .Y(_05532_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30325_ ( .A({ _21229_, _06930_, _07066_, _21261_ }), .Y(_05533_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30326_ ( .A({ _21228_, _06930_, _07066_, _21260_ }), .Y(_05534_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30327_ ( .A({ _21227_, _06930_, _07066_, _21259_ }), .Y(_05535_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30328_ ( .A({ _21226_, _06930_, _07066_, _21258_ }), .Y(_05536_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30329_ ( .A({ _21225_, _06930_, _07066_, _21257_ }), .Y(_05537_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30330_ ( .A({ _21224_, _06930_, _07066_, _21256_ }), .Y(_05538_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30331_ ( .A({ _21254_, _06930_, _07066_, _21286_ }), .Y(_05539_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30332_ ( .A({ _21253_, _06930_, _07066_, _21285_ }), .Y(_05540_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30333_ ( .A({ _21252_, _06930_, _07066_, _21284_ }), .Y(_05541_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30334_ ( .A({ _21251_, _06930_, _07066_, _21283_ }), .Y(_05542_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30335_ ( .A({ _21250_, _06930_, _07066_, _21282_ }), .Y(_05543_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30336_ ( .A({ _21249_, _06930_, _07066_, _21281_ }), .Y(_05544_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30337_ ( .A({ _21248_, _06930_, _07066_, _21280_ }), .Y(_05545_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30338_ ( .A({ _21245_, _06930_, _07066_, _21277_ }), .Y(_05546_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30339_ ( .A({ _21234_, _06930_, _07066_, _21266_ }), .Y(_05547_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _30340_ ( .A({ _21223_, _06930_, _07066_, _21255_ }), .Y(_05548_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30341_ ( .A({ _05945_, _07085_ }), .Y(_24045_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30342_ ( .A({ _05945_, _15810_, _07085_ }), .Y(_15811_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _30343_ ( .A({ _05937_, _07372_ }), .Y(_24043_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30344_ ( .A({ _07373_, max_pool_serial_18_comp_fsm[2], max_pool_serial_18_comp_fsm[3] }), .Y(_07372_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30345_ ( .A({ max_pool_serial_18_comp_fsm[1], _07379_, _07374_ }), .Y(_07373_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30346_ ( .A({ max_pool_serial_18_comp_fsm[0], _07378_, _07375_ }), .Y(_07374_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30347_ ( .A({ _07377_, _07376_ }), .Y(_07375_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30348_ ( .A(max_pool_serial_18_comp_fsm[15:12]), .Y(_07376_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30349_ ( .A(max_pool_serial_18_comp_fsm[11:8]), .Y(_07377_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30350_ ( .A(max_pool_serial_18_comp_fsm[7:4]), .Y(_07378_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30351_ ( .A({ _07383_, _07382_, _07381_, _07380_ }), .Y(_07379_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30352_ ( .A(max_pool_serial_18_comp_fsm[23:20]), .Y(_07380_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30353_ ( .A(max_pool_serial_18_comp_fsm[19:16]), .Y(_07381_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30354_ ( .A(max_pool_serial_18_comp_fsm[31:28]), .Y(_07382_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30355_ ( .A(max_pool_serial_18_comp_fsm[27:24]), .Y(_07383_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _30356_ ( .A({ _07384_, max_pool_serial_18_comp_fsm[0], _07379_, max_pool_serial_18_comp_fsm[1] }), .Y(_05937_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30357_ ( .A({ _07378_, _07375_, max_pool_serial_18_comp_fsm[3:2] }), .Y(_07384_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30358_ ( .A({ _07391_, _07388_, _07385_ }), .Y(_24042_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30359_ ( .A({ _05726_, _05937_, _07386_, _07372_ }), .Y(_07385_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30360_ ( .A({ _07373_, max_pool_serial_18_comp_fsm[3:2] }), .Y(_07386_) );
  \$lut  #( .LUT(16'hefff), .WIDTH(4) ) _30361_ ( .A({ _07378_, _07387_, max_pool_serial_18_comp_fsm[3:2] }), .Y(_05726_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30362_ ( .A({ _07375_, _07379_, max_pool_serial_18_comp_fsm[1:0] }), .Y(_07387_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30363_ ( .A({ _05935_, _07389_ }), .Y(_07388_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _30364_ ( .A({ _07387_, max_pool_serial_18_comp_fsm[2], _07378_, max_pool_serial_18_comp_fsm[3] }), .Y(_05935_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30365_ ( .A({ max_pool_serial_18_comp_fsm[1], _07390_, _07379_, max_pool_serial_18_comp_fsm[0] }), .Y(_07389_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30366_ ( .A({ _07375_, max_pool_serial_18_comp_fsm[2], _07378_, max_pool_serial_18_comp_fsm[3] }), .Y(_07390_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30367_ ( .A({ _05936_, _05934_ }), .Y(_07391_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _30368_ ( .A({ max_pool_serial_18_comp_fsm[1], _07384_, _07379_, max_pool_serial_18_comp_fsm[0] }), .Y(_05934_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _30369_ ( .A({ _07390_, max_pool_serial_18_comp_fsm[0], _07379_, max_pool_serial_18_comp_fsm[1] }), .Y(_05936_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30370_ ( .A({ _07393_, _07392_ }), .Y(_15512_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _30371_ ( .A({ _07388_, _05936_, _05726_, _15576_ }), .Y(_07392_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30372_ ( .A({ _15480_, _07372_, _15544_, _07386_ }), .Y(_07393_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30373_ ( .A({ _07394_, _15487_, _07372_ }), .Y(_15519_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30374_ ( .A({ _15551_, _07386_, _15583_, _05726_ }), .Y(_07394_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _30375_ ( .A({ _07396_, _07395_ }), .Y(_15490_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _30376_ ( .A({ _07388_, _05934_, _05726_, _15554_ }), .Y(_07395_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30377_ ( .A({ _15458_, _07372_, _15522_, _07386_ }), .Y(_07396_) );
  \$lut  #( .LUT(16'h8fff), .WIDTH(4) ) _30378_ ( .A({ _07397_, _07398_, _07386_, _15533_ }), .Y(_15501_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _30379_ ( .A({ _07391_, _07372_, _15469_ }), .Y(_07397_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _30380_ ( .A({ _05937_, _07389_, _05726_, _15565_ }), .Y(_07398_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30381_ ( .A({ _07399_, _15547_, _07386_ }), .Y(_15515_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30382_ ( .A({ _15483_, _07372_, _15579_, _05726_ }), .Y(_07399_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30383_ ( .A({ _07400_, _15484_, _07372_ }), .Y(_15516_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30384_ ( .A({ _15548_, _07386_, _15580_, _05726_ }), .Y(_07400_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30385_ ( .A({ _07401_, _15525_, _07386_ }), .Y(_15493_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30386_ ( .A({ _15461_, _07372_, _15557_, _05726_ }), .Y(_07401_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30387_ ( .A({ _07402_, _15485_, _07372_ }), .Y(_15517_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30388_ ( .A({ _15549_, _07386_, _15581_, _05726_ }), .Y(_07402_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30389_ ( .A({ _07403_, _15550_, _07386_ }), .Y(_15518_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30390_ ( .A({ _15486_, _07372_, _15582_, _05726_ }), .Y(_07403_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30391_ ( .A({ _07404_, _15552_, _07386_ }), .Y(_15520_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30392_ ( .A({ _15488_, _07372_, _15584_, _05726_ }), .Y(_07404_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30393_ ( .A({ _07405_, _15553_, _07386_ }), .Y(_15521_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30394_ ( .A({ _15489_, _07372_, _15585_, _05726_ }), .Y(_07405_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30395_ ( .A({ _07406_, _15464_, _07372_ }), .Y(_15496_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30396_ ( .A({ _15528_, _07386_, _15560_, _05726_ }), .Y(_07406_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30397_ ( .A({ _07407_, _15523_, _07386_ }), .Y(_15491_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30398_ ( .A({ _15459_, _07372_, _15555_, _05726_ }), .Y(_07407_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30399_ ( .A({ _07408_, _15460_, _07372_ }), .Y(_15492_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30400_ ( .A({ _15524_, _07386_, _15556_, _05726_ }), .Y(_07408_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30401_ ( .A({ _07409_, _15462_, _07372_ }), .Y(_15494_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30402_ ( .A({ _15526_, _07386_, _15558_, _05726_ }), .Y(_07409_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30403_ ( .A({ _07410_, _15463_, _07372_ }), .Y(_15495_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30404_ ( .A({ _15527_, _07386_, _15559_, _05726_ }), .Y(_07410_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30405_ ( .A({ _07411_, _15471_, _07372_ }), .Y(_15503_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30406_ ( .A({ _15535_, _07386_, _15567_, _05726_ }), .Y(_07411_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30407_ ( .A({ _07412_, _15529_, _07386_ }), .Y(_15497_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30408_ ( .A({ _15465_, _07372_, _15561_, _05726_ }), .Y(_07412_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30409_ ( .A({ _07413_, _15530_, _07386_ }), .Y(_15498_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30410_ ( .A({ _15466_, _07372_, _15562_, _05726_ }), .Y(_07413_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30411_ ( .A({ _07414_, _15476_, _07372_ }), .Y(_15508_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30412_ ( .A({ _15540_, _07386_, _15572_, _05726_ }), .Y(_07414_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30413_ ( .A({ _07415_, _15467_, _07372_ }), .Y(_15499_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30414_ ( .A({ _15531_, _07386_, _15563_, _05726_ }), .Y(_07415_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30415_ ( .A({ _07416_, _15532_, _07386_ }), .Y(_15500_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30416_ ( .A({ _15468_, _07372_, _15564_, _05726_ }), .Y(_07416_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30417_ ( .A({ _07417_, _15470_, _07372_ }), .Y(_15502_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30418_ ( .A({ _15534_, _07386_, _15566_, _05726_ }), .Y(_07417_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30419_ ( .A({ _07418_, _15536_, _07386_ }), .Y(_15504_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30420_ ( .A({ _15472_, _07372_, _15568_, _05726_ }), .Y(_07418_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30421_ ( .A({ _07419_, _15537_, _07386_ }), .Y(_15505_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30422_ ( .A({ _15473_, _07372_, _15569_, _05726_ }), .Y(_07419_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30423_ ( .A({ _07420_, _15538_, _07386_ }), .Y(_15506_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30424_ ( .A({ _15474_, _07372_, _15570_, _05726_ }), .Y(_07420_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30425_ ( .A({ _07421_, _15475_, _07372_ }), .Y(_15507_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30426_ ( .A({ _15539_, _07386_, _15571_, _05726_ }), .Y(_07421_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30427_ ( .A({ _07422_, _15477_, _07372_ }), .Y(_15509_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30428_ ( .A({ _15541_, _07386_, _15573_, _05726_ }), .Y(_07422_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30429_ ( .A({ _07423_, _15542_, _07386_ }), .Y(_15510_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30430_ ( .A({ _15478_, _07372_, _15574_, _05726_ }), .Y(_07423_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30431_ ( .A({ _07424_, _15479_, _07372_ }), .Y(_15511_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30432_ ( .A({ _15543_, _07386_, _15575_, _05726_ }), .Y(_07424_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30433_ ( .A({ _07425_, _15545_, _07386_ }), .Y(_15513_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30434_ ( .A({ _15481_, _07372_, _15577_, _05726_ }), .Y(_07425_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30435_ ( .A({ _07426_, _15482_, _07372_ }), .Y(_15514_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30436_ ( .A({ _15546_, _07386_, _15578_, _05726_ }), .Y(_07426_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30437_ ( .A({ _15416_, _05932_, _15448_, _07438_ }), .Y(_15384_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30438_ ( .A({ _stream_max_pool_serial_18_source_1_source_pat_fsm_0[0], _07436_, _07427_ }), .Y(_05932_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30439_ ( .A({ _07428_, _stream_max_pool_serial_18_source_1_source_pat_fsm_0[1] }), .Y(_07427_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30440_ ( .A({ _07435_, _07434_, _07429_ }), .Y(_07428_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30441_ ( .A({ _07433_, _07432_, _07431_, _07430_ }), .Y(_07429_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30442_ ( .A(_stream_max_pool_serial_18_source_1_source_pat_fsm_0[23:20]), .Y(_07430_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30443_ ( .A(_stream_max_pool_serial_18_source_1_source_pat_fsm_0[19:16]), .Y(_07431_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30444_ ( .A(_stream_max_pool_serial_18_source_1_source_pat_fsm_0[31:28]), .Y(_07432_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30445_ ( .A(_stream_max_pool_serial_18_source_1_source_pat_fsm_0[27:24]), .Y(_07433_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30446_ ( .A(_stream_max_pool_serial_18_source_1_source_pat_fsm_0[15:12]), .Y(_07434_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30447_ ( .A(_stream_max_pool_serial_18_source_1_source_pat_fsm_0[11:8]), .Y(_07435_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30448_ ( .A({ _07437_, _stream_max_pool_serial_18_source_1_source_pat_fsm_0[3:2] }), .Y(_07436_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30449_ ( .A(_stream_max_pool_serial_18_source_1_source_pat_fsm_0[7:4]), .Y(_07437_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30450_ ( .A({ _07439_, _07427_ }), .Y(_07438_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30451_ ( .A({ _07436_, _stream_max_pool_serial_18_source_1_source_pat_fsm_0[0] }), .Y(_07439_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _30452_ ( .A({ _05933_, _05932_, _07438_ }), .Y(_24041_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _30453_ ( .A({ _stream_max_pool_serial_18_source_1_source_pat_fsm_0[1], _07439_, _07428_ }), .Y(_05933_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30454_ ( .A({ _15421_, _05932_, _15453_, _07438_ }), .Y(_15389_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30455_ ( .A({ _15394_, _05932_, _15426_, _07438_ }), .Y(_15362_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30456_ ( .A({ _15405_, _05932_, _15437_, _07438_ }), .Y(_15373_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30457_ ( .A({ _15419_, _05932_, _15451_, _07438_ }), .Y(_15387_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30458_ ( .A({ _15420_, _05932_, _15452_, _07438_ }), .Y(_15388_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30459_ ( .A({ _15396_, _05932_, _15428_, _07438_ }), .Y(_15364_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30460_ ( .A({ _15422_, _05932_, _15454_, _07438_ }), .Y(_15390_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30461_ ( .A({ _15423_, _05932_, _15455_, _07438_ }), .Y(_15391_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30462_ ( .A({ _15401_, _05932_, _15433_, _07438_ }), .Y(_15369_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30463_ ( .A({ _15424_, _05932_, _15456_, _07438_ }), .Y(_15392_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30464_ ( .A({ _15425_, _05932_, _15457_, _07438_ }), .Y(_15393_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30465_ ( .A({ _15395_, _05932_, _15427_, _07438_ }), .Y(_15363_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30466_ ( .A({ _15397_, _05932_, _15429_, _07438_ }), .Y(_15365_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30467_ ( .A({ _15398_, _05932_, _15430_, _07438_ }), .Y(_15366_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30468_ ( .A({ _15399_, _05932_, _15431_, _07438_ }), .Y(_15367_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30469_ ( .A({ _15410_, _05932_, _15442_, _07438_ }), .Y(_15378_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30470_ ( .A({ _15400_, _05932_, _15432_, _07438_ }), .Y(_15368_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30471_ ( .A({ _15402_, _05932_, _15434_, _07438_ }), .Y(_15370_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30472_ ( .A({ _15403_, _05932_, _15435_, _07438_ }), .Y(_15371_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30473_ ( .A({ _15404_, _05932_, _15436_, _07438_ }), .Y(_15372_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30474_ ( .A({ _15406_, _05932_, _15438_, _07438_ }), .Y(_15374_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30475_ ( .A({ _15407_, _05932_, _15439_, _07438_ }), .Y(_15375_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30476_ ( .A({ _15408_, _05932_, _15440_, _07438_ }), .Y(_15376_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30477_ ( .A({ _15409_, _05932_, _15441_, _07438_ }), .Y(_15377_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30478_ ( .A({ _15411_, _05932_, _15443_, _07438_ }), .Y(_15379_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30479_ ( .A({ _15412_, _05932_, _15444_, _07438_ }), .Y(_15380_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30480_ ( .A({ _15413_, _05932_, _15445_, _07438_ }), .Y(_15381_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30481_ ( .A({ _15414_, _05932_, _15446_, _07438_ }), .Y(_15382_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30482_ ( .A({ _15415_, _05932_, _15447_, _07438_ }), .Y(_15383_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30483_ ( .A({ _15417_, _05932_, _15449_, _07438_ }), .Y(_15385_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _30484_ ( .A({ _15418_, _05932_, _15450_, _07438_ }), .Y(_15386_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30485_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15288_, _15352_ }), .Y(_15320_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30486_ ( .A({ _07448_, _07447_, _07442_, _07440_ }), .Y(_24040_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30487_ ( .A({ _07441_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[31:29] }), .Y(_07440_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30488_ ( .A(_stream_max_pool_serial_18_sink_3_sink_fsm_1[28:25]), .Y(_07441_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30489_ ( .A({ _07446_, _07445_, _07444_, _07443_ }), .Y(_07442_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30490_ ( .A(_stream_max_pool_serial_18_sink_3_sink_fsm_1[8:5]), .Y(_07443_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30491_ ( .A(_stream_max_pool_serial_18_sink_3_sink_fsm_1[4:1]), .Y(_07444_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30492_ ( .A(_stream_max_pool_serial_18_sink_3_sink_fsm_1[16:13]), .Y(_07445_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30493_ ( .A(_stream_max_pool_serial_18_sink_3_sink_fsm_1[12:9]), .Y(_07446_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30494_ ( .A(_stream_max_pool_serial_18_sink_3_sink_fsm_1[24:21]), .Y(_07447_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30495_ ( .A(_stream_max_pool_serial_18_sink_3_sink_fsm_1[20:17]), .Y(_07448_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30496_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15266_, _15330_ }), .Y(_15298_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30497_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15277_, _15341_ }), .Y(_15309_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30498_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15293_, _15357_ }), .Y(_15325_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30499_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15291_, _15355_ }), .Y(_15323_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30500_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15292_, _15356_ }), .Y(_15324_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30501_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15294_, _15358_ }), .Y(_15326_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30502_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15295_, _15359_ }), .Y(_15327_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30503_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15296_, _15360_ }), .Y(_15328_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30504_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15268_, _15332_ }), .Y(_15300_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30505_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15269_, _15333_ }), .Y(_15301_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30506_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15297_, _15361_ }), .Y(_15329_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30507_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15267_, _15331_ }), .Y(_15299_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30508_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15270_, _15334_ }), .Y(_15302_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30509_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15271_, _15335_ }), .Y(_15303_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30510_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15272_, _15336_ }), .Y(_15304_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30511_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15275_, _15339_ }), .Y(_15307_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30512_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15276_, _15340_ }), .Y(_15308_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30513_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15281_, _15345_ }), .Y(_15313_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30514_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15273_, _15337_ }), .Y(_15305_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30515_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15274_, _15338_ }), .Y(_15306_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30516_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15278_, _15342_ }), .Y(_15310_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30517_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15279_, _15343_ }), .Y(_15311_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30518_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15280_, _15344_ }), .Y(_15312_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30519_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15284_, _15348_ }), .Y(_15316_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30520_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15282_, _15346_ }), .Y(_15314_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30521_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15283_, _15347_ }), .Y(_15315_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30522_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15285_, _15349_ }), .Y(_15317_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30523_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15286_, _15350_ }), .Y(_15318_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30524_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15287_, _15351_ }), .Y(_15319_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30525_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15289_, _15353_ }), .Y(_15321_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30526_ ( .A({ _24040_, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _15290_, _15354_ }), .Y(_15322_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30527_ ( .A({ _07449_, _04736_, _07453_ }), .Y(_22821_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30528_ ( .A({ _04640_, _07450_, _07452_, _04512_ }), .Y(_07449_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30529_ ( .A({ _06887_, _07451_, _06891_, main_fsm[4] }), .Y(_07450_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _30530_ ( .A({ main_fsm[3], main_fsm[0], main_fsm[2:1] }), .Y(_07451_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30531_ ( .A({ main_fsm[4], _06914_, _06898_, _06891_ }), .Y(_07452_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30532_ ( .A({ main_fsm[4], _06911_, _06891_, _06887_ }), .Y(_07453_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30533_ ( .A({ _07454_, _04511_, _07452_ }), .Y(_22820_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30534_ ( .A({ _04735_, _07453_, _07450_, _04639_ }), .Y(_07454_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30535_ ( .A({ _07499_, _07496_, _07481_, _07455_ }), .Y(_22085_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30536_ ( .A({ _07475_, _07456_, _07479_, _22245_ }), .Y(_07455_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30537_ ( .A({ _07469_, _07467_, _07462_, _07457_ }), .Y(_07456_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30538_ ( .A({ _22341_, _07458_, _07460_, _22373_ }), .Y(_07457_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30539_ ( .A({ _07067_, _07459_, _06923_, _06920_ }), .Y(_07458_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30540_ ( .A({ _06932_, control_conv2d_16[4] }), .Y(_07459_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30541_ ( .A({ _07461_, _07459_, _06923_, _06920_ }), .Y(_07460_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30542_ ( .A({ control_conv2d_16[1:0], _06919_ }), .Y(_07461_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30543_ ( .A({ _22117_, _07463_, _07465_, _22277_ }), .Y(_07462_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30544_ ( .A({ _07464_, _06931_, _06923_, _06920_ }), .Y(_07463_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30545_ ( .A({ control_conv2d_16[1], control_conv2d_16[2], control_conv2d_16[0], control_conv2d_16[3] }), .Y(_07464_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30546_ ( .A({ _07466_, _07459_, _06923_, _06920_ }), .Y(_07465_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _30547_ ( .A(control_conv2d_16[3:0]), .Y(_07466_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30548_ ( .A({ _22149_, _06930_, _22053_, _06008_ }), .Y(_07467_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30549_ ( .A({ _07468_, _06931_, _06923_, _06920_ }), .Y(_06008_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30550_ ( .A({ control_conv2d_16[1:0], control_conv2d_16[2], control_conv2d_16[3] }), .Y(_07468_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30551_ ( .A({ _22181_, _07470_, _07472_, _22309_ }), .Y(_07469_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30552_ ( .A({ _07471_, _07459_, _06923_, _06920_ }), .Y(_07470_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30553_ ( .A({ control_conv2d_16[1:0], control_conv2d_16[3:2] }), .Y(_07471_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30554_ ( .A({ _07473_, _07459_, _06923_, _06920_ }), .Y(_07472_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30555_ ( .A({ _07474_, control_conv2d_16[0], control_conv2d_16[1] }), .Y(_07473_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _30556_ ( .A(control_conv2d_16[3:2]), .Y(_07474_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30557_ ( .A({ _22213_, _07476_, _07478_, _22405_ }), .Y(_07475_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30558_ ( .A({ _07477_, _07459_, _06923_, _06920_ }), .Y(_07476_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30559_ ( .A({ control_conv2d_16[1], control_conv2d_16[2], control_conv2d_16[3], control_conv2d_16[0] }), .Y(_07477_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30560_ ( .A({ _07459_, _06923_, _06920_, _06918_ }), .Y(_07478_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30561_ ( .A({ _07480_, _07459_, _06923_, _06920_ }), .Y(_07479_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _30562_ ( .A({ control_conv2d_16[2], control_conv2d_16[0], control_conv2d_16[3], control_conv2d_16[1] }), .Y(_07480_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30563_ ( .A({ _07494_, _07491_, _07487_, _07482_ }), .Y(_07481_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30564_ ( .A({ _22437_, _07483_, _07485_, _22789_ }), .Y(_07482_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30565_ ( .A({ _07480_, _07484_ }), .Y(_07483_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30566_ ( .A({ control_conv2d_16[4], _06929_, _06923_, _06920_ }), .Y(_07484_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30567_ ( .A({ _07486_, _06928_, _06923_, _06920_ }), .Y(_07485_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30568_ ( .A({ _06919_, control_conv2d_16[1:0] }), .Y(_07486_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30569_ ( .A({ _22597_, _07488_, _22501_, _07489_ }), .Y(_07487_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30570_ ( .A({ _06918_, _07484_ }), .Y(_07488_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30571_ ( .A({ _07490_, _07484_ }), .Y(_07489_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30572_ ( .A({ control_conv2d_16[1:0], _07474_ }), .Y(_07490_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30573_ ( .A({ _22693_, _07492_, _22661_, _07493_ }), .Y(_07491_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30574_ ( .A({ _07468_, _06928_, _06923_, _06920_ }), .Y(_07492_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30575_ ( .A({ _07490_, _06928_, _06923_, _06920_ }), .Y(_07493_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30576_ ( .A({ _22757_, _06021_, _22725_, _07495_ }), .Y(_07494_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30577_ ( .A({ _07464_, _06928_, _06923_, _06920_ }), .Y(_07495_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30578_ ( .A({ _22469_, _07497_, _07498_, _22629_ }), .Y(_07496_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30579_ ( .A({ _07466_, _07484_ }), .Y(_07497_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30580_ ( .A({ _07480_, _06928_, _06923_, _06920_ }), .Y(_07498_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30581_ ( .A({ _22565_, _07500_, _22533_, _07501_ }), .Y(_07499_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30582_ ( .A({ _06933_, _07484_ }), .Y(_07500_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _30583_ ( .A({ _07464_, _07484_ }), .Y(_07501_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30584_ ( .A({ _07502_, _04733_, _07453_ }), .Y(_22818_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30585_ ( .A({ _04637_, _07450_, _07452_, _04509_ }), .Y(_07502_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30586_ ( .A({ _07503_, _04732_, _07453_ }), .Y(_22817_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30587_ ( .A({ _04636_, _07450_, _07452_, _04508_ }), .Y(_07503_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30588_ ( .A({ _07517_, _07516_, _07511_, _07504_ }), .Y(_22084_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30589_ ( .A({ _07510_, _07505_, _07478_, _22404_ }), .Y(_07504_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30590_ ( .A({ _07509_, _07508_, _07507_, _07506_ }), .Y(_07505_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30591_ ( .A({ _22148_, _06930_, _22052_, _06008_ }), .Y(_07506_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30592_ ( .A({ _22372_, _07460_, _22308_, _07472_ }), .Y(_07507_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30593_ ( .A({ _22340_, _07458_, _22116_, _07463_ }), .Y(_07508_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30594_ ( .A({ _22244_, _07479_, _22180_, _07470_ }), .Y(_07509_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30595_ ( .A({ _22212_, _07476_, _07465_, _22276_ }), .Y(_07510_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30596_ ( .A({ _07515_, _07514_, _07513_, _07512_ }), .Y(_07511_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30597_ ( .A({ _22500_, _07489_, _07498_, _22628_ }), .Y(_07512_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30598_ ( .A({ _22564_, _07500_, _07493_, _22660_ }), .Y(_07513_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30599_ ( .A({ _22596_, _07488_, _07495_, _22724_ }), .Y(_07514_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30600_ ( .A({ _22468_, _07497_, _22436_, _07483_ }), .Y(_07515_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30601_ ( .A({ _22532_, _07501_, _07492_, _22692_ }), .Y(_07516_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30602_ ( .A({ _22756_, _06021_, _07485_, _22788_ }), .Y(_07517_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30603_ ( .A({ _07518_, _04507_, _07452_ }), .Y(_22816_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30604_ ( .A({ _04731_, _07453_, _07450_, _04635_ }), .Y(_07518_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30605_ ( .A({ _07532_, _07531_, _07526_, _07519_ }), .Y(_22082_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30606_ ( .A({ _07525_, _07520_, _06930_, _22146_ }), .Y(_07519_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30607_ ( .A({ _07524_, _07523_, _07522_, _07521_ }), .Y(_07520_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30608_ ( .A({ _22370_, _07460_, _22274_, _07465_ }), .Y(_07521_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30609_ ( .A({ _22050_, _06008_, _07470_, _22178_ }), .Y(_07522_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30610_ ( .A({ _22242_, _07479_, _07478_, _22402_ }), .Y(_07523_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30611_ ( .A({ _22210_, _07476_, _07472_, _22306_ }), .Y(_07524_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30612_ ( .A({ _22338_, _07458_, _22114_, _07463_ }), .Y(_07525_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30613_ ( .A({ _07530_, _07529_, _07528_, _07527_ }), .Y(_07526_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30614_ ( .A({ _22466_, _07497_, _22434_, _07483_ }), .Y(_07527_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30615_ ( .A({ _22498_, _07489_, _07492_, _22690_ }), .Y(_07528_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30616_ ( .A({ _22722_, _07495_, _07485_, _22786_ }), .Y(_07529_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30617_ ( .A({ _22754_, _06021_, _22658_, _07493_ }), .Y(_07530_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30618_ ( .A({ _22562_, _07500_, _07498_, _22626_ }), .Y(_07531_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30619_ ( .A({ _22530_, _07501_, _07488_, _22594_ }), .Y(_07532_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30620_ ( .A({ _07533_, _04506_, _07452_ }), .Y(_22815_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30621_ ( .A({ _04730_, _07453_, _07450_, _04634_ }), .Y(_07533_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30622_ ( .A({ _07547_, _07546_, _07541_, _07534_ }), .Y(_22081_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30623_ ( .A({ _07540_, _07535_, _06930_, _22145_ }), .Y(_07534_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30624_ ( .A({ _07539_, _07538_, _07537_, _07536_ }), .Y(_07535_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30625_ ( .A({ _22241_, _07479_, _22209_, _07476_ }), .Y(_07536_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30626_ ( .A({ _22273_, _07465_, _22177_, _07470_ }), .Y(_07537_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30627_ ( .A({ _22401_, _07478_, _22305_, _07472_ }), .Y(_07538_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30628_ ( .A({ _22369_, _07460_, _22113_, _07463_ }), .Y(_07539_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30629_ ( .A({ _22337_, _07458_, _22049_, _06008_ }), .Y(_07540_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30630_ ( .A({ _07545_, _07544_, _07543_, _07542_ }), .Y(_07541_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30631_ ( .A({ _22433_, _07483_, _07489_, _22497_ }), .Y(_07542_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30632_ ( .A({ _22593_, _07488_, _07485_, _22785_ }), .Y(_07543_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30633_ ( .A({ _22753_, _06021_, _22721_, _07495_ }), .Y(_07544_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30634_ ( .A({ _22689_, _07492_, _22657_, _07493_ }), .Y(_07545_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30635_ ( .A({ _22529_, _07501_, _07498_, _22625_ }), .Y(_07546_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30636_ ( .A({ _22465_, _07497_, _07500_, _22561_ }), .Y(_07547_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30637_ ( .A({ _07548_, _04729_, _07453_ }), .Y(_22814_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30638_ ( .A({ _04633_, _07450_, _07452_, _04505_ }), .Y(_07548_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30639_ ( .A({ _07562_, _07561_, _07556_, _07549_ }), .Y(_22080_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _30640_ ( .A({ _07555_, _07550_, _06008_, _22048_ }), .Y(_07549_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30641_ ( .A({ _07554_, _07553_, _07552_, _07551_ }), .Y(_07550_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30642_ ( .A({ _22208_, _07476_, _07465_, _22272_ }), .Y(_07551_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30643_ ( .A({ _22240_, _07479_, _22176_, _07470_ }), .Y(_07552_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30644_ ( .A({ _22336_, _07458_, _22304_, _07472_ }), .Y(_07553_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30645_ ( .A({ _22400_, _07478_, _22368_, _07460_ }), .Y(_07554_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30646_ ( .A({ _22144_, _06930_, _22112_, _07463_ }), .Y(_07555_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30647_ ( .A({ _07560_, _07559_, _07558_, _07557_ }), .Y(_07556_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30648_ ( .A({ _22464_, _07497_, _07489_, _22496_ }), .Y(_07557_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30649_ ( .A({ _22432_, _07483_, _22752_, _06021_ }), .Y(_07558_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30650_ ( .A({ _22688_, _07492_, _22656_, _07493_ }), .Y(_07559_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30651_ ( .A({ _22624_, _07498_, _07485_, _22784_ }), .Y(_07560_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30652_ ( .A({ _22560_, _07500_, _07488_, _22592_ }), .Y(_07561_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30653_ ( .A({ _22528_, _07501_, _07495_, _22720_ }), .Y(_07562_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30654_ ( .A({ _07563_, _04503_, _07452_ }), .Y(_22812_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30655_ ( .A({ _04727_, _07453_, _07450_, _04631_ }), .Y(_07563_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30656_ ( .A({ _07564_, _04728_, _07453_ }), .Y(_22813_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30657_ ( .A({ _04632_, _07450_, _07452_, _04504_ }), .Y(_07564_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30658_ ( .A({ _07578_, _07577_, _07572_, _07565_ }), .Y(_22079_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30659_ ( .A({ _07571_, _07566_, _07458_, _22335_ }), .Y(_07565_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30660_ ( .A({ _07570_, _07569_, _07568_, _07567_ }), .Y(_07566_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30661_ ( .A({ _22399_, _07478_, _22111_, _07463_ }), .Y(_07567_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30662_ ( .A({ _22143_, _06930_, _07476_, _22207_ }), .Y(_07568_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30663_ ( .A({ _22239_, _07479_, _22047_, _06008_ }), .Y(_07569_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30664_ ( .A({ _22271_, _07465_, _22175_, _07470_ }), .Y(_07570_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30665_ ( .A({ _22367_, _07460_, _22303_, _07472_ }), .Y(_07571_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30666_ ( .A({ _07576_, _07575_, _07574_, _07573_ }), .Y(_07572_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30667_ ( .A({ _22495_, _07489_, _07495_, _22719_ }), .Y(_07573_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30668_ ( .A({ _22591_, _07488_, _07492_, _22687_ }), .Y(_07574_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30669_ ( .A({ _22431_, _07483_, _22751_, _06021_ }), .Y(_07575_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30670_ ( .A({ _22559_, _07500_, _22527_, _07501_ }), .Y(_07576_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30671_ ( .A({ _22463_, _07497_, _07493_, _22655_ }), .Y(_07577_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30672_ ( .A({ _22623_, _07498_, _07485_, _22783_ }), .Y(_07578_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30673_ ( .A({ _07579_, _04726_, _07453_ }), .Y(_22811_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30674_ ( .A({ _04630_, _07450_, _07452_, _04502_ }), .Y(_07579_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30675_ ( .A({ _07593_, _07592_, _07587_, _07580_ }), .Y(_22078_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30676_ ( .A({ _07586_, _07581_, _07478_, _22398_ }), .Y(_07580_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30677_ ( .A({ _07585_, _07584_, _07583_, _07582_ }), .Y(_07581_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30678_ ( .A({ _22366_, _07460_, _22302_, _07472_ }), .Y(_07582_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30679_ ( .A({ _22142_, _06930_, _07465_, _22270_ }), .Y(_07583_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30680_ ( .A({ _22206_, _07476_, _07458_, _22334_ }), .Y(_07584_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30681_ ( .A({ _22238_, _07479_, _22174_, _07470_ }), .Y(_07585_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30682_ ( .A({ _22110_, _07463_, _22046_, _06008_ }), .Y(_07586_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30683_ ( .A({ _07591_, _07590_, _07589_, _07588_ }), .Y(_07587_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30684_ ( .A({ _22526_, _07501_, _22430_, _07483_ }), .Y(_07588_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30685_ ( .A({ _22462_, _07497_, _22750_, _06021_ }), .Y(_07589_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30686_ ( .A({ _22686_, _07492_, _22654_, _07493_ }), .Y(_07590_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30687_ ( .A({ _22622_, _07498_, _07485_, _22782_ }), .Y(_07591_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30688_ ( .A({ _22558_, _07500_, _22494_, _07489_ }), .Y(_07592_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30689_ ( .A({ _22590_, _07488_, _07495_, _22718_ }), .Y(_07593_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30690_ ( .A({ _07594_, _04725_, _07453_ }), .Y(_22810_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30691_ ( .A({ _04629_, _07450_, _07452_, _04501_ }), .Y(_07594_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30692_ ( .A({ _07608_, _07607_, _07602_, _07595_ }), .Y(_22077_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30693_ ( .A({ _07601_, _07596_, _06930_, _22141_ }), .Y(_07595_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30694_ ( .A({ _07600_, _07599_, _07598_, _07597_ }), .Y(_07596_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30695_ ( .A({ _22237_, _07479_, _22109_, _07463_ }), .Y(_07597_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30696_ ( .A({ _22205_, _07476_, _07458_, _22333_ }), .Y(_07598_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30697_ ( .A({ _22269_, _07465_, _07472_, _22301_ }), .Y(_07599_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30698_ ( .A({ _22397_, _07478_, _22365_, _07460_ }), .Y(_07600_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30699_ ( .A({ _22045_, _06008_, _07470_, _22173_ }), .Y(_07601_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30700_ ( .A({ _07606_, _07605_, _07604_, _07603_ }), .Y(_07602_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30701_ ( .A({ _22493_, _07489_, _07495_, _22717_ }), .Y(_07603_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30702_ ( .A({ _22429_, _07483_, _07485_, _22781_ }), .Y(_07604_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30703_ ( .A({ _22557_, _07500_, _07493_, _22653_ }), .Y(_07605_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30704_ ( .A({ _22749_, _06021_, _22685_, _07492_ }), .Y(_07606_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30705_ ( .A({ _22525_, _07501_, _07498_, _22621_ }), .Y(_07607_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30706_ ( .A({ _22461_, _07497_, _07488_, _22589_ }), .Y(_07608_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30707_ ( .A({ _07609_, _04500_, _07452_ }), .Y(_22809_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30708_ ( .A({ _04724_, _07453_, _07450_, _04628_ }), .Y(_07609_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30709_ ( .A({ _07623_, _07622_, _07617_, _07610_ }), .Y(_22076_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30710_ ( .A({ _07616_, _07611_, _07463_, _22108_ }), .Y(_07610_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30711_ ( .A({ _07615_, _07614_, _07613_, _07612_ }), .Y(_07611_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30712_ ( .A({ _22268_, _07465_, _22044_, _06008_ }), .Y(_07612_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30713_ ( .A({ _22332_, _07458_, _07460_, _22364_ }), .Y(_07613_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30714_ ( .A({ _22236_, _07479_, _07472_, _22300_ }), .Y(_07614_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30715_ ( .A({ _22204_, _07476_, _22172_, _07470_ }), .Y(_07615_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30716_ ( .A({ _22140_, _06930_, _07478_, _22396_ }), .Y(_07616_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30717_ ( .A({ _07621_, _07620_, _07619_, _07618_ }), .Y(_07617_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30718_ ( .A({ _22492_, _07489_, _07485_, _22780_ }), .Y(_07618_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30719_ ( .A({ _22428_, _07483_, _07488_, _22588_ }), .Y(_07619_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30720_ ( .A({ _22620_, _07498_, _07493_, _22652_ }), .Y(_07620_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30721_ ( .A({ _22684_, _07492_, _07495_, _22716_ }), .Y(_07621_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30722_ ( .A({ _22524_, _07501_, _22748_, _06021_ }), .Y(_07622_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30723_ ( .A({ _22460_, _07497_, _07500_, _22556_ }), .Y(_07623_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30724_ ( .A({ _07624_, _04722_, _07453_ }), .Y(_22807_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30725_ ( .A({ _04626_, _07450_, _07452_, _04498_ }), .Y(_07624_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30726_ ( .A({ _07638_, _07637_, _07632_, _07625_ }), .Y(_22075_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _30727_ ( .A({ _07631_, _07626_, _06008_, _22043_ }), .Y(_07625_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30728_ ( .A({ _07630_, _07629_, _07628_, _07627_ }), .Y(_07626_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30729_ ( .A({ _22363_, _07460_, _22299_, _07472_ }), .Y(_07627_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30730_ ( .A({ _22331_, _07458_, _22171_, _07470_ }), .Y(_07628_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30731_ ( .A({ _22139_, _06930_, _07479_, _22235_ }), .Y(_07629_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30732_ ( .A({ _22107_, _07463_, _07465_, _22267_ }), .Y(_07630_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30733_ ( .A({ _22203_, _07476_, _07478_, _22395_ }), .Y(_07631_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30734_ ( .A({ _07636_, _07635_, _07634_, _07633_ }), .Y(_07632_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30735_ ( .A({ _22459_, _07497_, _07495_, _22715_ }), .Y(_07633_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30736_ ( .A({ _22587_, _07488_, _07485_, _22779_ }), .Y(_07634_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30737_ ( .A({ _22555_, _07500_, _22523_, _07501_ }), .Y(_07635_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30738_ ( .A({ _22747_, _06021_, _22683_, _07492_ }), .Y(_07636_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30739_ ( .A({ _22491_, _07489_, _07498_, _22619_ }), .Y(_07637_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30740_ ( .A({ _22427_, _07483_, _07493_, _22651_ }), .Y(_07638_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30741_ ( .A({ _07639_, _04720_, _07453_ }), .Y(_22805_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30742_ ( .A({ _04624_, _07450_, _07452_, _04496_ }), .Y(_07639_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30743_ ( .A({ _07640_, _04721_, _07453_ }), .Y(_22806_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30744_ ( .A({ _04625_, _07450_, _07452_, _04497_ }), .Y(_07640_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30745_ ( .A({ _07654_, _07653_, _07648_, _07641_ }), .Y(_22074_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30746_ ( .A({ _07647_, _07642_, _07458_, _22330_ }), .Y(_07641_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30747_ ( .A({ _07646_, _07645_, _07644_, _07643_ }), .Y(_07642_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30748_ ( .A({ _22234_, _07479_, _07465_, _22266_ }), .Y(_07643_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30749_ ( .A({ _22138_, _06930_, _22106_, _07463_ }), .Y(_07644_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30750_ ( .A({ _22170_, _07470_, _07472_, _22298_ }), .Y(_07645_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30751_ ( .A({ _22202_, _07476_, _22042_, _06008_ }), .Y(_07646_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30752_ ( .A({ _22394_, _07478_, _22362_, _07460_ }), .Y(_07647_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30753_ ( .A({ _07652_, _07651_, _07650_, _07649_ }), .Y(_07648_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30754_ ( .A({ _22522_, _07501_, _07492_, _22682_ }), .Y(_07649_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30755_ ( .A({ _22554_, _07500_, _07493_, _22650_ }), .Y(_07650_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30756_ ( .A({ _22426_, _07483_, _07488_, _22586_ }), .Y(_07651_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30757_ ( .A({ _22458_, _07497_, _07498_, _22618_ }), .Y(_07652_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30758_ ( .A({ _22490_, _07489_, _07495_, _22714_ }), .Y(_07653_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30759_ ( .A({ _22746_, _06021_, _07485_, _22778_ }), .Y(_07654_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30760_ ( .A({ _07655_, _04719_, _07453_ }), .Y(_22804_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30761_ ( .A({ _04623_, _07450_, _07452_, _04495_ }), .Y(_07655_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30762_ ( .A({ _07669_, _07668_, _07663_, _07656_ }), .Y(_22073_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30763_ ( .A({ _07662_, _07657_, _07463_, _22105_ }), .Y(_07656_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30764_ ( .A({ _07661_, _07660_, _07659_, _07658_ }), .Y(_07657_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30765_ ( .A({ _22265_, _07465_, _22041_, _06008_ }), .Y(_07658_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30766_ ( .A({ _22329_, _07458_, _22169_, _07470_ }), .Y(_07659_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30767_ ( .A({ _22233_, _07479_, _07460_, _22361_ }), .Y(_07660_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30768_ ( .A({ _22201_, _07476_, _07472_, _22297_ }), .Y(_07661_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30769_ ( .A({ _22137_, _06930_, _07478_, _22393_ }), .Y(_07662_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30770_ ( .A({ _07667_, _07666_, _07665_, _07664_ }), .Y(_07663_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30771_ ( .A({ _22553_, _07500_, _22489_, _07489_ }), .Y(_07664_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30772_ ( .A({ _22585_, _07488_, _07492_, _22681_ }), .Y(_07665_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30773_ ( .A({ _22745_, _06021_, _22649_, _07493_ }), .Y(_07666_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30774_ ( .A({ _22617_, _07498_, _07485_, _22777_ }), .Y(_07667_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30775_ ( .A({ _22457_, _07497_, _07501_, _22521_ }), .Y(_07668_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30776_ ( .A({ _22425_, _07483_, _07495_, _22713_ }), .Y(_07669_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30777_ ( .A({ _07670_, _04718_, _07453_ }), .Y(_22803_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30778_ ( .A({ _04622_, _07450_, _07452_, _04494_ }), .Y(_07670_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30779_ ( .A({ _07684_, _07683_, _07678_, _07671_ }), .Y(_22071_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30780_ ( .A({ _07677_, _07672_, _06930_, _22135_ }), .Y(_07671_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30781_ ( .A({ _07676_, _07675_, _07674_, _07673_ }), .Y(_07672_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30782_ ( .A({ _22231_, _07479_, _07478_, _22391_ }), .Y(_07673_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30783_ ( .A({ _22327_, _07458_, _22103_, _07463_ }), .Y(_07674_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30784_ ( .A({ _22263_, _07465_, _22039_, _06008_ }), .Y(_07675_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30785_ ( .A({ _22167_, _07470_, _07472_, _22295_ }), .Y(_07676_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30786_ ( .A({ _22199_, _07476_, _07460_, _22359_ }), .Y(_07677_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30787_ ( .A({ _07682_, _07681_, _07680_, _07679_ }), .Y(_07678_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30788_ ( .A({ _22455_, _07497_, _07500_, _22551_ }), .Y(_07679_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30789_ ( .A({ _22423_, _07483_, _07489_, _22487_ }), .Y(_07680_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30790_ ( .A({ _22583_, _07488_, _07498_, _22615_ }), .Y(_07681_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30791_ ( .A({ _22743_, _06021_, _22647_, _07493_ }), .Y(_07682_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30792_ ( .A({ _22519_, _07501_, _07492_, _22679_ }), .Y(_07683_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30793_ ( .A({ _22711_, _07495_, _07485_, _22775_ }), .Y(_07684_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30794_ ( .A({ _07685_, _04717_, _07453_ }), .Y(_22802_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30795_ ( .A({ _04621_, _07450_, _07452_, _04493_ }), .Y(_07685_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30796_ ( .A({ _07699_, _07698_, _07693_, _07686_ }), .Y(_22070_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30797_ ( .A({ _07692_, _07687_, _07479_, _22230_ }), .Y(_07686_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30798_ ( .A({ _07691_, _07690_, _07689_, _07688_ }), .Y(_07687_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30799_ ( .A({ _22134_, _06930_, _07465_, _22262_ }), .Y(_07688_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30800_ ( .A({ _22390_, _07478_, _22038_, _06008_ }), .Y(_07689_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30801_ ( .A({ _22198_, _07476_, _22166_, _07470_ }), .Y(_07690_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30802_ ( .A({ _22102_, _07463_, _07472_, _22294_ }), .Y(_07691_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30803_ ( .A({ _22326_, _07458_, _07460_, _22358_ }), .Y(_07692_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30804_ ( .A({ _07697_, _07696_, _07695_, _07694_ }), .Y(_07693_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30805_ ( .A({ _22518_, _07501_, _07498_, _22614_ }), .Y(_07694_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30806_ ( .A({ _22422_, _07483_, _07488_, _22582_ }), .Y(_07695_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30807_ ( .A({ _22646_, _07493_, _07485_, _22774_ }), .Y(_07696_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30808_ ( .A({ _22742_, _06021_, _22678_, _07492_ }), .Y(_07697_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30809_ ( .A({ _22550_, _07500_, _07495_, _22710_ }), .Y(_07698_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30810_ ( .A({ _22454_, _07497_, _07489_, _22486_ }), .Y(_07699_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30811_ ( .A({ _07700_, _04492_, _07452_ }), .Y(_22801_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30812_ ( .A({ _04716_, _07453_, _07450_, _04620_ }), .Y(_07700_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30813_ ( .A({ _07714_, _07713_, _07708_, _07701_ }), .Y(_22069_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30814_ ( .A({ _07707_, _07702_, _06930_, _22133_ }), .Y(_07701_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30815_ ( .A({ _07706_, _07705_, _07704_, _07703_ }), .Y(_07702_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30816_ ( .A({ _22229_, _07479_, _07460_, _22357_ }), .Y(_07703_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30817_ ( .A({ _22389_, _07478_, _22165_, _07470_ }), .Y(_07704_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30818_ ( .A({ _22325_, _07458_, _22261_, _07465_ }), .Y(_07705_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30819_ ( .A({ _22197_, _07476_, _07472_, _22293_ }), .Y(_07706_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30820_ ( .A({ _22101_, _07463_, _22037_, _06008_ }), .Y(_07707_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30821_ ( .A({ _07712_, _07711_, _07710_, _07709_ }), .Y(_07708_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30822_ ( .A({ _22549_, _07500_, _07488_, _22581_ }), .Y(_07709_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30823_ ( .A({ _22517_, _07501_, _07492_, _22677_ }), .Y(_07710_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30824_ ( .A({ _22741_, _06021_, _22613_, _07498_ }), .Y(_07711_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30825_ ( .A({ _22709_, _07495_, _07485_, _22773_ }), .Y(_07712_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30826_ ( .A({ _22453_, _07497_, _22421_, _07483_ }), .Y(_07713_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30827_ ( .A({ _22485_, _07489_, _07493_, _22645_ }), .Y(_07714_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30828_ ( .A({ _07715_, _04490_, _07452_ }), .Y(_22799_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30829_ ( .A({ _04714_, _07453_, _07450_, _04618_ }), .Y(_07715_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30830_ ( .A({ _07716_, _04713_, _07453_ }), .Y(_22798_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30831_ ( .A({ _04617_, _07450_, _07452_, _04489_ }), .Y(_07716_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30832_ ( .A({ _07717_, _04491_, _07452_ }), .Y(_22800_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30833_ ( .A({ _04715_, _07453_, _07450_, _04619_ }), .Y(_07717_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30834_ ( .A({ _07731_, _07730_, _07725_, _07718_ }), .Y(_22068_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30835_ ( .A({ _07724_, _07719_, _07463_, _22100_ }), .Y(_07718_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30836_ ( .A({ _07723_, _07722_, _07721_, _07720_ }), .Y(_07719_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30837_ ( .A({ _22164_, _07470_, _07472_, _22292_ }), .Y(_07720_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30838_ ( .A({ _22196_, _07476_, _22036_, _06008_ }), .Y(_07721_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30839_ ( .A({ _22324_, _07458_, _07460_, _22356_ }), .Y(_07722_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30840_ ( .A({ _22228_, _07479_, _07478_, _22388_ }), .Y(_07723_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30841_ ( .A({ _22132_, _06930_, _07465_, _22260_ }), .Y(_07724_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30842_ ( .A({ _07729_, _07728_, _07727_, _07726_ }), .Y(_07725_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30843_ ( .A({ _22452_, _07497_, _07500_, _22548_ }), .Y(_07726_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30844_ ( .A({ _22484_, _07489_, _07492_, _22676_ }), .Y(_07727_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30845_ ( .A({ _22740_, _06021_, _22708_, _07495_ }), .Y(_07728_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30846_ ( .A({ _22612_, _07498_, _07485_, _22772_ }), .Y(_07729_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30847_ ( .A({ _22420_, _07483_, _07493_, _22644_ }), .Y(_07730_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30848_ ( .A({ _22516_, _07501_, _07488_, _22580_ }), .Y(_07731_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30849_ ( .A({ _07732_, _04743_, _07453_ }), .Y(_22828_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30850_ ( .A({ _04647_, _07450_, _07452_, _04519_ }), .Y(_07732_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30851_ ( .A({ _07746_, _07745_, _07740_, _07733_ }), .Y(_22067_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30852_ ( .A({ _07739_, _07734_, _07460_, _22355_ }), .Y(_07733_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30853_ ( .A({ _07738_, _07737_, _07736_, _07735_ }), .Y(_07734_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30854_ ( .A({ _22131_, _06930_, _07479_, _22227_ }), .Y(_07735_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30855_ ( .A({ _22099_, _07463_, _07470_, _22163_ }), .Y(_07736_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30856_ ( .A({ _22387_, _07478_, _22035_, _06008_ }), .Y(_07737_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30857_ ( .A({ _22195_, _07476_, _07472_, _22291_ }), .Y(_07738_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30858_ ( .A({ _22323_, _07458_, _22259_, _07465_ }), .Y(_07739_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30859_ ( .A({ _07744_, _07743_, _07742_, _07741_ }), .Y(_07740_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30860_ ( .A({ _22579_, _07488_, _22739_, _06021_ }), .Y(_07741_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30861_ ( .A({ _22451_, _07497_, _07498_, _22611_ }), .Y(_07742_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30862_ ( .A({ _22547_, _07500_, _07493_, _22643_ }), .Y(_07743_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30863_ ( .A({ _22707_, _07495_, _07485_, _22771_ }), .Y(_07744_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30864_ ( .A({ _22483_, _07489_, _07492_, _22675_ }), .Y(_07745_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30865_ ( .A({ _22515_, _07501_, _22419_, _07483_ }), .Y(_07746_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30866_ ( .A({ _07747_, _04742_, _07453_ }), .Y(_22827_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30867_ ( .A({ _04646_, _07450_, _07452_, _04518_ }), .Y(_07747_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30868_ ( .A({ _07761_, _07760_, _07755_, _07748_ }), .Y(_22066_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30869_ ( .A({ _07754_, _07749_, _07463_, _22098_ }), .Y(_07748_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30870_ ( .A({ _07753_, _07752_, _07751_, _07750_ }), .Y(_07749_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30871_ ( .A({ _22386_, _07478_, _22034_, _06008_ }), .Y(_07750_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30872_ ( .A({ _22162_, _07470_, _07472_, _22290_ }), .Y(_07751_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30873_ ( .A({ _22226_, _07479_, _07458_, _22322_ }), .Y(_07752_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30874_ ( .A({ _22354_, _07460_, _22258_, _07465_ }), .Y(_07753_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30875_ ( .A({ _22130_, _06930_, _07476_, _22194_ }), .Y(_07754_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30876_ ( .A({ _07759_, _07758_, _07757_, _07756_ }), .Y(_07755_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30877_ ( .A({ _22514_, _07501_, _07498_, _22610_ }), .Y(_07756_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30878_ ( .A({ _22546_, _07500_, _07488_, _22578_ }), .Y(_07757_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30879_ ( .A({ _22674_, _07492_, _07495_, _22706_ }), .Y(_07758_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30880_ ( .A({ _22738_, _06021_, _07485_, _22770_ }), .Y(_07759_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30881_ ( .A({ _22450_, _07497_, _07489_, _22482_ }), .Y(_07760_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30882_ ( .A({ _22418_, _07483_, _07493_, _22642_ }), .Y(_07761_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30883_ ( .A({ _07762_, _04517_, _07452_ }), .Y(_22826_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30884_ ( .A({ _04741_, _07453_, _07450_, _04645_ }), .Y(_07762_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30885_ ( .A({ _07776_, _07775_, _07770_, _07763_ }), .Y(_22065_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30886_ ( .A({ _07769_, _07764_, _07460_, _22353_ }), .Y(_07763_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30887_ ( .A({ _07768_, _07767_, _07766_, _07765_ }), .Y(_07764_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30888_ ( .A({ _22225_, _07479_, _22033_, _06008_ }), .Y(_07765_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30889_ ( .A({ _22257_, _07465_, _22161_, _07470_ }), .Y(_07766_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30890_ ( .A({ _22129_, _06930_, _07478_, _22385_ }), .Y(_07767_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30891_ ( .A({ _22321_, _07458_, _22097_, _07463_ }), .Y(_07768_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30892_ ( .A({ _22193_, _07476_, _07472_, _22289_ }), .Y(_07769_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30893_ ( .A({ _07774_, _07773_, _07772_, _07771_ }), .Y(_07770_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30894_ ( .A({ _22513_, _07501_, _22417_, _07483_ }), .Y(_07771_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30895_ ( .A({ _22545_, _07500_, _07495_, _22705_ }), .Y(_07772_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30896_ ( .A({ _22449_, _07497_, _07485_, _22769_ }), .Y(_07773_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30897_ ( .A({ _22609_, _07498_, _07493_, _22641_ }), .Y(_07774_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30898_ ( .A({ _22577_, _07488_, _22737_, _06021_ }), .Y(_07775_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30899_ ( .A({ _22481_, _07489_, _07492_, _22673_ }), .Y(_07776_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30900_ ( .A({ _07777_, _04740_, _07453_ }), .Y(_22825_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30901_ ( .A({ _04644_, _07450_, _07452_, _04516_ }), .Y(_07777_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30902_ ( .A({ _07778_, _04739_, _07453_ }), .Y(_22824_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30903_ ( .A({ _04643_, _07450_, _07452_, _04515_ }), .Y(_07778_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30904_ ( .A({ _07792_, _07791_, _07786_, _07779_ }), .Y(_22064_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _30905_ ( .A({ _07785_, _07780_, _06008_, _22032_ }), .Y(_07779_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30906_ ( .A({ _07784_, _07783_, _07782_, _07781_ }), .Y(_07780_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30907_ ( .A({ _22224_, _07479_, _07460_, _22352_ }), .Y(_07781_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30908_ ( .A({ _22192_, _07476_, _07465_, _22256_ }), .Y(_07782_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30909_ ( .A({ _22128_, _06930_, _07470_, _22160_ }), .Y(_07783_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30910_ ( .A({ _22384_, _07478_, _22320_, _07458_ }), .Y(_07784_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30911_ ( .A({ _22096_, _07463_, _07472_, _22288_ }), .Y(_07785_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30912_ ( .A({ _07790_, _07789_, _07788_, _07787_ }), .Y(_07786_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30913_ ( .A({ _22512_, _07501_, _07492_, _22672_ }), .Y(_07787_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30914_ ( .A({ _22544_, _07500_, _07493_, _22640_ }), .Y(_07788_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30915_ ( .A({ _22416_, _07483_, _07485_, _22768_ }), .Y(_07789_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30916_ ( .A({ _22448_, _07497_, _07488_, _22576_ }), .Y(_07790_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30917_ ( .A({ _22480_, _07489_, _07498_, _22608_ }), .Y(_07791_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30918_ ( .A({ _22736_, _06021_, _22704_, _07495_ }), .Y(_07792_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _30919_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18705_, _18737_ }), .Y(_18673_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _30920_ ( .A({ _07794_, _07802_, _stream_conv2d_16_source_22_source_pat_fsm_5[1] }), .Y(_07793_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _30921_ ( .A({ _07801_, _07800_, _07795_ }), .Y(_07794_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30922_ ( .A({ _07799_, _07798_, _07797_, _07796_ }), .Y(_07795_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30923_ ( .A(_stream_conv2d_16_source_22_source_pat_fsm_5[23:20]), .Y(_07796_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30924_ ( .A(_stream_conv2d_16_source_22_source_pat_fsm_5[19:16]), .Y(_07797_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30925_ ( .A(_stream_conv2d_16_source_22_source_pat_fsm_5[31:28]), .Y(_07798_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30926_ ( .A(_stream_conv2d_16_source_22_source_pat_fsm_5[27:24]), .Y(_07799_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30927_ ( .A(_stream_conv2d_16_source_22_source_pat_fsm_5[15:12]), .Y(_07800_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30928_ ( .A(_stream_conv2d_16_source_22_source_pat_fsm_5[11:8]), .Y(_07801_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _30929_ ( .A({ _07803_, _stream_conv2d_16_source_22_source_pat_fsm_5[3:2] }), .Y(_07802_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _30930_ ( .A(_stream_conv2d_16_source_22_source_pat_fsm_5[7:4]), .Y(_07803_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30931_ ( .A({ _07804_, _04738_, _07453_ }), .Y(_22823_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30932_ ( .A({ _04642_, _07450_, _07452_, _04514_ }), .Y(_07804_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30933_ ( .A({ _07805_, _04737_, _07453_ }), .Y(_22822_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30934_ ( .A({ _04641_, _07450_, _07452_, _04513_ }), .Y(_07805_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30935_ ( .A({ _07819_, _07818_, _07813_, _07806_ }), .Y(_22063_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30936_ ( .A({ _07812_, _07807_, _07472_, _22287_ }), .Y(_07806_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30937_ ( .A({ _07811_, _07810_, _07809_, _07808_ }), .Y(_07807_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30938_ ( .A({ _22191_, _07476_, _22159_, _07470_ }), .Y(_07808_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30939_ ( .A({ _22319_, _07458_, _07460_, _22351_ }), .Y(_07809_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30940_ ( .A({ _22127_, _06930_, _22095_, _07463_ }), .Y(_07810_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30941_ ( .A({ _22223_, _07479_, _07478_, _22383_ }), .Y(_07811_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30942_ ( .A({ _22255_, _07465_, _22031_, _06008_ }), .Y(_07812_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30943_ ( .A({ _07817_, _07816_, _07815_, _07814_ }), .Y(_07813_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30944_ ( .A({ _22447_, _07497_, _07485_, _22767_ }), .Y(_07814_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30945_ ( .A({ _22479_, _07489_, _07495_, _22703_ }), .Y(_07815_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30946_ ( .A({ _22415_, _07483_, _07488_, _22575_ }), .Y(_07816_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30947_ ( .A({ _22543_, _07500_, _22511_, _07501_ }), .Y(_07817_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30948_ ( .A({ _22671_, _07492_, _22639_, _07493_ }), .Y(_07818_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30949_ ( .A({ _22735_, _06021_, _22607_, _07498_ }), .Y(_07819_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30950_ ( .A({ _07820_, _04734_, _07453_ }), .Y(_22819_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30951_ ( .A({ _04638_, _07450_, _07452_, _04510_ }), .Y(_07820_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30952_ ( .A({ _07821_, _04499_, _07452_ }), .Y(_22808_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30953_ ( .A({ _04723_, _07453_, _07450_, _04627_ }), .Y(_07821_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30954_ ( .A({ _07835_, _07834_, _07829_, _07822_ }), .Y(_22062_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _30955_ ( .A({ _07828_, _07823_, _06008_, _22030_ }), .Y(_07822_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30956_ ( .A({ _07827_, _07826_, _07825_, _07824_ }), .Y(_07823_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30957_ ( .A({ _22318_, _07458_, _07460_, _22350_ }), .Y(_07824_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30958_ ( .A({ _22190_, _07476_, _22158_, _07470_ }), .Y(_07825_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30959_ ( .A({ _22382_, _07478_, _22286_, _07472_ }), .Y(_07826_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30960_ ( .A({ _22222_, _07479_, _22094_, _07463_ }), .Y(_07827_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30961_ ( .A({ _22126_, _06930_, _07465_, _22254_ }), .Y(_07828_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30962_ ( .A({ _07833_, _07832_, _07831_, _07830_ }), .Y(_07829_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30963_ ( .A({ _22414_, _07483_, _07493_, _22638_ }), .Y(_07830_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30964_ ( .A({ _22478_, _07489_, _22734_, _06021_ }), .Y(_07831_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30965_ ( .A({ _22574_, _07488_, _07492_, _22670_ }), .Y(_07832_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30966_ ( .A({ _22606_, _07498_, _07495_, _22702_ }), .Y(_07833_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30967_ ( .A({ _22446_, _07497_, _07500_, _22542_ }), .Y(_07834_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30968_ ( .A({ _22510_, _07501_, _07485_, _22766_ }), .Y(_07835_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _30969_ ( .A({ _07836_, _04712_, _07453_ }), .Y(_22797_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30970_ ( .A({ _04616_, _07450_, _07452_, _04488_ }), .Y(_07836_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30971_ ( .A({ _07850_, _07849_, _07844_, _07837_ }), .Y(_22092_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30972_ ( .A({ _07843_, _07838_, _07458_, _22348_ }), .Y(_07837_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30973_ ( .A({ _07842_, _07841_, _07840_, _07839_ }), .Y(_07838_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30974_ ( .A({ _22252_, _07479_, _22220_, _07476_ }), .Y(_07839_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30975_ ( .A({ _22156_, _06930_, _07465_, _22284_ }), .Y(_07840_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30976_ ( .A({ _22060_, _06008_, _07472_, _22316_ }), .Y(_07841_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30977_ ( .A({ _22124_, _07463_, _07470_, _22188_ }), .Y(_07842_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30978_ ( .A({ _22412_, _07478_, _22380_, _07460_ }), .Y(_07843_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30979_ ( .A({ _07848_, _07847_, _07846_, _07845_ }), .Y(_07844_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30980_ ( .A({ _22572_, _07500_, _22540_, _07501_ }), .Y(_07845_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30981_ ( .A({ _22444_, _07483_, _07488_, _22604_ }), .Y(_07846_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30982_ ( .A({ _22508_, _07489_, _07498_, _22636_ }), .Y(_07847_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30983_ ( .A({ _22700_, _07492_, _22668_, _07493_ }), .Y(_07848_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30984_ ( .A({ _22476_, _07497_, _07495_, _22732_ }), .Y(_07849_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30985_ ( .A({ _22764_, _06021_, _07485_, _22796_ }), .Y(_07850_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _30986_ ( .A({ _07864_, _07863_, _07858_, _07851_ }), .Y(_22091_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _30987_ ( .A({ _07857_, _07852_, _06930_, _22155_ }), .Y(_07851_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30988_ ( .A({ _07856_, _07855_, _07854_, _07853_ }), .Y(_07852_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30989_ ( .A({ _22251_, _07479_, _07460_, _22379_ }), .Y(_07853_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30990_ ( .A({ _22411_, _07478_, _22283_, _07465_ }), .Y(_07854_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30991_ ( .A({ _22219_, _07476_, _07458_, _22347_ }), .Y(_07855_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30992_ ( .A({ _22187_, _07470_, _07472_, _22315_ }), .Y(_07856_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _30993_ ( .A({ _22123_, _07463_, _22059_, _06008_ }), .Y(_07857_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _30994_ ( .A({ _07862_, _07861_, _07860_, _07859_ }), .Y(_07858_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30995_ ( .A({ _22507_, _07489_, _07485_, _22795_ }), .Y(_07859_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30996_ ( .A({ _22539_, _07501_, _07488_, _22603_ }), .Y(_07860_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _30997_ ( .A({ _22763_, _06021_, _22731_, _07495_ }), .Y(_07861_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30998_ ( .A({ _22699_, _07492_, _22667_, _07493_ }), .Y(_07862_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _30999_ ( .A({ _22571_, _07500_, _22443_, _07483_ }), .Y(_07863_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31000_ ( .A({ _22475_, _07497_, _07498_, _22635_ }), .Y(_07864_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31001_ ( .A({ _07878_, _07877_, _07872_, _07865_ }), .Y(_22090_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _31002_ ( .A({ _07871_, _07866_, _07463_, _22122_ }), .Y(_07865_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31003_ ( .A({ _07870_, _07869_, _07868_, _07867_ }), .Y(_07866_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31004_ ( .A({ _22058_, _06008_, _07470_, _22186_ }), .Y(_07867_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31005_ ( .A({ _22218_, _07476_, _07465_, _22282_ }), .Y(_07868_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31006_ ( .A({ _22346_, _07458_, _22314_, _07472_ }), .Y(_07869_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31007_ ( .A({ _22410_, _07478_, _22378_, _07460_ }), .Y(_07870_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31008_ ( .A({ _22154_, _06930_, _07479_, _22250_ }), .Y(_07871_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31009_ ( .A({ _07876_, _07875_, _07874_, _07873_ }), .Y(_07872_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31010_ ( .A({ _22602_, _07488_, _22506_, _07489_ }), .Y(_07873_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31011_ ( .A({ _22538_, _07501_, _07493_, _22666_ }), .Y(_07874_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31012_ ( .A({ _22442_, _07483_, _07492_, _22698_ }), .Y(_07875_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31013_ ( .A({ _22762_, _06021_, _22634_, _07498_ }), .Y(_07876_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31014_ ( .A({ _22474_, _07497_, _07495_, _22730_ }), .Y(_07877_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31015_ ( .A({ _22570_, _07500_, _07485_, _22794_ }), .Y(_07878_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _31016_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18799_, _18831_ }), .Y(_18767_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31017_ ( .A({ _07880_, _07888_, _stream_conv2d_16_source_21_source_pat_fsm_4[1] }), .Y(_07879_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31018_ ( .A({ _07887_, _07886_, _07881_ }), .Y(_07880_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31019_ ( .A({ _07885_, _07884_, _07883_, _07882_ }), .Y(_07881_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31020_ ( .A(_stream_conv2d_16_source_21_source_pat_fsm_4[23:20]), .Y(_07882_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31021_ ( .A(_stream_conv2d_16_source_21_source_pat_fsm_4[19:16]), .Y(_07883_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31022_ ( .A(_stream_conv2d_16_source_21_source_pat_fsm_4[31:28]), .Y(_07884_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31023_ ( .A(_stream_conv2d_16_source_21_source_pat_fsm_4[27:24]), .Y(_07885_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31024_ ( .A(_stream_conv2d_16_source_21_source_pat_fsm_4[15:12]), .Y(_07886_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31025_ ( .A(_stream_conv2d_16_source_21_source_pat_fsm_4[11:8]), .Y(_07887_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _31026_ ( .A({ _07889_, _stream_conv2d_16_source_21_source_pat_fsm_4[3:2] }), .Y(_07888_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31027_ ( .A(_stream_conv2d_16_source_21_source_pat_fsm_4[7:4]), .Y(_07889_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _31028_ ( .A({ _07452_, _07450_, _07453_ }), .Y(_24077_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31029_ ( .A({ _07903_, _07902_, _07897_, _07890_ }), .Y(_22089_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _31030_ ( .A({ _07896_, _07891_, _06008_, _22057_ }), .Y(_07890_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31031_ ( .A({ _07895_, _07894_, _07893_, _07892_ }), .Y(_07891_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31032_ ( .A({ _22153_, _06930_, _07472_, _22313_ }), .Y(_07892_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31033_ ( .A({ _22249_, _07479_, _22217_, _07476_ }), .Y(_07893_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31034_ ( .A({ _22345_, _07458_, _07460_, _22377_ }), .Y(_07894_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31035_ ( .A({ _22409_, _07478_, _22281_, _07465_ }), .Y(_07895_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31036_ ( .A({ _22121_, _07463_, _07470_, _22185_ }), .Y(_07896_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31037_ ( .A({ _07901_, _07900_, _07899_, _07898_ }), .Y(_07897_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31038_ ( .A({ _22473_, _07497_, _07501_, _22537_ }), .Y(_07898_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31039_ ( .A({ _22569_, _07500_, _07493_, _22665_ }), .Y(_07899_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31040_ ( .A({ _22761_, _06021_, _22633_, _07498_ }), .Y(_07900_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31041_ ( .A({ _22729_, _07495_, _07485_, _22793_ }), .Y(_07901_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31042_ ( .A({ _22601_, _07488_, _07492_, _22697_ }), .Y(_07902_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31043_ ( .A({ _22441_, _07483_, _07489_, _22505_ }), .Y(_07903_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31044_ ( .A({ _07471_, _07484_ }), .Y(_06012_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _31045_ ( .A({ _07905_, _07464_, _06933_ }), .Y(_07904_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31046_ ( .A({ _07459_, _06923_, _06920_ }), .Y(_07905_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _31047_ ( .A({ _07907_, _06008_, _22056_ }), .Y(_07906_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _31048_ ( .A({ _07066_, _07905_, _07908_ }), .Y(_07907_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _31049_ ( .A({ _07474_, control_conv2d_16[1:0] }), .Y(_07908_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31050_ ( .A({ control_conv2d_16[1], _07474_, control_conv2d_16[0] }), .Y(_07909_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31051_ ( .A({ _22344_, _07458_, _22120_, _07463_ }), .Y(_07910_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31052_ ( .A({ _22152_, _06930_, _07479_, _22248_ }), .Y(_07911_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31053_ ( .A({ _07921_, _07914_, _07913_ }), .Y(_07912_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31054_ ( .A({ _22536_, _07501_, _07493_, _22664_ }), .Y(_07913_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31055_ ( .A({ _07919_, _07917_, _07916_, _07915_ }), .Y(_07914_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31056_ ( .A({ _22408_, _07478_, _22312_, _07472_ }), .Y(_07915_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31057_ ( .A({ _22216_, _07476_, _07465_, _22280_ }), .Y(_07916_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31058_ ( .A({ _06919_, _07918_ }), .Y(_07917_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31059_ ( .A({ _06931_, _06923_, _06920_ }), .Y(_07918_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31060_ ( .A({ _07920_, _07905_, _22184_, _07470_ }), .Y(_07919_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31061_ ( .A({ _06919_, control_conv2d_16[1] }), .Y(_07920_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31062_ ( .A({ _22632_, _07498_, _07495_, _22728_ }), .Y(_07921_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31063_ ( .A({ _07926_, _07925_, _07924_, _07923_ }), .Y(_07922_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31064_ ( .A({ _22440_, _07483_, _07485_, _22792_ }), .Y(_07923_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31065_ ( .A({ _22472_, _07497_, _07489_, _22504_ }), .Y(_07924_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31066_ ( .A({ _22568_, _07500_, _07488_, _22600_ }), .Y(_07925_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31067_ ( .A({ _22760_, _06021_, _22696_, _07492_ }), .Y(_07926_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31068_ ( .A({ _07940_, _07937_, _07934_, _13052_ }), .Y(_22087_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31069_ ( .A({ _22343_, _07458_, _07460_, _22375_ }), .Y(_07927_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31070_ ( .A({ _22247_, _07479_, _22183_, _07470_ }), .Y(_07928_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31071_ ( .A({ _22055_, _06008_, _07472_, _22311_ }), .Y(_07929_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31072_ ( .A({ _07471_, _07930_ }), .Y(_06016_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31073_ ( .A({ _06928_, _06923_, _06920_ }), .Y(_07930_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31074_ ( .A({ _07067_, _07461_ }), .Y(_07931_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31075_ ( .A({ _07909_, _07484_ }), .Y(_07932_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31076_ ( .A({ _22215_, _07476_, _07465_, _22279_ }), .Y(_07933_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _31077_ ( .A({ _07935_, _07936_, _07497_, _22471_ }), .Y(_07934_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _31078_ ( .A({ _06013_, _07066_, _07500_, _22567_ }), .Y(_07935_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31079_ ( .A({ _07477_, _07484_ }), .Y(_06013_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _31080_ ( .A({ _07484_, _07908_, _07473_ }), .Y(_07936_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _31081_ ( .A({ _07938_, _07939_, _07488_, _22599_ }), .Y(_07937_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31082_ ( .A({ _22535_, _07501_, _22439_, _07483_ }), .Y(_07938_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31083_ ( .A({ _22151_, _06930_, _22119_, _07463_ }), .Y(_07939_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _31084_ ( .A({ _07942_, _07941_, _07498_, _22631_ }), .Y(_07940_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31085_ ( .A({ _22503_, _07489_, _07495_, _22727_ }), .Y(_07941_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31086_ ( .A({ _07944_, _07943_ }), .Y(_07942_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31087_ ( .A({ _22695_, _07492_, _07485_, _22791_ }), .Y(_07943_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31088_ ( .A({ _22759_, _06021_, _22663_, _07493_ }), .Y(_07944_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31089_ ( .A({ _07949_, _07948_, _07947_, _07946_ }), .Y(_07945_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31090_ ( .A({ _22246_, _07479_, _07460_, _22374_ }), .Y(_07946_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31091_ ( .A({ _22214_, _07476_, _07472_, _22310_ }), .Y(_07947_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31092_ ( .A({ _22054_, _06008_, _07484_, _07909_ }), .Y(_07948_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31093_ ( .A({ _22150_, _06930_, _07458_, _22342_ }), .Y(_07949_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31094_ ( .A({ _07468_, _07484_ }), .Y(_06015_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31095_ ( .A({ _07909_, _07930_ }), .Y(_07950_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31096_ ( .A({ _22278_, _07465_, _22182_, _07470_ }), .Y(_07951_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31097_ ( .A({ _22406_, _07478_, _22118_, _07463_ }), .Y(_07952_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31098_ ( .A({ _07954_, _07493_, _22662_ }), .Y(_07953_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _31099_ ( .A({ _07930_, _07466_, _07477_ }), .Y(_07954_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31100_ ( .A({ _22470_, _07497_, _22438_, _07483_ }), .Y(_07955_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31101_ ( .A({ _22630_, _07498_ }), .Y(_07956_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _31102_ ( .A({ _07959_, _07958_, _07488_, _22598_ }), .Y(_07957_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31103_ ( .A({ _22726_, _07495_ }), .Y(_07958_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31104_ ( .A({ _22694_, _07492_, _07485_, _22790_ }), .Y(_07959_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31105_ ( .A({ _22566_, _07500_, _22534_, _07501_ }), .Y(_07960_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31106_ ( .A({ _07979_, _07977_, _07972_, _07961_ }), .Y(_22083_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31107_ ( .A({ _07971_, _07970_, _07965_, _07962_ }), .Y(_07961_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31108_ ( .A({ _07964_, _07963_, _07904_ }), .Y(_07962_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31109_ ( .A({ _07461_, _07918_, _07490_, _07905_ }), .Y(_07963_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31110_ ( .A({ _22211_, _07476_, _07484_, _07931_ }), .Y(_07964_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31111_ ( .A({ _07969_, _07968_, _07967_, _07966_ }), .Y(_07965_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31112_ ( .A({ _22051_, _06008_ }), .Y(_07966_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31113_ ( .A({ _22339_, _07458_, _22115_, _07463_ }), .Y(_07967_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31114_ ( .A({ _07461_, _07930_, _22243_, _07479_ }), .Y(_07968_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31115_ ( .A({ _22275_, _07465_, _07472_, _22307_ }), .Y(_07969_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31116_ ( .A({ _22371_, _07460_, _22179_, _07470_ }), .Y(_07970_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31117_ ( .A({ _22147_, _06930_, _07478_, _22403_ }), .Y(_07971_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31118_ ( .A({ _07976_, _07975_, _07973_ }), .Y(_07972_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31119_ ( .A({ _06013_, _07974_, _07954_, _07066_ }), .Y(_07973_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31120_ ( .A({ _22755_, _06021_, _22659_, _07493_ }), .Y(_07974_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31121_ ( .A({ _22627_, _07498_, _07495_, _22723_ }), .Y(_07975_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31122_ ( .A({ _22691_, _07492_, _07485_, _22787_ }), .Y(_07976_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31123_ ( .A({ _07978_, _07501_, _22531_ }), .Y(_07977_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31124_ ( .A({ _22595_, _07488_, _22499_, _07489_ }), .Y(_07978_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _31125_ ( .A({ _07980_, _07981_, _07497_, _22467_ }), .Y(_07979_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31126_ ( .A({ _22563_, _07500_, _22435_, _07483_ }), .Y(_07980_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _31127_ ( .A({ _07930_, _07067_, _06933_ }), .Y(_07981_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _31128_ ( .A({ _07984_, _07983_, _07458_, _22328_ }), .Y(_07982_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _31129_ ( .A({ _07905_, _07464_, _07909_ }), .Y(_07983_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31130_ ( .A({ _22136_, _06930_, _22104_, _07463_ }), .Y(_07984_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31131_ ( .A({ _07477_, _07930_ }), .Y(_06017_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _31132_ ( .A({ _07950_, _07478_, _22392_ }), .Y(_07985_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31133_ ( .A({ _07991_, _07989_, _07988_, _07987_ }), .Y(_07986_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31134_ ( .A({ _22200_, _07476_, _07460_, _22360_ }), .Y(_07987_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31135_ ( .A({ _22264_, _07465_, _07472_, _22296_ }), .Y(_07988_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31136_ ( .A({ _07990_, _07930_, _22040_, _06008_ }), .Y(_07989_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _31137_ ( .A({ control_conv2d_16[0], control_conv2d_16[1], control_conv2d_16[2], control_conv2d_16[3] }), .Y(_07990_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31138_ ( .A({ _22232_, _07479_, _22168_, _07470_ }), .Y(_07991_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31139_ ( .A({ _22520_, _07501_, _07488_, _22584_ }), .Y(_07992_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _31140_ ( .A({ _06013_, _07932_, _07500_, _22552_ }), .Y(_07993_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31141_ ( .A({ _22648_, _07493_ }), .Y(_07994_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31142_ ( .A({ _22456_, _07497_, _07485_, _22776_ }), .Y(_07995_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31143_ ( .A({ _08000_, _07997_, _07998_, _07999_ }), .Y(_07996_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31144_ ( .A({ _22424_, _07483_, _07492_, _22680_ }), .Y(_07997_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31145_ ( .A({ _22488_, _07489_, _22744_, _06021_ }), .Y(_07998_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31146_ ( .A({ control_conv2d_16[0], _07920_, _07484_ }), .Y(_07999_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31147_ ( .A({ _22616_, _07498_, _07495_, _22712_ }), .Y(_08000_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31148_ ( .A({ _08005_, _08004_, _08003_, _08002_ }), .Y(_08001_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31149_ ( .A({ _22189_, _07476_ }), .Y(_08002_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31150_ ( .A({ _22125_, _06930_, _22029_, _06008_ }), .Y(_08003_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31151_ ( .A({ _22093_, _07463_, _07472_, _22285_ }), .Y(_08004_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31152_ ( .A({ _22317_, _07458_, _07460_, _22349_ }), .Y(_08005_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31153_ ( .A({ _22221_, _07479_, _07478_, _22381_ }), .Y(_08006_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31154_ ( .A({ _22253_, _07465_, _22157_, _07470_ }), .Y(_08007_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31155_ ( .A({ _08013_, _08012_, _08010_, _08009_ }), .Y(_08008_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31156_ ( .A({ _22413_, _07483_, _07492_, _22669_ }), .Y(_08009_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31157_ ( .A({ _08011_, _07907_, _06014_, _07950_ }), .Y(_08010_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31158_ ( .A({ _07908_, _07484_ }), .Y(_06014_) );
  \$lut  #( .LUT(16'h035f), .WIDTH(4) ) _31159_ ( .A({ _07486_, _07918_, _07905_, _06918_ }), .Y(_08011_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31160_ ( .A({ _07954_, _06013_, _07932_ }), .Y(_08012_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31161_ ( .A({ _22733_, _06021_, _22605_, _07498_ }), .Y(_08013_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31162_ ( .A({ _08018_, _08017_, _08016_, _08015_ }), .Y(_08014_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31163_ ( .A({ _22477_, _07489_, _07495_, _22701_ }), .Y(_08015_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31164_ ( .A({ _22541_, _07500_, _22509_, _07501_ }), .Y(_08016_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31165_ ( .A({ _22445_, _07497_, _07488_, _22573_ }), .Y(_08017_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31166_ ( .A({ _22637_, _07493_, _07485_, _22765_ }), .Y(_08018_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _31167_ ( .A({ _05978_, _07879_ }), .Y(_24065_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _31168_ ( .A({ _stream_conv2d_16_source_21_source_pat_fsm_4[1], _07880_, _07888_, _stream_conv2d_16_source_21_source_pat_fsm_4[0] }), .Y(_05978_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _31169_ ( .A({ _05924_, _08019_, _08045_, _08048_ }), .Y(_24039_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31170_ ( .A({ _08039_, _08037_, _24037_ }), .Y(_08019_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _31171_ ( .A({ _13755_, _24038_ }), .Y(_24037_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _31172_ ( .A({ _05929_, _08032_ }), .Y(_24038_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _31173_ ( .A({ _08020_, _08029_, _08025_, control_matmul_29[4] }), .Y(_05929_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31174_ ( .A({ _08024_, _08023_, _08022_, _08021_ }), .Y(_08020_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31175_ ( .A(control_matmul_29[23:20]), .Y(_08021_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31176_ ( .A(control_matmul_29[19:16]), .Y(_08022_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31177_ ( .A(control_matmul_29[31:28]), .Y(_08023_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31178_ ( .A(control_matmul_29[27:24]), .Y(_08024_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31179_ ( .A({ _08026_, _08028_, _08027_, control_matmul_29[5] }), .Y(_08025_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31180_ ( .A(control_matmul_29[15:12]), .Y(_08026_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31181_ ( .A(control_matmul_29[7:6]), .Y(_08027_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31182_ ( .A(control_matmul_29[11:8]), .Y(_08028_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31183_ ( .A({ _08031_, _08030_ }), .Y(_08029_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _31184_ ( .A(control_matmul_29[3:2]), .Y(_08030_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31185_ ( .A(control_matmul_29[1:0]), .Y(_08031_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31186_ ( .A({ _08020_, _08034_, _08033_, control_matmul_29[4] }), .Y(_08032_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31187_ ( .A({ control_matmul_29[5], _08028_, _08027_, _08026_ }), .Y(_08033_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31188_ ( .A({ control_matmul_29[2], control_matmul_29[3], control_matmul_29[0], control_matmul_29[1] }), .Y(_08034_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31189_ ( .A({ _08035_, _08033_, _08020_, control_matmul_29[4] }), .Y(_13755_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31190_ ( .A({ _08036_, control_matmul_29[2], control_matmul_29[3] }), .Y(_08035_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31191_ ( .A({ control_matmul_29[0], control_matmul_29[1] }), .Y(_08036_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31192_ ( .A({ _08030_, _08038_ }), .Y(_08037_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31193_ ( .A({ _08020_, _08033_, control_matmul_29[4] }), .Y(_08038_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31194_ ( .A({ _05926_, _05928_, _08041_, _08040_ }), .Y(_08039_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31195_ ( .A({ _08020_, _08034_, _08025_, control_matmul_29[4] }), .Y(_08040_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31196_ ( .A({ control_matmul_29[4], _08029_, _08025_, _08020_ }), .Y(_08041_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _31197_ ( .A({ _08020_, _08042_, _08025_, control_matmul_29[4] }), .Y(_05928_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _31198_ ( .A({ _08043_, control_matmul_29[0], control_matmul_29[1] }), .Y(_08042_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31199_ ( .A(control_matmul_29[3:2]), .Y(_08043_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31200_ ( .A({ control_matmul_29[4], _08044_, _08025_, _08020_ }), .Y(_05926_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31201_ ( .A({ _08031_, control_matmul_29[2], control_matmul_29[3] }), .Y(_08044_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _31202_ ( .A({ _08046_, _08051_, _08058_ }), .Y(_08045_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _31203_ ( .A({ _08055_, _08052_, _08050_, _08047_ }), .Y(_08046_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31204_ ( .A({ _08049_, _08048_ }), .Y(_08047_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31205_ ( .A({ _08020_, _08025_, control_matmul_29[4] }), .Y(_08048_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31206_ ( .A({ _08030_, _08036_ }), .Y(_08049_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31207_ ( .A({ _08043_, _08031_, _08051_ }), .Y(_08050_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31208_ ( .A({ control_matmul_29[4], _08025_, _08020_ }), .Y(_08051_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31209_ ( .A({ _08020_, _08053_, _08025_, control_matmul_29[4] }), .Y(_08052_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31210_ ( .A({ _08043_, _08054_ }), .Y(_08053_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31211_ ( .A({ control_matmul_29[0], control_matmul_29[1] }), .Y(_08054_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31212_ ( .A({ _08020_, _08044_, _08033_, control_matmul_29[4] }), .Y(_08055_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _31213_ ( .A({ _08030_, control_matmul_29[0], control_matmul_29[1] }), .Y(_08056_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31214_ ( .A({ _08054_, _08030_ }), .Y(_08057_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31215_ ( .A({ _08020_, _08056_, _08025_, control_matmul_29[4] }), .Y(_08058_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31216_ ( .A({ _08060_, _08048_ }), .Y(_08059_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31217_ ( .A({ _08054_, control_matmul_29[2], control_matmul_29[3] }), .Y(_08060_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31218_ ( .A({ _08043_, _08031_, _08048_ }), .Y(_08061_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31219_ ( .A({ control_matmul_29[4], _08034_, _08025_, _08020_ }), .Y(_08062_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31220_ ( .A({ control_matmul_29[4], _08049_, _08025_, _08020_ }), .Y(_08063_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _31221_ ( .A({ _08057_, _08048_ }), .Y(_05931_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31222_ ( .A({ _08020_, _08044_, _08025_, control_matmul_29[4] }), .Y(_08064_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31223_ ( .A({ control_matmul_29[4], _08025_, _08020_, _08035_ }), .Y(_08065_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _31224_ ( .A({ _08020_, _08060_, _08033_, control_matmul_29[4] }), .Y(_05924_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31225_ ( .A(control_matmul_29[3:2]), .Y(_08066_) );
  \$lut  #( .LUT(16'h9fff), .WIDTH(4) ) _31226_ ( .A({ _08036_, _08048_, control_matmul_29[3:2] }), .Y(_08067_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31227_ ( .A({ _08066_, _08051_, control_matmul_29[0], control_matmul_29[1] }), .Y(_08068_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31228_ ( .A({ _08066_, _08036_, _08051_ }), .Y(_08069_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31229_ ( .A({ _08066_, _08031_, _08051_ }), .Y(_08070_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31230_ ( .A({ _08066_, _08054_, _08051_ }), .Y(_08071_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _31231_ ( .A({ _08084_, _08079_, _08072_ }), .Y(_14722_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31232_ ( .A({ _08078_, _08076_, _08073_ }), .Y(_08072_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _31233_ ( .A({ _08075_, _08074_, _08064_, _15170_ }), .Y(_08073_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31234_ ( .A({ _15202_, _05929_, _15234_, _08058_ }), .Y(_08074_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _31235_ ( .A({ _08051_, _08043_, control_matmul_29[0] }), .Y(_08075_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31236_ ( .A({ _14946_, _08077_, _15042_, _08063_ }), .Y(_08076_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31237_ ( .A({ _08043_, _08036_, _08051_ }), .Y(_08077_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31238_ ( .A({ _15138_, _08059_, _08062_, _15010_ }), .Y(_08078_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _31239_ ( .A({ _08083_, _08080_, _13755_, _14786_ }), .Y(_08079_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _31240_ ( .A({ _08082_, _08081_, _08065_, _14978_ }), .Y(_08080_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31241_ ( .A({ _08048_, _08066_, control_matmul_29[0] }), .Y(_08081_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31242_ ( .A({ _15106_, _08052_, _14690_, _05924_ }), .Y(_08082_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31243_ ( .A({ 1'h1, _08032_, _08055_, _14754_ }), .Y(_08083_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31244_ ( .A({ _08091_, _08088_, _08087_, _08085_ }), .Y(_08084_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31245_ ( .A({ _15074_, _08086_ }), .Y(_08085_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31246_ ( .A({ _08066_, _08036_, _08048_ }), .Y(_08086_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31247_ ( .A({ _14850_, _08070_, _08071_, _14818_ }), .Y(_08087_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _31248_ ( .A({ _08089_, _08039_, _08061_ }), .Y(_08088_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _31249_ ( .A({ _08090_, _08038_, _08051_ }), .Y(_08089_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _31250_ ( .A({ _08030_, control_matmul_29[0] }), .Y(_08090_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31251_ ( .A({ _14882_, _08069_, _14914_, _08068_ }), .Y(_08091_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _31252_ ( .A({ _08105_, _08103_, _08092_ }), .Y(_14733_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31253_ ( .A({ _08098_, _08095_, _08094_, _08093_ }), .Y(_08092_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31254_ ( .A({ _15149_, _08059_, _08062_, _15021_ }), .Y(_08093_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31255_ ( .A({ _14957_, _08077_, _15053_, _08063_ }), .Y(_08094_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31256_ ( .A({ _08097_, _08096_, _08067_ }), .Y(_08095_) );
  \$lut  #( .LUT(16'h035f), .WIDTH(4) ) _31257_ ( .A({ _08029_, _08038_, _08051_, _08049_ }), .Y(_08096_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31258_ ( .A({ 1'h0, _08032_, _15117_, _08052_ }), .Y(_08097_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31259_ ( .A({ _08102_, _08101_, _08100_, _08099_ }), .Y(_08098_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31260_ ( .A({ _15181_, _08064_ }), .Y(_08099_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31261_ ( .A({ _14765_, _08055_, _14701_, _05924_ }), .Y(_08100_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31262_ ( .A({ _14797_, _13755_, _15245_, _08058_ }), .Y(_08101_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31263_ ( .A({ _15213_, _05929_, _08065_, _14989_ }), .Y(_08102_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31264_ ( .A({ _08104_, _08068_, _14925_ }), .Y(_08103_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31265_ ( .A({ _14829_, _08071_, _15085_, _08086_ }), .Y(_08104_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _31266_ ( .A({ _08107_, _08106_, _08070_, _14861_ }), .Y(_08105_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31267_ ( .A({ _05926_, _08061_, _08050_, _08047_ }), .Y(_08106_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31268_ ( .A({ _14893_, _08069_, _08081_, control_matmul_29[1] }), .Y(_08107_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31269_ ( .A({ _08112_, _08111_, _08110_, _08109_ }), .Y(_08108_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31270_ ( .A({ _15160_, _08059_, _08032_, 1'h1 }), .Y(_08109_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31271_ ( .A({ _14968_, _08077_, _15000_, _08065_ }), .Y(_08110_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31272_ ( .A({ _14808_, _13755_, _15256_, _08058_ }), .Y(_08111_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31273_ ( .A({ _15128_, _08052_, _14712_, _05924_ }), .Y(_08112_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31274_ ( .A({ _08115_, _08114_ }), .Y(_08113_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31275_ ( .A({ _14904_, _08069_, _08071_, _14840_ }), .Y(_08114_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31276_ ( .A({ _14936_, _08068_, _15096_, _08086_ }), .Y(_08115_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31277_ ( .A({ _05926_, _08048_, _08035_ }), .Y(_08116_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _31278_ ( .A({ _08081_, _08064_, _15192_ }), .Y(_08117_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31279_ ( .A({ _08120_, _08119_ }), .Y(_08118_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31280_ ( .A({ _15032_, _08062_, _15064_, _08063_ }), .Y(_08119_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31281_ ( .A({ _15224_, _05929_, _08055_, _14776_ }), .Y(_08120_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _31282_ ( .A({ _08123_, _08122_, _08064_, _15195_ }), .Y(_08121_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31283_ ( .A({ _14971_, _08077_, _08032_, 1'h0 }), .Y(_08122_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31284_ ( .A({ _08127_, _08126_, _08125_, _08124_ }), .Y(_08123_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31285_ ( .A({ _14811_, _13755_, _15067_, _08063_ }), .Y(_08124_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _31286_ ( .A({ _15227_, _05929_, _14715_, _05924_ }), .Y(_08125_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31287_ ( .A({ _15131_, _08052_, _08065_, _15003_ }), .Y(_08126_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31288_ ( .A({ _14779_, _08055_, _15035_, _08062_ }), .Y(_08127_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _31289_ ( .A({ _08081_, _08058_, _15259_ }), .Y(_08128_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _31290_ ( .A({ _08051_, _08060_, _08053_ }), .Y(_08129_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31291_ ( .A({ _14875_, _08070_, _08071_, _14843_ }), .Y(_08130_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31292_ ( .A({ _14939_, _08068_, _15099_, _08086_ }), .Y(_08131_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31293_ ( .A({ _08146_, _08145_, _08138_, _08132_ }), .Y(_14748_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31294_ ( .A({ _08137_, _08136_, _08134_, _08133_ }), .Y(_08132_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31295_ ( .A({ _15164_, _08059_, _08062_, _15036_ }), .Y(_08133_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _31296_ ( .A({ _08135_, _08064_, _15196_ }), .Y(_08134_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31297_ ( .A({ _08066_, _08054_, _08048_ }), .Y(_08135_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31298_ ( .A({ _14972_, _08077_, _13755_, _14812_ }), .Y(_08136_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31299_ ( .A({ _15228_, _05929_, _08055_, _14780_ }), .Y(_08137_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31300_ ( .A({ _08143_, _08141_, _08140_, _08139_ }), .Y(_08138_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31301_ ( .A({ _14876_, _08070_, _08071_, _14844_ }), .Y(_08139_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31302_ ( .A({ _14908_, _08069_, _15100_, _08086_ }), .Y(_08140_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31303_ ( .A({ _08142_, _08129_, _08075_ }), .Y(_08141_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31304_ ( .A({ _15004_, _08065_, _15068_, _08063_ }), .Y(_08142_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31305_ ( .A({ _08144_, _08068_, _14940_ }), .Y(_08143_) );
  \$lut  #( .LUT(16'h01ff), .WIDTH(4) ) _31306_ ( .A({ _08051_, _08057_, _08090_, _08044_ }), .Y(_08144_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31307_ ( .A({ _15260_, _08058_, _08052_, _15132_ }), .Y(_08145_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31308_ ( .A({ 1'h0, _08032_, _14716_, _05924_ }), .Y(_08146_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31309_ ( .A({ _08157_, _08154_, _08152_, _08147_ }), .Y(_14749_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31310_ ( .A({ _08151_, _08150_, _08149_, _08148_ }), .Y(_08147_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31311_ ( .A({ _15165_, _08059_, _13755_, _14813_ }), .Y(_08148_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31312_ ( .A({ _14973_, _08077_, _15133_, _08052_ }), .Y(_08149_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31313_ ( .A({ _15197_, _08064_, _14717_, _05924_ }), .Y(_08150_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31314_ ( .A({ _15229_, _05929_, _08032_, 1'h1 }), .Y(_08151_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31315_ ( .A({ _08153_, _08070_, _14877_ }), .Y(_08152_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31316_ ( .A({ _14941_, _08068_, _15101_, _08086_ }), .Y(_08153_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31317_ ( .A({ _08156_, _08037_, _08155_ }), .Y(_08154_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31318_ ( .A({ _14909_, _08069_, _08071_, _14845_ }), .Y(_08155_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31319_ ( .A({ _15261_, _08058_, _08055_, _14781_ }), .Y(_08156_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31320_ ( .A({ _08158_, _08065_, _15005_ }), .Y(_08157_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31321_ ( .A({ _15037_, _08062_, _15069_, _08063_ }), .Y(_08158_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31322_ ( .A({ _08170_, _08169_, _08164_, _08159_ }), .Y(_14750_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31323_ ( .A({ _08163_, _08162_, _08161_, _08160_ }), .Y(_08159_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31324_ ( .A({ _14942_, _08068_ }), .Y(_08160_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31325_ ( .A({ _14974_, _08077_, _15038_, _08062_ }), .Y(_08161_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31326_ ( .A({ _14782_, _08055_, _14718_, _05924_ }), .Y(_08162_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31327_ ( .A({ 1'h0, _08032_, _15134_, _08052_ }), .Y(_08163_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31328_ ( .A({ _08168_, _08167_, _08165_ }), .Y(_08164_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31329_ ( .A({ _08166_, _08063_, _15070_ }), .Y(_08165_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31330_ ( .A({ _15006_, _08065_, _15198_, _08064_ }), .Y(_08166_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31331_ ( .A({ _15166_, _08059_, _15230_, _05929_ }), .Y(_08167_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31332_ ( .A({ _14814_, _13755_, _15262_, _08058_ }), .Y(_08168_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31333_ ( .A({ _14910_, _08069_, _08071_, _14846_ }), .Y(_08169_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31334_ ( .A({ _14878_, _08070_, _15102_, _08086_ }), .Y(_08170_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31335_ ( .A({ _08182_, _08181_, _08176_, _08171_ }), .Y(_14751_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31336_ ( .A({ _08175_, _08173_, _08172_ }), .Y(_08171_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31337_ ( .A({ _14975_, _08077_, _15071_, _08063_ }), .Y(_08172_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31338_ ( .A({ _08174_, _08068_, _14943_ }), .Y(_08173_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31339_ ( .A({ _14815_, _13755_, _15007_, _08065_ }), .Y(_08174_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31340_ ( .A({ _14783_, _08055_, _14719_, _05924_ }), .Y(_08175_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31341_ ( .A({ _08180_, _08179_, _08177_, _08178_ }), .Y(_08176_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31342_ ( .A({ _15167_, _08059_, _08032_, 1'h0 }), .Y(_08177_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31343_ ( .A({ _15135_, _08052_ }), .Y(_08178_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31344_ ( .A({ _15231_, _05929_, _08064_, _15199_ }), .Y(_08179_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31345_ ( .A({ _15263_, _08058_, _08062_, _15039_ }), .Y(_08180_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31346_ ( .A({ _14911_, _08069_, _15103_, _08086_ }), .Y(_08181_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31347_ ( .A({ _14879_, _08070_, _08071_, _14847_ }), .Y(_08182_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31348_ ( .A({ _08194_, _08193_, _08188_, _08183_ }), .Y(_14752_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31349_ ( .A({ _08187_, _08186_, _08185_, _08184_ }), .Y(_08183_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31350_ ( .A({ _14944_, _08068_ }), .Y(_08184_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31351_ ( .A({ _14976_, _08077_, _15040_, _08062_ }), .Y(_08185_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31352_ ( .A({ _14784_, _08055_, _14720_, _05924_ }), .Y(_08186_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31353_ ( .A({ 1'h0, _08032_, _15136_, _08052_ }), .Y(_08187_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31354_ ( .A({ _08192_, _08191_, _08189_ }), .Y(_08188_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31355_ ( .A({ _08190_, _08063_, _15072_ }), .Y(_08189_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31356_ ( .A({ _15008_, _08065_, _15200_, _08064_ }), .Y(_08190_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31357_ ( .A({ _15168_, _08059_, _15232_, _05929_ }), .Y(_08191_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31358_ ( .A({ _14816_, _13755_, _15264_, _08058_ }), .Y(_08192_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31359_ ( .A({ _14912_, _08069_, _08071_, _14848_ }), .Y(_08193_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31360_ ( .A({ _14880_, _08070_, _15104_, _08086_ }), .Y(_08194_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31361_ ( .A({ _08206_, _08205_, _08200_, _08195_ }), .Y(_14753_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31362_ ( .A({ _08199_, _08197_, _08196_ }), .Y(_08195_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31363_ ( .A({ _15169_, _08059_, _08065_, _15009_ }), .Y(_08196_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31364_ ( .A({ _08198_, _08069_, _14913_ }), .Y(_08197_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31365_ ( .A({ _15233_, _05929_, _08032_, 1'h0 }), .Y(_08198_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31366_ ( .A({ _15265_, _08058_, _14721_, _05924_ }), .Y(_08199_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31367_ ( .A({ _08204_, _08203_, _08201_ }), .Y(_08200_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31368_ ( .A({ _08202_, _08077_, _14977_ }), .Y(_08201_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31369_ ( .A({ _15137_, _08052_, _08063_, _15073_ }), .Y(_08202_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31370_ ( .A({ _14785_, _08055_, _15201_, _08064_ }), .Y(_08203_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31371_ ( .A({ _14817_, _13755_, _15041_, _08062_ }), .Y(_08204_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31372_ ( .A({ _14849_, _08071_, _15105_, _08086_ }), .Y(_08205_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31373_ ( .A({ _14881_, _08070_, _14945_, _08068_ }), .Y(_08206_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31374_ ( .A({ _08218_, _08217_, _08212_, _08207_ }), .Y(_14723_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31375_ ( .A({ _08211_, _08210_, _08209_, _08208_ }), .Y(_08207_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31376_ ( .A({ _14915_, _08068_ }), .Y(_08208_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31377_ ( .A({ _14947_, _08077_, _15011_, _08062_ }), .Y(_08209_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31378_ ( .A({ _14755_, _08055_, _14691_, _05924_ }), .Y(_08210_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31379_ ( .A({ 1'h0, _08032_, _15107_, _08052_ }), .Y(_08211_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31380_ ( .A({ _08216_, _08215_, _08213_ }), .Y(_08212_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31381_ ( .A({ _08214_, _08063_, _15043_ }), .Y(_08213_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31382_ ( .A({ _14979_, _08065_, _15171_, _08064_ }), .Y(_08214_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31383_ ( .A({ _15139_, _08059_, _15203_, _05929_ }), .Y(_08215_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31384_ ( .A({ _14787_, _13755_, _15235_, _08058_ }), .Y(_08216_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31385_ ( .A({ _14883_, _08069_, _08071_, _14819_ }), .Y(_08217_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31386_ ( .A({ _14851_, _08070_, _15075_, _08086_ }), .Y(_08218_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31387_ ( .A({ _08230_, _08229_, _08224_, _08219_ }), .Y(_14724_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31388_ ( .A({ _08223_, _08222_, _08220_ }), .Y(_08219_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31389_ ( .A({ _08221_, _08071_, _14820_ }), .Y(_08220_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31390_ ( .A({ _15236_, _08058_, _08065_, _14980_ }), .Y(_08221_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31391_ ( .A({ _14788_, _13755_, _15204_, _05929_ }), .Y(_08222_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31392_ ( .A({ _14756_, _08055_, _14692_, _05924_ }), .Y(_08223_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31393_ ( .A({ _08228_, _08225_, _08226_, _08227_ }), .Y(_08224_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31394_ ( .A({ _14948_, _08077_, _15012_, _08062_ }), .Y(_08225_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31395_ ( .A({ _15140_, _08059_, _08032_, 1'h0 }), .Y(_08226_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31396_ ( .A({ _15108_, _08052_ }), .Y(_08227_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31397_ ( .A({ _15172_, _08064_, _08063_, _15044_ }), .Y(_08228_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31398_ ( .A({ _14884_, _08069_, _08070_, _14852_ }), .Y(_08229_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31399_ ( .A({ _14916_, _08068_, _15076_, _08086_ }), .Y(_08230_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31400_ ( .A({ _08242_, _08241_, _08236_, _08231_ }), .Y(_14725_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31401_ ( .A({ _08235_, _08234_, _08232_ }), .Y(_08231_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31402_ ( .A({ _08233_, _08069_, _14885_ }), .Y(_08232_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31403_ ( .A({ _14789_, _13755_, _14981_, _08065_ }), .Y(_08233_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31404_ ( .A({ _15013_, _08062_, _14693_, _05924_ }), .Y(_08234_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31405_ ( .A({ _15237_, _08058_, _08064_, _15173_ }), .Y(_08235_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31406_ ( .A({ _08240_, _08237_, _08238_, _08239_ }), .Y(_08236_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31407_ ( .A({ _15141_, _08059_, _08032_, 1'h0 }), .Y(_08237_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31408_ ( .A({ _14949_, _08077_, _15045_, _08063_ }), .Y(_08238_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31409_ ( .A({ _15109_, _08052_ }), .Y(_08239_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31410_ ( .A({ _15205_, _05929_, _08055_, _14757_ }), .Y(_08240_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31411_ ( .A({ _14853_, _08070_, _08071_, _14821_ }), .Y(_08241_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31412_ ( .A({ _14917_, _08068_, _15077_, _08086_ }), .Y(_08242_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31413_ ( .A({ _08254_, _08253_, _08248_, _08243_ }), .Y(_14726_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31414_ ( .A({ _08247_, _08246_, _08245_, _08244_ }), .Y(_08243_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31415_ ( .A({ _15078_, _08086_ }), .Y(_08244_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31416_ ( .A({ _14950_, _08077_, _15046_, _08063_ }), .Y(_08245_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31417_ ( .A({ _15238_, _08058_, _08065_, _14982_ }), .Y(_08246_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31418_ ( .A({ _14758_, _08055_, _15174_, _08064_ }), .Y(_08247_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31419_ ( .A({ _08252_, _08251_, _08249_, _08250_ }), .Y(_08248_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31420_ ( .A({ _15142_, _08059_, _15206_, _05929_ }), .Y(_08249_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31421_ ( .A({ _14790_, _13755_ }), .Y(_08250_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31422_ ( .A({ _15014_, _08062_, _14694_, _05924_ }), .Y(_08251_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31423_ ( .A({ 1'h0, _08032_, _15110_, _08052_ }), .Y(_08252_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31424_ ( .A({ _14822_, _08071_, _14918_, _08068_ }), .Y(_08253_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31425_ ( .A({ _14886_, _08069_, _08070_, _14854_ }), .Y(_08254_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31426_ ( .A({ _08266_, _08265_, _08260_, _08255_ }), .Y(_14727_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31427_ ( .A({ _08259_, _08257_, _08256_ }), .Y(_08255_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31428_ ( .A({ _15143_, _08059_, _08065_, _14983_ }), .Y(_08256_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31429_ ( .A({ _08258_, _08069_, _14887_ }), .Y(_08257_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31430_ ( .A({ _15207_, _05929_, _08032_, 1'h0 }), .Y(_08258_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31431_ ( .A({ _15175_, _08064_, _14695_, _05924_ }), .Y(_08259_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31432_ ( .A({ _08264_, _08263_, _08261_ }), .Y(_08260_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31433_ ( .A({ _08262_, _08077_, _14951_ }), .Y(_08261_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31434_ ( .A({ _15111_, _08052_, _08063_, _15047_ }), .Y(_08262_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31435_ ( .A({ _15239_, _08058_, _08055_, _14759_ }), .Y(_08263_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31436_ ( .A({ _14791_, _13755_, _15015_, _08062_ }), .Y(_08264_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31437_ ( .A({ _14823_, _08071_, _15079_, _08086_ }), .Y(_08265_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31438_ ( .A({ _14855_, _08070_, _14919_, _08068_ }), .Y(_08266_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31439_ ( .A({ _08278_, _08277_, _08272_, _08267_ }), .Y(_14728_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31440_ ( .A({ _08271_, _08270_, _08269_, _08268_ }), .Y(_08267_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31441_ ( .A({ _15080_, _08086_ }), .Y(_08268_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31442_ ( .A({ _14952_, _08077_, _15048_, _08063_ }), .Y(_08269_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31443_ ( .A({ _14984_, _08065_, _15176_, _08064_ }), .Y(_08270_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31444_ ( .A({ _15240_, _08058_, _08055_, _14760_ }), .Y(_08271_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31445_ ( .A({ _08276_, _08275_, _08273_, _08274_ }), .Y(_08272_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31446_ ( .A({ _15144_, _08059_, _15208_, _05929_ }), .Y(_08273_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31447_ ( .A({ _14792_, _13755_ }), .Y(_08274_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31448_ ( .A({ _15016_, _08062_, _14696_, _05924_ }), .Y(_08275_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31449_ ( .A({ 1'h0, _08032_, _15112_, _08052_ }), .Y(_08276_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31450_ ( .A({ _14824_, _08071_, _14920_, _08068_ }), .Y(_08277_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31451_ ( .A({ _14888_, _08069_, _08070_, _14856_ }), .Y(_08278_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31452_ ( .A({ _08290_, _08289_, _08284_, _08279_ }), .Y(_14729_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31453_ ( .A({ _08283_, _08282_, _08281_, _08280_ }), .Y(_08279_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31454_ ( .A({ _14921_, _08068_ }), .Y(_08280_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31455_ ( .A({ _14953_, _08077_, _15017_, _08062_ }), .Y(_08281_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31456_ ( .A({ _14761_, _08055_, _14697_, _05924_ }), .Y(_08282_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31457_ ( .A({ 1'h0, _08032_, _15113_, _08052_ }), .Y(_08283_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31458_ ( .A({ _08288_, _08287_, _08285_ }), .Y(_08284_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31459_ ( .A({ _08286_, _08063_, _15049_ }), .Y(_08285_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31460_ ( .A({ _15241_, _08058_, _08065_, _14985_ }), .Y(_08286_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31461_ ( .A({ _15145_, _08059_, _15209_, _05929_ }), .Y(_08287_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31462_ ( .A({ _14793_, _13755_, _15177_, _08064_ }), .Y(_08288_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31463_ ( .A({ _14889_, _08069_, _08071_, _14825_ }), .Y(_08289_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31464_ ( .A({ _14857_, _08070_, _15081_, _08086_ }), .Y(_08290_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31465_ ( .A({ _08302_, _08301_, _08296_, _08291_ }), .Y(_14730_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31466_ ( .A({ _08295_, _08293_, _08292_ }), .Y(_08291_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31467_ ( .A({ _15146_, _08059_, _08065_, _14986_ }), .Y(_08292_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31468_ ( .A({ _08294_, _08069_, _14890_ }), .Y(_08293_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31469_ ( .A({ _15210_, _05929_, _08032_, 1'h0 }), .Y(_08294_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31470_ ( .A({ _15242_, _08058_, _14698_, _05924_ }), .Y(_08295_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31471_ ( .A({ _08300_, _08299_, _08297_ }), .Y(_08296_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31472_ ( .A({ _08298_, _08077_, _14954_ }), .Y(_08297_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31473_ ( .A({ _15114_, _08052_, _08063_, _15050_ }), .Y(_08298_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31474_ ( .A({ _14762_, _08055_, _15178_, _08064_ }), .Y(_08299_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31475_ ( .A({ _14794_, _13755_, _15018_, _08062_ }), .Y(_08300_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31476_ ( .A({ _14826_, _08071_, _15082_, _08086_ }), .Y(_08301_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31477_ ( .A({ _14858_, _08070_, _14922_, _08068_ }), .Y(_08302_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31478_ ( .A({ _08314_, _08313_, _08308_, _08303_ }), .Y(_14731_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31479_ ( .A({ _08307_, _08306_, _08304_ }), .Y(_08303_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31480_ ( .A({ _08305_, _08069_, _14891_ }), .Y(_08304_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31481_ ( .A({ _14795_, _13755_, _14987_, _08065_ }), .Y(_08305_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31482_ ( .A({ _15019_, _08062_, _14699_, _05924_ }), .Y(_08306_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31483_ ( .A({ _15243_, _08058_, _08064_, _15179_ }), .Y(_08307_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31484_ ( .A({ _08312_, _08309_, _08310_, _08311_ }), .Y(_08308_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31485_ ( .A({ _15147_, _08059_, _08032_, 1'h0 }), .Y(_08309_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31486_ ( .A({ _14955_, _08077_, _15051_, _08063_ }), .Y(_08310_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31487_ ( .A({ _15115_, _08052_ }), .Y(_08311_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31488_ ( .A({ _15211_, _05929_, _08055_, _14763_ }), .Y(_08312_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31489_ ( .A({ _14859_, _08070_, _08071_, _14827_ }), .Y(_08313_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31490_ ( .A({ _14923_, _08068_, _15083_, _08086_ }), .Y(_08314_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31491_ ( .A({ _08326_, _08325_, _08320_, _08315_ }), .Y(_14732_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31492_ ( .A({ _08319_, _08318_, _08316_ }), .Y(_08315_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31493_ ( .A({ _08317_, _08086_, _15084_ }), .Y(_08316_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31494_ ( .A({ _15244_, _08058_, _08062_, _15020_ }), .Y(_08317_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31495_ ( .A({ _14796_, _13755_, _15212_, _05929_ }), .Y(_08318_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31496_ ( .A({ 1'h0, _08032_, _15116_, _08052_ }), .Y(_08319_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31497_ ( .A({ _08324_, _08321_, _08322_, _08323_ }), .Y(_08320_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31498_ ( .A({ _14956_, _08077_, _14700_, _05924_ }), .Y(_08321_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31499_ ( .A({ _15148_, _08059_, _15180_, _08064_ }), .Y(_08322_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31500_ ( .A({ _14764_, _08055_ }), .Y(_08323_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31501_ ( .A({ _14988_, _08065_, _15052_, _08063_ }), .Y(_08324_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31502_ ( .A({ _14828_, _08071_, _14924_, _08068_ }), .Y(_08325_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31503_ ( .A({ _14892_, _08069_, _08070_, _14860_ }), .Y(_08326_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31504_ ( .A({ _08338_, _08337_, _08332_, _08327_ }), .Y(_14734_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31505_ ( .A({ _08331_, _08330_, _08329_, _08328_ }), .Y(_08327_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31506_ ( .A({ _15086_, _08086_ }), .Y(_08328_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31507_ ( .A({ _14958_, _08077_, _15054_, _08063_ }), .Y(_08329_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31508_ ( .A({ _14990_, _08065_, _15182_, _08064_ }), .Y(_08330_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31509_ ( .A({ _15246_, _08058_, _08055_, _14766_ }), .Y(_08331_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31510_ ( .A({ _08336_, _08335_, _08333_, _08334_ }), .Y(_08332_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31511_ ( .A({ _15150_, _08059_, _15214_, _05929_ }), .Y(_08333_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31512_ ( .A({ _14798_, _13755_ }), .Y(_08334_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31513_ ( .A({ _15022_, _08062_, _14702_, _05924_ }), .Y(_08335_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31514_ ( .A({ 1'h0, _08032_, _15118_, _08052_ }), .Y(_08336_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31515_ ( .A({ _14830_, _08071_, _14926_, _08068_ }), .Y(_08337_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31516_ ( .A({ _14894_, _08069_, _08070_, _14862_ }), .Y(_08338_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31517_ ( .A({ _08350_, _08349_, _08344_, _08339_ }), .Y(_14735_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31518_ ( .A({ _08343_, _08342_, _08341_, _08340_ }), .Y(_08339_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31519_ ( .A({ _14927_, _08068_ }), .Y(_08340_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31520_ ( .A({ _14959_, _08077_, _15023_, _08062_ }), .Y(_08341_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31521_ ( .A({ _14767_, _08055_, _14703_, _05924_ }), .Y(_08342_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31522_ ( .A({ 1'h0, _08032_, _15119_, _08052_ }), .Y(_08343_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31523_ ( .A({ _08348_, _08347_, _08345_ }), .Y(_08344_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31524_ ( .A({ _08346_, _08063_, _15055_ }), .Y(_08345_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31525_ ( .A({ _14991_, _08065_, _15183_, _08064_ }), .Y(_08346_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31526_ ( .A({ _15151_, _08059_, _15215_, _05929_ }), .Y(_08347_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31527_ ( .A({ _14799_, _13755_, _15247_, _08058_ }), .Y(_08348_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31528_ ( .A({ _14895_, _08069_, _08071_, _14831_ }), .Y(_08349_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31529_ ( .A({ _14863_, _08070_, _15087_, _08086_ }), .Y(_08350_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31530_ ( .A({ _08362_, _08361_, _08356_, _08351_ }), .Y(_14736_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31531_ ( .A({ _08355_, _08354_, _08353_, _08352_ }), .Y(_08351_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31532_ ( .A({ _14928_, _08068_ }), .Y(_08352_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31533_ ( .A({ _14960_, _08077_, _15024_, _08062_ }), .Y(_08353_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31534_ ( .A({ _14768_, _08055_, _14704_, _05924_ }), .Y(_08354_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31535_ ( .A({ 1'h0, _08032_, _15120_, _08052_ }), .Y(_08355_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31536_ ( .A({ _08360_, _08359_, _08357_ }), .Y(_08356_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31537_ ( .A({ _08358_, _08063_, _15056_ }), .Y(_08357_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31538_ ( .A({ _14992_, _08065_, _15184_, _08064_ }), .Y(_08358_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31539_ ( .A({ _15152_, _08059_, _15216_, _05929_ }), .Y(_08359_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31540_ ( .A({ _14800_, _13755_, _15248_, _08058_ }), .Y(_08360_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31541_ ( .A({ _14896_, _08069_, _08071_, _14832_ }), .Y(_08361_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31542_ ( .A({ _14864_, _08070_, _15088_, _08086_ }), .Y(_08362_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31543_ ( .A({ _08374_, _08373_, _08368_, _08363_ }), .Y(_14737_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31544_ ( .A({ _08367_, _08366_, _08364_ }), .Y(_08363_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31545_ ( .A({ _08365_, _08086_, _15089_ }), .Y(_08364_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31546_ ( .A({ _15185_, _08064_, _08062_, _15025_ }), .Y(_08365_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31547_ ( .A({ _14801_, _13755_, _15217_, _05929_ }), .Y(_08366_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31548_ ( .A({ 1'h0, _08032_, _15121_, _08052_ }), .Y(_08367_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31549_ ( .A({ _08372_, _08369_, _08370_, _08371_ }), .Y(_08368_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31550_ ( .A({ _14961_, _08077_, _14705_, _05924_ }), .Y(_08369_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31551_ ( .A({ _15153_, _08059_, _15249_, _08058_ }), .Y(_08370_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31552_ ( .A({ _14769_, _08055_ }), .Y(_08371_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31553_ ( .A({ _14993_, _08065_, _15057_, _08063_ }), .Y(_08372_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31554_ ( .A({ _14833_, _08071_, _14929_, _08068_ }), .Y(_08373_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31555_ ( .A({ _14897_, _08069_, _08070_, _14865_ }), .Y(_08374_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31556_ ( .A({ _08386_, _08385_, _08380_, _08375_ }), .Y(_14738_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31557_ ( .A({ _08379_, _08378_, _08377_, _08376_ }), .Y(_08375_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31558_ ( .A({ _15090_, _08086_ }), .Y(_08376_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31559_ ( .A({ _14962_, _08077_, _15058_, _08063_ }), .Y(_08377_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31560_ ( .A({ _15250_, _08058_, _08065_, _14994_ }), .Y(_08378_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31561_ ( .A({ _14770_, _08055_, _15186_, _08064_ }), .Y(_08379_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31562_ ( .A({ _08384_, _08383_, _08381_, _08382_ }), .Y(_08380_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31563_ ( .A({ _15154_, _08059_, _15218_, _05929_ }), .Y(_08381_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31564_ ( .A({ _14802_, _13755_ }), .Y(_08382_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31565_ ( .A({ _15026_, _08062_, _14706_, _05924_ }), .Y(_08383_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31566_ ( .A({ 1'h0, _08032_, _15122_, _08052_ }), .Y(_08384_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31567_ ( .A({ _14834_, _08071_, _14930_, _08068_ }), .Y(_08385_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31568_ ( .A({ _14898_, _08069_, _08070_, _14866_ }), .Y(_08386_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31569_ ( .A({ _08398_, _08397_, _08392_, _08387_ }), .Y(_14739_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31570_ ( .A({ _08391_, _08390_, _08388_ }), .Y(_08387_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31571_ ( .A({ _08389_, _08086_, _15091_ }), .Y(_08388_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31572_ ( .A({ _15187_, _08064_, _08062_, _15027_ }), .Y(_08389_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31573_ ( .A({ _14803_, _13755_, _15219_, _05929_ }), .Y(_08390_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31574_ ( .A({ 1'h0, _08032_, _15123_, _08052_ }), .Y(_08391_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31575_ ( .A({ _08396_, _08393_, _08394_, _08395_ }), .Y(_08392_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31576_ ( .A({ _14963_, _08077_, _14707_, _05924_ }), .Y(_08393_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31577_ ( .A({ _15155_, _08059_, _15251_, _08058_ }), .Y(_08394_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31578_ ( .A({ _14771_, _08055_ }), .Y(_08395_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31579_ ( .A({ _14995_, _08065_, _15059_, _08063_ }), .Y(_08396_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31580_ ( .A({ _14835_, _08071_, _14931_, _08068_ }), .Y(_08397_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31581_ ( .A({ _14899_, _08069_, _08070_, _14867_ }), .Y(_08398_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31582_ ( .A({ _08410_, _08409_, _08404_, _08399_ }), .Y(_14740_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31583_ ( .A({ _08403_, _08402_, _08401_, _08400_ }), .Y(_08399_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31584_ ( .A({ _14932_, _08068_ }), .Y(_08400_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31585_ ( .A({ _14964_, _08077_, _15028_, _08062_ }), .Y(_08401_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31586_ ( .A({ _14772_, _08055_, _14708_, _05924_ }), .Y(_08402_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31587_ ( .A({ 1'h0, _08032_, _15124_, _08052_ }), .Y(_08403_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31588_ ( .A({ _08408_, _08407_, _08405_ }), .Y(_08404_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31589_ ( .A({ _08406_, _08063_, _15060_ }), .Y(_08405_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31590_ ( .A({ _15252_, _08058_, _08065_, _14996_ }), .Y(_08406_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31591_ ( .A({ _15156_, _08059_, _15220_, _05929_ }), .Y(_08407_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31592_ ( .A({ _14804_, _13755_, _15188_, _08064_ }), .Y(_08408_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31593_ ( .A({ _14900_, _08069_, _08071_, _14836_ }), .Y(_08409_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31594_ ( .A({ _14868_, _08070_, _15092_, _08086_ }), .Y(_08410_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31595_ ( .A({ _08422_, _08421_, _08416_, _08411_ }), .Y(_14741_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31596_ ( .A({ _08415_, _08414_, _08413_, _08412_ }), .Y(_08411_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31597_ ( .A({ _15093_, _08086_ }), .Y(_08412_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31598_ ( .A({ _14965_, _08077_, _15061_, _08063_ }), .Y(_08413_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31599_ ( .A({ _14997_, _08065_, _15189_, _08064_ }), .Y(_08414_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31600_ ( .A({ _15253_, _08058_, _08055_, _14773_ }), .Y(_08415_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31601_ ( .A({ _08420_, _08419_, _08417_, _08418_ }), .Y(_08416_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31602_ ( .A({ _15157_, _08059_, _15221_, _05929_ }), .Y(_08417_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31603_ ( .A({ _14805_, _13755_ }), .Y(_08418_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31604_ ( .A({ _15029_, _08062_, _14709_, _05924_ }), .Y(_08419_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31605_ ( .A({ 1'h0, _08032_, _15125_, _08052_ }), .Y(_08420_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31606_ ( .A({ _14837_, _08071_, _14933_, _08068_ }), .Y(_08421_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31607_ ( .A({ _14901_, _08069_, _08070_, _14869_ }), .Y(_08422_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31608_ ( .A({ _08434_, _08433_, _08428_, _08423_ }), .Y(_14742_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31609_ ( .A({ _08427_, _08425_, _08424_ }), .Y(_08423_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31610_ ( .A({ _14966_, _08077_, _15062_, _08063_ }), .Y(_08424_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31611_ ( .A({ _08426_, _08068_, _14934_ }), .Y(_08425_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31612_ ( .A({ _14806_, _13755_, _14998_, _08065_ }), .Y(_08426_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31613_ ( .A({ _14774_, _08055_, _14710_, _05924_ }), .Y(_08427_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31614_ ( .A({ _08432_, _08431_, _08429_, _08430_ }), .Y(_08428_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31615_ ( .A({ _15158_, _08059_, _08032_, 1'h0 }), .Y(_08429_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31616_ ( .A({ _15126_, _08052_ }), .Y(_08430_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _31617_ ( .A({ _15222_, _05929_, _15254_, _08058_ }), .Y(_08431_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31618_ ( .A({ _15190_, _08064_, _08062_, _15030_ }), .Y(_08432_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31619_ ( .A({ _14902_, _08069_, _15094_, _08086_ }), .Y(_08433_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31620_ ( .A({ _14870_, _08070_, _08071_, _14838_ }), .Y(_08434_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31621_ ( .A({ _08446_, _08445_, _08440_, _08435_ }), .Y(_14743_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31622_ ( .A({ _08439_, _08438_, _08436_ }), .Y(_08435_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31623_ ( .A({ _08437_, _08071_, _14839_ }), .Y(_08436_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31624_ ( .A({ _15255_, _08058_, _08065_, _14999_ }), .Y(_08437_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31625_ ( .A({ _14807_, _13755_, _15223_, _05929_ }), .Y(_08438_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31626_ ( .A({ _14775_, _08055_, _14711_, _05924_ }), .Y(_08439_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31627_ ( .A({ _08444_, _08441_, _08442_, _08443_ }), .Y(_08440_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31628_ ( .A({ _14967_, _08077_, _15031_, _08062_ }), .Y(_08441_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31629_ ( .A({ _15159_, _08059_, _08032_, 1'h0 }), .Y(_08442_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31630_ ( .A({ _15127_, _08052_ }), .Y(_08443_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31631_ ( .A({ _15191_, _08064_, _08063_, _15063_ }), .Y(_08444_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31632_ ( .A({ _14903_, _08069_, _08070_, _14871_ }), .Y(_08445_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31633_ ( .A({ _14935_, _08068_, _15095_, _08086_ }), .Y(_08446_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31634_ ( .A({ _08458_, _08457_, _08452_, _08447_ }), .Y(_14745_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31635_ ( .A({ _08451_, _08450_, _08449_, _08448_ }), .Y(_08447_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31636_ ( .A({ _14937_, _08068_ }), .Y(_08448_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31637_ ( .A({ _14969_, _08077_, _15033_, _08062_ }), .Y(_08449_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31638_ ( .A({ _14777_, _08055_, _14713_, _05924_ }), .Y(_08450_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31639_ ( .A({ 1'h0, _08032_, _15129_, _08052_ }), .Y(_08451_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _31640_ ( .A({ _08456_, _08455_, _08453_ }), .Y(_08452_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _31641_ ( .A({ _08454_, _08063_, _15065_ }), .Y(_08453_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31642_ ( .A({ _15001_, _08065_, _15193_, _08064_ }), .Y(_08454_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31643_ ( .A({ _15161_, _08059_, _15225_, _05929_ }), .Y(_08455_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31644_ ( .A({ _14809_, _13755_, _15257_, _08058_ }), .Y(_08456_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31645_ ( .A({ _14905_, _08069_, _08071_, _14841_ }), .Y(_08457_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31646_ ( .A({ _14873_, _08070_, _15097_, _08086_ }), .Y(_08458_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _31647_ ( .A({ _08470_, _08469_, _08464_, _08459_ }), .Y(_14746_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31648_ ( .A({ _08463_, _08462_, _08461_, _08460_ }), .Y(_08459_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31649_ ( .A({ _15098_, _08086_ }), .Y(_08460_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31650_ ( .A({ _14970_, _08077_, _15066_, _08063_ }), .Y(_08461_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31651_ ( .A({ _15258_, _08058_, _08065_, _15002_ }), .Y(_08462_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31652_ ( .A({ _14778_, _08055_, _15194_, _08064_ }), .Y(_08463_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31653_ ( .A({ _08468_, _08467_, _08465_, _08466_ }), .Y(_08464_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31654_ ( .A({ _15162_, _08059_, _15226_, _05929_ }), .Y(_08465_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31655_ ( .A({ _14810_, _13755_ }), .Y(_08466_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _31656_ ( .A({ _15034_, _08062_, _14714_, _05924_ }), .Y(_08467_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31657_ ( .A({ 1'h0, _08032_, _15130_, _08052_ }), .Y(_08468_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31658_ ( .A({ _14842_, _08071_, _14938_, _08068_ }), .Y(_08469_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31659_ ( .A({ _14906_, _08069_, _08070_, _14874_ }), .Y(_08470_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31660_ ( .A({ _14594_, _13755_, _14626_, _08032_ }), .Y(_05549_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31661_ ( .A({ _14605_, _13755_, _14637_, _08032_ }), .Y(_05550_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31662_ ( .A({ _14616_, _13755_, _14648_, _08032_ }), .Y(_05551_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31663_ ( .A({ _14619_, _13755_, _14651_, _08032_ }), .Y(_05552_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31664_ ( .A({ _14620_, _13755_, _14652_, _08032_ }), .Y(_05553_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31665_ ( .A({ _14621_, _13755_, _14653_, _08032_ }), .Y(_05554_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31666_ ( .A({ _14622_, _13755_, _14654_, _08032_ }), .Y(_05555_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31667_ ( .A({ _14623_, _13755_, _14655_, _08032_ }), .Y(_05556_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31668_ ( .A({ _14624_, _13755_, _14656_, _08032_ }), .Y(_05557_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31669_ ( .A({ _14625_, _13755_, _14657_, _08032_ }), .Y(_05558_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31670_ ( .A({ _14595_, _13755_, _14627_, _08032_ }), .Y(_05559_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31671_ ( .A({ _14596_, _13755_, _14628_, _08032_ }), .Y(_05560_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31672_ ( .A({ _14597_, _13755_, _14629_, _08032_ }), .Y(_05561_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31673_ ( .A({ _14598_, _13755_, _14630_, _08032_ }), .Y(_05562_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31674_ ( .A({ _14599_, _13755_, _14631_, _08032_ }), .Y(_05563_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31675_ ( .A({ _14600_, _13755_, _14632_, _08032_ }), .Y(_05564_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31676_ ( .A({ _14601_, _13755_, _14633_, _08032_ }), .Y(_05565_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31677_ ( .A({ _14602_, _13755_, _14634_, _08032_ }), .Y(_05566_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31678_ ( .A({ _14603_, _13755_, _14635_, _08032_ }), .Y(_05567_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31679_ ( .A({ _14604_, _13755_, _14636_, _08032_ }), .Y(_05568_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31680_ ( .A({ _14606_, _13755_, _14638_, _08032_ }), .Y(_05569_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31681_ ( .A({ _14607_, _13755_, _14639_, _08032_ }), .Y(_05570_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31682_ ( .A({ _14608_, _13755_, _14640_, _08032_ }), .Y(_05571_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31683_ ( .A({ _14609_, _13755_, _14641_, _08032_ }), .Y(_05572_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31684_ ( .A({ _14610_, _13755_, _14642_, _08032_ }), .Y(_05573_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31685_ ( .A({ _14611_, _13755_, _14643_, _08032_ }), .Y(_05574_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31686_ ( .A({ _14612_, _13755_, _14644_, _08032_ }), .Y(_05575_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31687_ ( .A({ _14613_, _13755_, _14645_, _08032_ }), .Y(_05576_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31688_ ( .A({ _14614_, _13755_, _14646_, _08032_ }), .Y(_05577_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31689_ ( .A({ _14615_, _13755_, _14647_, _08032_ }), .Y(_05578_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31690_ ( .A({ _14617_, _13755_, _14649_, _08032_ }), .Y(_05579_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _31691_ ( .A({ _14618_, _13755_, _14650_, _08032_ }), .Y(_05580_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31692_ ( .A({ _08471_, _04701_, _08474_ }), .Y(_22850_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31693_ ( .A({ _04605_, _08472_, _08473_, _04477_ }), .Y(_08471_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31694_ ( .A({ _06887_, _06900_, _06891_, main_fsm[4] }), .Y(_08472_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31695_ ( .A({ main_fsm[4], _06904_, _06898_, _06891_ }), .Y(_08473_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31696_ ( .A({ main_fsm[4], _06917_, _06891_, _06887_ }), .Y(_08474_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31697_ ( .A({ _08475_, _04700_, _08474_ }), .Y(_22849_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31698_ ( .A({ _04604_, _08472_, _08473_, _04476_ }), .Y(_08475_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31699_ ( .A({ _08476_, _04475_, _08473_ }), .Y(_22848_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31700_ ( .A({ _04699_, _08474_, _08472_, _04603_ }), .Y(_08476_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31701_ ( .A({ _08477_, _04474_, _08473_ }), .Y(_22847_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31702_ ( .A({ _04698_, _08474_, _08472_, _04602_ }), .Y(_08477_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31703_ ( .A({ _08478_, _04473_, _08473_ }), .Y(_22846_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31704_ ( .A({ _04697_, _08474_, _08472_, _04601_ }), .Y(_08478_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31705_ ( .A({ _08479_, _04472_, _08473_ }), .Y(_22845_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31706_ ( .A({ _04696_, _08474_, _08472_, _04600_ }), .Y(_08479_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31707_ ( .A({ _08480_, _04695_, _08474_ }), .Y(_22844_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31708_ ( .A({ _04599_, _08472_, _08473_, _04471_ }), .Y(_08480_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31709_ ( .A({ _08481_, _04694_, _08474_ }), .Y(_22843_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31710_ ( .A({ _04598_, _08472_, _08473_, _04470_ }), .Y(_08481_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31711_ ( .A({ _08482_, _04693_, _08474_ }), .Y(_22842_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31712_ ( .A({ _04597_, _08472_, _08473_, _04469_ }), .Y(_08482_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31713_ ( .A({ _08483_, _04692_, _08474_ }), .Y(_22841_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31714_ ( .A({ _04596_, _08472_, _08473_, _04468_ }), .Y(_08483_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31715_ ( .A({ _08484_, _04690_, _08474_ }), .Y(_22839_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31716_ ( .A({ _04594_, _08472_, _08473_, _04466_ }), .Y(_08484_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31717_ ( .A({ _08485_, _04689_, _08474_ }), .Y(_22838_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31718_ ( .A({ _04593_, _08472_, _08473_, _04465_ }), .Y(_08485_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31719_ ( .A({ _08486_, _04464_, _08473_ }), .Y(_22837_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31720_ ( .A({ _04688_, _08474_, _08472_, _04592_ }), .Y(_08486_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31721_ ( .A({ _08487_, _04687_, _08474_ }), .Y(_22836_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31722_ ( .A({ _04591_, _08472_, _08473_, _04463_ }), .Y(_08487_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31723_ ( .A({ _08488_, _04686_, _08474_ }), .Y(_22835_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31724_ ( .A({ _04590_, _08472_, _08473_, _04462_ }), .Y(_08488_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31725_ ( .A({ _08489_, _04685_, _08474_ }), .Y(_22834_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31726_ ( .A({ _04589_, _08472_, _08473_, _04461_ }), .Y(_08489_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31727_ ( .A({ _08490_, _04684_, _08474_ }), .Y(_22833_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31728_ ( .A({ _04588_, _08472_, _08473_, _04460_ }), .Y(_08490_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31729_ ( .A({ _08491_, _04459_, _08473_ }), .Y(_22832_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31730_ ( .A({ _04683_, _08474_, _08472_, _04587_ }), .Y(_08491_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31731_ ( .A({ _08492_, _04458_, _08473_ }), .Y(_22831_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31732_ ( .A({ _04682_, _08474_, _08472_, _04586_ }), .Y(_08492_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31733_ ( .A({ _08493_, _04457_, _08473_ }), .Y(_22830_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31734_ ( .A({ _04681_, _08474_, _08472_, _04585_ }), .Y(_08493_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31735_ ( .A({ _08494_, _04711_, _08474_ }), .Y(_22860_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31736_ ( .A({ _04615_, _08472_, _08473_, _04487_ }), .Y(_08494_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31737_ ( .A({ _08495_, _04710_, _08474_ }), .Y(_22859_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31738_ ( .A({ _04614_, _08472_, _08473_, _04486_ }), .Y(_08495_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31739_ ( .A({ _08496_, _04485_, _08473_ }), .Y(_22858_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31740_ ( .A({ _04709_, _08474_, _08472_, _04613_ }), .Y(_08496_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31741_ ( .A({ _08497_, _04484_, _08473_ }), .Y(_22857_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31742_ ( .A({ _04708_, _08474_, _08472_, _04612_ }), .Y(_08497_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31743_ ( .A({ _08498_, _04707_, _08474_ }), .Y(_22856_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31744_ ( .A({ _04611_, _08472_, _08473_, _04483_ }), .Y(_08498_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31745_ ( .A({ _08499_, _04482_, _08473_ }), .Y(_22855_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31746_ ( .A({ _04706_, _08474_, _08472_, _04610_ }), .Y(_08499_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31747_ ( .A({ _08500_, _04705_, _08474_ }), .Y(_22854_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31748_ ( .A({ _04609_, _08472_, _08473_, _04481_ }), .Y(_08500_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31749_ ( .A({ _08501_, _04702_, _08474_ }), .Y(_22851_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31750_ ( .A({ _04606_, _08472_, _08473_, _04478_ }), .Y(_08501_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31751_ ( .A({ _08502_, _04467_, _08473_ }), .Y(_22840_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31752_ ( .A({ _04691_, _08474_, _08472_, _04595_ }), .Y(_08502_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31753_ ( .A({ _08503_, _04680_, _08474_ }), .Y(_22829_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31754_ ( .A({ _04584_, _08472_, _08473_, _04456_ }), .Y(_08503_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _31755_ ( .A({ _08473_, _08472_, _08474_ }), .Y(_24078_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _31756_ ( .A({ _08505_, _07463_, _06930_ }), .Y(_08504_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _31757_ ( .A({ _06008_, _07472_, _07470_, _07066_ }), .Y(_08505_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31758_ ( .A({ _08506_, _04448_, _08509_ }), .Y(_22885_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31759_ ( .A({ _04576_, _08507_, _04672_, _08508_ }), .Y(_08506_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31760_ ( .A({ _06905_, _06886_ }), .Y(_08507_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31761_ ( .A({ main_fsm[4], _06897_, _06891_, _06887_ }), .Y(_08508_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31762_ ( .A({ main_fsm[4], _06909_, _06898_, _06891_ }), .Y(_08509_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31763_ ( .A({ _08510_, _04447_, _08509_ }), .Y(_22884_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31764_ ( .A({ _04575_, _08507_, _04671_, _08508_ }), .Y(_08510_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31765_ ( .A({ _08511_, _04669_, _08508_ }), .Y(_22882_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31766_ ( .A({ _04573_, _08507_, _08509_, _04445_ }), .Y(_08511_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31767_ ( .A({ _08512_, _04668_, _08508_ }), .Y(_22881_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31768_ ( .A({ _04572_, _08507_, _08509_, _04444_ }), .Y(_08512_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31769_ ( .A({ _08513_, _04665_, _08508_ }), .Y(_22878_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31770_ ( .A({ _04569_, _08507_, _08509_, _04441_ }), .Y(_08513_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31771_ ( .A({ _08514_, _04664_, _08508_ }), .Y(_22877_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31772_ ( .A({ _04568_, _08507_, _08509_, _04440_ }), .Y(_08514_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31773_ ( .A({ _08515_, _04663_, _08508_ }), .Y(_22876_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31774_ ( .A({ _04567_, _08507_, _08509_, _04439_ }), .Y(_08515_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31775_ ( .A({ _08516_, _04438_, _08509_ }), .Y(_22875_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31776_ ( .A({ _04566_, _08507_, _04662_, _08508_ }), .Y(_08516_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31777_ ( .A({ _08517_, _04661_, _08508_ }), .Y(_22874_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31778_ ( .A({ _04565_, _08507_, _08509_, _04437_ }), .Y(_08517_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31779_ ( .A({ _08518_, _04660_, _08508_ }), .Y(_22873_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31780_ ( .A({ _04564_, _08507_, _08509_, _04436_ }), .Y(_08518_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31781_ ( .A({ _08519_, _04658_, _08508_ }), .Y(_22871_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31782_ ( .A({ _04562_, _08507_, _08509_, _04434_ }), .Y(_08519_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31783_ ( .A({ _08520_, _04433_, _08509_ }), .Y(_22870_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31784_ ( .A({ _04561_, _08507_, _04657_, _08508_ }), .Y(_08520_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31785_ ( .A({ _08521_, _04656_, _08508_ }), .Y(_22869_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31786_ ( .A({ _04560_, _08507_, _08509_, _04432_ }), .Y(_08521_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31787_ ( .A({ _08522_, _04655_, _08508_ }), .Y(_22868_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31788_ ( .A({ _04559_, _08507_, _08509_, _04431_ }), .Y(_08522_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31789_ ( .A({ _08523_, _04654_, _08508_ }), .Y(_22867_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31790_ ( .A({ _04558_, _08507_, _08509_, _04430_ }), .Y(_08523_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31791_ ( .A({ _08524_, _04429_, _08509_ }), .Y(_22866_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31792_ ( .A({ _04557_, _08507_, _04653_, _08508_ }), .Y(_08524_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31793_ ( .A({ _08525_, _04652_, _08508_ }), .Y(_22865_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31794_ ( .A({ _04556_, _08507_, _08509_, _04428_ }), .Y(_08525_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31795_ ( .A({ _08526_, _04427_, _08509_ }), .Y(_22864_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31796_ ( .A({ _04555_, _08507_, _04651_, _08508_ }), .Y(_08526_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31797_ ( .A({ _08527_, _04426_, _08509_ }), .Y(_22863_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31798_ ( .A({ _04554_, _08507_, _04650_, _08508_ }), .Y(_08527_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31799_ ( .A({ _08528_, _04425_, _08509_ }), .Y(_22862_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31800_ ( .A({ _04553_, _08507_, _04649_, _08508_ }), .Y(_08528_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31801_ ( .A({ _08529_, _04679_, _08508_ }), .Y(_22892_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31802_ ( .A({ _04583_, _08507_, _08509_, _04455_ }), .Y(_08529_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31803_ ( .A({ _08530_, _04678_, _08508_ }), .Y(_22891_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31804_ ( .A({ _04582_, _08507_, _08509_, _04454_ }), .Y(_08530_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31805_ ( .A({ _08531_, _04677_, _08508_ }), .Y(_22890_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31806_ ( .A({ _04581_, _08507_, _08509_, _04453_ }), .Y(_08531_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31807_ ( .A({ _08532_, _04676_, _08508_ }), .Y(_22889_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31808_ ( .A({ _04580_, _08507_, _08509_, _04452_ }), .Y(_08532_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31809_ ( .A({ _08533_, _04675_, _08508_ }), .Y(_22888_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31810_ ( .A({ _04579_, _08507_, _08509_, _04451_ }), .Y(_08533_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31811_ ( .A({ _08534_, _04674_, _08508_ }), .Y(_22887_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31812_ ( .A({ _04578_, _08507_, _08509_, _04450_ }), .Y(_08534_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31813_ ( .A({ _08535_, _04673_, _08508_ }), .Y(_22886_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31814_ ( .A({ _04577_, _08507_, _08509_, _04449_ }), .Y(_08535_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31815_ ( .A({ _08536_, _04446_, _08509_ }), .Y(_22883_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31816_ ( .A({ _04574_, _08507_, _04670_, _08508_ }), .Y(_08536_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31817_ ( .A({ _08537_, _04659_, _08508_ }), .Y(_22872_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31818_ ( .A({ _04563_, _08507_, _08509_, _04435_ }), .Y(_08537_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31819_ ( .A({ _08538_, _04648_, _08508_ }), .Y(_22861_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31820_ ( .A({ _04552_, _08507_, _08509_, _04424_ }), .Y(_08538_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _31821_ ( .A({ _08508_, _08509_, _08507_ }), .Y(_24079_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31822_ ( .A({ _08540_, _04416_, _08539_ }), .Y(_22917_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31823_ ( .A({ _06910_, _06886_ }), .Y(_08539_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31824_ ( .A({ _04544_, _08541_, _08542_, _04384_ }), .Y(_08540_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31825_ ( .A({ _06887_, _06907_, _06891_, main_fsm[4] }), .Y(_08541_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31826_ ( .A({ main_fsm[4], _06916_, _06898_, _06891_ }), .Y(_08542_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31827_ ( .A({ _08543_, _04415_, _08539_ }), .Y(_22916_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31828_ ( .A({ _04543_, _08541_, _08542_, _04383_ }), .Y(_08543_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31829_ ( .A({ _08544_, _04541_, _08541_ }), .Y(_22914_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31830_ ( .A({ _04413_, _08539_, _08542_, _04381_ }), .Y(_08544_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31831_ ( .A({ _08545_, _04540_, _08541_ }), .Y(_22913_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31832_ ( .A({ _04412_, _08539_, _08542_, _04380_ }), .Y(_08545_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31833_ ( .A({ _08546_, _04411_, _08539_ }), .Y(_22912_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31834_ ( .A({ _04539_, _08541_, _08542_, _04379_ }), .Y(_08546_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31835_ ( .A({ _08547_, _04538_, _08541_ }), .Y(_22911_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31836_ ( .A({ _04410_, _08539_, _08542_, _04378_ }), .Y(_08547_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31837_ ( .A({ _08548_, _04409_, _08539_ }), .Y(_22910_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31838_ ( .A({ _04537_, _08541_, _08542_, _04377_ }), .Y(_08548_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31839_ ( .A({ _08549_, _04536_, _08541_ }), .Y(_22909_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31840_ ( .A({ _04408_, _08539_, _08542_, _04376_ }), .Y(_08549_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31841_ ( .A({ _08550_, _04535_, _08541_ }), .Y(_22908_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31842_ ( .A({ _04407_, _08539_, _08542_, _04375_ }), .Y(_08550_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31843_ ( .A({ _08551_, _04406_, _08539_ }), .Y(_22907_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31844_ ( .A({ _04534_, _08541_, _08542_, _04374_ }), .Y(_08551_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31845_ ( .A({ _08552_, _04405_, _08539_ }), .Y(_22906_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31846_ ( .A({ _04533_, _08541_, _08542_, _04373_ }), .Y(_08552_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31847_ ( .A({ _08553_, _04404_, _08539_ }), .Y(_22905_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31848_ ( .A({ _04532_, _08541_, _08542_, _04372_ }), .Y(_08553_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31849_ ( .A({ _08554_, _04530_, _08541_ }), .Y(_22903_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31850_ ( .A({ _04402_, _08539_, _08542_, _04370_ }), .Y(_08554_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31851_ ( .A({ _08555_, _04401_, _08539_ }), .Y(_22902_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31852_ ( .A({ _04529_, _08541_, _08542_, _04369_ }), .Y(_08555_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31853_ ( .A({ _08556_, _04528_, _08541_ }), .Y(_22901_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31854_ ( .A({ _04400_, _08539_, _08542_, _04368_ }), .Y(_08556_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31855_ ( .A({ _08557_, _04527_, _08541_ }), .Y(_22900_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31856_ ( .A({ _04399_, _08539_, _08542_, _04367_ }), .Y(_08557_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31857_ ( .A({ _08558_, _04526_, _08541_ }), .Y(_22899_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31858_ ( .A({ _04398_, _08539_, _08542_, _04366_ }), .Y(_08558_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31859_ ( .A({ _08559_, _04525_, _08541_ }), .Y(_22898_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31860_ ( .A({ _04397_, _08539_, _08542_, _04365_ }), .Y(_08559_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31861_ ( .A({ _08560_, _04396_, _08539_ }), .Y(_22897_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31862_ ( .A({ _04524_, _08541_, _08542_, _04364_ }), .Y(_08560_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31863_ ( .A({ _08561_, _04395_, _08539_ }), .Y(_22896_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31864_ ( .A({ _04523_, _08541_, _08542_, _04363_ }), .Y(_08561_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31865_ ( .A({ _08562_, _04394_, _08539_ }), .Y(_22895_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31866_ ( .A({ _04522_, _08541_, _08542_, _04362_ }), .Y(_08562_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31867_ ( .A({ _08563_, _04393_, _08539_ }), .Y(_22894_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31868_ ( .A({ _04521_, _08541_, _08542_, _04361_ }), .Y(_08563_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31869_ ( .A({ _08564_, _04423_, _08539_ }), .Y(_22924_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31870_ ( .A({ _04551_, _08541_, _08542_, _04391_ }), .Y(_08564_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31871_ ( .A({ _08565_, _04550_, _08541_ }), .Y(_22923_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31872_ ( .A({ _04422_, _08539_, _08542_, _04390_ }), .Y(_08565_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31873_ ( .A({ _08566_, _04421_, _08539_ }), .Y(_22922_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31874_ ( .A({ _04549_, _08541_, _08542_, _04389_ }), .Y(_08566_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31875_ ( .A({ _08567_, _04420_, _08539_ }), .Y(_22921_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31876_ ( .A({ _04548_, _08541_, _08542_, _04388_ }), .Y(_08567_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31877_ ( .A({ _08568_, _04547_, _08541_ }), .Y(_22920_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31878_ ( .A({ _04419_, _08539_, _08542_, _04387_ }), .Y(_08568_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31879_ ( .A({ _08569_, _04418_, _08539_ }), .Y(_22919_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31880_ ( .A({ _04546_, _08541_, _08542_, _04386_ }), .Y(_08569_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31881_ ( .A({ _08570_, _04545_, _08541_ }), .Y(_22918_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31882_ ( .A({ _04417_, _08539_, _08542_, _04385_ }), .Y(_08570_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31883_ ( .A({ _08571_, _04414_, _08539_ }), .Y(_22915_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31884_ ( .A({ _04542_, _08541_, _08542_, _04382_ }), .Y(_08571_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31885_ ( .A({ _08572_, _04403_, _08539_ }), .Y(_22904_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31886_ ( .A({ _04531_, _08541_, _08542_, _04371_ }), .Y(_08572_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31887_ ( .A({ _08573_, _04520_, _08541_ }), .Y(_22893_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31888_ ( .A({ _04392_, _08539_, _08542_, _04360_ }), .Y(_08573_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _31889_ ( .A({ _08542_, _08541_, _08539_ }), .Y(_24080_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31890_ ( .A({ _08574_, _04544_, _08578_ }), .Y(_22949_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31891_ ( .A({ _04416_, _08575_, _saxi_register_11[31], _08577_ }), .Y(_08574_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _31892_ ( .A({ main_fsm[4], _08576_, _06898_, _06891_ }), .Y(_08575_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _31893_ ( .A({ main_fsm[1], main_fsm[3], main_fsm[0], main_fsm[2] }), .Y(_08576_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31894_ ( .A({ _06887_, _06914_, _06891_, main_fsm[4] }), .Y(_08577_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31895_ ( .A({ _06887_, _06902_, _06891_, main_fsm[4] }), .Y(_08578_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31896_ ( .A({ _08579_, _04543_, _08578_ }), .Y(_22948_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31897_ ( .A({ _04415_, _08575_, _saxi_register_11[30], _08577_ }), .Y(_08579_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31898_ ( .A({ _08580_, _saxi_register_11[29], _08577_ }), .Y(_22946_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31899_ ( .A({ _04541_, _08578_, _08575_, _04413_ }), .Y(_08580_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31900_ ( .A({ _08581_, _04540_, _08578_ }), .Y(_22945_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31901_ ( .A({ _04412_, _08575_, _saxi_register_11[28], _08577_ }), .Y(_08581_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31902_ ( .A({ _08582_, _04539_, _08578_ }), .Y(_22944_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31903_ ( .A({ _04411_, _08575_, _saxi_register_11[27], _08577_ }), .Y(_08582_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31904_ ( .A({ _08583_, _04538_, _08578_ }), .Y(_22943_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31905_ ( .A({ _04410_, _08575_, _saxi_register_11[26], _08577_ }), .Y(_08583_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31906_ ( .A({ _08584_, _04537_, _08578_ }), .Y(_22942_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31907_ ( .A({ _04409_, _08575_, _saxi_register_11[25], _08577_ }), .Y(_08584_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31908_ ( .A({ _08585_, _04536_, _08578_ }), .Y(_22941_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31909_ ( .A({ _04408_, _08575_, _saxi_register_11[24], _08577_ }), .Y(_08585_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31910_ ( .A({ _08586_, _saxi_register_11[23], _08577_ }), .Y(_22940_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31911_ ( .A({ _04535_, _08578_, _08575_, _04407_ }), .Y(_08586_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31912_ ( .A({ _08587_, _saxi_register_11[22], _08577_ }), .Y(_22939_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31913_ ( .A({ _04534_, _08578_, _08575_, _04406_ }), .Y(_08587_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31914_ ( .A({ _08588_, _saxi_register_11[21], _08577_ }), .Y(_22938_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31915_ ( .A({ _04533_, _08578_, _08575_, _04405_ }), .Y(_08588_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31916_ ( .A({ _08589_, _04532_, _08578_ }), .Y(_22937_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31917_ ( .A({ _04404_, _08575_, _saxi_register_11[20], _08577_ }), .Y(_08589_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31918_ ( .A({ _08590_, _saxi_register_11[19], _08577_ }), .Y(_22935_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31919_ ( .A({ _04530_, _08578_, _08575_, _04402_ }), .Y(_08590_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31920_ ( .A({ _08591_, _04529_, _08578_ }), .Y(_22934_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31921_ ( .A({ _04401_, _08575_, _saxi_register_11[18], _08577_ }), .Y(_08591_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31922_ ( .A({ _08592_, _saxi_register_11[17], _08577_ }), .Y(_22933_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31923_ ( .A({ _04528_, _08578_, _08575_, _04400_ }), .Y(_08592_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31924_ ( .A({ _08593_, _saxi_register_11[16], _08577_ }), .Y(_22932_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31925_ ( .A({ _04527_, _08578_, _08575_, _04399_ }), .Y(_08593_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31926_ ( .A({ _08594_, _04526_, _08578_ }), .Y(_22931_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31927_ ( .A({ _04398_, _08575_, _saxi_register_11[15], _08577_ }), .Y(_08594_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31928_ ( .A({ _08595_, _04525_, _08578_ }), .Y(_22930_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31929_ ( .A({ _04397_, _08575_, _saxi_register_11[14], _08577_ }), .Y(_08595_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31930_ ( .A({ _08596_, _saxi_register_11[13], _08577_ }), .Y(_22929_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31931_ ( .A({ _04524_, _08578_, _08575_, _04396_ }), .Y(_08596_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31932_ ( .A({ _08597_, _04523_, _08578_ }), .Y(_22928_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31933_ ( .A({ _04395_, _08575_, _saxi_register_11[12], _08577_ }), .Y(_08597_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31934_ ( .A({ _08598_, _saxi_register_11[11], _08577_ }), .Y(_22927_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31935_ ( .A({ _04522_, _08578_, _08575_, _04394_ }), .Y(_08598_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31936_ ( .A({ _08599_, _saxi_register_11[10], _08577_ }), .Y(_22926_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31937_ ( .A({ _04521_, _08578_, _08575_, _04393_ }), .Y(_08599_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31938_ ( .A({ _08600_, _04551_, _08578_ }), .Y(_22956_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31939_ ( .A({ _04423_, _08575_, _saxi_register_11[9], _08577_ }), .Y(_08600_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31940_ ( .A({ _08601_, _saxi_register_11[8], _08577_ }), .Y(_22955_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31941_ ( .A({ _04550_, _08578_, _08575_, _04422_ }), .Y(_08601_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31942_ ( .A({ _08602_, _saxi_register_11[7], _08577_ }), .Y(_22954_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31943_ ( .A({ _04549_, _08578_, _08575_, _04421_ }), .Y(_08602_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31944_ ( .A({ _08603_, _04548_, _08578_ }), .Y(_22953_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31945_ ( .A({ _04420_, _08575_, _saxi_register_11[6], _08577_ }), .Y(_08603_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31946_ ( .A({ _08604_, _saxi_register_11[5], _08577_ }), .Y(_22952_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31947_ ( .A({ _04547_, _08578_, _08575_, _04419_ }), .Y(_08604_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31948_ ( .A({ _08605_, _04546_, _08578_ }), .Y(_22951_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31949_ ( .A({ _04418_, _08575_, _saxi_register_11[4], _08577_ }), .Y(_08605_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31950_ ( .A({ _08606_, _saxi_register_11[3], _08577_ }), .Y(_22950_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31951_ ( .A({ _04545_, _08578_, _08575_, _04417_ }), .Y(_08606_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31952_ ( .A({ _08607_, _04542_, _08578_ }), .Y(_22947_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31953_ ( .A({ _04414_, _08575_, _saxi_register_11[2], _08577_ }), .Y(_08607_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31954_ ( .A({ _08608_, _saxi_register_11[1], _08577_ }), .Y(_22936_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31955_ ( .A({ _04531_, _08578_, _08575_, _04403_ }), .Y(_08608_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31956_ ( .A({ _08609_, _saxi_register_11[0], _08577_ }), .Y(_22925_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31957_ ( .A({ _04520_, _08578_, _08575_, _04392_ }), .Y(_08609_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _31958_ ( .A({ _08577_, _08575_, _08578_ }), .Y(_24081_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31959_ ( .A({ _08610_, _04096_, _08613_ }), .Y(_22981_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31960_ ( .A({ _saxi_register_10[31], _08611_, _04256_, _08612_ }), .Y(_08610_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31961_ ( .A({ _06897_, _06908_ }), .Y(_08611_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _31962_ ( .A({ _06911_, _06901_ }), .Y(_08612_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _31963_ ( .A({ _06891_, _06917_, _06898_, main_fsm[4] }), .Y(_08613_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31964_ ( .A({ _08614_, _04095_, _08613_ }), .Y(_22980_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31965_ ( .A({ _saxi_register_10[30], _08611_, _04255_, _08612_ }), .Y(_08614_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31966_ ( .A({ _08615_, _04093_, _08613_ }), .Y(_22978_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31967_ ( .A({ _saxi_register_10[29], _08611_, _04253_, _08612_ }), .Y(_08615_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31968_ ( .A({ _08616_, _04092_, _08613_ }), .Y(_22977_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31969_ ( .A({ _saxi_register_10[28], _08611_, _04252_, _08612_ }), .Y(_08616_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31970_ ( .A({ _08617_, _04091_, _08613_ }), .Y(_22976_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31971_ ( .A({ _saxi_register_10[27], _08611_, _04251_, _08612_ }), .Y(_08617_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31972_ ( .A({ _08618_, _04090_, _08613_ }), .Y(_22975_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31973_ ( .A({ _saxi_register_10[26], _08611_, _04250_, _08612_ }), .Y(_08618_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31974_ ( .A({ _08619_, _04089_, _08613_ }), .Y(_22974_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31975_ ( .A({ _saxi_register_10[25], _08611_, _04249_, _08612_ }), .Y(_08619_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31976_ ( .A({ _08620_, _04088_, _08613_ }), .Y(_22973_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31977_ ( .A({ _saxi_register_10[24], _08611_, _04248_, _08612_ }), .Y(_08620_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31978_ ( .A({ _08621_, _04087_, _08613_ }), .Y(_22972_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31979_ ( .A({ _saxi_register_10[23], _08611_, _04247_, _08612_ }), .Y(_08621_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31980_ ( .A({ _08622_, _04086_, _08613_ }), .Y(_22971_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31981_ ( .A({ _saxi_register_10[22], _08611_, _04246_, _08612_ }), .Y(_08622_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31982_ ( .A({ _08623_, _04085_, _08613_ }), .Y(_22970_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31983_ ( .A({ _saxi_register_10[21], _08611_, _04245_, _08612_ }), .Y(_08623_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31984_ ( .A({ _08624_, _04084_, _08613_ }), .Y(_22969_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31985_ ( .A({ _saxi_register_10[20], _08611_, _04244_, _08612_ }), .Y(_08624_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31986_ ( .A({ _08625_, _04082_, _08613_ }), .Y(_22967_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31987_ ( .A({ _saxi_register_10[19], _08611_, _04242_, _08612_ }), .Y(_08625_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31988_ ( .A({ _08626_, _04081_, _08613_ }), .Y(_22966_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31989_ ( .A({ _saxi_register_10[18], _08611_, _04241_, _08612_ }), .Y(_08626_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31990_ ( .A({ _08627_, _04080_, _08613_ }), .Y(_22965_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31991_ ( .A({ _saxi_register_10[17], _08611_, _04240_, _08612_ }), .Y(_08627_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31992_ ( .A({ _08628_, _04079_, _08613_ }), .Y(_22964_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31993_ ( .A({ _saxi_register_10[16], _08611_, _04239_, _08612_ }), .Y(_08628_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31994_ ( .A({ _08629_, _04078_, _08613_ }), .Y(_22963_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31995_ ( .A({ _saxi_register_10[15], _08611_, _04238_, _08612_ }), .Y(_08629_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31996_ ( .A({ _08630_, _04077_, _08613_ }), .Y(_22962_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31997_ ( .A({ _saxi_register_10[14], _08611_, _04237_, _08612_ }), .Y(_08630_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _31998_ ( .A({ _08631_, _04076_, _08613_ }), .Y(_22961_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _31999_ ( .A({ _saxi_register_10[13], _08611_, _04236_, _08612_ }), .Y(_08631_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32000_ ( .A({ _08632_, _04075_, _08613_ }), .Y(_22960_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32001_ ( .A({ _saxi_register_10[12], _08611_, _04235_, _08612_ }), .Y(_08632_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32002_ ( .A({ _08633_, _04074_, _08613_ }), .Y(_22959_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32003_ ( .A({ _saxi_register_10[11], _08611_, _04234_, _08612_ }), .Y(_08633_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32004_ ( .A({ _08634_, _04073_, _08613_ }), .Y(_22958_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32005_ ( .A({ _saxi_register_10[10], _08611_, _04233_, _08612_ }), .Y(_08634_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32006_ ( .A({ _08635_, _04103_, _08613_ }), .Y(_22988_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32007_ ( .A({ _saxi_register_10[9], _08611_, _04263_, _08612_ }), .Y(_08635_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32008_ ( .A({ _08636_, _04102_, _08613_ }), .Y(_22987_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32009_ ( .A({ _saxi_register_10[8], _08611_, _04262_, _08612_ }), .Y(_08636_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32010_ ( .A({ _08637_, _04101_, _08613_ }), .Y(_22986_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32011_ ( .A({ _saxi_register_10[7], _08611_, _04261_, _08612_ }), .Y(_08637_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32012_ ( .A({ _08638_, _04100_, _08613_ }), .Y(_22985_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32013_ ( .A({ _saxi_register_10[6], _08611_, _04260_, _08612_ }), .Y(_08638_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32014_ ( .A({ _08639_, _04099_, _08613_ }), .Y(_22984_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32015_ ( .A({ _saxi_register_10[5], _08611_, _04259_, _08612_ }), .Y(_08639_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32016_ ( .A({ _08640_, _04098_, _08613_ }), .Y(_22983_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32017_ ( .A({ _saxi_register_10[4], _08611_, _04258_, _08612_ }), .Y(_08640_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32018_ ( .A({ _08641_, _04097_, _08613_ }), .Y(_22982_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32019_ ( .A({ _saxi_register_10[3], _08611_, _04257_, _08612_ }), .Y(_08641_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32020_ ( .A({ _08642_, _04094_, _08613_ }), .Y(_22979_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32021_ ( .A({ _saxi_register_10[2], _08611_, _04254_, _08612_ }), .Y(_08642_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32022_ ( .A({ _08643_, _04083_, _08613_ }), .Y(_22968_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32023_ ( .A({ _saxi_register_10[1], _08611_, _04243_, _08612_ }), .Y(_08643_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32024_ ( .A({ _08644_, _04072_, _08613_ }), .Y(_22957_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32025_ ( .A({ _saxi_register_10[0], _08611_, _04232_, _08612_ }), .Y(_08644_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _32026_ ( .A({ _08613_, _08612_, _08611_ }), .Y(_24082_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32027_ ( .A({ _08645_, _04384_, _08648_ }), .Y(_23013_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32028_ ( .A({ _04064_, _08646_, _04224_, _08647_ }), .Y(_08645_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32029_ ( .A({ _06907_, _06915_ }), .Y(_08646_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _32030_ ( .A({ _06891_, _06897_, _06898_, main_fsm[4] }), .Y(_08647_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32031_ ( .A({ _06917_, _06901_ }), .Y(_08648_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32032_ ( .A({ _08649_, _04223_, _08647_ }), .Y(_23012_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32033_ ( .A({ _04383_, _08648_, _04063_, _08646_ }), .Y(_08649_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32034_ ( .A({ _08650_, _04221_, _08647_ }), .Y(_23010_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32035_ ( .A({ _04381_, _08648_, _04061_, _08646_ }), .Y(_08650_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32036_ ( .A({ _08651_, _04220_, _08647_ }), .Y(_23009_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32037_ ( .A({ _04380_, _08648_, _04060_, _08646_ }), .Y(_08651_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32038_ ( .A({ _08652_, _04219_, _08647_ }), .Y(_23008_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32039_ ( .A({ _04379_, _08648_, _04059_, _08646_ }), .Y(_08652_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32040_ ( .A({ _08653_, _04218_, _08647_ }), .Y(_23007_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32041_ ( .A({ _04378_, _08648_, _04058_, _08646_ }), .Y(_08653_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32042_ ( .A({ _08654_, _04217_, _08647_ }), .Y(_23006_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32043_ ( .A({ _04377_, _08648_, _04057_, _08646_ }), .Y(_08654_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32044_ ( .A({ _08655_, _04376_, _08648_ }), .Y(_23005_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32045_ ( .A({ _04056_, _08646_, _04216_, _08647_ }), .Y(_08655_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32046_ ( .A({ _08656_, _04215_, _08647_ }), .Y(_23004_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32047_ ( .A({ _04375_, _08648_, _04055_, _08646_ }), .Y(_08656_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32048_ ( .A({ _08657_, _04214_, _08647_ }), .Y(_23003_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32049_ ( .A({ _04374_, _08648_, _04054_, _08646_ }), .Y(_08657_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32050_ ( .A({ _08658_, _04213_, _08647_ }), .Y(_23002_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32051_ ( .A({ _04373_, _08648_, _04053_, _08646_ }), .Y(_08658_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32052_ ( .A({ _08659_, _04212_, _08647_ }), .Y(_23001_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32053_ ( .A({ _04372_, _08648_, _04052_, _08646_ }), .Y(_08659_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32054_ ( .A({ _08660_, _04210_, _08647_ }), .Y(_22999_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32055_ ( .A({ _04370_, _08648_, _04050_, _08646_ }), .Y(_08660_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32056_ ( .A({ _08661_, _04369_, _08648_ }), .Y(_22998_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32057_ ( .A({ _04049_, _08646_, _04209_, _08647_ }), .Y(_08661_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32058_ ( .A({ _08662_, _04208_, _08647_ }), .Y(_22997_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32059_ ( .A({ _04368_, _08648_, _04048_, _08646_ }), .Y(_08662_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32060_ ( .A({ _08663_, _04367_, _08648_ }), .Y(_22996_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32061_ ( .A({ _04047_, _08646_, _04207_, _08647_ }), .Y(_08663_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32062_ ( .A({ _08664_, _04206_, _08647_ }), .Y(_22995_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32063_ ( .A({ _04366_, _08648_, _04046_, _08646_ }), .Y(_08664_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32064_ ( .A({ _08665_, _04205_, _08647_ }), .Y(_22994_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32065_ ( .A({ _04365_, _08648_, _04045_, _08646_ }), .Y(_08665_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32066_ ( .A({ _08666_, _04204_, _08647_ }), .Y(_22993_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32067_ ( .A({ _04364_, _08648_, _04044_, _08646_ }), .Y(_08666_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32068_ ( .A({ _08667_, _04203_, _08647_ }), .Y(_22992_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32069_ ( .A({ _04363_, _08648_, _04043_, _08646_ }), .Y(_08667_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32070_ ( .A({ _08668_, _04202_, _08647_ }), .Y(_22991_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32071_ ( .A({ _04362_, _08648_, _04042_, _08646_ }), .Y(_08668_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32072_ ( .A({ _08669_, _04201_, _08647_ }), .Y(_22990_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32073_ ( .A({ _04361_, _08648_, _04041_, _08646_ }), .Y(_08669_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32074_ ( .A({ _08670_, _04231_, _08647_ }), .Y(_23020_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32075_ ( .A({ _04391_, _08648_, _04071_, _08646_ }), .Y(_08670_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32076_ ( .A({ _08671_, _04390_, _08648_ }), .Y(_23019_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32077_ ( .A({ _04070_, _08646_, _04230_, _08647_ }), .Y(_08671_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32078_ ( .A({ _08672_, _04229_, _08647_ }), .Y(_23018_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32079_ ( .A({ _04389_, _08648_, _04069_, _08646_ }), .Y(_08672_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32080_ ( .A({ _08673_, _04228_, _08647_ }), .Y(_23017_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32081_ ( .A({ _04388_, _08648_, _04068_, _08646_ }), .Y(_08673_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32082_ ( .A({ _08674_, _04227_, _08647_ }), .Y(_23016_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32083_ ( .A({ _04387_, _08648_, _04067_, _08646_ }), .Y(_08674_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32084_ ( .A({ _08675_, _04386_, _08648_ }), .Y(_23015_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32085_ ( .A({ _04066_, _08646_, _04226_, _08647_ }), .Y(_08675_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32086_ ( .A({ _08676_, _04225_, _08647_ }), .Y(_23014_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32087_ ( .A({ _04385_, _08648_, _04065_, _08646_ }), .Y(_08676_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32088_ ( .A({ _08677_, _04222_, _08647_ }), .Y(_23011_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32089_ ( .A({ _04382_, _08648_, _04062_, _08646_ }), .Y(_08677_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32090_ ( .A({ _08678_, _04211_, _08647_ }), .Y(_23000_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32091_ ( .A({ _04371_, _08648_, _04051_, _08646_ }), .Y(_08678_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32092_ ( .A({ _08679_, _04360_, _08648_ }), .Y(_22989_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32093_ ( .A({ _04040_, _08646_, _04200_, _08647_ }), .Y(_08679_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _32094_ ( .A({ _08647_, _08646_, _08648_ }), .Y(_24083_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32095_ ( .A({ _08680_, _04192_, _08684_ }), .Y(_23045_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32096_ ( .A({ _04032_, _08681_, _04352_, _08683_ }), .Y(_08680_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32097_ ( .A({ _08682_, _06915_ }), .Y(_08681_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _32098_ ( .A({ main_fsm[0], main_fsm[3:1] }), .Y(_08682_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32099_ ( .A({ _06916_, _06903_ }), .Y(_08683_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32100_ ( .A({ _08576_, _06908_ }), .Y(_08684_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32101_ ( .A({ _08685_, _04191_, _08684_ }), .Y(_23044_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32102_ ( .A({ _04031_, _08681_, _04351_, _08683_ }), .Y(_08685_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32103_ ( .A({ _08686_, _04349_, _08683_ }), .Y(_23042_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32104_ ( .A({ _04189_, _08684_, _08681_, _04029_ }), .Y(_08686_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32105_ ( .A({ _08687_, _04348_, _08683_ }), .Y(_23041_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32106_ ( .A({ _04188_, _08684_, _08681_, _04028_ }), .Y(_08687_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32107_ ( .A({ _08688_, _04347_, _08683_ }), .Y(_23040_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32108_ ( .A({ _04187_, _08684_, _08681_, _04027_ }), .Y(_08688_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32109_ ( .A({ _08689_, _04346_, _08683_ }), .Y(_23039_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32110_ ( .A({ _04186_, _08684_, _08681_, _04026_ }), .Y(_08689_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32111_ ( .A({ _08690_, _04185_, _08684_ }), .Y(_23038_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32112_ ( .A({ _04025_, _08681_, _04345_, _08683_ }), .Y(_08690_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32113_ ( .A({ _08691_, _04344_, _08683_ }), .Y(_23037_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32114_ ( .A({ _04184_, _08684_, _08681_, _04024_ }), .Y(_08691_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32115_ ( .A({ _08692_, _04183_, _08684_ }), .Y(_23036_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32116_ ( .A({ _04023_, _08681_, _04343_, _08683_ }), .Y(_08692_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32117_ ( .A({ _08693_, _04182_, _08684_ }), .Y(_23035_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32118_ ( .A({ _04022_, _08681_, _04342_, _08683_ }), .Y(_08693_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32119_ ( .A({ _08694_, _04181_, _08684_ }), .Y(_23034_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32120_ ( .A({ _04021_, _08681_, _04341_, _08683_ }), .Y(_08694_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32121_ ( .A({ _08695_, _04340_, _08683_ }), .Y(_23033_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32122_ ( .A({ _04180_, _08684_, _08681_, _04020_ }), .Y(_08695_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32123_ ( .A({ _08696_, _04338_, _08683_ }), .Y(_23031_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32124_ ( .A({ _04178_, _08684_, _08681_, _04018_ }), .Y(_08696_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32125_ ( .A({ _08697_, _04177_, _08684_ }), .Y(_23030_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32126_ ( .A({ _04017_, _08681_, _04337_, _08683_ }), .Y(_08697_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32127_ ( .A({ _08698_, _04336_, _08683_ }), .Y(_23029_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32128_ ( .A({ _04176_, _08684_, _08681_, _04016_ }), .Y(_08698_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32129_ ( .A({ _08699_, _04335_, _08683_ }), .Y(_23028_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32130_ ( .A({ _04175_, _08684_, _08681_, _04015_ }), .Y(_08699_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32131_ ( .A({ _08700_, _04334_, _08683_ }), .Y(_23027_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32132_ ( .A({ _04174_, _08684_, _08681_, _04014_ }), .Y(_08700_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32133_ ( .A({ _08701_, _04173_, _08684_ }), .Y(_23026_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32134_ ( .A({ _04013_, _08681_, _04333_, _08683_ }), .Y(_08701_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32135_ ( .A({ _08702_, _04332_, _08683_ }), .Y(_23025_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32136_ ( .A({ _04172_, _08684_, _08681_, _04012_ }), .Y(_08702_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32137_ ( .A({ _08703_, _04331_, _08683_ }), .Y(_23024_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32138_ ( .A({ _04171_, _08684_, _08681_, _04011_ }), .Y(_08703_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32139_ ( .A({ _08704_, _04330_, _08683_ }), .Y(_23023_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32140_ ( .A({ _04170_, _08684_, _08681_, _04010_ }), .Y(_08704_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32141_ ( .A({ _08705_, _04169_, _08684_ }), .Y(_23022_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32142_ ( .A({ _04009_, _08681_, _04329_, _08683_ }), .Y(_08705_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32143_ ( .A({ _08706_, _04359_, _08683_ }), .Y(_23052_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32144_ ( .A({ _04199_, _08684_, _08681_, _04039_ }), .Y(_08706_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32145_ ( .A({ _08707_, _04358_, _08683_ }), .Y(_23051_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32146_ ( .A({ _04198_, _08684_, _08681_, _04038_ }), .Y(_08707_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32147_ ( .A({ _08708_, _04357_, _08683_ }), .Y(_23050_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32148_ ( .A({ _04197_, _08684_, _08681_, _04037_ }), .Y(_08708_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32149_ ( .A({ _08709_, _04356_, _08683_ }), .Y(_23049_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32150_ ( .A({ _04196_, _08684_, _08681_, _04036_ }), .Y(_08709_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32151_ ( .A({ _08710_, _04195_, _08684_ }), .Y(_23048_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32152_ ( .A({ _04035_, _08681_, _04355_, _08683_ }), .Y(_08710_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32153_ ( .A({ _08711_, _04354_, _08683_ }), .Y(_23047_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32154_ ( .A({ _04194_, _08684_, _08681_, _04034_ }), .Y(_08711_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32155_ ( .A({ _08712_, _04353_, _08683_ }), .Y(_23046_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32156_ ( .A({ _04193_, _08684_, _08681_, _04033_ }), .Y(_08712_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32157_ ( .A({ _08713_, _04190_, _08684_ }), .Y(_23043_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32158_ ( .A({ _04030_, _08681_, _04350_, _08683_ }), .Y(_08713_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32159_ ( .A({ _08714_, _04339_, _08683_ }), .Y(_23032_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32160_ ( .A({ _04179_, _08684_, _08681_, _04019_ }), .Y(_08714_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32161_ ( .A({ _08715_, _04328_, _08683_ }), .Y(_23021_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32162_ ( .A({ _04168_, _08684_, _08681_, _04008_ }), .Y(_08715_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _32163_ ( .A({ _08683_, _08681_, _08684_ }), .Y(_24084_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32164_ ( .A({ _14204_, _13755_, _14236_, _08032_ }), .Y(_05581_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32165_ ( .A({ _14178_, _13755_, _14210_, _08032_ }), .Y(_05582_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32166_ ( .A({ _14189_, _13755_, _14221_, _08032_ }), .Y(_05583_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32167_ ( .A({ _14200_, _13755_, _14232_, _08032_ }), .Y(_05584_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32168_ ( .A({ _14203_, _13755_, _14235_, _08032_ }), .Y(_05585_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32169_ ( .A({ _14205_, _13755_, _14237_, _08032_ }), .Y(_05586_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32170_ ( .A({ _14206_, _13755_, _14238_, _08032_ }), .Y(_05587_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32171_ ( .A({ _14207_, _13755_, _14239_, _08032_ }), .Y(_05588_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32172_ ( .A({ _14208_, _13755_, _14240_, _08032_ }), .Y(_05589_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32173_ ( .A({ _14182_, _13755_, _14214_, _08032_ }), .Y(_05590_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32174_ ( .A({ _14209_, _13755_, _14241_, _08032_ }), .Y(_05591_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32175_ ( .A({ _14186_, _13755_, _14218_, _08032_ }), .Y(_05592_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32176_ ( .A({ _14179_, _13755_, _14211_, _08032_ }), .Y(_05593_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32177_ ( .A({ _14180_, _13755_, _14212_, _08032_ }), .Y(_05594_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32178_ ( .A({ _14181_, _13755_, _14213_, _08032_ }), .Y(_05595_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32179_ ( .A({ _14190_, _13755_, _14222_, _08032_ }), .Y(_05596_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32180_ ( .A({ _14183_, _13755_, _14215_, _08032_ }), .Y(_05597_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32181_ ( .A({ _14184_, _13755_, _14216_, _08032_ }), .Y(_05598_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32182_ ( .A({ _14185_, _13755_, _14217_, _08032_ }), .Y(_05599_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32183_ ( .A({ _14187_, _13755_, _14219_, _08032_ }), .Y(_05600_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32184_ ( .A({ _14188_, _13755_, _14220_, _08032_ }), .Y(_05601_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32185_ ( .A({ _14191_, _13755_, _14223_, _08032_ }), .Y(_05602_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32186_ ( .A({ _14194_, _13755_, _14226_, _08032_ }), .Y(_05603_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32187_ ( .A({ _14192_, _13755_, _14224_, _08032_ }), .Y(_05604_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32188_ ( .A({ _14193_, _13755_, _14225_, _08032_ }), .Y(_05605_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32189_ ( .A({ _14196_, _13755_, _14228_, _08032_ }), .Y(_05606_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32190_ ( .A({ _14195_, _13755_, _14227_, _08032_ }), .Y(_05607_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32191_ ( .A({ _14199_, _13755_, _14231_, _08032_ }), .Y(_05608_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32192_ ( .A({ _14197_, _13755_, _14229_, _08032_ }), .Y(_05609_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32193_ ( .A({ _14202_, _13755_, _14234_, _08032_ }), .Y(_05610_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32194_ ( .A({ _14198_, _13755_, _14230_, _08032_ }), .Y(_05611_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32195_ ( .A({ _14201_, _13755_, _14233_, _08032_ }), .Y(_05612_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32196_ ( .A({ _08716_, _04320_, _08719_ }), .Y(_23077_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32197_ ( .A({ _04000_, _08717_, _04160_, _08718_ }), .Y(_08716_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32198_ ( .A({ _07451_, _06915_ }), .Y(_08717_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32199_ ( .A({ _08682_, _06908_ }), .Y(_08718_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32200_ ( .A({ _08576_, _06903_ }), .Y(_08719_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32201_ ( .A({ _08720_, _04319_, _08719_ }), .Y(_23076_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32202_ ( .A({ _03999_, _08717_, _04159_, _08718_ }), .Y(_08720_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32203_ ( .A({ _08721_, _04317_, _08719_ }), .Y(_23074_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32204_ ( .A({ _03997_, _08717_, _04157_, _08718_ }), .Y(_08721_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32205_ ( .A({ _08722_, _04156_, _08718_ }), .Y(_23073_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32206_ ( .A({ _04316_, _08719_, _08717_, _03996_ }), .Y(_08722_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32207_ ( .A({ _08723_, _04155_, _08718_ }), .Y(_23072_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32208_ ( .A({ _04315_, _08719_, _08717_, _03995_ }), .Y(_08723_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32209_ ( .A({ _08724_, _04314_, _08719_ }), .Y(_23071_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32210_ ( .A({ _03994_, _08717_, _04154_, _08718_ }), .Y(_08724_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32211_ ( .A({ _08725_, _04153_, _08718_ }), .Y(_23070_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32212_ ( .A({ _04313_, _08719_, _08717_, _03993_ }), .Y(_08725_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32213_ ( .A({ _08726_, _04152_, _08718_ }), .Y(_23069_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32214_ ( .A({ _04312_, _08719_, _08717_, _03992_ }), .Y(_08726_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32215_ ( .A({ _08727_, _04311_, _08719_ }), .Y(_23068_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32216_ ( .A({ _03991_, _08717_, _04151_, _08718_ }), .Y(_08727_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32217_ ( .A({ _08728_, _04150_, _08718_ }), .Y(_23067_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32218_ ( .A({ _04310_, _08719_, _08717_, _03990_ }), .Y(_08728_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32219_ ( .A({ _08729_, _04149_, _08718_ }), .Y(_23066_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32220_ ( .A({ _04309_, _08719_, _08717_, _03989_ }), .Y(_08729_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32221_ ( .A({ _08730_, _04308_, _08719_ }), .Y(_23065_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32222_ ( .A({ _03988_, _08717_, _04148_, _08718_ }), .Y(_08730_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32223_ ( .A({ _08731_, _04306_, _08719_ }), .Y(_23063_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32224_ ( .A({ _03986_, _08717_, _04146_, _08718_ }), .Y(_08731_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32225_ ( .A({ _08732_, _04305_, _08719_ }), .Y(_23062_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32226_ ( .A({ _03985_, _08717_, _04145_, _08718_ }), .Y(_08732_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32227_ ( .A({ _08733_, _04304_, _08719_ }), .Y(_23061_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32228_ ( .A({ _03984_, _08717_, _04144_, _08718_ }), .Y(_08733_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32229_ ( .A({ _08734_, _04143_, _08718_ }), .Y(_23060_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32230_ ( .A({ _04303_, _08719_, _08717_, _03983_ }), .Y(_08734_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32231_ ( .A({ _08735_, _04142_, _08718_ }), .Y(_23059_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32232_ ( .A({ _04302_, _08719_, _08717_, _03982_ }), .Y(_08735_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32233_ ( .A({ _08736_, _04301_, _08719_ }), .Y(_23058_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32234_ ( .A({ _03981_, _08717_, _04141_, _08718_ }), .Y(_08736_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32235_ ( .A({ _08737_, _04140_, _08718_ }), .Y(_23057_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32236_ ( .A({ _04300_, _08719_, _08717_, _03980_ }), .Y(_08737_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32237_ ( .A({ _08738_, _04299_, _08719_ }), .Y(_23056_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32238_ ( .A({ _03979_, _08717_, _04139_, _08718_ }), .Y(_08738_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32239_ ( .A({ _08739_, _04298_, _08719_ }), .Y(_23055_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32240_ ( .A({ _03978_, _08717_, _04138_, _08718_ }), .Y(_08739_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32241_ ( .A({ _08740_, _04137_, _08718_ }), .Y(_23054_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32242_ ( .A({ _04297_, _08719_, _08717_, _03977_ }), .Y(_08740_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32243_ ( .A({ _08741_, _04167_, _08718_ }), .Y(_23084_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32244_ ( .A({ _04327_, _08719_, _08717_, _04007_ }), .Y(_08741_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32245_ ( .A({ _08742_, _04326_, _08719_ }), .Y(_23083_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32246_ ( .A({ _04006_, _08717_, _04166_, _08718_ }), .Y(_08742_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32247_ ( .A({ _08743_, _04325_, _08719_ }), .Y(_23082_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32248_ ( .A({ _04005_, _08717_, _04165_, _08718_ }), .Y(_08743_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32249_ ( .A({ _08744_, _04324_, _08719_ }), .Y(_23081_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32250_ ( .A({ _04004_, _08717_, _04164_, _08718_ }), .Y(_08744_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32251_ ( .A({ _08745_, _04323_, _08719_ }), .Y(_23080_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32252_ ( .A({ _04003_, _08717_, _04163_, _08718_ }), .Y(_08745_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32253_ ( .A({ _08746_, _04162_, _08718_ }), .Y(_23079_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32254_ ( .A({ _04322_, _08719_, _08717_, _04002_ }), .Y(_08746_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32255_ ( .A({ _08747_, _04161_, _08718_ }), .Y(_23078_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32256_ ( .A({ _04321_, _08719_, _08717_, _04001_ }), .Y(_08747_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32257_ ( .A({ _08748_, _04318_, _08719_ }), .Y(_23075_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32258_ ( .A({ _03998_, _08717_, _04158_, _08718_ }), .Y(_08748_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32259_ ( .A({ _08749_, _04147_, _08718_ }), .Y(_23064_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32260_ ( .A({ _04307_, _08719_, _08717_, _03987_ }), .Y(_08749_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32261_ ( .A({ _08750_, _04136_, _08718_ }), .Y(_23053_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32262_ ( .A({ _04296_, _08719_, _08717_, _03976_ }), .Y(_08750_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _32263_ ( .A({ _08718_, _08717_, _08719_ }), .Y(_24085_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32264_ ( .A({ _08751_, _04128_, _08754_ }), .Y(_23109_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32265_ ( .A({ _04288_, _08752_, _08753_, _saxi_register_13[31] }), .Y(_08751_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32266_ ( .A({ _08682_, _06903_ }), .Y(_08752_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32267_ ( .A({ _06900_, _06915_ }), .Y(_08753_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32268_ ( .A({ main_fsm[4], _07451_, _06906_, _06891_ }), .Y(_08754_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32269_ ( .A({ _08755_, _04287_, _08752_ }), .Y(_23108_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32270_ ( .A({ _saxi_register_13[30], _08753_, _04127_, _08754_ }), .Y(_08755_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32271_ ( .A({ _08756_, _04285_, _08752_ }), .Y(_23106_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32272_ ( .A({ _saxi_register_13[29], _08753_, _04125_, _08754_ }), .Y(_08756_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32273_ ( .A({ _08757_, _04284_, _08752_ }), .Y(_23105_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32274_ ( .A({ _saxi_register_13[28], _08753_, _04124_, _08754_ }), .Y(_08757_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32275_ ( .A({ _08758_, _04123_, _08754_ }), .Y(_23104_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32276_ ( .A({ _04283_, _08752_, _08753_, _saxi_register_13[27] }), .Y(_08758_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32277_ ( .A({ _08759_, _04122_, _08754_ }), .Y(_23103_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32278_ ( .A({ _04282_, _08752_, _08753_, _saxi_register_13[26] }), .Y(_08759_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32279_ ( .A({ _08760_, _04121_, _08754_ }), .Y(_23102_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32280_ ( .A({ _04281_, _08752_, _08753_, _saxi_register_13[25] }), .Y(_08760_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32281_ ( .A({ _08761_, _04120_, _08754_ }), .Y(_23101_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32282_ ( .A({ _04280_, _08752_, _08753_, _saxi_register_13[24] }), .Y(_08761_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32283_ ( .A({ _08762_, _04119_, _08754_ }), .Y(_23100_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32284_ ( .A({ _04279_, _08752_, _08753_, _saxi_register_13[23] }), .Y(_08762_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32285_ ( .A({ _08763_, _04118_, _08754_ }), .Y(_23099_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32286_ ( .A({ _04278_, _08752_, _08753_, _saxi_register_13[22] }), .Y(_08763_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32287_ ( .A({ _08764_, _04277_, _08752_ }), .Y(_23098_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32288_ ( .A({ _saxi_register_13[21], _08753_, _04117_, _08754_ }), .Y(_08764_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32289_ ( .A({ _08765_, _04276_, _08752_ }), .Y(_23097_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32290_ ( .A({ _saxi_register_13[20], _08753_, _04116_, _08754_ }), .Y(_08765_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32291_ ( .A({ _08766_, _04274_, _08752_ }), .Y(_23095_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32292_ ( .A({ _saxi_register_13[19], _08753_, _04114_, _08754_ }), .Y(_08766_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32293_ ( .A({ _08767_, _04273_, _08752_ }), .Y(_23094_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32294_ ( .A({ _saxi_register_13[18], _08753_, _04113_, _08754_ }), .Y(_08767_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32295_ ( .A({ _08768_, _04272_, _08752_ }), .Y(_23093_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32296_ ( .A({ _saxi_register_13[17], _08753_, _04112_, _08754_ }), .Y(_08768_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32297_ ( .A({ _08769_, _04271_, _08752_ }), .Y(_23092_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32298_ ( .A({ _saxi_register_13[16], _08753_, _04111_, _08754_ }), .Y(_08769_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32299_ ( .A({ _08770_, _04270_, _08752_ }), .Y(_23091_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32300_ ( .A({ _saxi_register_13[15], _08753_, _04110_, _08754_ }), .Y(_08770_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32301_ ( .A({ _08771_, _04269_, _08752_ }), .Y(_23090_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32302_ ( .A({ _saxi_register_13[14], _08753_, _04109_, _08754_ }), .Y(_08771_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32303_ ( .A({ _08772_, _04268_, _08752_ }), .Y(_23089_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32304_ ( .A({ _saxi_register_13[13], _08753_, _04108_, _08754_ }), .Y(_08772_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32305_ ( .A({ _08773_, _04267_, _08752_ }), .Y(_23088_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32306_ ( .A({ _saxi_register_13[12], _08753_, _04107_, _08754_ }), .Y(_08773_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32307_ ( .A({ _08774_, _04106_, _08754_ }), .Y(_23087_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32308_ ( .A({ _04266_, _08752_, _08753_, _saxi_register_13[11] }), .Y(_08774_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32309_ ( .A({ _08775_, _04105_, _08754_ }), .Y(_23086_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32310_ ( .A({ _04265_, _08752_, _08753_, _saxi_register_13[10] }), .Y(_08775_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32311_ ( .A({ _08776_, _04295_, _08752_ }), .Y(_23116_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32312_ ( .A({ _saxi_register_13[9], _08753_, _04135_, _08754_ }), .Y(_08776_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32313_ ( .A({ _08777_, _04294_, _08752_ }), .Y(_23115_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32314_ ( .A({ _saxi_register_13[8], _08753_, _04134_, _08754_ }), .Y(_08777_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32315_ ( .A({ _08778_, _04133_, _08754_ }), .Y(_23114_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32316_ ( .A({ _04293_, _08752_, _08753_, _saxi_register_13[7] }), .Y(_08778_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32317_ ( .A({ _08779_, _04132_, _08754_ }), .Y(_23113_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32318_ ( .A({ _04292_, _08752_, _08753_, _saxi_register_13[6] }), .Y(_08779_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32319_ ( .A({ _08780_, _04291_, _08752_ }), .Y(_23112_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32320_ ( .A({ _saxi_register_13[5], _08753_, _04131_, _08754_ }), .Y(_08780_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32321_ ( .A({ _08781_, _04290_, _08752_ }), .Y(_23111_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32322_ ( .A({ _saxi_register_13[4], _08753_, _04130_, _08754_ }), .Y(_08781_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32323_ ( .A({ _08782_, _04289_, _08752_ }), .Y(_23110_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32324_ ( .A({ _saxi_register_13[3], _08753_, _04129_, _08754_ }), .Y(_08782_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32325_ ( .A({ _08783_, _04126_, _08754_ }), .Y(_23107_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32326_ ( .A({ _04286_, _08752_, _08753_, _saxi_register_13[2] }), .Y(_08783_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32327_ ( .A({ _08784_, _04275_, _08752_ }), .Y(_23096_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32328_ ( .A({ _saxi_register_13[1], _08753_, _04115_, _08754_ }), .Y(_08784_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32329_ ( .A({ _08785_, _04264_, _08752_ }), .Y(_23085_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32330_ ( .A({ _saxi_register_13[0], _08753_, _04104_, _08754_ }), .Y(_08785_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _32331_ ( .A({ _08754_, _08753_, _08752_ }), .Y(_24086_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32332_ ( .A({ _08786_, _04064_, _08789_ }), .Y(_23141_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32333_ ( .A({ _saxi_register_12[31], _08787_, _08788_, _04224_ }), .Y(_08786_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32334_ ( .A({ _06905_, _06915_ }), .Y(_08787_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _32335_ ( .A({ _06891_, _07451_, _06898_, main_fsm[4] }), .Y(_08788_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32336_ ( .A({ main_fsm[4], _06900_, _06906_, _06891_ }), .Y(_08789_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32337_ ( .A({ _08790_, _04223_, _08788_ }), .Y(_23140_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32338_ ( .A({ _saxi_register_12[30], _08787_, _08789_, _04063_ }), .Y(_08790_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32339_ ( .A({ _08791_, _04221_, _08788_ }), .Y(_23138_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32340_ ( .A({ _saxi_register_12[29], _08787_, _08789_, _04061_ }), .Y(_08791_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32341_ ( .A({ _08792_, _04220_, _08788_ }), .Y(_23137_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32342_ ( .A({ _saxi_register_12[28], _08787_, _08789_, _04060_ }), .Y(_08792_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32343_ ( .A({ _08793_, _04219_, _08788_ }), .Y(_23136_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32344_ ( .A({ _saxi_register_12[27], _08787_, _08789_, _04059_ }), .Y(_08793_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32345_ ( .A({ _08794_, _04058_, _08789_ }), .Y(_23135_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32346_ ( .A({ _saxi_register_12[26], _08787_, _08788_, _04218_ }), .Y(_08794_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32347_ ( .A({ _08795_, _04217_, _08788_ }), .Y(_23134_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32348_ ( .A({ _saxi_register_12[25], _08787_, _08789_, _04057_ }), .Y(_08795_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32349_ ( .A({ _08796_, _04056_, _08789_ }), .Y(_23133_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32350_ ( .A({ _saxi_register_12[24], _08787_, _08788_, _04216_ }), .Y(_08796_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32351_ ( .A({ _08797_, _04055_, _08789_ }), .Y(_23132_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32352_ ( .A({ _saxi_register_12[23], _08787_, _08788_, _04215_ }), .Y(_08797_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32353_ ( .A({ _08798_, _04214_, _08788_ }), .Y(_23131_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32354_ ( .A({ _saxi_register_12[22], _08787_, _08789_, _04054_ }), .Y(_08798_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32355_ ( .A({ _08799_, _04053_, _08789_ }), .Y(_23130_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32356_ ( .A({ _saxi_register_12[21], _08787_, _08788_, _04213_ }), .Y(_08799_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32357_ ( .A({ _08800_, _04212_, _08788_ }), .Y(_23129_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32358_ ( .A({ _saxi_register_12[20], _08787_, _08789_, _04052_ }), .Y(_08800_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32359_ ( .A({ _08801_, _04210_, _08788_ }), .Y(_23127_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32360_ ( .A({ _saxi_register_12[19], _08787_, _08789_, _04050_ }), .Y(_08801_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32361_ ( .A({ _08802_, _04209_, _08788_ }), .Y(_23126_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32362_ ( .A({ _saxi_register_12[18], _08787_, _08789_, _04049_ }), .Y(_08802_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32363_ ( .A({ _08803_, _04048_, _08789_ }), .Y(_23125_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32364_ ( .A({ _saxi_register_12[17], _08787_, _08788_, _04208_ }), .Y(_08803_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32365_ ( .A({ _08804_, _04207_, _08788_ }), .Y(_23124_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32366_ ( .A({ _saxi_register_12[16], _08787_, _08789_, _04047_ }), .Y(_08804_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32367_ ( .A({ _08805_, _04206_, _08788_ }), .Y(_23123_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32368_ ( .A({ _saxi_register_12[15], _08787_, _08789_, _04046_ }), .Y(_08805_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32369_ ( .A({ _08806_, _04205_, _08788_ }), .Y(_23122_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32370_ ( .A({ _saxi_register_12[14], _08787_, _08789_, _04045_ }), .Y(_08806_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32371_ ( .A({ _08807_, _04044_, _08789_ }), .Y(_23121_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32372_ ( .A({ _saxi_register_12[13], _08787_, _08788_, _04204_ }), .Y(_08807_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32373_ ( .A({ _08808_, _04203_, _08788_ }), .Y(_23120_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32374_ ( .A({ _saxi_register_12[12], _08787_, _08789_, _04043_ }), .Y(_08808_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32375_ ( .A({ _08809_, _04202_, _08788_ }), .Y(_23119_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32376_ ( .A({ _saxi_register_12[11], _08787_, _08789_, _04042_ }), .Y(_08809_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32377_ ( .A({ _08810_, _04041_, _08789_ }), .Y(_23118_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32378_ ( .A({ _saxi_register_12[10], _08787_, _08788_, _04201_ }), .Y(_08810_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32379_ ( .A({ _08811_, _04071_, _08789_ }), .Y(_23148_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32380_ ( .A({ _saxi_register_12[9], _08787_, _08788_, _04231_ }), .Y(_08811_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32381_ ( .A({ _08812_, _04070_, _08789_ }), .Y(_23147_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32382_ ( .A({ _saxi_register_12[8], _08787_, _08788_, _04230_ }), .Y(_08812_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32383_ ( .A({ _08813_, _04069_, _08789_ }), .Y(_23146_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32384_ ( .A({ _saxi_register_12[7], _08787_, _08788_, _04229_ }), .Y(_08813_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32385_ ( .A({ _08814_, _04228_, _08788_ }), .Y(_23145_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32386_ ( .A({ _saxi_register_12[6], _08787_, _08789_, _04068_ }), .Y(_08814_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32387_ ( .A({ _08815_, _04067_, _08789_ }), .Y(_23144_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32388_ ( .A({ _saxi_register_12[5], _08787_, _08788_, _04227_ }), .Y(_08815_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32389_ ( .A({ _08816_, _04226_, _08788_ }), .Y(_23143_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32390_ ( .A({ _saxi_register_12[4], _08787_, _08789_, _04066_ }), .Y(_08816_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32391_ ( .A({ _13760_, _13755_, _13792_, _08032_ }), .Y(_05613_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32392_ ( .A({ _13771_, _13755_, _13803_, _08032_ }), .Y(_05614_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32393_ ( .A({ _13782_, _13755_, _13814_, _08032_ }), .Y(_05615_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32394_ ( .A({ _13785_, _13755_, _13817_, _08032_ }), .Y(_05616_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32395_ ( .A({ _13786_, _13755_, _13818_, _08032_ }), .Y(_05617_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32396_ ( .A({ _13787_, _13755_, _13819_, _08032_ }), .Y(_05618_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32397_ ( .A({ _13788_, _13755_, _13820_, _08032_ }), .Y(_05619_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32398_ ( .A({ _13789_, _13755_, _13821_, _08032_ }), .Y(_05620_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32399_ ( .A({ _13790_, _13755_, _13822_, _08032_ }), .Y(_05621_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32400_ ( .A({ _13791_, _13755_, _13823_, _08032_ }), .Y(_05622_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32401_ ( .A({ _13761_, _13755_, _13793_, _08032_ }), .Y(_05623_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32402_ ( .A({ _13762_, _13755_, _13794_, _08032_ }), .Y(_05624_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32403_ ( .A({ _13763_, _13755_, _13795_, _08032_ }), .Y(_05625_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32404_ ( .A({ _13764_, _13755_, _13796_, _08032_ }), .Y(_05626_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32405_ ( .A({ _13765_, _13755_, _13797_, _08032_ }), .Y(_05627_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32406_ ( .A({ _13766_, _13755_, _13798_, _08032_ }), .Y(_05628_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32407_ ( .A({ _13767_, _13755_, _13799_, _08032_ }), .Y(_05629_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32408_ ( .A({ _13768_, _13755_, _13800_, _08032_ }), .Y(_05630_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32409_ ( .A({ _13769_, _13755_, _13801_, _08032_ }), .Y(_05631_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32410_ ( .A({ _13770_, _13755_, _13802_, _08032_ }), .Y(_05632_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32411_ ( .A({ _13772_, _13755_, _13804_, _08032_ }), .Y(_05633_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32412_ ( .A({ _13773_, _13755_, _13805_, _08032_ }), .Y(_05634_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32413_ ( .A({ _13774_, _13755_, _13806_, _08032_ }), .Y(_05635_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32414_ ( .A({ _13775_, _13755_, _13807_, _08032_ }), .Y(_05636_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32415_ ( .A({ _13776_, _13755_, _13808_, _08032_ }), .Y(_05637_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32416_ ( .A({ _13777_, _13755_, _13809_, _08032_ }), .Y(_05638_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32417_ ( .A({ _13780_, _13755_, _13812_, _08032_ }), .Y(_05639_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32418_ ( .A({ _13781_, _13755_, _13813_, _08032_ }), .Y(_05640_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32419_ ( .A({ _13778_, _13755_, _13810_, _08032_ }), .Y(_05641_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32420_ ( .A({ _13779_, _13755_, _13811_, _08032_ }), .Y(_05642_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32421_ ( .A({ _13783_, _13755_, _13815_, _08032_ }), .Y(_05643_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _32422_ ( .A({ _13784_, _13755_, _13816_, _08032_ }), .Y(_05644_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32423_ ( .A({ _08817_, _04065_, _08789_ }), .Y(_23142_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32424_ ( .A({ _saxi_register_12[3], _08787_, _08788_, _04225_ }), .Y(_08817_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32425_ ( .A({ _08818_, _04062_, _08789_ }), .Y(_23139_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32426_ ( .A({ _saxi_register_12[2], _08787_, _08788_, _04222_ }), .Y(_08818_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32427_ ( .A({ _08819_, _04211_, _08788_ }), .Y(_23128_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32428_ ( .A({ _saxi_register_12[1], _08787_, _08789_, _04051_ }), .Y(_08819_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32429_ ( .A({ _08820_, _04040_, _08789_ }), .Y(_23117_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32430_ ( .A({ _saxi_register_12[0], _08787_, _08788_, _04200_ }), .Y(_08820_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _32431_ ( .A({ _08788_, _08789_, _08787_ }), .Y(_24087_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32432_ ( .A({ _08821_, _04256_, _08824_ }), .Y(_23173_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32433_ ( .A({ _saxi_register_10[31], _08822_, _04096_, _08823_ }), .Y(_08821_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32434_ ( .A({ _06910_, _06915_ }), .Y(_08822_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32435_ ( .A({ main_fsm[4], _06905_, _06906_, _06891_ }), .Y(_08823_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _32436_ ( .A({ _06891_, _06900_, _06898_, main_fsm[4] }), .Y(_08824_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32437_ ( .A({ _08825_, _04255_, _08824_ }), .Y(_23172_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32438_ ( .A({ _saxi_register_10[30], _08822_, _04095_, _08823_ }), .Y(_08825_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32439_ ( .A({ _08826_, _04253_, _08824_ }), .Y(_23170_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32440_ ( .A({ _saxi_register_10[29], _08822_, _04093_, _08823_ }), .Y(_08826_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32441_ ( .A({ _08827_, _04092_, _08823_ }), .Y(_23169_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32442_ ( .A({ _saxi_register_10[28], _08822_, _04252_, _08824_ }), .Y(_08827_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32443_ ( .A({ _08828_, _04251_, _08824_ }), .Y(_23168_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32444_ ( .A({ _saxi_register_10[27], _08822_, _04091_, _08823_ }), .Y(_08828_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32445_ ( .A({ _08829_, _04250_, _08824_ }), .Y(_23167_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32446_ ( .A({ _saxi_register_10[26], _08822_, _04090_, _08823_ }), .Y(_08829_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32447_ ( .A({ _08830_, _04249_, _08824_ }), .Y(_23166_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32448_ ( .A({ _saxi_register_10[25], _08822_, _04089_, _08823_ }), .Y(_08830_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32449_ ( .A({ _08831_, _04088_, _08823_ }), .Y(_23165_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32450_ ( .A({ _saxi_register_10[24], _08822_, _04248_, _08824_ }), .Y(_08831_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32451_ ( .A({ _08832_, _04087_, _08823_ }), .Y(_23164_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32452_ ( .A({ _saxi_register_10[23], _08822_, _04247_, _08824_ }), .Y(_08832_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32453_ ( .A({ _08833_, _04086_, _08823_ }), .Y(_23163_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32454_ ( .A({ _saxi_register_10[22], _08822_, _04246_, _08824_ }), .Y(_08833_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32455_ ( .A({ _08834_, _04245_, _08824_ }), .Y(_23162_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32456_ ( .A({ _saxi_register_10[21], _08822_, _04085_, _08823_ }), .Y(_08834_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32457_ ( .A({ _08835_, _04244_, _08824_ }), .Y(_23161_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32458_ ( .A({ _saxi_register_10[20], _08822_, _04084_, _08823_ }), .Y(_08835_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32459_ ( .A({ _08836_, _04242_, _08824_ }), .Y(_23159_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32460_ ( .A({ _saxi_register_10[19], _08822_, _04082_, _08823_ }), .Y(_08836_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32461_ ( .A({ _08837_, _04241_, _08824_ }), .Y(_23158_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32462_ ( .A({ _saxi_register_10[18], _08822_, _04081_, _08823_ }), .Y(_08837_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32463_ ( .A({ _08838_, _04080_, _08823_ }), .Y(_23157_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32464_ ( .A({ _saxi_register_10[17], _08822_, _04240_, _08824_ }), .Y(_08838_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32465_ ( .A({ _08839_, _04239_, _08824_ }), .Y(_23156_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32466_ ( .A({ _saxi_register_10[16], _08822_, _04079_, _08823_ }), .Y(_08839_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32467_ ( .A({ _08840_, _04238_, _08824_ }), .Y(_23155_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32468_ ( .A({ _saxi_register_10[15], _08822_, _04078_, _08823_ }), .Y(_08840_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32469_ ( .A({ _08841_, _04237_, _08824_ }), .Y(_23154_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32470_ ( .A({ _saxi_register_10[14], _08822_, _04077_, _08823_ }), .Y(_08841_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32471_ ( .A({ _08842_, _04236_, _08824_ }), .Y(_23153_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32472_ ( .A({ _saxi_register_10[13], _08822_, _04076_, _08823_ }), .Y(_08842_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32473_ ( .A({ _08843_, _04235_, _08824_ }), .Y(_23152_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32474_ ( .A({ _saxi_register_10[12], _08822_, _04075_, _08823_ }), .Y(_08843_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32475_ ( .A({ _08844_, _04234_, _08824_ }), .Y(_23151_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32476_ ( .A({ _saxi_register_10[11], _08822_, _04074_, _08823_ }), .Y(_08844_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32477_ ( .A({ _08845_, _04233_, _08824_ }), .Y(_23150_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32478_ ( .A({ _saxi_register_10[10], _08822_, _04073_, _08823_ }), .Y(_08845_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32479_ ( .A({ _08846_, _04263_, _08824_ }), .Y(_23180_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32480_ ( .A({ _saxi_register_10[9], _08822_, _04103_, _08823_ }), .Y(_08846_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32481_ ( .A({ _08847_, _04102_, _08823_ }), .Y(_23179_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32482_ ( .A({ _saxi_register_10[8], _08822_, _04262_, _08824_ }), .Y(_08847_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32483_ ( .A({ _08848_, _04101_, _08823_ }), .Y(_23178_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32484_ ( .A({ _saxi_register_10[7], _08822_, _04261_, _08824_ }), .Y(_08848_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32485_ ( .A({ _08849_, _04260_, _08824_ }), .Y(_23177_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32486_ ( .A({ _saxi_register_10[6], _08822_, _04100_, _08823_ }), .Y(_08849_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32487_ ( .A({ _08850_, _04259_, _08824_ }), .Y(_23176_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32488_ ( .A({ _saxi_register_10[5], _08822_, _04099_, _08823_ }), .Y(_08850_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32489_ ( .A({ _08851_, _04258_, _08824_ }), .Y(_23175_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32490_ ( .A({ _saxi_register_10[4], _08822_, _04098_, _08823_ }), .Y(_08851_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32491_ ( .A({ _08852_, _04257_, _08824_ }), .Y(_23174_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32492_ ( .A({ _saxi_register_10[3], _08822_, _04097_, _08823_ }), .Y(_08852_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32493_ ( .A({ _08853_, _04094_, _08823_ }), .Y(_23171_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32494_ ( .A({ _saxi_register_10[2], _08822_, _04254_, _08824_ }), .Y(_08853_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32495_ ( .A({ _08854_, _04083_, _08823_ }), .Y(_23160_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32496_ ( .A({ _saxi_register_10[1], _08822_, _04243_, _08824_ }), .Y(_08854_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32497_ ( .A({ _08855_, _04232_, _08824_ }), .Y(_23149_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32498_ ( .A({ _saxi_register_10[0], _08822_, _04072_, _08823_ }), .Y(_08855_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _32499_ ( .A({ _08823_, _08824_, _08822_ }), .Y(_24088_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32500_ ( .A({ _05929_, _13753_, _13755_ }), .Y(_13754_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32501_ ( .A({ _05920_, _08856_ }), .Y(_24036_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32502_ ( .A({ _08862_, _08857_ }), .Y(_08856_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32503_ ( .A({ matmul_29_comp_fsm[2], _08858_, matmul_29_comp_fsm[3] }), .Y(_08857_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32504_ ( .A({ _08861_, _08860_, _08859_ }), .Y(_08858_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32505_ ( .A(matmul_29_comp_fsm[15:12]), .Y(_08859_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32506_ ( .A(matmul_29_comp_fsm[7:4]), .Y(_08860_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32507_ ( .A(matmul_29_comp_fsm[11:8]), .Y(_08861_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32508_ ( .A({ matmul_29_comp_fsm[1], _08863_, matmul_29_comp_fsm[0] }), .Y(_08862_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32509_ ( .A({ _08867_, _08866_, _08865_, _08864_ }), .Y(_08863_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32510_ ( .A(matmul_29_comp_fsm[23:20]), .Y(_08864_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32511_ ( .A(matmul_29_comp_fsm[19:16]), .Y(_08865_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32512_ ( .A(matmul_29_comp_fsm[31:28]), .Y(_08866_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32513_ ( .A(matmul_29_comp_fsm[27:24]), .Y(_08867_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _32514_ ( .A({ _08868_, _08869_, matmul_29_comp_fsm[1] }), .Y(_05920_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32515_ ( .A({ matmul_29_comp_fsm[0], _08863_ }), .Y(_08868_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _32516_ ( .A({ _08858_, matmul_29_comp_fsm[2], matmul_29_comp_fsm[3] }), .Y(_08869_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32517_ ( .A({ _08873_, _08870_ }), .Y(_24035_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _32518_ ( .A({ _05917_, _05725_, _08872_, _08856_ }), .Y(_08870_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32519_ ( .A({ matmul_29_comp_fsm[1], _08869_, _08868_ }), .Y(_05917_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32520_ ( .A({ _08871_, _08869_ }), .Y(_05725_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _32521_ ( .A({ _08863_, matmul_29_comp_fsm[1:0] }), .Y(_08871_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32522_ ( .A({ _08871_, _08857_ }), .Y(_08872_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32523_ ( .A({ _05916_, _05920_, _08874_ }), .Y(_08873_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32524_ ( .A({ _08857_, _08868_, matmul_29_comp_fsm[1] }), .Y(_08874_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32525_ ( .A({ _08869_, _08862_ }), .Y(_05916_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _32526_ ( .A({ _08875_, _05917_, _08874_ }), .Y(_13679_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32527_ ( .A({ _13743_, _05725_, _08872_, _13711_ }), .Y(_08875_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _32528_ ( .A({ _08876_, _13689_, _08872_ }), .Y(_13657_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _32529_ ( .A({ _05916_, _05725_, _13721_ }), .Y(_08876_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _32530_ ( .A({ _08877_, _08873_ }), .Y(_13668_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32531_ ( .A({ _13732_, _05725_, _08872_, _13700_ }), .Y(_08877_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32532_ ( .A({ _13746_, _05725_, _08872_, _13714_ }), .Y(_13682_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32533_ ( .A({ _13749_, _05725_, _08872_, _13717_ }), .Y(_13685_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32534_ ( .A({ _13751_, _05725_, _08872_, _13719_ }), .Y(_13687_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32535_ ( .A({ _13747_, _05725_, _08872_, _13715_ }), .Y(_13683_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32536_ ( .A({ _13748_, _05725_, _08872_, _13716_ }), .Y(_13684_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32537_ ( .A({ _13750_, _05725_, _08872_, _13718_ }), .Y(_13686_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32538_ ( .A({ _13722_, _05725_, _08872_, _13690_ }), .Y(_13658_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32539_ ( .A({ _13727_, _05725_, _08872_, _13695_ }), .Y(_13663_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32540_ ( .A({ _13752_, _05725_, _08872_, _13720_ }), .Y(_13688_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32541_ ( .A({ _13723_, _05725_, _08872_, _13691_ }), .Y(_13659_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32542_ ( .A({ _13724_, _05725_, _08872_, _13692_ }), .Y(_13660_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32543_ ( .A({ _13728_, _05725_, _08872_, _13696_ }), .Y(_13664_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32544_ ( .A({ _13725_, _05725_, _08872_, _13693_ }), .Y(_13661_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32545_ ( .A({ _13726_, _05725_, _08872_, _13694_ }), .Y(_13662_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32546_ ( .A({ _13731_, _05725_, _08872_, _13699_ }), .Y(_13667_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32547_ ( .A({ _13729_, _05725_, _08872_, _13697_ }), .Y(_13665_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32548_ ( .A({ _13734_, _05725_, _08872_, _13702_ }), .Y(_13670_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32549_ ( .A({ _13730_, _05725_, _08872_, _13698_ }), .Y(_13666_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32550_ ( .A({ _13733_, _05725_, _08872_, _13701_ }), .Y(_13669_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32551_ ( .A({ _13737_, _05725_, _08872_, _13705_ }), .Y(_13673_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32552_ ( .A({ _13735_, _05725_, _08872_, _13703_ }), .Y(_13671_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32553_ ( .A({ _13739_, _05725_, _08872_, _13707_ }), .Y(_13675_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32554_ ( .A({ _13736_, _05725_, _08872_, _13704_ }), .Y(_13672_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32555_ ( .A({ _13738_, _05725_, _08872_, _13706_ }), .Y(_13674_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32556_ ( .A({ _13742_, _05725_, _08872_, _13710_ }), .Y(_13678_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32557_ ( .A({ _13744_, _05725_, _08872_, _13712_ }), .Y(_13680_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32558_ ( .A({ _13740_, _05725_, _08872_, _13708_ }), .Y(_13676_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32559_ ( .A({ _13741_, _05725_, _08872_, _13709_ }), .Y(_13677_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _32560_ ( .A({ _13745_, _05725_, _08872_, _13713_ }), .Y(_13681_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _32561_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18343_, _18375_ }), .Y(_18311_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32562_ ( .A({ _08879_, _08887_, _stream_conv2d_16_source_26_source_pat_fsm_9[1] }), .Y(_08878_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32563_ ( .A({ _08886_, _08885_, _08880_ }), .Y(_08879_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32564_ ( .A({ _08884_, _08883_, _08882_, _08881_ }), .Y(_08880_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32565_ ( .A(_stream_conv2d_16_source_26_source_pat_fsm_9[23:20]), .Y(_08881_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32566_ ( .A(_stream_conv2d_16_source_26_source_pat_fsm_9[19:16]), .Y(_08882_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32567_ ( .A(_stream_conv2d_16_source_26_source_pat_fsm_9[31:28]), .Y(_08883_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32568_ ( .A(_stream_conv2d_16_source_26_source_pat_fsm_9[27:24]), .Y(_08884_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32569_ ( .A(_stream_conv2d_16_source_26_source_pat_fsm_9[15:12]), .Y(_08885_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32570_ ( .A(_stream_conv2d_16_source_26_source_pat_fsm_9[11:8]), .Y(_08886_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _32571_ ( .A({ _08888_, _stream_conv2d_16_source_26_source_pat_fsm_9[3:2] }), .Y(_08887_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32572_ ( .A(_stream_conv2d_16_source_26_source_pat_fsm_9[7:4]), .Y(_08888_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _32573_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18342_, _18374_ }), .Y(_18310_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _32574_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18338_, _18370_ }), .Y(_18306_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _32575_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18337_, _18369_ }), .Y(_18305_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _32576_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18336_, _18368_ }), .Y(_18304_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _32577_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18335_, _18367_ }), .Y(_18303_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _32578_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18334_, _18366_ }), .Y(_18302_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _32579_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18333_, _18365_ }), .Y(_18301_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _32580_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18332_, _18364_ }), .Y(_18300_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _32581_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18331_, _18363_ }), .Y(_18299_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32582_ ( .A({ _08901_, _08898_, _08889_ }), .Y(_23205_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32583_ ( .A({ _08896_, _08893_, _08890_ }), .Y(_08889_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32584_ ( .A({ _23269_, _08891_, _08892_, _23493_ }), .Y(_08890_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _32585_ ( .A({ _06887_, _06909_, _06891_, main_fsm[4] }), .Y(_08891_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32586_ ( .A({ _06904_, _06912_, _06891_ }), .Y(_08892_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32587_ ( .A({ _23365_, _08894_, _08895_, _23461_ }), .Y(_08893_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _32588_ ( .A({ _06891_, _06907_, _06898_, main_fsm[4] }), .Y(_08894_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32589_ ( .A({ main_fsm[4], _06902_, _06906_, _06891_ }), .Y(_08895_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32590_ ( .A({ _23525_, _05684_, _23397_, _08897_ }), .Y(_08896_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32591_ ( .A({ _06897_, _06912_, _06891_ }), .Y(_05684_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _32592_ ( .A({ _06891_, _06910_, _06898_, main_fsm[4] }), .Y(_08897_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32593_ ( .A({ _23301_, _08899_, _23237_, _08900_ }), .Y(_08898_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _32594_ ( .A({ _06887_, _06911_, _06891_, main_fsm[4] }), .Y(_08899_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32595_ ( .A({ main_fsm[4], _06905_, _06891_, _06887_ }), .Y(_08900_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32596_ ( .A({ _23333_, _08902_, _23429_, _08903_ }), .Y(_08901_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32597_ ( .A({ main_fsm[4], _06905_, _06898_, _06891_ }), .Y(_08902_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32598_ ( .A({ main_fsm[4], _06914_, _06906_, _06891_ }), .Y(_08903_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32599_ ( .A({ _08909_, _08908_, _08904_ }), .Y(_23204_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32600_ ( .A({ _08907_, _08906_, _08905_ }), .Y(_08904_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32601_ ( .A({ _23492_, _08892_, _23460_, _08895_ }), .Y(_08905_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32602_ ( .A({ _23236_, _08900_, _08897_, _23396_ }), .Y(_08906_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32603_ ( .A({ _23428_, _08903_, _08891_, _23268_ }), .Y(_08907_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32604_ ( .A({ _23332_, _08902_, _08894_, _23364_ }), .Y(_08908_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32605_ ( .A({ _23300_, _08899_, _23524_, _05684_ }), .Y(_08909_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32606_ ( .A({ _08915_, _08914_, _08910_ }), .Y(_23200_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32607_ ( .A({ _08913_, _08912_, _08911_ }), .Y(_08910_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32608_ ( .A({ _23232_, _08900_, _08892_, _23488_ }), .Y(_08911_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32609_ ( .A({ _23296_, _08899_, _08895_, _23456_ }), .Y(_08912_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32610_ ( .A({ _23328_, _08902_, _23264_, _08891_ }), .Y(_08913_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32611_ ( .A({ _23520_, _05684_, _23392_, _08897_ }), .Y(_08914_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32612_ ( .A({ _23424_, _08903_, _08894_, _23360_ }), .Y(_08915_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32613_ ( .A({ _08921_, _08920_, _08916_ }), .Y(_23201_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32614_ ( .A({ _08919_, _08918_, _08917_ }), .Y(_08916_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32615_ ( .A({ _23425_, _08903_, _08891_, _23265_ }), .Y(_08917_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32616_ ( .A({ _23297_, _08899_, _08897_, _23393_ }), .Y(_08918_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32617_ ( .A({ _23233_, _08900_, _08894_, _23361_ }), .Y(_08919_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32618_ ( .A({ _23329_, _08902_, _23521_, _05684_ }), .Y(_08920_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32619_ ( .A({ _23489_, _08892_, _23457_, _08895_ }), .Y(_08921_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32620_ ( .A({ _08927_, _08926_, _08922_ }), .Y(_23202_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32621_ ( .A({ _08925_, _08924_, _08923_ }), .Y(_08922_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32622_ ( .A({ _23490_, _08892_, _23458_, _08895_ }), .Y(_08923_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32623_ ( .A({ _23234_, _08900_, _08897_, _23394_ }), .Y(_08924_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32624_ ( .A({ _23426_, _08903_, _08891_, _23266_ }), .Y(_08925_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32625_ ( .A({ _23330_, _08902_, _08894_, _23362_ }), .Y(_08926_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32626_ ( .A({ _23298_, _08899_, _23522_, _05684_ }), .Y(_08927_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32627_ ( .A({ _08933_, _08932_, _08928_ }), .Y(_23198_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32628_ ( .A({ _08931_, _08930_, _08929_ }), .Y(_08928_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32629_ ( .A({ _23230_, _08900_, _08897_, _23390_ }), .Y(_08929_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32630_ ( .A({ _23294_, _08899_, _23518_, _05684_ }), .Y(_08930_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32631_ ( .A({ _23262_, _08891_, _08894_, _23358_ }), .Y(_08931_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32632_ ( .A({ _23326_, _08902_, _08895_, _23454_ }), .Y(_08932_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32633_ ( .A({ _23422_, _08903_, _08892_, _23486_ }), .Y(_08933_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32634_ ( .A({ _08939_, _08938_, _08934_ }), .Y(_23199_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32635_ ( .A({ _08937_, _08936_, _08935_ }), .Y(_08934_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32636_ ( .A({ _23263_, _08891_, _08892_, _23487_ }), .Y(_08935_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32637_ ( .A({ _23359_, _08894_, _08895_, _23455_ }), .Y(_08936_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32638_ ( .A({ _23519_, _05684_, _23391_, _08897_ }), .Y(_08937_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32639_ ( .A({ _23295_, _08899_, _23231_, _08900_ }), .Y(_08938_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32640_ ( .A({ _23327_, _08902_, _23423_, _08903_ }), .Y(_08939_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32641_ ( .A({ _08945_, _08944_, _08940_ }), .Y(_23197_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32642_ ( .A({ _08943_, _08942_, _08941_ }), .Y(_08940_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32643_ ( .A({ _23261_, _08891_, _08892_, _23485_ }), .Y(_08941_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32644_ ( .A({ _23293_, _08899_, _23229_, _08900_ }), .Y(_08942_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32645_ ( .A({ _23453_, _08895_, _23517_, _05684_ }), .Y(_08943_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32646_ ( .A({ _23357_, _08894_, _08897_, _23389_ }), .Y(_08944_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32647_ ( .A({ _23325_, _08902_, _23421_, _08903_ }), .Y(_08945_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32648_ ( .A({ _08951_, _08950_, _08946_ }), .Y(_23195_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32649_ ( .A({ _08949_, _08948_, _08947_ }), .Y(_08946_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32650_ ( .A({ _23259_, _08891_, _08892_, _23483_ }), .Y(_08947_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32651_ ( .A({ _23355_, _08894_, _08895_, _23451_ }), .Y(_08948_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32652_ ( .A({ _23515_, _05684_, _23387_, _08897_ }), .Y(_08949_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32653_ ( .A({ _23291_, _08899_, _23227_, _08900_ }), .Y(_08950_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32654_ ( .A({ _23323_, _08902_, _23419_, _08903_ }), .Y(_08951_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32655_ ( .A({ _08957_, _08956_, _08952_ }), .Y(_23196_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32656_ ( .A({ _08955_, _08954_, _08953_ }), .Y(_08952_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32657_ ( .A({ _23260_, _08891_, _08892_, _23484_ }), .Y(_08953_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32658_ ( .A({ _23452_, _08895_, _23516_, _05684_ }), .Y(_08954_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32659_ ( .A({ _23420_, _08903_, _08894_, _23356_ }), .Y(_08955_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32660_ ( .A({ _23292_, _08899_, _23228_, _08900_ }), .Y(_08956_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32661_ ( .A({ _23324_, _08902_, _08897_, _23388_ }), .Y(_08957_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32662_ ( .A({ _08963_, _08962_, _08958_ }), .Y(_23190_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32663_ ( .A({ _08961_, _08960_, _08959_ }), .Y(_08958_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32664_ ( .A({ _23222_, _08900_, _08892_, _23478_ }), .Y(_08959_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32665_ ( .A({ _23286_, _08899_, _08895_, _23446_ }), .Y(_08960_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32666_ ( .A({ _23318_, _08902_, _23254_, _08891_ }), .Y(_08961_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32667_ ( .A({ _23510_, _05684_, _23382_, _08897_ }), .Y(_08962_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32668_ ( .A({ _23414_, _08903_, _08894_, _23350_ }), .Y(_08963_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32669_ ( .A({ _08969_, _08968_, _08964_ }), .Y(_23191_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32670_ ( .A({ _08967_, _08966_, _08965_ }), .Y(_08964_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32671_ ( .A({ _23223_, _08900_, _23415_, _08903_ }), .Y(_08965_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32672_ ( .A({ _23287_, _08899_, _08897_, _23383_ }), .Y(_08966_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32673_ ( .A({ _23255_, _08891_, _08892_, _23479_ }), .Y(_08967_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32674_ ( .A({ _23319_, _08902_, _08895_, _23447_ }), .Y(_08968_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32675_ ( .A({ _23351_, _08894_, _23511_, _05684_ }), .Y(_08969_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32676_ ( .A({ _08975_, _08974_, _08970_ }), .Y(_23185_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32677_ ( .A({ _08973_, _08972_, _08971_ }), .Y(_08970_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32678_ ( .A({ _23473_, _08892_, _23441_, _08895_ }), .Y(_08971_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32679_ ( .A({ _23217_, _08900_, _08897_, _23377_ }), .Y(_08972_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32680_ ( .A({ _23409_, _08903_, _08891_, _23249_ }), .Y(_08973_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32681_ ( .A({ _23313_, _08902_, _08894_, _23345_ }), .Y(_08974_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32682_ ( .A({ _23281_, _08899_, _23505_, _05684_ }), .Y(_08975_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32683_ ( .A({ _08981_, _08980_, _08976_ }), .Y(_23188_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32684_ ( .A({ _08979_, _08978_, _08977_ }), .Y(_08976_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32685_ ( .A({ _23252_, _08891_, _08892_, _23476_ }), .Y(_08977_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32686_ ( .A({ _23444_, _08895_, _23508_, _05684_ }), .Y(_08978_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32687_ ( .A({ _23412_, _08903_, _08894_, _23348_ }), .Y(_08979_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32688_ ( .A({ _23284_, _08899_, _23220_, _08900_ }), .Y(_08980_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32689_ ( .A({ _23316_, _08902_, _08897_, _23380_ }), .Y(_08981_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32690_ ( .A({ _08987_, _08986_, _08982_ }), .Y(_23193_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32691_ ( .A({ _08985_, _08984_, _08983_ }), .Y(_08982_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32692_ ( .A({ _23225_, _08900_, _08891_, _23257_ }), .Y(_08983_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32693_ ( .A({ _23289_, _08899_, _08894_, _23353_ }), .Y(_08984_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32694_ ( .A({ _23417_, _08903_, _08892_, _23481_ }), .Y(_08985_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32695_ ( .A({ _23449_, _08895_, _23513_, _05684_ }), .Y(_08986_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32696_ ( .A({ _23321_, _08902_, _08897_, _23385_ }), .Y(_08987_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32697_ ( .A({ _08993_, _08992_, _08988_ }), .Y(_23186_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32698_ ( .A({ _08991_, _08990_, _08989_ }), .Y(_08988_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32699_ ( .A({ _23474_, _08892_, _23442_, _08895_ }), .Y(_08989_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32700_ ( .A({ _23218_, _08900_, _08897_, _23378_ }), .Y(_08990_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32701_ ( .A({ _23410_, _08903_, _08891_, _23250_ }), .Y(_08991_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32702_ ( .A({ _23314_, _08902_, _08894_, _23346_ }), .Y(_08992_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32703_ ( .A({ _23282_, _08899_, _23506_, _05684_ }), .Y(_08993_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32704_ ( .A({ _08999_, _08998_, _08994_ }), .Y(_23194_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32705_ ( .A({ _08997_, _08996_, _08995_ }), .Y(_08994_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32706_ ( .A({ _23258_, _08891_, _08892_, _23482_ }), .Y(_08995_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32707_ ( .A({ _23354_, _08894_, _08895_, _23450_ }), .Y(_08996_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32708_ ( .A({ _23514_, _05684_, _23386_, _08897_ }), .Y(_08997_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32709_ ( .A({ _23290_, _08899_, _23226_, _08900_ }), .Y(_08998_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32710_ ( .A({ _23322_, _08902_, _23418_, _08903_ }), .Y(_08999_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32711_ ( .A({ _09005_, _09004_, _09000_ }), .Y(_23189_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32712_ ( .A({ _09003_, _09002_, _09001_ }), .Y(_09000_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32713_ ( .A({ _23253_, _08891_, _08892_, _23477_ }), .Y(_09001_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32714_ ( .A({ _23285_, _08899_, _23221_, _08900_ }), .Y(_09002_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32715_ ( .A({ _23445_, _08895_, _23509_, _05684_ }), .Y(_09003_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32716_ ( .A({ _23349_, _08894_, _08897_, _23381_ }), .Y(_09004_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32717_ ( .A({ _23317_, _08902_, _23413_, _08903_ }), .Y(_09005_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32718_ ( .A({ _09011_, _09010_, _09006_ }), .Y(_23187_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32719_ ( .A({ _09009_, _09008_, _09007_ }), .Y(_09006_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32720_ ( .A({ _23315_, _08902_, _08894_, _23347_ }), .Y(_09007_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32721_ ( .A({ _23219_, _08900_, _08895_, _23443_ }), .Y(_09008_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32722_ ( .A({ _23251_, _08891_, _23507_, _05684_ }), .Y(_09009_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32723_ ( .A({ _23283_, _08899_, _23411_, _08903_ }), .Y(_09010_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32724_ ( .A({ _23475_, _08892_, _23379_, _08897_ }), .Y(_09011_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32725_ ( .A({ _09017_, _09016_, _09012_ }), .Y(_23182_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32726_ ( .A({ _09015_, _09014_, _09013_ }), .Y(_09012_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32727_ ( .A({ _23246_, _08891_, _08892_, _23470_ }), .Y(_09013_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32728_ ( .A({ _23342_, _08894_, _08895_, _23438_ }), .Y(_09014_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32729_ ( .A({ _23502_, _05684_, _23374_, _08897_ }), .Y(_09015_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32730_ ( .A({ _23278_, _08899_, _23214_, _08900_ }), .Y(_09016_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32731_ ( .A({ _23310_, _08902_, _23406_, _08903_ }), .Y(_09017_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32732_ ( .A({ _09023_, _09022_, _09018_ }), .Y(_23184_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32733_ ( .A({ _09021_, _09020_, _09019_ }), .Y(_09018_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32734_ ( .A({ _23248_, _08891_, _08892_, _23472_ }), .Y(_09019_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32735_ ( .A({ _23344_, _08894_, _08895_, _23440_ }), .Y(_09020_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32736_ ( .A({ _23504_, _05684_, _23376_, _08897_ }), .Y(_09021_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32737_ ( .A({ _23280_, _08899_, _23216_, _08900_ }), .Y(_09022_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32738_ ( .A({ _23312_, _08902_, _23408_, _08903_ }), .Y(_09023_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32739_ ( .A({ _09029_, _09028_, _09024_ }), .Y(_23183_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32740_ ( .A({ _09027_, _09026_, _09025_ }), .Y(_09024_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32741_ ( .A({ _23407_, _08903_, _08891_, _23247_ }), .Y(_09025_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32742_ ( .A({ _23503_, _05684_, _23375_, _08897_ }), .Y(_09026_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32743_ ( .A({ _23471_, _08892_, _23439_, _08895_ }), .Y(_09027_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32744_ ( .A({ _23279_, _08899_, _08902_, _23311_ }), .Y(_09028_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32745_ ( .A({ _23215_, _08900_, _08894_, _23343_ }), .Y(_09029_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32746_ ( .A({ _09035_, _09034_, _09030_ }), .Y(_23211_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32747_ ( .A({ _09033_, _09032_, _09031_ }), .Y(_09030_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32748_ ( .A({ _23275_, _08891_, _08892_, _23499_ }), .Y(_09031_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32749_ ( .A({ _23371_, _08894_, _08895_, _23467_ }), .Y(_09032_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32750_ ( .A({ _23531_, _05684_, _23403_, _08897_ }), .Y(_09033_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32751_ ( .A({ _23307_, _08899_, _23243_, _08900_ }), .Y(_09034_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32752_ ( .A({ _23339_, _08902_, _23435_, _08903_ }), .Y(_09035_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _32753_ ( .A({ _09056_, _09053_, _09045_, _09036_ }), .Y(_23209_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32754_ ( .A({ _09042_, _09040_, _09037_ }), .Y(_09036_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _32755_ ( .A({ _09038_, _08902_, _23337_ }), .Y(_09037_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32756_ ( .A({ _06917_, _06886_, _09039_, _06910_ }), .Y(_09038_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32757_ ( .A({ main_fsm[4], _06891_, _06887_ }), .Y(_09039_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _32758_ ( .A({ _09041_, _08891_, _23273_ }), .Y(_09040_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32759_ ( .A({ _06897_, _06886_, _06907_, _06901_ }), .Y(_09041_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _32760_ ( .A({ _09044_, _09043_, _08897_, _23401_ }), .Y(_09042_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32761_ ( .A({ _23305_, _08899_, _08892_, _23497_ }), .Y(_09043_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _32762_ ( .A({ _09039_, _07451_, _06900_ }), .Y(_09044_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _32763_ ( .A({ _09050_, _09046_, _08895_, _23465_ }), .Y(_09045_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32764_ ( .A({ _09049_, _09048_, _09047_ }), .Y(_09046_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _32765_ ( .A({ _08577_, _06886_, _06904_ }), .Y(_09047_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _32766_ ( .A({ _09039_, _06902_, _06896_ }), .Y(_09048_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32767_ ( .A({ _08541_, _08508_, _08474_, _07453_ }), .Y(_09049_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _32768_ ( .A({ _09051_, _08894_, _23369_ }), .Y(_09050_) );
  \$lut  #( .LUT(8'h4f), .WIDTH(3) ) _32769_ ( .A({ _09039_, _09052_, _06916_ }), .Y(_09051_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32770_ ( .A({ _08682_, _08576_ }), .Y(_09052_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32771_ ( .A({ _09055_, _09054_ }), .Y(_09053_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32772_ ( .A({ _06916_, _06886_, _23433_, _08903_ }), .Y(_09054_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32773_ ( .A({ _23241_, _08900_, _23529_, _05684_ }), .Y(_09055_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _32774_ ( .A({ _09058_, _09057_, _08539_, _08507_ }), .Y(_09056_) );
  \$lut  #( .LUT(16'h004f), .WIDTH(4) ) _32775_ ( .A({ _08578_, _06886_, _09052_, _06896_ }), .Y(_09057_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32776_ ( .A({ _08472_, _07450_ }), .Y(_09058_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32777_ ( .A({ _09064_, _09063_, _09059_ }), .Y(_23212_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32778_ ( .A({ _09062_, _09061_, _09060_ }), .Y(_09059_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32779_ ( .A({ _23276_, _08891_, _08892_, _23500_ }), .Y(_09060_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32780_ ( .A({ _23372_, _08894_, _08895_, _23468_ }), .Y(_09061_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32781_ ( .A({ _23532_, _05684_, _23404_, _08897_ }), .Y(_09062_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32782_ ( .A({ _23308_, _08899_, _23244_, _08900_ }), .Y(_09063_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32783_ ( .A({ _23340_, _08902_, _23436_, _08903_ }), .Y(_09064_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32784_ ( .A({ _09070_, _09069_, _09065_ }), .Y(_23210_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32785_ ( .A({ _09068_, _09067_, _09066_ }), .Y(_09065_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32786_ ( .A({ _23434_, _08903_, _08891_, _23274_ }), .Y(_09066_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32787_ ( .A({ _23306_, _08899_, _08897_, _23402_ }), .Y(_09067_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32788_ ( .A({ _23242_, _08900_, _08894_, _23370_ }), .Y(_09068_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32789_ ( .A({ _23338_, _08902_, _23530_, _05684_ }), .Y(_09069_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32790_ ( .A({ _23498_, _08892_, _23466_, _08895_ }), .Y(_09070_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _32791_ ( .A({ _09087_, _09082_, _09080_, _13067_ }), .Y(_23207_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32792_ ( .A({ _09075_, _09073_, _09072_, _09049_ }), .Y(_09071_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _32793_ ( .A({ _05732_, _09039_, _07451_, _06900_ }), .Y(_09072_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32794_ ( .A({ _05730_, _09074_, _08473_, _07452_ }), .Y(_09073_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32795_ ( .A({ main_fsm[4], _07451_, _06898_, _06891_ }), .Y(_09074_) );
  \$lut  #( .LUT(16'h001f), .WIDTH(4) ) _32796_ ( .A({ _09076_, _06908_, _06904_, _06896_ }), .Y(_09075_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32797_ ( .A({ main_fsm[4], _06910_, _06898_, _06891_ }), .Y(_09076_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _32798_ ( .A({ _08648_, _08612_, _08895_, _23463_ }), .Y(_09077_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _32799_ ( .A({ _08646_, _08611_, _08892_, _23495_ }), .Y(_09078_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _32800_ ( .A({ _06908_, _06917_, _06911_ }), .Y(_09079_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32801_ ( .A({ _09081_, _09051_ }), .Y(_09080_) );
  \$lut  #( .LUT(16'h000b), .WIDTH(4) ) _32802_ ( .A({ _08509_, _08542_, _06901_, _09052_ }), .Y(_09081_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32803_ ( .A({ _09086_, _09085_, _09084_, _09083_ }), .Y(_09082_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32804_ ( .A({ _23335_, _08902_, _23431_, _08903_ }), .Y(_09083_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32805_ ( .A({ _23239_, _08900_, _08897_, _23399_ }), .Y(_09084_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32806_ ( .A({ _23303_, _08899_, _23527_, _05684_ }), .Y(_09085_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32807_ ( .A({ _23271_, _08891_, _08894_, _23367_ }), .Y(_09086_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32808_ ( .A({ _09090_, _09089_, _09088_ }), .Y(_09087_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _32809_ ( .A({ _08823_, _06908_, _06910_ }), .Y(_09088_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _32810_ ( .A({ _06908_, _06916_, _06909_ }), .Y(_09089_) );
  \$lut  #( .LUT(16'h000b), .WIDTH(4) ) _32811_ ( .A({ _08754_, _08789_, _06908_, _09052_ }), .Y(_09090_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32812_ ( .A({ _09099_, _09098_, _09095_, _09092_ }), .Y(_09091_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _32813_ ( .A({ _09094_, _09093_, _08902_, _23320_ }), .Y(_09092_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _32814_ ( .A({ _08613_, _06903_, _06911_ }), .Y(_09093_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32815_ ( .A({ _23288_, _08899_, _23512_, _05684_ }), .Y(_09094_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _32816_ ( .A({ _09097_, _09096_, _08892_, _23480_ }), .Y(_09095_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32817_ ( .A({ _23416_, _08903_, _08895_, _23448_ }), .Y(_09096_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _32818_ ( .A({ _06915_, _08682_, _08576_ }), .Y(_09097_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32819_ ( .A({ _23224_, _08900_, _08891_, _23256_ }), .Y(_09098_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32820_ ( .A({ _23352_, _08894_, _08897_, _23384_ }), .Y(_09099_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32821_ ( .A({ _09106_, _09105_, _09103_, _09101_ }), .Y(_09100_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32822_ ( .A({ _05742_, _09102_, _05743_ }), .Y(_09101_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _32823_ ( .A({ _06915_, _06910_, _06905_ }), .Y(_09102_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32824_ ( .A({ _05740_, _05734_, _09104_ }), .Y(_09103_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _32825_ ( .A({ _06903_, _06914_, _06904_ }), .Y(_09104_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32826_ ( .A({ _08473_, _07452_, _08539_, _08507_ }), .Y(_09105_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32827_ ( .A({ _09079_, _09038_ }), .Y(_09106_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _32828_ ( .A({ _09109_, _09108_, _08474_, _07453_ }), .Y(_09107_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32829_ ( .A({ _08648_, _08612_ }), .Y(_09108_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _32830_ ( .A({ _09088_, _09076_, _06908_, _06904_ }), .Y(_09109_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32831_ ( .A({ _06911_, _06903_ }), .Y(_05646_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32832_ ( .A({ _09121_, _09118_, _09110_ }), .Y(_23208_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32833_ ( .A({ _09117_, _09116_, _09113_, _09111_ }), .Y(_09110_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _32834_ ( .A({ _09112_, _08891_, _23272_ }), .Y(_09111_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32835_ ( .A({ _23496_, _08892_, _23368_, _08894_ }), .Y(_09112_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _32836_ ( .A({ _09115_, _09114_, _05684_, _23528_ }), .Y(_09113_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32837_ ( .A({ _23240_, _08900_, _08895_, _23464_ }), .Y(_09114_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32838_ ( .A({ _05734_, _05732_ }), .Y(_09115_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32839_ ( .A({ _23304_, _08899_, _08902_, _23336_ }), .Y(_09116_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32840_ ( .A({ _23432_, _08903_, _08897_, _23400_ }), .Y(_09117_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32841_ ( .A({ _09120_, _09119_, _09093_, _09108_ }), .Y(_09118_) );
  \$lut  #( .LUT(16'h111f), .WIDTH(4) ) _32842_ ( .A({ _06903_, _06901_, _06902_, _06896_ }), .Y(_09119_) );
  \$lut  #( .LUT(16'h10ff), .WIDTH(4) ) _32843_ ( .A({ _06903_, _09052_, _06916_, _06909_ }), .Y(_09120_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32844_ ( .A({ _09123_, _09073_, _09122_ }), .Y(_09121_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _32845_ ( .A({ _09081_, _09104_, _09076_ }), .Y(_09122_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32846_ ( .A({ _05736_, _08824_, _08788_, _08647_ }), .Y(_09123_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32847_ ( .A({ _08682_, _06886_ }), .Y(_05681_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _32848_ ( .A({ _09138_, _09127_, _09124_ }), .Y(_23206_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32849_ ( .A({ _09090_, _09089_, _09125_, _09080_ }), .Y(_09124_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _32850_ ( .A({ _09126_, _09097_, _08753_, _08717_ }), .Y(_09125_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _32851_ ( .A({ _06915_, _06916_, _06909_ }), .Y(_09126_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32852_ ( .A({ _09135_, _09133_, _09131_, _09128_ }), .Y(_09127_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32853_ ( .A({ _09130_, _09129_ }), .Y(_09128_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32854_ ( .A({ _23238_, _08900_, _08902_, _23334_ }), .Y(_09129_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32855_ ( .A({ _23430_, _08903_, _08895_, _23462_ }), .Y(_09130_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32856_ ( .A({ _09132_, _09104_, _09047_, _09058_ }), .Y(_09131_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _32857_ ( .A({ _08824_, _08788_ }), .Y(_09132_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _32858_ ( .A({ _09134_, _08891_, _23270_ }), .Y(_09133_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32859_ ( .A({ _23302_, _08899_, _08897_, _23398_ }), .Y(_09134_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _32860_ ( .A({ _09137_, _09136_, _05684_, _23526_ }), .Y(_09135_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32861_ ( .A({ _23494_, _08892_, _23366_, _08894_ }), .Y(_09136_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _32862_ ( .A({ _05740_, _06886_, _06916_ }), .Y(_09137_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32863_ ( .A({ _09139_, _09120_, _09073_, _09044_ }), .Y(_09138_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _32864_ ( .A({ _06886_, _09052_, _06904_, _06908_ }), .Y(_09139_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32865_ ( .A({ _06909_, _06903_ }), .Y(_05645_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _32866_ ( .A({ _09152_, _13073_, _09143_, _09140_ }), .Y(_23181_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _32867_ ( .A({ _09115_, _09141_, _08894_, _23341_ }), .Y(_09140_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _32868_ ( .A({ _09142_, _08903_, _23405_ }), .Y(_09141_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32869_ ( .A({ _06909_, _06903_, _08576_, _06915_ }), .Y(_09142_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32870_ ( .A({ _09145_, _09144_ }), .Y(_09143_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32871_ ( .A({ _08508_, _08612_, _08611_, _08507_ }), .Y(_09144_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32872_ ( .A({ _08788_, _08787_, _08717_, _08719_ }), .Y(_09145_) );
  \$lut  #( .LUT(16'h1fff), .WIDTH(4) ) _32873_ ( .A({ _06912_, _06891_, _06902_, _06909_ }), .Y(_09146_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32874_ ( .A({ _09149_, _09148_, _05737_, _05731_ }), .Y(_09147_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _32875_ ( .A({ _05739_, _05742_, _05740_, _08509_ }), .Y(_09148_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _32876_ ( .A({ _09150_, _06886_, _06897_ }), .Y(_09149_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32877_ ( .A({ _08576_, _06891_, _06887_ }), .Y(_09150_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32878_ ( .A({ _08823_, _08754_, _08647_, _08684_ }), .Y(_09151_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32879_ ( .A({ _09156_, _09155_, _09154_, _09153_ }), .Y(_09152_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32880_ ( .A({ _23309_, _08902_, _08892_, _23469_ }), .Y(_09153_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32881_ ( .A({ _23245_, _08891_, _23501_, _05684_ }), .Y(_09154_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32882_ ( .A({ _23277_, _08899_, _08897_, _23373_ }), .Y(_09155_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32883_ ( .A({ _23213_, _08900_, _08895_, _23437_ }), .Y(_09156_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32884_ ( .A({ _06896_, _09039_ }), .Y(_05680_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32885_ ( .A({ _06896_, _06901_ }), .Y(_05682_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32886_ ( .A({ _06916_, _06908_ }), .Y(_05683_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _32887_ ( .A({ _09167_, _09163_, _09162_, _09157_ }), .Y(_23203_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32888_ ( .A({ _09089_, _09088_, _09161_, _09158_ }), .Y(_09157_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _32889_ ( .A({ _09159_, _09126_, _08894_, _23363_ }), .Y(_09158_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _32890_ ( .A({ _09160_, _08891_, _23267_ }), .Y(_09159_) );
  \$lut  #( .LUT(16'h1fff), .WIDTH(4) ) _32891_ ( .A({ _06912_, _06891_, _06896_, _06902_ }), .Y(_09160_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _32892_ ( .A({ _09102_, _05645_, _08683_ }), .Y(_09161_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32893_ ( .A({ _09119_, _09105_, _09103_ }), .Y(_09162_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32894_ ( .A({ _09075_, _09048_, _09047_, _09164_ }), .Y(_09163_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _32895_ ( .A({ _09166_, _09165_, _08542_, _08509_ }), .Y(_09164_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _32896_ ( .A({ _08578_, _06886_, _06896_ }), .Y(_09165_) );
  \$lut  #( .LUT(16'h035f), .WIDTH(4) ) _32897_ ( .A({ _06916_, _09039_, _06886_, _06910_ }), .Y(_09166_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32898_ ( .A({ _09171_, _09170_, _09169_, _09168_ }), .Y(_09167_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32899_ ( .A({ _23491_, _08892_, _23459_, _08895_ }), .Y(_09168_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32900_ ( .A({ _23299_, _08899_, _08902_, _23331_ }), .Y(_09169_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _32901_ ( .A({ _23427_, _08903_, _08897_, _23395_ }), .Y(_09170_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _32902_ ( .A({ _23235_, _08900_, _23523_, _05684_ }), .Y(_09171_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32903_ ( .A({ _05912_, _09172_ }), .Y(_24034_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32904_ ( .A({ _09181_, _09178_, _09173_ }), .Y(_09172_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32905_ ( .A({ _09177_, _09176_, _09175_, _09174_ }), .Y(_09173_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32906_ ( .A(_stream_matmul_29_source_6_source_pat_fsm_0[23:20]), .Y(_09174_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32907_ ( .A(_stream_matmul_29_source_6_source_pat_fsm_0[19:16]), .Y(_09175_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32908_ ( .A(_stream_matmul_29_source_6_source_pat_fsm_0[31:28]), .Y(_09176_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32909_ ( .A(_stream_matmul_29_source_6_source_pat_fsm_0[27:24]), .Y(_09177_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32910_ ( .A({ _09180_, _09179_ }), .Y(_09178_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32911_ ( .A(_stream_matmul_29_source_6_source_pat_fsm_0[15:12]), .Y(_09179_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32912_ ( .A(_stream_matmul_29_source_6_source_pat_fsm_0[11:8]), .Y(_09180_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32913_ ( .A({ _09182_, _stream_matmul_29_source_6_source_pat_fsm_0[3:2], _stream_matmul_29_source_6_source_pat_fsm_0[0] }), .Y(_09181_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32914_ ( .A(_stream_matmul_29_source_6_source_pat_fsm_0[7:4]), .Y(_09182_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _32915_ ( .A({ _09183_, _09182_, _09178_, _09173_ }), .Y(_05912_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32916_ ( .A({ _stream_matmul_29_source_6_source_pat_fsm_0[0], _stream_matmul_29_source_6_source_pat_fsm_0[3:1] }), .Y(_09183_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32917_ ( .A({ _13653_, _09184_, _13621_, _05912_ }), .Y(_13589_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32918_ ( .A({ _09172_, _stream_matmul_29_source_6_source_pat_fsm_0[1] }), .Y(_09184_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32919_ ( .A({ _13652_, _09184_, _13620_, _05912_ }), .Y(_13588_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32920_ ( .A({ _13651_, _09184_, _13619_, _05912_ }), .Y(_13587_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32921_ ( .A({ _13626_, _09184_, _13594_, _05912_ }), .Y(_13562_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32922_ ( .A({ _13654_, _09184_, _13622_, _05912_ }), .Y(_13590_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32923_ ( .A({ _13632_, _09184_, _13600_, _05912_ }), .Y(_13568_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32924_ ( .A({ _13650_, _09184_, _13618_, _05912_ }), .Y(_13586_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32925_ ( .A({ _13636_, _09184_, _13604_, _05912_ }), .Y(_13572_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32926_ ( .A({ _13625_, _09184_, _13593_, _05912_ }), .Y(_13561_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32927_ ( .A({ _13647_, _09184_, _13615_, _05912_ }), .Y(_13583_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32928_ ( .A({ _13631_, _09184_, _13599_, _05912_ }), .Y(_13567_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32929_ ( .A({ _13630_, _09184_, _13598_, _05912_ }), .Y(_13566_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32930_ ( .A({ _13656_, _09184_, _13624_, _05912_ }), .Y(_13592_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32931_ ( .A({ _13655_, _09184_, _13623_, _05912_ }), .Y(_13591_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32932_ ( .A({ _13637_, _09184_, _13605_, _05912_ }), .Y(_13573_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32933_ ( .A({ _13633_, _09184_, _13601_, _05912_ }), .Y(_13569_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32934_ ( .A({ _13629_, _09184_, _13597_, _05912_ }), .Y(_13565_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32935_ ( .A({ _13628_, _09184_, _13596_, _05912_ }), .Y(_13564_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32936_ ( .A({ _13627_, _09184_, _13595_, _05912_ }), .Y(_13563_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32937_ ( .A({ _13644_, _09184_, _13612_, _05912_ }), .Y(_13580_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32938_ ( .A({ _13635_, _09184_, _13603_, _05912_ }), .Y(_13571_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32939_ ( .A({ _13643_, _09184_, _13611_, _05912_ }), .Y(_13579_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32940_ ( .A({ _13642_, _09184_, _13610_, _05912_ }), .Y(_13578_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32941_ ( .A({ _13634_, _09184_, _13602_, _05912_ }), .Y(_13570_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32942_ ( .A({ _13648_, _09184_, _13616_, _05912_ }), .Y(_13584_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32943_ ( .A({ _13645_, _09184_, _13613_, _05912_ }), .Y(_13581_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32944_ ( .A({ _13641_, _09184_, _13609_, _05912_ }), .Y(_13577_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32945_ ( .A({ _13639_, _09184_, _13607_, _05912_ }), .Y(_13575_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32946_ ( .A({ _13638_, _09184_, _13606_, _05912_ }), .Y(_13574_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32947_ ( .A({ _13640_, _09184_, _13608_, _05912_ }), .Y(_13576_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32948_ ( .A({ _13646_, _09184_, _13614_, _05912_ }), .Y(_13582_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32949_ ( .A({ _13649_, _09184_, _13617_, _05912_ }), .Y(_13585_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _32950_ ( .A({ _05911_, _09185_ }), .Y(_24033_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32951_ ( .A({ _09194_, _09191_, _09186_ }), .Y(_09185_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32952_ ( .A({ _09190_, _09189_, _09188_, _09187_ }), .Y(_09186_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32953_ ( .A(_stream_matmul_29_source_8_source_pat_fsm_1[23:20]), .Y(_09187_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32954_ ( .A(_stream_matmul_29_source_8_source_pat_fsm_1[19:16]), .Y(_09188_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32955_ ( .A(_stream_matmul_29_source_8_source_pat_fsm_1[31:28]), .Y(_09189_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32956_ ( .A(_stream_matmul_29_source_8_source_pat_fsm_1[27:24]), .Y(_09190_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _32957_ ( .A({ _09193_, _09192_ }), .Y(_09191_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32958_ ( .A(_stream_matmul_29_source_8_source_pat_fsm_1[15:12]), .Y(_09192_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32959_ ( .A(_stream_matmul_29_source_8_source_pat_fsm_1[11:8]), .Y(_09193_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32960_ ( .A({ _09195_, _stream_matmul_29_source_8_source_pat_fsm_1[3:2], _stream_matmul_29_source_8_source_pat_fsm_1[0] }), .Y(_09194_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _32961_ ( .A(_stream_matmul_29_source_8_source_pat_fsm_1[7:4]), .Y(_09195_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _32962_ ( .A({ _09196_, _09195_, _09191_, _09186_ }), .Y(_05911_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _32963_ ( .A({ _stream_matmul_29_source_8_source_pat_fsm_1[0], _stream_matmul_29_source_8_source_pat_fsm_1[3:1] }), .Y(_09196_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32964_ ( .A({ _13540_, _09197_, _13508_, _05911_ }), .Y(_13476_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _32965_ ( .A({ _09185_, _stream_matmul_29_source_8_source_pat_fsm_1[1] }), .Y(_09197_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32966_ ( .A({ _13551_, _09197_, _13519_, _05911_ }), .Y(_13487_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32967_ ( .A({ _13529_, _09197_, _13497_, _05911_ }), .Y(_13465_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32968_ ( .A({ _13555_, _09197_, _13523_, _05911_ }), .Y(_13491_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32969_ ( .A({ _13530_, _09197_, _13498_, _05911_ }), .Y(_13466_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32970_ ( .A({ _13554_, _09197_, _13522_, _05911_ }), .Y(_13490_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32971_ ( .A({ _13557_, _09197_, _13525_, _05911_ }), .Y(_13493_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32972_ ( .A({ _13531_, _09197_, _13499_, _05911_ }), .Y(_13467_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32973_ ( .A({ _13560_, _09197_, _13528_, _05911_ }), .Y(_13496_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32974_ ( .A({ _13559_, _09197_, _13527_, _05911_ }), .Y(_13495_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32975_ ( .A({ _13558_, _09197_, _13526_, _05911_ }), .Y(_13494_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32976_ ( .A({ _13556_, _09197_, _13524_, _05911_ }), .Y(_13492_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32977_ ( .A({ _13538_, _09197_, _13506_, _05911_ }), .Y(_13474_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32978_ ( .A({ _13532_, _09197_, _13500_, _05911_ }), .Y(_13468_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32979_ ( .A({ _13533_, _09197_, _13501_, _05911_ }), .Y(_13469_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32980_ ( .A({ _13539_, _09197_, _13507_, _05911_ }), .Y(_13475_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32981_ ( .A({ _13537_, _09197_, _13505_, _05911_ }), .Y(_13473_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32982_ ( .A({ _13536_, _09197_, _13504_, _05911_ }), .Y(_13472_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32983_ ( .A({ _13548_, _09197_, _13516_, _05911_ }), .Y(_13484_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32984_ ( .A({ _13541_, _09197_, _13509_, _05911_ }), .Y(_13477_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32985_ ( .A({ _13542_, _09197_, _13510_, _05911_ }), .Y(_13478_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32986_ ( .A({ _13535_, _09197_, _13503_, _05911_ }), .Y(_13471_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32987_ ( .A({ _13547_, _09197_, _13515_, _05911_ }), .Y(_13483_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32988_ ( .A({ _13546_, _09197_, _13514_, _05911_ }), .Y(_13482_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32989_ ( .A({ _13534_, _09197_, _13502_, _05911_ }), .Y(_13470_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32990_ ( .A({ _13549_, _09197_, _13517_, _05911_ }), .Y(_13485_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32991_ ( .A({ _13545_, _09197_, _13513_, _05911_ }), .Y(_13481_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32992_ ( .A({ _13543_, _09197_, _13511_, _05911_ }), .Y(_13479_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32993_ ( .A({ _13552_, _09197_, _13520_, _05911_ }), .Y(_13488_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32994_ ( .A({ _13544_, _09197_, _13512_, _05911_ }), .Y(_13480_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32995_ ( .A({ _13550_, _09197_, _13518_, _05911_ }), .Y(_13486_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _32996_ ( .A({ _13553_, _09197_, _13521_, _05911_ }), .Y(_13489_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _32997_ ( .A({ _09202_, _09200_, _09198_, _09118_ }), .Y(_24089_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _32998_ ( .A({ _09075_, _09199_, _09101_, _09087_ }), .Y(_09198_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _32999_ ( .A({ _09123_, _09079_, _09038_ }), .Y(_09199_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33000_ ( .A({ _09201_, _09125_, _09080_, _09046_ }), .Y(_09200_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33001_ ( .A({ _09160_, _09137_, _09104_ }), .Y(_09201_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33002_ ( .A({ _09206_, _09204_, _09203_, _09056_ }), .Y(_09202_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33003_ ( .A({ _09073_, _09072_ }), .Y(_09203_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33004_ ( .A({ _09205_, _09041_, _08646_, _08611_ }), .Y(_09204_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33005_ ( .A({ _05734_, _08894_, _08892_, _08891_ }), .Y(_09205_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33006_ ( .A({ _09208_, _09207_, _08902_, _08900_ }), .Y(_09206_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _33007_ ( .A({ _08903_, _09039_, _06909_ }), .Y(_09207_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33008_ ( .A({ _05684_, _08897_, _08895_, _08899_ }), .Y(_09208_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33009_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13331_, _13363_ }), .Y(_13299_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33010_ ( .A({ _09210_, _09218_, _stream_matmul_29_source_20_source_pat_fsm_3[1] }), .Y(_09209_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33011_ ( .A({ _09217_, _09216_, _09211_ }), .Y(_09210_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33012_ ( .A({ _09215_, _09214_, _09213_, _09212_ }), .Y(_09211_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33013_ ( .A(_stream_matmul_29_source_20_source_pat_fsm_3[23:20]), .Y(_09212_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33014_ ( .A(_stream_matmul_29_source_20_source_pat_fsm_3[19:16]), .Y(_09213_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33015_ ( .A(_stream_matmul_29_source_20_source_pat_fsm_3[31:28]), .Y(_09214_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33016_ ( .A(_stream_matmul_29_source_20_source_pat_fsm_3[27:24]), .Y(_09215_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33017_ ( .A(_stream_matmul_29_source_20_source_pat_fsm_3[15:12]), .Y(_09216_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33018_ ( .A(_stream_matmul_29_source_20_source_pat_fsm_3[11:8]), .Y(_09217_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33019_ ( .A({ _09219_, _stream_matmul_29_source_20_source_pat_fsm_3[3:2] }), .Y(_09218_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33020_ ( .A(_stream_matmul_29_source_20_source_pat_fsm_3[7:4]), .Y(_09219_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33021_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13330_, _13362_ }), .Y(_13298_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33022_ ( .A({ _05908_, _09209_ }), .Y(_24031_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _33023_ ( .A({ _stream_matmul_29_source_20_source_pat_fsm_3[1], _09210_, _09218_, _stream_matmul_29_source_20_source_pat_fsm_3[0] }), .Y(_05908_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33024_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13335_, _13367_ }), .Y(_13303_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33025_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13332_, _13364_ }), .Y(_13300_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33026_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13310_, _13342_ }), .Y(_13278_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33027_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13327_, _13359_ }), .Y(_13295_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33028_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13316_, _13348_ }), .Y(_13284_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33029_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13334_, _13366_ }), .Y(_13302_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33030_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13305_, _13337_ }), .Y(_13273_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33031_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13309_, _13341_ }), .Y(_13277_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33032_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13333_, _13365_ }), .Y(_13301_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33033_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13311_, _13343_ }), .Y(_13279_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33034_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13308_, _13340_ }), .Y(_13276_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33035_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13336_, _13368_ }), .Y(_13304_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33036_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13319_, _13351_ }), .Y(_13287_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33037_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13307_, _13339_ }), .Y(_13275_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33038_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13314_, _13346_ }), .Y(_13282_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33039_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13306_, _13338_ }), .Y(_13274_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33040_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13318_, _13350_ }), .Y(_13286_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33041_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13317_, _13349_ }), .Y(_13285_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33042_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13313_, _13345_ }), .Y(_13281_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33043_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13312_, _13344_ }), .Y(_13280_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33044_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13323_, _13355_ }), .Y(_13291_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33045_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13320_, _13352_ }), .Y(_13288_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33046_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13315_, _13347_ }), .Y(_13283_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33047_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13322_, _13354_ }), .Y(_13290_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33048_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13321_, _13353_ }), .Y(_13289_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33049_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13329_, _13361_ }), .Y(_13297_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33050_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13326_, _13358_ }), .Y(_13294_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33051_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13325_, _13357_ }), .Y(_13293_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33052_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13328_, _13360_ }), .Y(_13296_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33053_ ( .A({ _09209_, _stream_matmul_29_source_20_source_pat_fsm_3[0], _13324_, _13356_ }), .Y(_13292_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33054_ ( .A({ _05913_, _09220_ }), .Y(_24032_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33055_ ( .A({ _09221_, _09226_, _stream_matmul_29_source_19_source_pat_fsm_2[0] }), .Y(_09220_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33056_ ( .A({ _09225_, _09224_, _09222_ }), .Y(_09221_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33057_ ( .A({ _09223_, _stream_matmul_29_source_19_source_pat_fsm_2[3:2] }), .Y(_09222_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33058_ ( .A(_stream_matmul_29_source_19_source_pat_fsm_2[7:4]), .Y(_09223_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33059_ ( .A(_stream_matmul_29_source_19_source_pat_fsm_2[15:12]), .Y(_09224_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33060_ ( .A(_stream_matmul_29_source_19_source_pat_fsm_2[11:8]), .Y(_09225_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33061_ ( .A({ _09230_, _09229_, _09228_, _09227_ }), .Y(_09226_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33062_ ( .A(_stream_matmul_29_source_19_source_pat_fsm_2[23:20]), .Y(_09227_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33063_ ( .A(_stream_matmul_29_source_19_source_pat_fsm_2[19:16]), .Y(_09228_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33064_ ( .A(_stream_matmul_29_source_19_source_pat_fsm_2[31:28]), .Y(_09229_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33065_ ( .A(_stream_matmul_29_source_19_source_pat_fsm_2[27:24]), .Y(_09230_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _33066_ ( .A({ _09221_, _stream_matmul_29_source_19_source_pat_fsm_2[0], _09226_, _stream_matmul_29_source_19_source_pat_fsm_2[1] }), .Y(_05913_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33067_ ( .A({ _13433_, _09231_, _13401_, _05913_ }), .Y(_13369_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33068_ ( .A({ _09220_, _stream_matmul_29_source_19_source_pat_fsm_2[1] }), .Y(_09231_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33069_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18339_, _18371_ }), .Y(_18307_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33070_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18340_, _18372_ }), .Y(_18308_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33071_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18329_, _18361_ }), .Y(_18297_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33072_ ( .A({ _13455_, _09231_, _13423_, _05913_ }), .Y(_13391_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33073_ ( .A({ _13444_, _09231_, _13412_, _05913_ }), .Y(_13380_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33074_ ( .A({ _13458_, _09231_, _13426_, _05913_ }), .Y(_13394_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33075_ ( .A({ _13459_, _09231_, _13427_, _05913_ }), .Y(_13395_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33076_ ( .A({ _13460_, _09231_, _13428_, _05913_ }), .Y(_13396_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33077_ ( .A({ _13461_, _09231_, _13429_, _05913_ }), .Y(_13397_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33078_ ( .A({ _13462_, _09231_, _13430_, _05913_ }), .Y(_13398_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33079_ ( .A({ _13463_, _09231_, _13431_, _05913_ }), .Y(_13399_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33080_ ( .A({ _13464_, _09231_, _13432_, _05913_ }), .Y(_13400_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33081_ ( .A({ _13434_, _09231_, _13402_, _05913_ }), .Y(_13370_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33082_ ( .A({ _13435_, _09231_, _13403_, _05913_ }), .Y(_13371_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33083_ ( .A({ _13436_, _09231_, _13404_, _05913_ }), .Y(_13372_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33084_ ( .A({ _13437_, _09231_, _13405_, _05913_ }), .Y(_13373_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33085_ ( .A({ _13438_, _09231_, _13406_, _05913_ }), .Y(_13374_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33086_ ( .A({ _13439_, _09231_, _13407_, _05913_ }), .Y(_13375_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33087_ ( .A({ _13440_, _09231_, _13408_, _05913_ }), .Y(_13376_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33088_ ( .A({ _13441_, _09231_, _13409_, _05913_ }), .Y(_13377_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33089_ ( .A({ _13442_, _09231_, _13410_, _05913_ }), .Y(_13378_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33090_ ( .A({ _13443_, _09231_, _13411_, _05913_ }), .Y(_13379_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33091_ ( .A({ _13445_, _09231_, _13413_, _05913_ }), .Y(_13381_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33092_ ( .A({ _13446_, _09231_, _13414_, _05913_ }), .Y(_13382_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33093_ ( .A({ _13447_, _09231_, _13415_, _05913_ }), .Y(_13383_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33094_ ( .A({ _13448_, _09231_, _13416_, _05913_ }), .Y(_13384_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33095_ ( .A({ _13449_, _09231_, _13417_, _05913_ }), .Y(_13385_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33096_ ( .A({ _13450_, _09231_, _13418_, _05913_ }), .Y(_13386_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33097_ ( .A({ _13451_, _09231_, _13419_, _05913_ }), .Y(_13387_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33098_ ( .A({ _13452_, _09231_, _13420_, _05913_ }), .Y(_13388_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33099_ ( .A({ _13453_, _09231_, _13421_, _05913_ }), .Y(_13389_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33100_ ( .A({ _13454_, _09231_, _13422_, _05913_ }), .Y(_13390_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33101_ ( .A({ _13456_, _09231_, _13424_, _05913_ }), .Y(_13392_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33102_ ( .A({ _13457_, _09231_, _13425_, _05913_ }), .Y(_13393_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33103_ ( .A({ _09240_, _09239_, _09234_, _09232_ }), .Y(_24030_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33104_ ( .A({ _09233_, _stream_matmul_29_sink_21_sink_fsm_4[31:29] }), .Y(_09232_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33105_ ( .A(_stream_matmul_29_sink_21_sink_fsm_4[28:25]), .Y(_09233_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33106_ ( .A({ _09238_, _09237_, _09236_, _09235_ }), .Y(_09234_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33107_ ( .A(_stream_matmul_29_sink_21_sink_fsm_4[8:5]), .Y(_09235_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33108_ ( .A(_stream_matmul_29_sink_21_sink_fsm_4[4:1]), .Y(_09236_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33109_ ( .A(_stream_matmul_29_sink_21_sink_fsm_4[16:13]), .Y(_09237_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33110_ ( .A(_stream_matmul_29_sink_21_sink_fsm_4[12:9]), .Y(_09238_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33111_ ( .A(_stream_matmul_29_sink_21_sink_fsm_4[24:21]), .Y(_09239_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33112_ ( .A(_stream_matmul_29_sink_21_sink_fsm_4[20:17]), .Y(_09240_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33113_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13177_, _13241_ }), .Y(_13209_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33114_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13188_, _13252_ }), .Y(_13220_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33115_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13199_, _13263_ }), .Y(_13231_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33116_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13202_, _13266_ }), .Y(_13234_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33117_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13203_, _13267_ }), .Y(_13235_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33118_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13204_, _13268_ }), .Y(_13236_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33119_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13205_, _13269_ }), .Y(_13237_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33120_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13206_, _13270_ }), .Y(_13238_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33121_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13207_, _13271_ }), .Y(_13239_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33122_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13208_, _13272_ }), .Y(_13240_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33123_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13178_, _13242_ }), .Y(_13210_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33124_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13179_, _13243_ }), .Y(_13211_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33125_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13180_, _13244_ }), .Y(_13212_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33126_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13181_, _13245_ }), .Y(_13213_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33127_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13182_, _13246_ }), .Y(_13214_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33128_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13183_, _13247_ }), .Y(_13215_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33129_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13184_, _13248_ }), .Y(_13216_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33130_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13185_, _13249_ }), .Y(_13217_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33131_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13186_, _13250_ }), .Y(_13218_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33132_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13187_, _13251_ }), .Y(_13219_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33133_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13189_, _13253_ }), .Y(_13221_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33134_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13190_, _13254_ }), .Y(_13222_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33135_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13191_, _13255_ }), .Y(_13223_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33136_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13192_, _13256_ }), .Y(_13224_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33137_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13193_, _13257_ }), .Y(_13225_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33138_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13194_, _13258_ }), .Y(_13226_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33139_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13195_, _13259_ }), .Y(_13227_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33140_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13196_, _13260_ }), .Y(_13228_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33141_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13197_, _13261_ }), .Y(_13229_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33142_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13198_, _13262_ }), .Y(_13230_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33143_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13200_, _13264_ }), .Y(_13232_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33144_ ( .A({ _24030_, _stream_matmul_29_sink_21_sink_fsm_4[0], _13201_, _13265_ }), .Y(_13233_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33145_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18421_, _18453_ }), .Y(_18389_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33146_ ( .A({ _09242_, _09250_, _stream_conv2d_16_source_25_source_pat_fsm_8[1] }), .Y(_09241_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33147_ ( .A({ _09249_, _09248_, _09243_ }), .Y(_09242_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33148_ ( .A({ _09247_, _09246_, _09245_, _09244_ }), .Y(_09243_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33149_ ( .A(_stream_conv2d_16_source_25_source_pat_fsm_8[23:20]), .Y(_09244_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33150_ ( .A(_stream_conv2d_16_source_25_source_pat_fsm_8[19:16]), .Y(_09245_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33151_ ( .A(_stream_conv2d_16_source_25_source_pat_fsm_8[31:28]), .Y(_09246_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33152_ ( .A(_stream_conv2d_16_source_25_source_pat_fsm_8[27:24]), .Y(_09247_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33153_ ( .A(_stream_conv2d_16_source_25_source_pat_fsm_8[15:12]), .Y(_09248_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33154_ ( .A(_stream_conv2d_16_source_25_source_pat_fsm_8[11:8]), .Y(_09249_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33155_ ( .A({ _09251_, _stream_conv2d_16_source_25_source_pat_fsm_8[3:2] }), .Y(_09250_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33156_ ( .A(_stream_conv2d_16_source_25_source_pat_fsm_8[7:4]), .Y(_09251_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33157_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18530_, _18562_ }), .Y(_18498_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33158_ ( .A({ _09253_, _09261_, _stream_conv2d_16_source_24_source_pat_fsm_7[1] }), .Y(_09252_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33159_ ( .A({ _09260_, _09259_, _09254_ }), .Y(_09253_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33160_ ( .A({ _09258_, _09257_, _09256_, _09255_ }), .Y(_09254_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33161_ ( .A(_stream_conv2d_16_source_24_source_pat_fsm_7[23:20]), .Y(_09255_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33162_ ( .A(_stream_conv2d_16_source_24_source_pat_fsm_7[19:16]), .Y(_09256_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33163_ ( .A(_stream_conv2d_16_source_24_source_pat_fsm_7[31:28]), .Y(_09257_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33164_ ( .A(_stream_conv2d_16_source_24_source_pat_fsm_7[27:24]), .Y(_09258_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33165_ ( .A(_stream_conv2d_16_source_24_source_pat_fsm_7[15:12]), .Y(_09259_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33166_ ( .A(_stream_conv2d_16_source_24_source_pat_fsm_7[11:8]), .Y(_09260_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33167_ ( .A({ _09262_, _stream_conv2d_16_source_24_source_pat_fsm_7[3:2] }), .Y(_09261_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33168_ ( .A(_stream_conv2d_16_source_24_source_pat_fsm_7[7:4]), .Y(_09262_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33169_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18906_, _18938_ }), .Y(_18874_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33170_ ( .A({ _09264_, _09272_, _stream_conv2d_16_source_20_source_pat_fsm_3[1] }), .Y(_09263_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33171_ ( .A({ _09271_, _09270_, _09265_ }), .Y(_09264_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33172_ ( .A({ _09269_, _09268_, _09267_, _09266_ }), .Y(_09265_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33173_ ( .A(_stream_conv2d_16_source_20_source_pat_fsm_3[23:20]), .Y(_09266_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33174_ ( .A(_stream_conv2d_16_source_20_source_pat_fsm_3[19:16]), .Y(_09267_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33175_ ( .A(_stream_conv2d_16_source_20_source_pat_fsm_3[31:28]), .Y(_09268_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33176_ ( .A(_stream_conv2d_16_source_20_source_pat_fsm_3[27:24]), .Y(_09269_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33177_ ( .A(_stream_conv2d_16_source_20_source_pat_fsm_3[15:12]), .Y(_09270_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33178_ ( .A(_stream_conv2d_16_source_20_source_pat_fsm_3[11:8]), .Y(_09271_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33179_ ( .A({ _09273_, _stream_conv2d_16_source_20_source_pat_fsm_3[3:2] }), .Y(_09272_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33180_ ( .A(_stream_conv2d_16_source_20_source_pat_fsm_3[7:4]), .Y(_09273_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33181_ ( .A({ _20105_, _05996_, _09285_, _20171_ }), .Y(_20138_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _33182_ ( .A({ _maxi_read_fsm[0], _09283_, _09274_ }), .Y(_05996_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33183_ ( .A({ _09280_, _09275_ }), .Y(_09274_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33184_ ( .A({ _09279_, _09278_, _09277_, _09276_ }), .Y(_09275_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33185_ ( .A(_maxi_read_fsm[23:20]), .Y(_09276_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33186_ ( .A(_maxi_read_fsm[19:16]), .Y(_09277_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33187_ ( .A(_maxi_read_fsm[31:28]), .Y(_09278_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33188_ ( .A(_maxi_read_fsm[27:24]), .Y(_09279_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33189_ ( .A({ _09282_, _09281_ }), .Y(_09280_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33190_ ( .A(_maxi_read_fsm[15:12]), .Y(_09281_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33191_ ( .A(_maxi_read_fsm[11:8]), .Y(_09282_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33192_ ( .A({ _09284_, _maxi_read_fsm[2:1], _maxi_read_fsm[3] }), .Y(_09283_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33193_ ( .A(_maxi_read_fsm[7:4]), .Y(_09284_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33194_ ( .A({ _09275_, _09286_, _maxi_read_fsm[1:0] }), .Y(_09285_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33195_ ( .A({ _09284_, _09280_, _maxi_read_fsm[2], _maxi_read_fsm[3] }), .Y(_09286_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _33196_ ( .A({ _05991_, _20019_, _09298_ }), .Y(_20021_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _33197_ ( .A({ _09287_, _09293_, conv2d_16_comp_fsm[1] }), .Y(_05991_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33198_ ( .A({ conv2d_16_comp_fsm[0], _09288_ }), .Y(_09287_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33199_ ( .A({ _09292_, _09291_, _09290_, _09289_ }), .Y(_09288_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33200_ ( .A(conv2d_16_comp_fsm[23:20]), .Y(_09289_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33201_ ( .A(conv2d_16_comp_fsm[19:16]), .Y(_09290_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33202_ ( .A(conv2d_16_comp_fsm[31:28]), .Y(_09291_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33203_ ( .A(conv2d_16_comp_fsm[27:24]), .Y(_09292_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33204_ ( .A({ _09294_, conv2d_16_comp_fsm[2], conv2d_16_comp_fsm[3] }), .Y(_09293_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33205_ ( .A({ _09297_, _09296_, _09295_ }), .Y(_09294_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33206_ ( .A(conv2d_16_comp_fsm[15:12]), .Y(_09295_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33207_ ( .A(conv2d_16_comp_fsm[7:4]), .Y(_09296_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33208_ ( .A(conv2d_16_comp_fsm[11:8]), .Y(_09297_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33209_ ( .A({ _09300_, _09299_ }), .Y(_09298_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33210_ ( .A({ conv2d_16_comp_fsm[2], _09294_, conv2d_16_comp_fsm[3] }), .Y(_09299_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33211_ ( .A({ conv2d_16_comp_fsm[1], _09288_, conv2d_16_comp_fsm[0] }), .Y(_09300_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33212_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18420_, _18452_ }), .Y(_18388_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33213_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18529_, _18561_ }), .Y(_18497_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33214_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18895_, _18927_ }), .Y(_18863_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33215_ ( .A({ _20104_, _05996_, _09285_, _20170_ }), .Y(_20137_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33216_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18419_, _18451_ }), .Y(_18387_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33217_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18528_, _18560_ }), .Y(_18496_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33218_ ( .A({ _20103_, _05996_, _09285_, _20169_ }), .Y(_20136_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33219_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18418_, _18450_ }), .Y(_18386_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33220_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18527_, _18559_ }), .Y(_18495_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33221_ ( .A({ _20102_, _05996_, _09285_, _20168_ }), .Y(_20135_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33222_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18526_, _18558_ }), .Y(_18494_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33223_ ( .A({ _20101_, _05996_, _09285_, _20167_ }), .Y(_20134_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33224_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18525_, _18557_ }), .Y(_18493_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33225_ ( .A({ _20100_, _05996_, _09285_, _20166_ }), .Y(_20133_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33226_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18524_, _18556_ }), .Y(_18492_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33227_ ( .A({ _05980_, _09263_ }), .Y(_24066_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _33228_ ( .A({ _stream_conv2d_16_source_20_source_pat_fsm_3[1], _09264_, _09272_, _stream_conv2d_16_source_20_source_pat_fsm_3[0] }), .Y(_05980_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33229_ ( .A({ _20099_, _05996_, _09285_, _20165_ }), .Y(_20132_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _33230_ ( .A({ _09304_, _09301_ }), .Y(_24070_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33231_ ( .A({ _05989_, _05727_, _09303_, _09298_ }), .Y(_09301_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _33232_ ( .A({ conv2d_16_comp_fsm[1], _09293_, _09287_ }), .Y(_05989_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _33233_ ( .A({ _09302_, _09293_ }), .Y(_05727_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33234_ ( .A({ _09288_, conv2d_16_comp_fsm[1:0] }), .Y(_09302_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33235_ ( .A({ _09302_, _09299_ }), .Y(_09303_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33236_ ( .A({ _05990_, _05991_, _09305_ }), .Y(_09304_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33237_ ( .A({ _09287_, _09299_, conv2d_16_comp_fsm[1] }), .Y(_09305_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _33238_ ( .A({ _09300_, _09293_ }), .Y(_05990_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33239_ ( .A({ _20098_, _05996_, _09285_, _20164_ }), .Y(_20131_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33240_ ( .A({ _20096_, _05996_, _09285_, _20162_ }), .Y(_20129_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33241_ ( .A({ cparam_matmul_29_max_och_count[3], matmul_29_och_count[3], cparam_matmul_29_max_och_count[2], matmul_29_och_count[2] }), .Y(_09306_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _33242_ ( .A({ cparam_matmul_29_max_och_count[1], matmul_29_och_count[1:0], cparam_matmul_29_max_och_count[0] }), .Y(_09307_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33243_ ( .A({ cparam_matmul_29_max_och_count[2], cparam_matmul_29_max_och_count[3], matmul_29_och_count[2], matmul_29_och_count[3] }), .Y(_09308_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33244_ ( .A({ cparam_matmul_29_max_och_count[5], matmul_29_och_count[5] }), .Y(_09309_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33245_ ( .A({ cparam_matmul_29_max_och_count[6], matmul_29_och_count[6], cparam_matmul_29_max_och_count[7], matmul_29_och_count[7] }), .Y(_09310_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33246_ ( .A({ matmul_29_och_count[5], cparam_matmul_29_max_och_count[5], matmul_29_och_count[6], cparam_matmul_29_max_och_count[6] }), .Y(_09311_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33247_ ( .A({ _09306_, _09313_, matmul_29_och_count[0], cparam_matmul_29_max_och_count[0] }), .Y(_09312_) );
  \$lut  #( .LUT(16'h9000), .WIDTH(4) ) _33248_ ( .A({ _09315_, _09314_, cparam_matmul_29_max_och_count[6], matmul_29_och_count[6] }), .Y(_09313_) );
  \$lut  #( .LUT(8'h41), .WIDTH(3) ) _33249_ ( .A({ cparam_matmul_29_max_och_count[4], matmul_29_och_count[4], _09309_ }), .Y(_09314_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _33250_ ( .A({ cparam_matmul_29_max_och_count[7], matmul_29_och_count[7], matmul_29_och_count[5], cparam_matmul_29_max_och_count[5] }), .Y(_09315_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33251_ ( .A({ _09324_, _09323_, _09321_, _09317_ }), .Y(_09316_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33252_ ( .A({ _09320_, _09319_, _09318_ }), .Y(_09317_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33253_ ( .A(matmul_29_och_count[31:28]), .Y(_09318_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33254_ ( .A(matmul_29_och_count[27:24]), .Y(_09319_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33255_ ( .A(matmul_29_och_count[23:20]), .Y(_09320_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _33256_ ( .A({ _09322_, matmul_29_och_count[7], cparam_matmul_29_max_och_count[7] }), .Y(_09321_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33257_ ( .A(matmul_29_och_count[11:8]), .Y(_09322_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33258_ ( .A(matmul_29_och_count[19:16]), .Y(_09323_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33259_ ( .A(matmul_29_och_count[15:12]), .Y(_09324_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33260_ ( .A({ _20095_, _05996_, _09285_, _20161_ }), .Y(_20128_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33261_ ( .A({ _20094_, _05996_, _09285_, _20160_ }), .Y(_20127_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33262_ ( .A({ _20093_, _05996_, _09285_, _20159_ }), .Y(_20126_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33263_ ( .A({ _20092_, _05996_, _09285_, _20158_ }), .Y(_20125_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33264_ ( .A({ _20091_, _05996_, _09285_, _20157_ }), .Y(_20124_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33265_ ( .A({ _20090_, _05996_, _09285_, _20156_ }), .Y(_20123_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33266_ ( .A({ _20089_, _05996_, _09285_, _20155_ }), .Y(_20122_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33267_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18417_, _18449_ }), .Y(_18385_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33268_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18523_, _18555_ }), .Y(_18491_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33269_ ( .A({ _20088_, _05996_, _09285_, _20154_ }), .Y(_20121_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33270_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18416_, _18448_ }), .Y(_18384_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33271_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18521_, _18553_ }), .Y(_18489_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33272_ ( .A({ _20087_, _05996_, _09285_, _20153_ }), .Y(_20120_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _33273_ ( .A({ _09340_, _09335_, _09326_, _09338_ }), .Y(_09325_) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _33274_ ( .A({ matmul_29_sync_comp_count[7], _09327_, _09334_, _05191_ }), .Y(_09326_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _33275_ ( .A({ _09333_, _09332_, _09331_, _09328_ }), .Y(_09327_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _33276_ ( .A({ _09330_, matmul_29_sync_comp_count[2], _05184_, _09329_ }), .Y(_09328_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _33277_ ( .A({ _05162_, matmul_29_sync_comp_count[0], matmul_29_sync_comp_count[1], _05173_ }), .Y(_09329_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33278_ ( .A({ _05187_, matmul_29_sync_comp_count[3] }), .Y(_09330_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33279_ ( .A({ matmul_29_sync_comp_count[3], _05187_, matmul_29_sync_comp_count[4], _05188_ }), .Y(_09331_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33280_ ( .A({ _05188_, matmul_29_sync_comp_count[4], _05189_, matmul_29_sync_comp_count[5] }), .Y(_09332_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33281_ ( .A({ matmul_29_sync_comp_count[5], _05189_, matmul_29_sync_comp_count[6], _05190_ }), .Y(_09333_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33282_ ( .A({ _05190_, matmul_29_sync_comp_count[6] }), .Y(_09334_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _33283_ ( .A({ _09337_, _09336_, _05193_, matmul_29_sync_comp_count[9] }), .Y(_09335_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33284_ ( .A({ matmul_29_sync_comp_count[8], _05192_, matmul_29_sync_comp_count[9], _05193_ }), .Y(_09336_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33285_ ( .A({ matmul_29_sync_comp_count[11], _05164_, matmul_29_sync_comp_count[10], _05163_ }), .Y(_09337_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33286_ ( .A({ _09339_, _09337_, _09336_ }), .Y(_09338_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33287_ ( .A({ _05192_, matmul_29_sync_comp_count[8], _05193_, matmul_29_sync_comp_count[9] }), .Y(_09339_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33288_ ( .A({ matmul_29_sync_comp_count[10], matmul_29_sync_comp_count[11], _05163_, _05164_ }), .Y(_09340_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33289_ ( .A({ _09352_, _09348_, _09342_ }), .Y(_09341_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33290_ ( .A({ _09347_, _09346_, _09343_ }), .Y(_09342_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33291_ ( .A({ _09345_, _09344_ }), .Y(_09343_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33292_ ( .A({ matmul_29_sync_comp_count[31], _05186_, matmul_29_sync_comp_count[30], _05185_ }), .Y(_09344_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33293_ ( .A({ matmul_29_sync_comp_count[29], _05183_, matmul_29_sync_comp_count[28], _05182_ }), .Y(_09345_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33294_ ( .A({ matmul_29_sync_comp_count[27], _05181_, matmul_29_sync_comp_count[26], _05180_ }), .Y(_09346_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33295_ ( .A({ matmul_29_sync_comp_count[25], _05179_, matmul_29_sync_comp_count[24], _05178_ }), .Y(_09347_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _33296_ ( .A({ _09351_, _09349_, _05169_, matmul_29_sync_comp_count[16] }), .Y(_09348_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _33297_ ( .A({ _09350_, _05170_, matmul_29_sync_comp_count[17] }), .Y(_09349_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33298_ ( .A({ matmul_29_sync_comp_count[19], _05172_, matmul_29_sync_comp_count[18], _05171_ }), .Y(_09350_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33299_ ( .A({ matmul_29_sync_comp_count[16], _05169_, matmul_29_sync_comp_count[17], _05170_ }), .Y(_09351_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33300_ ( .A({ _09354_, _09353_ }), .Y(_09352_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33301_ ( .A({ matmul_29_sync_comp_count[23], _05177_, matmul_29_sync_comp_count[22], _05176_ }), .Y(_09353_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33302_ ( .A({ matmul_29_sync_comp_count[21], _05175_, matmul_29_sync_comp_count[20], _05174_ }), .Y(_09354_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33303_ ( .A({ matmul_29_sync_comp_count[15], _05168_, matmul_29_sync_comp_count[14], _05167_ }), .Y(_09355_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33304_ ( .A({ matmul_29_sync_comp_count[13], _05166_, matmul_29_sync_comp_count[12], _05165_ }), .Y(_09356_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33305_ ( .A({ matmul_29_sync_comp_count[14], matmul_29_sync_comp_count[15], _05167_, _05168_ }), .Y(_09357_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33306_ ( .A({ matmul_29_sync_comp_count[12], matmul_29_sync_comp_count[13], _05165_, _05166_ }), .Y(_09358_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _33307_ ( .A({ _09364_, _09362_, _09360_, _09352_ }), .Y(_09359_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _33308_ ( .A({ _09361_, _09349_, _09351_ }), .Y(_09360_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33309_ ( .A({ matmul_29_sync_comp_count[18], matmul_29_sync_comp_count[19], _05171_, _05172_ }), .Y(_09361_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _33310_ ( .A({ _09353_, matmul_29_sync_comp_count[21], _05175_, _09363_ }), .Y(_09362_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33311_ ( .A({ matmul_29_sync_comp_count[20], _05174_ }), .Y(_09363_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33312_ ( .A({ matmul_29_sync_comp_count[22], matmul_29_sync_comp_count[23], _05176_, _05177_ }), .Y(_09364_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _33313_ ( .A({ _09370_, _09366_, _09344_, _09369_ }), .Y(_09365_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _33314_ ( .A({ _09343_, _09367_, _09368_, _09346_ }), .Y(_09366_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33315_ ( .A({ matmul_29_sync_comp_count[26], matmul_29_sync_comp_count[27], _05180_, _05181_ }), .Y(_09367_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33316_ ( .A({ matmul_29_sync_comp_count[24], matmul_29_sync_comp_count[25], _05178_, _05179_ }), .Y(_09368_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33317_ ( .A({ matmul_29_sync_comp_count[28], matmul_29_sync_comp_count[29], _05182_, _05183_ }), .Y(_09369_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33318_ ( .A({ matmul_29_sync_comp_count[30], matmul_29_sync_comp_count[31], _05185_, _05186_ }), .Y(_09370_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33319_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18631_, _18663_ }), .Y(_18599_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33320_ ( .A({ _09372_, _09380_, _stream_conv2d_16_source_23_source_pat_fsm_6[1] }), .Y(_09371_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33321_ ( .A({ _09379_, _09378_, _09373_ }), .Y(_09372_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33322_ ( .A({ _09377_, _09376_, _09375_, _09374_ }), .Y(_09373_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33323_ ( .A(_stream_conv2d_16_source_23_source_pat_fsm_6[23:20]), .Y(_09374_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33324_ ( .A(_stream_conv2d_16_source_23_source_pat_fsm_6[19:16]), .Y(_09375_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33325_ ( .A(_stream_conv2d_16_source_23_source_pat_fsm_6[31:28]), .Y(_09376_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33326_ ( .A(_stream_conv2d_16_source_23_source_pat_fsm_6[27:24]), .Y(_09377_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33327_ ( .A(_stream_conv2d_16_source_23_source_pat_fsm_6[15:12]), .Y(_09378_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33328_ ( .A(_stream_conv2d_16_source_23_source_pat_fsm_6[11:8]), .Y(_09379_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33329_ ( .A({ _09381_, _stream_conv2d_16_source_23_source_pat_fsm_6[3:2] }), .Y(_09380_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33330_ ( .A(_stream_conv2d_16_source_23_source_pat_fsm_6[7:4]), .Y(_09381_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33331_ ( .A({ _20118_, _05996_, _09285_, _20184_ }), .Y(_20151_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33332_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18630_, _18662_ }), .Y(_18598_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33333_ ( .A({ _20117_, _05996_, _09285_, _20183_ }), .Y(_20150_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33334_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18628_, _18660_ }), .Y(_18596_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33335_ ( .A({ _20116_, _05996_, _09285_, _20182_ }), .Y(_20149_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33336_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18627_, _18659_ }), .Y(_18595_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33337_ ( .A({ _20115_, _05996_, _09285_, _20181_ }), .Y(_20148_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _33338_ ( .A({ _09383_, max_pool_serial_18_col_count[2], cparam_max_pool_serial_18_max_col_count[2], _09384_ }), .Y(_09382_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33339_ ( .A({ cparam_max_pool_serial_18_max_col_count[3], max_pool_serial_18_col_count[3] }), .Y(_09383_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33340_ ( .A({ max_pool_serial_18_col_count[1], cparam_max_pool_serial_18_max_col_count[1] }), .Y(_09384_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33341_ ( .A({ _09383_, max_pool_serial_18_col_count[1], cparam_max_pool_serial_18_max_col_count[1] }), .Y(_09385_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33342_ ( .A({ cparam_max_pool_serial_18_max_col_count[2], max_pool_serial_18_col_count[2], cparam_max_pool_serial_18_max_col_count[0], max_pool_serial_18_col_count[0] }), .Y(_09386_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33343_ ( .A({ _09390_, _09388_ }), .Y(_09387_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33344_ ( .A({ _09389_, max_pool_serial_18_col_count[18], max_pool_serial_18_col_count[9], max_pool_serial_18_col_count[21] }), .Y(_09388_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33345_ ( .A({ max_pool_serial_18_col_count[17:16], max_pool_serial_18_col_count[14], max_pool_serial_18_col_count[10] }), .Y(_09389_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33346_ ( .A({ max_pool_serial_18_col_count[20], max_pool_serial_18_col_count[15], max_pool_serial_18_col_count[13:12] }), .Y(_09390_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33347_ ( .A({ _09395_, _09394_, _09392_ }), .Y(_09391_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33348_ ( .A({ _09393_, max_pool_serial_18_col_count[31], max_pool_serial_18_col_count[8], max_pool_serial_18_col_count[30] }), .Y(_09392_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33349_ ( .A(max_pool_serial_18_col_count[29:26]), .Y(_09393_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33350_ ( .A(max_pool_serial_18_col_count[25:22]), .Y(_09394_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33351_ ( .A({ max_pool_serial_18_col_count[19], max_pool_serial_18_col_count[11], max_pool_serial_18_col_count[7:6] }), .Y(_09395_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33352_ ( .A({ _20114_, _05996_, _09285_, _20180_ }), .Y(_20147_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33353_ ( .A({ _20113_, _05996_, _09285_, _20179_ }), .Y(_20146_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33354_ ( .A({ _20112_, _05996_, _09285_, _20178_ }), .Y(_20145_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33355_ ( .A({ _20108_, _05996_, _09285_, _20174_ }), .Y(_20141_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33356_ ( .A({ _20097_, _05996_, _09285_, _20163_ }), .Y(_20130_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33357_ ( .A({ _09397_, max_pool_serial_18_row_count[18], max_pool_serial_18_row_count[15] }), .Y(_09396_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33358_ ( .A({ _09404_, _09403_, _09402_, _09398_ }), .Y(_09397_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33359_ ( .A({ _09401_, _09399_, max_pool_serial_18_row_count[19], max_pool_serial_18_row_count[14] }), .Y(_09398_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33360_ ( .A({ _09400_, max_pool_serial_18_row_count[7:6] }), .Y(_09399_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33361_ ( .A({ max_pool_serial_18_row_count[13:11], max_pool_serial_18_row_count[8] }), .Y(_09400_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33362_ ( .A({ max_pool_serial_18_row_count[31:29], max_pool_serial_18_row_count[25] }), .Y(_09401_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33363_ ( .A({ max_pool_serial_18_row_count[28:26], max_pool_serial_18_row_count[24] }), .Y(_09402_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33364_ ( .A(max_pool_serial_18_row_count[23:20]), .Y(_09403_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33365_ ( .A({ max_pool_serial_18_row_count[17:16], max_pool_serial_18_row_count[10:9] }), .Y(_09404_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _33366_ ( .A({ _09406_, max_pool_serial_18_row_count[2], cparam_max_pool_serial_18_max_col_count[2], _09407_ }), .Y(_09405_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33367_ ( .A({ cparam_max_pool_serial_18_max_col_count[3], max_pool_serial_18_row_count[3] }), .Y(_09406_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33368_ ( .A({ max_pool_serial_18_row_count[1], cparam_max_pool_serial_18_max_col_count[1] }), .Y(_09407_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _33369_ ( .A({ _09406_, max_pool_serial_18_row_count[1], cparam_max_pool_serial_18_max_col_count[1] }), .Y(_09408_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33370_ ( .A({ cparam_max_pool_serial_18_max_col_count[0], max_pool_serial_18_row_count[0], cparam_max_pool_serial_18_max_col_count[2], max_pool_serial_18_row_count[2] }), .Y(_09409_) );
  \$lut  #( .LUT(16'hbf00), .WIDTH(4) ) _33371_ ( .A({ _09428_, _09432_, _09430_, _09411_ }), .Y(_09410_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _33372_ ( .A({ _09424_, _09421_, _09427_, _09412_ }), .Y(_09411_) );
  \$lut  #( .LUT(16'h00f4), .WIDTH(4) ) _33373_ ( .A({ _09418_, _09419_, _09420_, _09413_ }), .Y(_09412_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _33374_ ( .A({ _09417_, _09416_, _09414_, _09415_ }), .Y(_09413_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _33375_ ( .A({ _05130_, max_pool_serial_18_comp_count[0], max_pool_serial_18_comp_count[1], _05141_ }), .Y(_09414_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _33376_ ( .A({ max_pool_serial_18_comp_count[2], _05152_, _05155_, max_pool_serial_18_comp_count[3] }), .Y(_09415_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _33377_ ( .A({ max_pool_serial_18_comp_count[2], _05152_, _05155_, max_pool_serial_18_comp_count[3] }), .Y(_09416_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33378_ ( .A({ max_pool_serial_18_comp_count[3], _05155_, max_pool_serial_18_comp_count[4], _05156_ }), .Y(_09417_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33379_ ( .A({ _05158_, max_pool_serial_18_comp_count[6] }), .Y(_09418_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33380_ ( .A({ max_pool_serial_18_comp_count[5], _05157_ }), .Y(_09419_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33381_ ( .A({ _05156_, max_pool_serial_18_comp_count[4], _05157_, max_pool_serial_18_comp_count[5] }), .Y(_09420_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _33382_ ( .A({ _09423_, _09422_, _05159_, max_pool_serial_18_comp_count[7] }), .Y(_09421_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33383_ ( .A({ max_pool_serial_18_comp_count[11], _05132_, max_pool_serial_18_comp_count[10], _05131_ }), .Y(_09422_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33384_ ( .A({ max_pool_serial_18_comp_count[9], _05161_, max_pool_serial_18_comp_count[8], _05160_ }), .Y(_09423_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _33385_ ( .A({ _09425_, _09422_, _09426_ }), .Y(_09424_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33386_ ( .A({ max_pool_serial_18_comp_count[10], max_pool_serial_18_comp_count[11], _05131_, _05132_ }), .Y(_09425_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33387_ ( .A({ max_pool_serial_18_comp_count[8], max_pool_serial_18_comp_count[9], _05160_, _05161_ }), .Y(_09426_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33388_ ( .A({ max_pool_serial_18_comp_count[6], _05158_, max_pool_serial_18_comp_count[7], _05159_ }), .Y(_09427_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _33389_ ( .A({ _09429_, _09430_, _09431_ }), .Y(_09428_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33390_ ( .A({ max_pool_serial_18_comp_count[14], max_pool_serial_18_comp_count[15], _05135_, _05136_ }), .Y(_09429_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33391_ ( .A({ max_pool_serial_18_comp_count[15], _05136_, max_pool_serial_18_comp_count[14], _05135_ }), .Y(_09430_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33392_ ( .A({ max_pool_serial_18_comp_count[12], max_pool_serial_18_comp_count[13], _05133_, _05134_ }), .Y(_09431_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33393_ ( .A({ max_pool_serial_18_comp_count[13], _05134_, max_pool_serial_18_comp_count[12], _05133_ }), .Y(_09432_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _33394_ ( .A({ _09441_, _09434_, _09435_, _09443_ }), .Y(_09433_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33395_ ( .A({ _09440_, _09439_, _09435_ }), .Y(_09434_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _33396_ ( .A({ _09438_, _09436_, _05142_, max_pool_serial_18_comp_count[20] }), .Y(_09435_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _33397_ ( .A({ _09437_, max_pool_serial_18_comp_count[22], _05144_ }), .Y(_09436_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _33398_ ( .A({ max_pool_serial_18_comp_count[23], _05145_, _05143_, max_pool_serial_18_comp_count[21] }), .Y(_09437_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33399_ ( .A({ max_pool_serial_18_comp_count[20], _05142_, max_pool_serial_18_comp_count[21], _05143_ }), .Y(_09438_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33400_ ( .A({ max_pool_serial_18_comp_count[19], _05140_, max_pool_serial_18_comp_count[18], _05139_ }), .Y(_09439_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33401_ ( .A({ max_pool_serial_18_comp_count[16], max_pool_serial_18_comp_count[17], _05137_, _05138_ }), .Y(_09440_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _33402_ ( .A({ _09442_, _09436_, _09438_ }), .Y(_09441_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33403_ ( .A({ max_pool_serial_18_comp_count[22], max_pool_serial_18_comp_count[23], _05144_, _05145_ }), .Y(_09442_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33404_ ( .A({ max_pool_serial_18_comp_count[18], max_pool_serial_18_comp_count[19], _05139_, _05140_ }), .Y(_09443_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33405_ ( .A({ _09445_, _09439_, _09435_ }), .Y(_09444_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33406_ ( .A({ max_pool_serial_18_comp_count[17], _05138_, max_pool_serial_18_comp_count[16], _05137_ }), .Y(_09445_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33407_ ( .A({ _09450_, _09447_ }), .Y(_09446_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33408_ ( .A({ _09449_, _09448_ }), .Y(_09447_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33409_ ( .A({ max_pool_serial_18_comp_count[31], _05154_, max_pool_serial_18_comp_count[30], _05153_ }), .Y(_09448_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33410_ ( .A({ max_pool_serial_18_comp_count[29], _05151_, max_pool_serial_18_comp_count[28], _05150_ }), .Y(_09449_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33411_ ( .A({ max_pool_serial_18_comp_count[27], _05149_, max_pool_serial_18_comp_count[26], _05148_ }), .Y(_09450_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33412_ ( .A({ max_pool_serial_18_comp_count[25], _05147_, max_pool_serial_18_comp_count[24], _05146_ }), .Y(_09451_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _33413_ ( .A({ _09456_, _09453_, _09447_, _09455_ }), .Y(_09452_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _33414_ ( .A({ _09448_, max_pool_serial_18_comp_count[29], _05151_, _09454_ }), .Y(_09453_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33415_ ( .A({ max_pool_serial_18_comp_count[28], _05150_ }), .Y(_09454_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33416_ ( .A({ max_pool_serial_18_comp_count[26], max_pool_serial_18_comp_count[27], _05148_, _05149_ }), .Y(_09455_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33417_ ( .A({ max_pool_serial_18_comp_count[30], max_pool_serial_18_comp_count[31], _05153_, _05154_ }), .Y(_09456_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33418_ ( .A({ max_pool_serial_18_comp_count[24], max_pool_serial_18_comp_count[25], _05146_, _05147_ }), .Y(_09457_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33419_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18446_, _18478_ }), .Y(_18414_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33420_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18520_, _18552_ }), .Y(_18488_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33421_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18626_, _18658_ }), .Y(_18594_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33422_ ( .A({ _20086_, _05996_, _09285_, _20152_ }), .Y(_20119_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _33423_ ( .A({ _09463_, _09458_ }), .Y(_06158_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33424_ ( .A({ _09462_, _09461_, _09460_, _09459_ }), .Y(_09458_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33425_ ( .A({ _05108_, _05107_, _05106_, _05105_ }), .Y(_09459_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33426_ ( .A({ _05104_, _05103_, _05102_, _05101_ }), .Y(_09460_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33427_ ( .A({ _05122_, _05121_, _05119_, _05118_ }), .Y(_09461_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33428_ ( .A({ _05116_, _05115_, _05113_, _05110_ }), .Y(_09462_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33429_ ( .A({ _05117_, _05114_, _05112_, _05111_ }), .Y(_09463_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33430_ ( .A({ _09464_, _09473_, _09470_, _maxi_write_rest_size[8] }), .Y(_06176_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33431_ ( .A({ _09469_, _09465_ }), .Y(_09464_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33432_ ( .A({ _09468_, _09466_, _maxi_write_rest_size[20:19] }), .Y(_09465_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33433_ ( .A({ _09467_, _maxi_write_rest_size[32:30] }), .Y(_09466_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33434_ ( .A({ _maxi_write_rest_size[28:27], _maxi_write_rest_size[25], _maxi_write_rest_size[22] }), .Y(_09467_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33435_ ( .A({ _maxi_write_rest_size[21], _maxi_write_rest_size[18:16] }), .Y(_09468_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33436_ ( .A({ _maxi_write_rest_size[29], _maxi_write_rest_size[26], _maxi_write_rest_size[24:23] }), .Y(_09469_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33437_ ( .A({ _09472_, _09471_ }), .Y(_09470_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33438_ ( .A(_maxi_write_rest_size[7:4]), .Y(_09471_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33439_ ( .A(_maxi_write_rest_size[3:0]), .Y(_09472_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33440_ ( .A({ _09474_, _maxi_write_rest_size[14], _maxi_write_rest_size[11:10] }), .Y(_09473_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33441_ ( .A({ _maxi_write_rest_size[15], _maxi_write_rest_size[13:12], _maxi_write_rest_size[9] }), .Y(_09474_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33442_ ( .A({ _05966_, _09475_ }), .Y(_24058_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33443_ ( .A({ _09476_, _09481_, _stream_conv2d_16_source_28_source_pat_fsm_11[0] }), .Y(_09475_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33444_ ( .A({ _09480_, _09479_, _09477_ }), .Y(_09476_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33445_ ( .A({ _09478_, _stream_conv2d_16_source_28_source_pat_fsm_11[3:2] }), .Y(_09477_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33446_ ( .A(_stream_conv2d_16_source_28_source_pat_fsm_11[7:4]), .Y(_09478_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33447_ ( .A(_stream_conv2d_16_source_28_source_pat_fsm_11[15:12]), .Y(_09479_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33448_ ( .A(_stream_conv2d_16_source_28_source_pat_fsm_11[11:8]), .Y(_09480_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33449_ ( .A({ _09485_, _09484_, _09483_, _09482_ }), .Y(_09481_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33450_ ( .A(_stream_conv2d_16_source_28_source_pat_fsm_11[23:20]), .Y(_09482_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33451_ ( .A(_stream_conv2d_16_source_28_source_pat_fsm_11[19:16]), .Y(_09483_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33452_ ( .A(_stream_conv2d_16_source_28_source_pat_fsm_11[31:28]), .Y(_09484_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33453_ ( .A(_stream_conv2d_16_source_28_source_pat_fsm_11[27:24]), .Y(_09485_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _33454_ ( .A({ _09476_, _stream_conv2d_16_source_28_source_pat_fsm_11[0], _09481_, _stream_conv2d_16_source_28_source_pat_fsm_11[1] }), .Y(_05966_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33455_ ( .A({ _18159_, _09486_, _18127_, _05966_ }), .Y(_18095_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33456_ ( .A({ _09475_, _stream_conv2d_16_source_28_source_pat_fsm_11[1] }), .Y(_09486_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33457_ ( .A({ _18170_, _09486_, _18138_, _05966_ }), .Y(_18106_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33458_ ( .A({ _18181_, _09486_, _18149_, _05966_ }), .Y(_18117_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33459_ ( .A({ _18184_, _09486_, _18152_, _05966_ }), .Y(_18120_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33460_ ( .A({ _18185_, _09486_, _18153_, _05966_ }), .Y(_18121_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33461_ ( .A({ _18186_, _09486_, _18154_, _05966_ }), .Y(_18122_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33462_ ( .A({ _18187_, _09486_, _18155_, _05966_ }), .Y(_18123_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33463_ ( .A({ _18188_, _09486_, _18156_, _05966_ }), .Y(_18124_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33464_ ( .A({ _18189_, _09486_, _18157_, _05966_ }), .Y(_18125_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33465_ ( .A({ _18190_, _09486_, _18158_, _05966_ }), .Y(_18126_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33466_ ( .A({ _18160_, _09486_, _18128_, _05966_ }), .Y(_18096_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33467_ ( .A({ _18161_, _09486_, _18129_, _05966_ }), .Y(_18097_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33468_ ( .A({ _18162_, _09486_, _18130_, _05966_ }), .Y(_18098_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33469_ ( .A({ _18163_, _09486_, _18131_, _05966_ }), .Y(_18099_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33470_ ( .A({ _18164_, _09486_, _18132_, _05966_ }), .Y(_18100_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33471_ ( .A({ _18165_, _09486_, _18133_, _05966_ }), .Y(_18101_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33472_ ( .A({ _18166_, _09486_, _18134_, _05966_ }), .Y(_18102_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33473_ ( .A({ _18167_, _09486_, _18135_, _05966_ }), .Y(_18103_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33474_ ( .A({ _18168_, _09486_, _18136_, _05966_ }), .Y(_18104_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33475_ ( .A({ _18169_, _09486_, _18137_, _05966_ }), .Y(_18105_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33476_ ( .A({ _18171_, _09486_, _18139_, _05966_ }), .Y(_18107_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33477_ ( .A({ _18172_, _09486_, _18140_, _05966_ }), .Y(_18108_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33478_ ( .A({ _18173_, _09486_, _18141_, _05966_ }), .Y(_18109_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33479_ ( .A({ _18174_, _09486_, _18142_, _05966_ }), .Y(_18110_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33480_ ( .A({ _18175_, _09486_, _18143_, _05966_ }), .Y(_18111_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33481_ ( .A({ _18176_, _09486_, _18144_, _05966_ }), .Y(_18112_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33482_ ( .A({ _18177_, _09486_, _18145_, _05966_ }), .Y(_18113_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33483_ ( .A({ _18178_, _09486_, _18146_, _05966_ }), .Y(_18114_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33484_ ( .A({ _18179_, _09486_, _18147_, _05966_ }), .Y(_18115_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33485_ ( .A({ _18180_, _09486_, _18148_, _05966_ }), .Y(_18116_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33486_ ( .A({ _18182_, _09486_, _18150_, _05966_ }), .Y(_18118_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33487_ ( .A({ _18183_, _09486_, _18151_, _05966_ }), .Y(_18119_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33488_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18445_, _18477_ }), .Y(_18413_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33489_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18519_, _18551_ }), .Y(_18487_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33490_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18625_, _18657_ }), .Y(_18593_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33491_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18324_, _18356_ }), .Y(_18292_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33492_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18347_, _18379_ }), .Y(_18315_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33493_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18444_, _18476_ }), .Y(_18412_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33494_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18518_, _18550_ }), .Y(_18486_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33495_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18624_, _18656_ }), .Y(_18592_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33496_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18346_, _18378_ }), .Y(_18314_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33497_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18323_, _18355_ }), .Y(_18291_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33498_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18443_, _18475_ }), .Y(_18411_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33499_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18517_, _18549_ }), .Y(_18485_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33500_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18623_, _18655_ }), .Y(_18591_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33501_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18322_, _18354_ }), .Y(_18290_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33502_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18345_, _18377_ }), .Y(_18313_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33503_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18442_, _18474_ }), .Y(_18410_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33504_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18516_, _18548_ }), .Y(_18484_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33505_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18622_, _18654_ }), .Y(_18590_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33506_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18441_, _18473_ }), .Y(_18409_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33507_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18515_, _18547_ }), .Y(_18483_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33508_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18621_, _18653_ }), .Y(_18589_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33509_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18440_, _18472_ }), .Y(_18408_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33510_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18514_, _18546_ }), .Y(_18482_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33511_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18620_, _18652_ }), .Y(_18588_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33512_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18437_, _18469_ }), .Y(_18405_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33513_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18513_, _18545_ }), .Y(_18481_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33514_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18619_, _18651_ }), .Y(_18587_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33515_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18512_, _18544_ }), .Y(_18480_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33516_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18617_, _18649_ }), .Y(_18585_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33517_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18616_, _18648_ }), .Y(_18584_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33518_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18615_, _18647_ }), .Y(_18583_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33519_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18614_, _18646_ }), .Y(_18582_) );
  \$lut  #( .LUT(16'h0bff), .WIDTH(4) ) _33520_ ( .A({ _09491_, _09487_, cparam_conv2d_16_max_col_count[4], conv2d_16_col_count[4] }), .Y(_06156_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _33521_ ( .A({ _09490_, cparam_conv2d_16_max_col_count[3], conv2d_16_col_count[3], _09488_ }), .Y(_09487_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _33522_ ( .A({ cparam_conv2d_16_max_col_count[2], conv2d_16_col_count[2], _09489_ }), .Y(_09488_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33523_ ( .A({ cparam_conv2d_16_max_col_count[0], cparam_conv2d_16_max_col_count[1], conv2d_16_col_count[0], conv2d_16_col_count[1] }), .Y(_09489_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33524_ ( .A({ conv2d_16_col_count[4], cparam_conv2d_16_max_col_count[4] }), .Y(_09490_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33525_ ( .A({ _09499_, _09498_, _09497_, _09492_ }), .Y(_09491_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33526_ ( .A({ _09496_, _09495_, _09494_, _09493_ }), .Y(_09492_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33527_ ( .A({ conv2d_16_col_count[14:13], conv2d_16_col_count[11:10] }), .Y(_09493_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33528_ ( .A({ conv2d_16_col_count[9:8], conv2d_16_col_count[6:5] }), .Y(_09494_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33529_ ( .A(conv2d_16_col_count[23:20]), .Y(_09495_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33530_ ( .A(conv2d_16_col_count[18:15]), .Y(_09496_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _33531_ ( .A({ conv2d_16_col_count[31:30], conv2d_16_col_count[28] }), .Y(_09497_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33532_ ( .A({ conv2d_16_col_count[24], conv2d_16_col_count[19], conv2d_16_col_count[12], conv2d_16_col_count[7] }), .Y(_09498_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33533_ ( .A({ conv2d_16_col_count[29], conv2d_16_col_count[27:25] }), .Y(_09499_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _33534_ ( .A({ _09505_, _09500_ }), .Y(_06157_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33535_ ( .A({ _09504_, _09503_, _09502_, _09501_ }), .Y(_09500_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33536_ ( .A({ _05048_, _05047_, _05046_, _05045_ }), .Y(_09501_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33537_ ( .A({ _05043_, _05042_, _05041_, _05040_ }), .Y(_09502_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33538_ ( .A({ _05057_, _05056_, _05054_, _05053_ }), .Y(_09503_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33539_ ( .A({ _05052_, _05051_, _05050_, _05049_ }), .Y(_09504_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33540_ ( .A({ _09509_, _09508_, _09507_, _09506_ }), .Y(_09505_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _33541_ ( .A({ _05058_, _05055_, _05044_, _05033_ }), .Y(_09506_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33542_ ( .A({ _05062_, _05061_, _05060_, _05059_ }), .Y(_09507_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33543_ ( .A({ _05039_, _05038_, _05037_, _05036_ }), .Y(_09508_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33544_ ( .A({ _05035_, _05034_, _05064_, _05063_ }), .Y(_09509_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33545_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18426_, _18458_ }), .Y(_18394_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33546_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18542_, _18574_ }), .Y(_18510_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33547_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18613_, _18645_ }), .Y(_18581_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33548_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18415_, _18447_ }), .Y(_18383_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33549_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18541_, _18573_ }), .Y(_18509_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33550_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18612_, _18644_ }), .Y(_18580_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33551_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18540_, _18572_ }), .Y(_18508_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _33552_ ( .A({ _09515_, _09510_ }), .Y(_06155_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33553_ ( .A({ _09514_, _09513_, _09512_, _09511_ }), .Y(_09510_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33554_ ( .A({ _05013_, _05011_, _05010_, _05009_ }), .Y(_09511_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33555_ ( .A({ _05008_, _05007_, _05006_, _05005_ }), .Y(_09512_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33556_ ( .A({ _05004_, _05025_, _05024_, _05022_ }), .Y(_09513_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33557_ ( .A({ _05020_, _05019_, _05017_, _05014_ }), .Y(_09514_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33558_ ( .A({ _05021_, _05018_, _05016_, _05015_ }), .Y(_09515_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33559_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18611_, _18643_ }), .Y(_18579_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _33560_ ( .A({ _09516_, _09525_, _09522_, _maxi_read_rest_size[8] }), .Y(_06175_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33561_ ( .A({ _09521_, _09517_ }), .Y(_09516_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33562_ ( .A({ _09520_, _09518_, _maxi_read_rest_size[20:19] }), .Y(_09517_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33563_ ( .A({ _09519_, _maxi_read_rest_size[32:30] }), .Y(_09518_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33564_ ( .A({ _maxi_read_rest_size[28:27], _maxi_read_rest_size[25], _maxi_read_rest_size[22] }), .Y(_09519_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33565_ ( .A({ _maxi_read_rest_size[21], _maxi_read_rest_size[18:16] }), .Y(_09520_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33566_ ( .A({ _maxi_read_rest_size[29], _maxi_read_rest_size[26], _maxi_read_rest_size[24:23] }), .Y(_09521_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33567_ ( .A({ _09524_, _09523_ }), .Y(_09522_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33568_ ( .A(_maxi_read_rest_size[7:4]), .Y(_09523_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33569_ ( .A(_maxi_read_rest_size[3:0]), .Y(_09524_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33570_ ( .A({ _09526_, _maxi_read_rest_size[14], _maxi_read_rest_size[11:10] }), .Y(_09525_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33571_ ( .A({ _maxi_read_rest_size[15], _maxi_read_rest_size[13:12], _maxi_read_rest_size[9] }), .Y(_09526_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33572_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18539_, _18571_ }), .Y(_18507_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33573_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18610_, _18642_ }), .Y(_18578_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33574_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18538_, _18570_ }), .Y(_18506_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33575_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18609_, _18641_ }), .Y(_18577_) );
  \$lut  #( .LUT(16'hf4ff), .WIDTH(4) ) _33576_ ( .A({ _09531_, _09527_, conv2d_16_row_count[4], cparam_conv2d_16_max_col_count[4] }), .Y(conv2d_16_update_filter) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _33577_ ( .A({ _09530_, conv2d_16_row_count[3], cparam_conv2d_16_max_col_count[3], _09528_ }), .Y(_09527_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _33578_ ( .A({ conv2d_16_row_count[2], cparam_conv2d_16_max_col_count[2], _09529_ }), .Y(_09528_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33579_ ( .A({ cparam_conv2d_16_max_col_count[0], cparam_conv2d_16_max_col_count[1], conv2d_16_row_count[0], conv2d_16_row_count[1] }), .Y(_09529_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33580_ ( .A({ cparam_conv2d_16_max_col_count[4], conv2d_16_row_count[4] }), .Y(_09530_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33581_ ( .A({ _09540_, _09539_, _09536_, _09532_ }), .Y(_09531_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33582_ ( .A({ _09535_, _09534_, _09533_ }), .Y(_09532_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _33583_ ( .A({ conv2d_16_row_count[30], conv2d_16_row_count[28], conv2d_16_row_count[22] }), .Y(_09533_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33584_ ( .A({ conv2d_16_row_count[20], conv2d_16_row_count[18], conv2d_16_row_count[16], conv2d_16_row_count[14] }), .Y(_09534_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33585_ ( .A({ conv2d_16_row_count[12], conv2d_16_row_count[10], conv2d_16_row_count[8], conv2d_16_row_count[6] }), .Y(_09535_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33586_ ( .A({ _09538_, _09537_ }), .Y(_09536_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33587_ ( .A({ conv2d_16_row_count[21], conv2d_16_row_count[19], conv2d_16_row_count[17], conv2d_16_row_count[15] }), .Y(_09537_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33588_ ( .A({ conv2d_16_row_count[13], conv2d_16_row_count[11], conv2d_16_row_count[9], conv2d_16_row_count[7] }), .Y(_09538_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33589_ ( .A({ conv2d_16_row_count[5], conv2d_16_row_count[31], conv2d_16_row_count[29], conv2d_16_row_count[27] }), .Y(_09539_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33590_ ( .A(conv2d_16_row_count[26:23]), .Y(_09540_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33591_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18537_, _18569_ }), .Y(_18505_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33592_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18608_, _18640_ }), .Y(_18576_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33593_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18433_, _18465_ }), .Y(_18401_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33594_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18638_, _18670_ }), .Y(_18606_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33595_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18637_, _18669_ }), .Y(_18605_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33596_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18636_, _18668_ }), .Y(_18604_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _33597_ ( .A({ _09546_, _09541_ }), .Y(_06154_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33598_ ( .A({ _09545_, _09544_, _09543_, _09542_ }), .Y(_09541_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33599_ ( .A({ _04855_, _04854_, _04853_, _04852_ }), .Y(_09542_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33600_ ( .A({ _04850_, _04849_, _04848_, _04847_ }), .Y(_09543_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33601_ ( .A({ _04864_, _04863_, _04861_, _04860_ }), .Y(_09544_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33602_ ( .A({ _04859_, _04858_, _04857_, _04856_ }), .Y(_09545_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33603_ ( .A({ _09550_, _09549_, _09548_, _09547_ }), .Y(_09546_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _33604_ ( .A({ _04865_, _04862_, _04851_, _04840_ }), .Y(_09547_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33605_ ( .A({ _04869_, _04868_, _04867_, _04866_ }), .Y(_09548_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33606_ ( .A({ _04846_, _04845_, _04844_, _04843_ }), .Y(_09549_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33607_ ( .A({ _04842_, _04841_, _04871_, _04870_ }), .Y(_09550_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33608_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18635_, _18667_ }), .Y(_18603_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _33609_ ( .A({ _09559_, _09563_, _09552_, _09562_ }), .Y(_09551_) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _33610_ ( .A({ conv2d_16_sync_comp_count[5], _09553_, _09558_, _04771_ }), .Y(_09552_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _33611_ ( .A({ _09554_, _09556_, _09555_, _09557_ }), .Y(_09553_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33612_ ( .A({ conv2d_16_sync_comp_count[3], _04769_, conv2d_16_sync_comp_count[4], _04770_ }), .Y(_09554_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _33613_ ( .A({ _04744_, conv2d_16_sync_comp_count[0], conv2d_16_sync_comp_count[1], _04755_ }), .Y(_09555_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _33614_ ( .A({ conv2d_16_sync_comp_count[2], _04766_, _04769_, conv2d_16_sync_comp_count[3] }), .Y(_09556_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _33615_ ( .A({ conv2d_16_sync_comp_count[2], _04766_, _04769_, conv2d_16_sync_comp_count[3] }), .Y(_09557_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33616_ ( .A({ _04770_, conv2d_16_sync_comp_count[4] }), .Y(_09558_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _33617_ ( .A({ _09561_, _09560_, _04773_, conv2d_16_sync_comp_count[7] }), .Y(_09559_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33618_ ( .A({ conv2d_16_sync_comp_count[11], _04746_, conv2d_16_sync_comp_count[10], _04745_ }), .Y(_09560_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33619_ ( .A({ conv2d_16_sync_comp_count[9], _04775_, conv2d_16_sync_comp_count[8], _04774_ }), .Y(_09561_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33620_ ( .A({ _04772_, conv2d_16_sync_comp_count[6] }), .Y(_09562_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33621_ ( .A({ conv2d_16_sync_comp_count[6], _04772_, conv2d_16_sync_comp_count[7], _04773_ }), .Y(_09563_) );
  \$lut  #( .LUT(16'h0071), .WIDTH(4) ) _33622_ ( .A({ _09565_, _04746_, conv2d_16_sync_comp_count[11], _09567_ }), .Y(_09564_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _33623_ ( .A({ _09560_, conv2d_16_sync_comp_count[9], _04775_, _09566_ }), .Y(_09565_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33624_ ( .A({ conv2d_16_sync_comp_count[8], _04774_ }), .Y(_09566_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33625_ ( .A({ conv2d_16_sync_comp_count[10], _04745_ }), .Y(_09567_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33626_ ( .A({ conv2d_16_sync_comp_count[15], _04750_, conv2d_16_sync_comp_count[14], _04749_ }), .Y(_09568_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33627_ ( .A({ conv2d_16_sync_comp_count[13], _04748_, conv2d_16_sync_comp_count[12], _04747_ }), .Y(_09569_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33628_ ( .A({ conv2d_16_sync_comp_count[12], conv2d_16_sync_comp_count[13], _04747_, _04748_ }), .Y(_09570_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33629_ ( .A({ conv2d_16_sync_comp_count[14], conv2d_16_sync_comp_count[15], _04749_, _04750_ }), .Y(_09571_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33630_ ( .A({ _09579_, _09573_ }), .Y(_09572_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33631_ ( .A({ _09578_, _09574_ }), .Y(_09573_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _33632_ ( .A({ _09577_, _09575_, _04756_, conv2d_16_sync_comp_count[20] }), .Y(_09574_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _33633_ ( .A({ _09576_, _04757_, conv2d_16_sync_comp_count[21] }), .Y(_09575_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33634_ ( .A({ conv2d_16_sync_comp_count[23], _04759_, conv2d_16_sync_comp_count[22], _04758_ }), .Y(_09576_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33635_ ( .A({ conv2d_16_sync_comp_count[20], _04756_, conv2d_16_sync_comp_count[21], _04757_ }), .Y(_09577_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33636_ ( .A({ conv2d_16_sync_comp_count[19], _04754_, conv2d_16_sync_comp_count[18], _04753_ }), .Y(_09578_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33637_ ( .A({ conv2d_16_sync_comp_count[17], _04752_, conv2d_16_sync_comp_count[16], _04751_ }), .Y(_09579_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _33638_ ( .A({ _09583_, _09581_, _09573_, _09585_ }), .Y(_09580_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33639_ ( .A({ _09582_, _09574_ }), .Y(_09581_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33640_ ( .A({ conv2d_16_sync_comp_count[18], conv2d_16_sync_comp_count[19], _04753_, _04754_ }), .Y(_09582_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _33641_ ( .A({ _09584_, _09575_, _09577_ }), .Y(_09583_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33642_ ( .A({ conv2d_16_sync_comp_count[22], conv2d_16_sync_comp_count[23], _04758_, _04759_ }), .Y(_09584_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33643_ ( .A({ conv2d_16_sync_comp_count[16], conv2d_16_sync_comp_count[17], _04751_, _04752_ }), .Y(_09585_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33644_ ( .A({ _09591_, _09590_, _09587_ }), .Y(_09586_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33645_ ( .A({ _09589_, _09588_ }), .Y(_09587_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33646_ ( .A({ conv2d_16_sync_comp_count[31], _04768_, conv2d_16_sync_comp_count[30], _04767_ }), .Y(_09588_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33647_ ( .A({ conv2d_16_sync_comp_count[29], _04765_, conv2d_16_sync_comp_count[28], _04764_ }), .Y(_09589_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33648_ ( .A({ conv2d_16_sync_comp_count[25], _04761_, conv2d_16_sync_comp_count[24], _04760_ }), .Y(_09590_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33649_ ( .A({ conv2d_16_sync_comp_count[27], _04763_, conv2d_16_sync_comp_count[26], _04762_ }), .Y(_09591_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _33650_ ( .A({ _09597_, _09593_, _09588_, _09596_ }), .Y(_09592_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _33651_ ( .A({ _09587_, _09594_, _09595_, _09591_ }), .Y(_09593_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33652_ ( .A({ conv2d_16_sync_comp_count[26], conv2d_16_sync_comp_count[27], _04762_, _04763_ }), .Y(_09594_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33653_ ( .A({ conv2d_16_sync_comp_count[24], conv2d_16_sync_comp_count[25], _04760_, _04761_ }), .Y(_09595_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33654_ ( .A({ conv2d_16_sync_comp_count[28], conv2d_16_sync_comp_count[29], _04764_, _04765_ }), .Y(_09596_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33655_ ( .A({ conv2d_16_sync_comp_count[30], conv2d_16_sync_comp_count[31], _04767_, _04768_ }), .Y(_09597_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33656_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18634_, _18666_ }), .Y(_18602_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33657_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18633_, _18665_ }), .Y(_18601_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33658_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18632_, _18664_ }), .Y(_18600_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _33659_ ( .A({ _09633_, _09643_, _09628_, _09598_ }), .Y(_06152_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _33660_ ( .A({ _09615_, _09625_, _09622_, _09599_ }), .Y(_09598_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _33661_ ( .A({ _09614_, _09609_, _09600_, _09612_ }), .Y(_09599_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _33662_ ( .A({ _09608_, _24016_, _counter_count_782[6], _09601_ }), .Y(_09600_) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _33663_ ( .A({ _counter_count_782[5], _09602_, _09607_, _24015_ }), .Y(_09601_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _33664_ ( .A({ _09606_, _09605_, _09604_, _09603_ }), .Y(_09602_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33665_ ( .A({ _23988_, _counter_count_782[0], _23999_, _counter_count_782[1] }), .Y(_09603_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33666_ ( .A({ _counter_count_782[1], _23999_, _counter_count_782[2], _24010_ }), .Y(_09604_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33667_ ( .A({ _24010_, _counter_count_782[2], _24013_, _counter_count_782[3] }), .Y(_09605_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33668_ ( .A({ _counter_count_782[3], _24013_, _counter_count_782[4], _24014_ }), .Y(_09606_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33669_ ( .A({ _24014_, _counter_count_782[4] }), .Y(_09607_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33670_ ( .A({ _counter_count_782[7], _24017_ }), .Y(_09608_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _33671_ ( .A({ _09610_, _counter_count_782[9], _24019_, _09611_ }), .Y(_09609_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33672_ ( .A({ _counter_count_782[11], _23990_, _counter_count_782[10], _23989_ }), .Y(_09610_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33673_ ( .A({ _counter_count_782[8], _24018_ }), .Y(_09611_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _33674_ ( .A({ _09613_, _09610_, _24017_, _counter_count_782[7] }), .Y(_09612_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33675_ ( .A({ _counter_count_782[9], _24019_, _counter_count_782[8], _24018_ }), .Y(_09613_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33676_ ( .A({ _counter_count_782[10], _counter_count_782[11], _23989_, _23990_ }), .Y(_09614_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33677_ ( .A({ _09621_, _09620_, _09616_ }), .Y(_09615_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _33678_ ( .A({ _09619_, _09617_, _24000_, _counter_count_782[20] }), .Y(_09616_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _33679_ ( .A({ _09618_, _24001_, _counter_count_782[21] }), .Y(_09617_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33680_ ( .A({ _counter_count_782[23], _24003_, _counter_count_782[22], _24002_ }), .Y(_09618_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33681_ ( .A({ _counter_count_782[20], _24000_, _counter_count_782[21], _24001_ }), .Y(_09619_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33682_ ( .A({ _counter_count_782[17], _23996_, _counter_count_782[16], _23995_ }), .Y(_09620_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33683_ ( .A({ _counter_count_782[19], _23998_, _counter_count_782[18], _23997_ }), .Y(_09621_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33684_ ( .A({ _09624_, _09623_ }), .Y(_09622_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33685_ ( .A({ _counter_count_782[15], _23994_, _counter_count_782[14], _23993_ }), .Y(_09623_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33686_ ( .A({ _counter_count_782[13], _23992_, _counter_count_782[12], _23991_ }), .Y(_09624_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _33687_ ( .A({ _09626_, _09623_, _09627_ }), .Y(_09625_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33688_ ( .A({ _counter_count_782[14], _counter_count_782[15], _23993_, _23994_ }), .Y(_09626_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33689_ ( .A({ _counter_count_782[12], _counter_count_782[13], _23991_, _23992_ }), .Y(_09627_) );
  \$lut  #( .LUT(16'h000b), .WIDTH(4) ) _33690_ ( .A({ _09632_, _09629_, _09617_, _09619_ }), .Y(_09628_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _33691_ ( .A({ _09616_, _09630_, _09631_, _09621_ }), .Y(_09629_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33692_ ( .A({ _counter_count_782[18], _counter_count_782[19], _23997_, _23998_ }), .Y(_09630_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33693_ ( .A({ _counter_count_782[16], _counter_count_782[17], _23995_, _23996_ }), .Y(_09631_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33694_ ( .A({ _counter_count_782[22], _counter_count_782[23], _24002_, _24003_ }), .Y(_09632_) );
  \$lut  #( .LUT(16'h000b), .WIDTH(4) ) _33695_ ( .A({ _09642_, _09634_, _09636_, _09638_ }), .Y(_09633_) );
  \$lut  #( .LUT(16'h8f00), .WIDTH(4) ) _33696_ ( .A({ _09635_, _09641_, _09640_, _09639_ }), .Y(_09634_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _33697_ ( .A({ _09638_, _09636_, _24008_, _counter_count_782[28] }), .Y(_09635_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _33698_ ( .A({ _09637_, _24009_, _counter_count_782[29] }), .Y(_09636_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33699_ ( .A({ _counter_count_782[31], _24012_, _counter_count_782[30], _24011_ }), .Y(_09637_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33700_ ( .A({ _counter_count_782[28], _24008_, _counter_count_782[29], _24009_ }), .Y(_09638_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33701_ ( .A({ _counter_count_782[27], _24007_, _counter_count_782[26], _24006_ }), .Y(_09639_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33702_ ( .A({ _counter_count_782[24], _counter_count_782[25], _24004_, _24005_ }), .Y(_09640_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33703_ ( .A({ _counter_count_782[26], _counter_count_782[27], _24006_, _24007_ }), .Y(_09641_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33704_ ( .A({ _counter_count_782[30], _counter_count_782[31], _24011_, _24012_ }), .Y(_09642_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33705_ ( .A({ _09644_, _09639_, _09635_ }), .Y(_09643_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33706_ ( .A({ _counter_count_782[25], _24005_, _counter_count_782[24], _24004_ }), .Y(_09644_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33707_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18629_, _18661_ }), .Y(_18597_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33708_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18618_, _18650_ }), .Y(_18586_) );
  \$lut  #( .LUT(16'h7100), .WIDTH(4) ) _33709_ ( .A({ _09651_, _pulse_count_213[8], _23986_, _13087_ }), .Y(_06151_) );
  \$lut  #( .LUT(16'h5701), .WIDTH(4) ) _33710_ ( .A({ _pulse_count_213[5], _09646_, _09650_, _23983_ }), .Y(_09645_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _33711_ ( .A({ _09649_, _23981_, _pulse_count_213[3], _09647_ }), .Y(_09646_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _33712_ ( .A({ _23978_, _pulse_count_213[2], _09648_ }), .Y(_09647_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _33713_ ( .A({ _23956_, _pulse_count_213[0], _pulse_count_213[1], _23967_ }), .Y(_09648_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33714_ ( .A({ _pulse_count_213[4], _23982_ }), .Y(_09649_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33715_ ( .A({ _23982_, _pulse_count_213[4] }), .Y(_09650_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33716_ ( .A({ _09654_, _09652_ }), .Y(_09651_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _33717_ ( .A({ _09653_, _23979_, _23971_, _23969_ }), .Y(_09652_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33718_ ( .A({ _23962_, _23960_, _23987_, _23974_ }), .Y(_09653_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33719_ ( .A({ _09658_, _09657_, _09656_, _09655_ }), .Y(_09654_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33720_ ( .A({ _23972_, _23970_, _23968_, _23965_ }), .Y(_09655_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33721_ ( .A({ _23963_, _23961_, _23959_, _23957_ }), .Y(_09656_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33722_ ( .A({ _23964_, _23958_, _23977_, _23976_ }), .Y(_09657_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33723_ ( .A({ _23980_, _23975_, _23973_, _23966_ }), .Y(_09658_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33724_ ( .A({ _20273_, _09285_, _20209_, maxi_rready }), .Y(_20241_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33725_ ( .A({ _maxi_read_fsm[0], _09659_, _09274_ }), .Y(maxi_rready) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _33726_ ( .A({ _09284_, _maxi_read_fsm[1], _maxi_read_fsm[2], _maxi_read_fsm[3] }), .Y(_09659_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _33727_ ( .A({ _09651_, _09660_, _reducemax_count_211[8], _23986_ }), .Y(_06150_) );
  \$lut  #( .LUT(16'hbbb0), .WIDTH(4) ) _33728_ ( .A({ _09669_, _09661_, _reducemax_count_211[8], _23986_ }), .Y(_09660_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _33729_ ( .A({ _09668_, _23984_, _reducemax_count_211[6], _09662_ }), .Y(_09661_) );
  \$lut  #( .LUT(8'h71), .WIDTH(3) ) _33730_ ( .A({ _23983_, _reducemax_count_211[5], _09663_ }), .Y(_09662_) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _33731_ ( .A({ _23982_, _09664_, _09667_, _reducemax_count_211[4] }), .Y(_09663_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _33732_ ( .A({ _09666_, _reducemax_count_211[2], _23978_, _09665_ }), .Y(_09664_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33733_ ( .A({ _23956_, _23967_, _reducemax_count_211[0], _reducemax_count_211[1] }), .Y(_09665_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33734_ ( .A({ _23981_, _reducemax_count_211[3] }), .Y(_09666_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33735_ ( .A({ _reducemax_count_211[3], _23981_ }), .Y(_09667_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33736_ ( .A({ _reducemax_count_211[7], _23985_ }), .Y(_09668_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33737_ ( .A({ _23985_, _reducemax_count_211[7] }), .Y(_09669_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33738_ ( .A({ _20272_, _09285_, _20208_, maxi_rready }), .Y(_20240_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33739_ ( .A({ _20270_, _09285_, _20206_, maxi_rready }), .Y(_20238_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33740_ ( .A({ _20269_, _09285_, _20205_, maxi_rready }), .Y(_20237_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33741_ ( .A({ _20268_, _09285_, _20204_, maxi_rready }), .Y(_20236_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33742_ ( .A({ _20267_, _09285_, _20203_, maxi_rready }), .Y(_20235_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33743_ ( .A({ _05991_, _09298_ }), .Y(_24071_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33744_ ( .A({ _20266_, _09285_, _20202_, maxi_rready }), .Y(_20234_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33745_ ( .A({ _20265_, _09285_, _20201_, maxi_rready }), .Y(_20233_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33746_ ( .A({ _20264_, _09285_, _20200_, maxi_rready }), .Y(_20232_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33747_ ( .A({ _20263_, _09285_, _20199_, maxi_rready }), .Y(_20231_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33748_ ( .A({ _20262_, _09285_, _20198_, maxi_rready }), .Y(_20230_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33749_ ( .A({ _20261_, _09285_, _20197_, maxi_rready }), .Y(_20229_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33750_ ( .A({ _09670_, _19850_, _09298_ }), .Y(_19882_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33751_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[6], _05991_ }), .Y(_09670_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33752_ ( .A({ _20259_, _09285_, _20195_, maxi_rready }), .Y(_20227_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33753_ ( .A({ _09670_, _19849_, _09298_ }), .Y(_19881_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33754_ ( .A({ _20258_, _09285_, _20194_, maxi_rready }), .Y(_20226_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33755_ ( .A({ _09670_, _19847_, _09298_ }), .Y(_19879_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33756_ ( .A({ _20257_, _09285_, _20193_, maxi_rready }), .Y(_20225_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33757_ ( .A({ _09670_, _19846_, _09298_ }), .Y(_19878_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33758_ ( .A({ _20256_, _09285_, _20192_, maxi_rready }), .Y(_20224_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33759_ ( .A({ _09670_, _19845_, _09298_ }), .Y(_19877_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33760_ ( .A({ _20255_, _09285_, _20191_, maxi_rready }), .Y(_20223_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33761_ ( .A({ _09670_, _19844_, _09298_ }), .Y(_19876_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33762_ ( .A({ _20254_, _09285_, _20190_, maxi_rready }), .Y(_20222_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33763_ ( .A({ _09670_, _19843_, _09298_ }), .Y(_19875_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33764_ ( .A({ _20253_, _09285_, _20189_, maxi_rready }), .Y(_20221_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33765_ ( .A({ _09670_, _19842_, _09298_ }), .Y(_19874_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33766_ ( .A({ _20252_, _09285_, _20188_, maxi_rready }), .Y(_20220_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33767_ ( .A({ _09670_, _19841_, _09298_ }), .Y(_19873_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33768_ ( .A({ _20251_, _09285_, _20187_, maxi_rready }), .Y(_20219_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33769_ ( .A({ _09670_, _19840_, _09298_ }), .Y(_19872_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33770_ ( .A({ _20250_, _09285_, _20186_, maxi_rready }), .Y(_20218_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33771_ ( .A({ _09670_, _19839_, _09298_ }), .Y(_19871_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33772_ ( .A({ _20280_, _09285_, _20216_, maxi_rready }), .Y(_20248_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33773_ ( .A({ _09670_, _19838_, _09298_ }), .Y(_19870_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33774_ ( .A({ _20279_, _09285_, _20215_, maxi_rready }), .Y(_20247_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33775_ ( .A({ _09670_, _19836_, _09298_ }), .Y(_19868_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33776_ ( .A({ _20278_, _09285_, _20214_, maxi_rready }), .Y(_20246_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33777_ ( .A({ _09670_, _19835_, _09298_ }), .Y(_19867_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33778_ ( .A({ _20277_, _09285_, _20213_, maxi_rready }), .Y(_20245_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33779_ ( .A({ _09670_, _19834_, _09298_ }), .Y(_19866_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33780_ ( .A({ _20276_, _09285_, _20212_, maxi_rready }), .Y(_20244_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33781_ ( .A({ _09670_, _19832_, _09298_ }), .Y(_19864_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33782_ ( .A({ _20275_, _09285_, _20211_, maxi_rready }), .Y(_20243_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _33783_ ( .A({ _09711_, _09671_, _pulse_count_19[32], _23948_ }), .Y(_06148_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _33784_ ( .A({ _09704_, _13091_, _09702_, _09672_ }), .Y(_09671_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _33785_ ( .A({ _09690_, _09686_, _09692_, _09673_ }), .Y(_09672_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _33786_ ( .A({ _09681_, _09685_, _09674_, _09684_ }), .Y(_09673_) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _33787_ ( .A({ _pulse_count_19[5], _09675_, _09680_, _23951_ }), .Y(_09674_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _33788_ ( .A({ _09679_, _09678_, _09676_, _09677_ }), .Y(_09675_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _33789_ ( .A({ _23923_, _pulse_count_19[0], _pulse_count_19[1], _23934_ }), .Y(_09676_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _33790_ ( .A({ _pulse_count_19[2], _23945_, _23949_, _pulse_count_19[3] }), .Y(_09677_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33791_ ( .A({ _pulse_count_19[4], _23950_ }), .Y(_09678_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33792_ ( .A({ _pulse_count_19[2], _pulse_count_19[3], _23945_, _23949_ }), .Y(_09679_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33793_ ( .A({ _23950_, _pulse_count_19[4] }), .Y(_09680_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _33794_ ( .A({ _09683_, _09682_, _23953_, _pulse_count_19[7] }), .Y(_09681_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33795_ ( .A({ _pulse_count_19[11], _23925_, _pulse_count_19[10], _23924_ }), .Y(_09682_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33796_ ( .A({ _pulse_count_19[9], _23955_, _pulse_count_19[8], _23954_ }), .Y(_09683_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33797_ ( .A({ _23952_, _pulse_count_19[6] }), .Y(_09684_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33798_ ( .A({ _pulse_count_19[6], _23952_, _pulse_count_19[7], _23953_ }), .Y(_09685_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _33799_ ( .A({ _09687_, _23926_, _pulse_count_19[12] }), .Y(_09686_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _33800_ ( .A({ _09688_, _23927_, _pulse_count_19[13] }), .Y(_09687_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33801_ ( .A({ _pulse_count_19[15], _23929_, _pulse_count_19[14], _23928_ }), .Y(_09688_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33802_ ( .A({ _pulse_count_19[12], _23926_, _pulse_count_19[13], _23927_ }), .Y(_09689_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _33803_ ( .A({ _09691_, _09687_, _09689_ }), .Y(_09690_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33804_ ( .A({ _pulse_count_19[14], _pulse_count_19[15], _23928_, _23929_ }), .Y(_09691_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _33805_ ( .A({ _09694_, _09682_, _09693_ }), .Y(_09692_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33806_ ( .A({ _pulse_count_19[8], _pulse_count_19[9], _23954_, _23955_ }), .Y(_09693_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33807_ ( .A({ _pulse_count_19[10], _pulse_count_19[11], _23924_, _23925_ }), .Y(_09694_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _33808_ ( .A({ _09698_, _09696_, _23935_, _pulse_count_19[20] }), .Y(_09695_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _33809_ ( .A({ _09697_, _pulse_count_19[22], _23937_ }), .Y(_09696_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _33810_ ( .A({ _pulse_count_19[23], _23938_, _23936_, _pulse_count_19[21] }), .Y(_09697_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33811_ ( .A({ _pulse_count_19[20], _23935_, _pulse_count_19[21], _23936_ }), .Y(_09698_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33812_ ( .A({ _pulse_count_19[19], _23933_, _pulse_count_19[18], _23932_ }), .Y(_09699_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33813_ ( .A({ _pulse_count_19[16], _pulse_count_19[17], _23930_, _23931_ }), .Y(_09700_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33814_ ( .A({ _pulse_count_19[22], _pulse_count_19[23], _23937_, _23938_ }), .Y(_09701_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33815_ ( .A({ _09703_, _09699_, _09695_ }), .Y(_09702_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33816_ ( .A({ _pulse_count_19[17], _23931_, _pulse_count_19[16], _23930_ }), .Y(_09703_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33817_ ( .A({ _09710_, _09705_ }), .Y(_09704_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33818_ ( .A({ _09709_, _09706_ }), .Y(_09705_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33819_ ( .A({ _09708_, _09707_ }), .Y(_09706_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33820_ ( .A({ _pulse_count_19[31], _23947_, _pulse_count_19[30], _23946_ }), .Y(_09707_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33821_ ( .A({ _pulse_count_19[29], _23944_, _pulse_count_19[28], _23943_ }), .Y(_09708_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33822_ ( .A({ _pulse_count_19[27], _23942_, _pulse_count_19[26], _23941_ }), .Y(_09709_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33823_ ( .A({ _pulse_count_19[25], _23940_, _pulse_count_19[24], _23939_ }), .Y(_09710_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _33824_ ( .A({ _09712_, _09705_, _09717_ }), .Y(_09711_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _33825_ ( .A({ _09716_, _09713_, _09706_, _09715_ }), .Y(_09712_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _33826_ ( .A({ _09707_, _pulse_count_19[29], _23944_, _09714_ }), .Y(_09713_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33827_ ( .A({ _pulse_count_19[28], _23943_ }), .Y(_09714_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33828_ ( .A({ _pulse_count_19[26], _pulse_count_19[27], _23941_, _23942_ }), .Y(_09715_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _33829_ ( .A({ _pulse_count_19[30], _pulse_count_19[31], _23946_, _23947_ }), .Y(_09716_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33830_ ( .A({ _pulse_count_19[24], _pulse_count_19[25], _23939_, _23940_ }), .Y(_09717_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33831_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18325_, _18357_ }), .Y(_18293_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33832_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18348_, _18380_ }), .Y(_18316_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _33833_ ( .A({ _09735_, _09751_, _09748_, _09719_ }), .Y(_09718_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _33834_ ( .A({ _09731_, _09728_, _09734_, _09720_ }), .Y(_09719_) );
  \$lut  #( .LUT(16'h00f4), .WIDTH(4) ) _33835_ ( .A({ _09725_, _09726_, _09727_, _09721_ }), .Y(_09720_) );
  \$lut  #( .LUT(16'h00b2), .WIDTH(4) ) _33836_ ( .A({ _09724_, _23949_, _reduceadd_count_17[3], _09722_ }), .Y(_09721_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _33837_ ( .A({ _23945_, _reduceadd_count_17[2], _09723_ }), .Y(_09722_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _33838_ ( .A({ _23923_, _23934_, _reduceadd_count_17[0], _reduceadd_count_17[1] }), .Y(_09723_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33839_ ( .A({ _reduceadd_count_17[4], _23950_ }), .Y(_09724_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33840_ ( .A({ _23952_, _reduceadd_count_17[6] }), .Y(_09725_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33841_ ( .A({ _reduceadd_count_17[5], _23951_ }), .Y(_09726_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33842_ ( .A({ _23950_, _reduceadd_count_17[4], _23951_, _reduceadd_count_17[5] }), .Y(_09727_) );
  \$lut  #( .LUT(16'h9000), .WIDTH(4) ) _33843_ ( .A({ _09730_, _09729_, _23955_, _reduceadd_count_17[9] }), .Y(_09728_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33844_ ( .A({ _23925_, _reduceadd_count_17[11], _23924_, _reduceadd_count_17[10] }), .Y(_09729_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _33845_ ( .A({ _23954_, _reduceadd_count_17[8], _23953_, _reduceadd_count_17[7] }), .Y(_09730_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _33846_ ( .A({ _09733_, _09729_, _09732_ }), .Y(_09731_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _33847_ ( .A({ _reduceadd_count_17[8], _23954_, _23955_, _reduceadd_count_17[9] }), .Y(_09732_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _33848_ ( .A({ _reduceadd_count_17[10], _23924_, _23925_, _reduceadd_count_17[11] }), .Y(_09733_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _33849_ ( .A({ _reduceadd_count_17[6], _23952_, _reduceadd_count_17[7], _23953_ }), .Y(_09734_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33850_ ( .A({ _09745_, _09742_, _09739_, _09736_ }), .Y(_09735_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _33851_ ( .A({ _09737_, _23930_, _reduceadd_count_17[16] }), .Y(_09736_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _33852_ ( .A({ _09738_, _23931_, _reduceadd_count_17[17] }), .Y(_09737_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33853_ ( .A({ _23933_, _reduceadd_count_17[19], _23932_, _reduceadd_count_17[18] }), .Y(_09738_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33854_ ( .A({ _09741_, _09740_ }), .Y(_09739_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33855_ ( .A({ _23947_, _reduceadd_count_17[31], _23946_, _reduceadd_count_17[30] }), .Y(_09740_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33856_ ( .A({ _23944_, _reduceadd_count_17[29], _23943_, _reduceadd_count_17[28] }), .Y(_09741_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33857_ ( .A({ _09744_, _09743_ }), .Y(_09742_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33858_ ( .A({ _23942_, _reduceadd_count_17[27], _23941_, _reduceadd_count_17[26] }), .Y(_09743_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33859_ ( .A({ _23940_, _reduceadd_count_17[25], _23939_, _reduceadd_count_17[24] }), .Y(_09744_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33860_ ( .A({ _09747_, _09746_ }), .Y(_09745_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33861_ ( .A({ _23938_, _reduceadd_count_17[23], _23937_, _reduceadd_count_17[22] }), .Y(_09746_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33862_ ( .A({ _23936_, _reduceadd_count_17[21], _23935_, _reduceadd_count_17[20] }), .Y(_09747_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33863_ ( .A({ _09750_, _09749_ }), .Y(_09748_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33864_ ( .A({ _23929_, _reduceadd_count_17[15], _23928_, _reduceadd_count_17[14] }), .Y(_09749_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _33865_ ( .A({ _23927_, _reduceadd_count_17[13], _23926_, _reduceadd_count_17[12] }), .Y(_09750_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _33866_ ( .A({ _09752_, _09749_, _09753_ }), .Y(_09751_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _33867_ ( .A({ _reduceadd_count_17[14], _23928_, _23929_, _reduceadd_count_17[15] }), .Y(_09752_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _33868_ ( .A({ _reduceadd_count_17[12], _23926_, _23927_, _reduceadd_count_17[13] }), .Y(_09753_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _33869_ ( .A({ _09739_, _09762_, _09742_, _09755_ }), .Y(_09754_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _33870_ ( .A({ _09761_, _09759_, _09756_, _09745_ }), .Y(_09755_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _33871_ ( .A({ _23933_, _reduceadd_count_17[19], _09757_ }), .Y(_09756_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _33872_ ( .A({ _23932_, _reduceadd_count_17[18], _09758_ }), .Y(_09757_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _33873_ ( .A({ _reduceadd_count_17[16], _23930_, _23931_, _reduceadd_count_17[17] }), .Y(_09758_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _33874_ ( .A({ _09746_, _reduceadd_count_17[21], _23936_, _09760_ }), .Y(_09759_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33875_ ( .A({ _reduceadd_count_17[20], _23935_ }), .Y(_09760_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _33876_ ( .A({ _reduceadd_count_17[22], _23937_, _23938_, _reduceadd_count_17[23] }), .Y(_09761_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _33877_ ( .A({ _09764_, _09743_, _09763_ }), .Y(_09762_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _33878_ ( .A({ _reduceadd_count_17[24], _23939_, _23940_, _reduceadd_count_17[25] }), .Y(_09763_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _33879_ ( .A({ _reduceadd_count_17[26], _23941_, _23942_, _reduceadd_count_17[27] }), .Y(_09764_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _33880_ ( .A({ _09740_, _reduceadd_count_17[29], _23944_, _09766_ }), .Y(_09765_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33881_ ( .A({ _reduceadd_count_17[28], _23943_ }), .Y(_09766_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _33882_ ( .A({ _reduceadd_count_17[30], _23946_, _23947_, _reduceadd_count_17[31] }), .Y(_09767_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33883_ ( .A({ _09670_, _19831_, _09298_ }), .Y(_19863_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33884_ ( .A({ _20274_, _09285_, _20210_, maxi_rready }), .Y(_20242_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33885_ ( .A({ _09670_, _19830_, _09298_ }), .Y(_19862_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33886_ ( .A({ _09670_, _19829_, _09298_ }), .Y(_19861_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33887_ ( .A({ _09670_, _19828_, _09298_ }), .Y(_19860_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33888_ ( .A({ _09670_, _19827_, _09298_ }), .Y(_19859_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33889_ ( .A({ _09670_, _19857_, _09298_ }), .Y(_19889_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33890_ ( .A({ _09670_, _19856_, _09298_ }), .Y(_19888_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33891_ ( .A({ _09670_, _19855_, _09298_ }), .Y(_19887_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33892_ ( .A({ _09670_, _19854_, _09298_ }), .Y(_19886_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33893_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[5], _05991_, _09298_, _19853_ }), .Y(_19885_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33894_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[4], _05991_, _09298_, _19852_ }), .Y(_19884_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33895_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[2], _05991_, _09298_, _19848_ }), .Y(_19880_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33896_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[3], _05991_, _09298_, _19851_ }), .Y(_19883_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33897_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[1], _05991_, _09298_, _19837_ }), .Y(_19869_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33898_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[0], _05991_, _09298_, _19826_ }), .Y(_19858_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33899_ ( .A({ _20271_, _09285_, _20207_, maxi_rready }), .Y(_20239_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33900_ ( .A({ _20260_, _09285_, _20196_, maxi_rready }), .Y(_20228_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _33901_ ( .A({ _20249_, _09285_, _20185_, maxi_rready }), .Y(_20217_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _33902_ ( .A({ maxi_rready, _09285_ }), .Y(_24072_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33903_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19013_, _19045_ }), .Y(_18981_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33904_ ( .A({ _09769_, _09777_, _stream_conv2d_16_source_19_source_pat_fsm_2[1] }), .Y(_09768_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33905_ ( .A({ _09776_, _09775_, _09770_ }), .Y(_09769_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33906_ ( .A({ _09774_, _09773_, _09772_, _09771_ }), .Y(_09770_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33907_ ( .A(_stream_conv2d_16_source_19_source_pat_fsm_2[23:20]), .Y(_09771_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33908_ ( .A(_stream_conv2d_16_source_19_source_pat_fsm_2[19:16]), .Y(_09772_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33909_ ( .A(_stream_conv2d_16_source_19_source_pat_fsm_2[31:28]), .Y(_09773_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33910_ ( .A(_stream_conv2d_16_source_19_source_pat_fsm_2[27:24]), .Y(_09774_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33911_ ( .A(_stream_conv2d_16_source_19_source_pat_fsm_2[15:12]), .Y(_09775_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33912_ ( .A(_stream_conv2d_16_source_19_source_pat_fsm_2[11:8]), .Y(_09776_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33913_ ( .A({ _09778_, _stream_conv2d_16_source_19_source_pat_fsm_2[3:2] }), .Y(_09777_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33914_ ( .A(_stream_conv2d_16_source_19_source_pat_fsm_2[7:4]), .Y(_09778_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33915_ ( .A({ _19199_, _05987_, _09790_, _19231_ }), .Y(_19167_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _33916_ ( .A({ _stream_conv2d_16_source_6_source_pat_fsm_0[0], _09788_, _09779_ }), .Y(_05987_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33917_ ( .A({ _09780_, _stream_conv2d_16_source_6_source_pat_fsm_0[1] }), .Y(_09779_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33918_ ( .A({ _09787_, _09786_, _09781_ }), .Y(_09780_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33919_ ( .A({ _09785_, _09784_, _09783_, _09782_ }), .Y(_09781_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33920_ ( .A(_stream_conv2d_16_source_6_source_pat_fsm_0[23:20]), .Y(_09782_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33921_ ( .A(_stream_conv2d_16_source_6_source_pat_fsm_0[19:16]), .Y(_09783_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33922_ ( .A(_stream_conv2d_16_source_6_source_pat_fsm_0[31:28]), .Y(_09784_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33923_ ( .A(_stream_conv2d_16_source_6_source_pat_fsm_0[27:24]), .Y(_09785_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33924_ ( .A(_stream_conv2d_16_source_6_source_pat_fsm_0[15:12]), .Y(_09786_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33925_ ( .A(_stream_conv2d_16_source_6_source_pat_fsm_0[11:8]), .Y(_09787_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33926_ ( .A({ _09789_, _stream_conv2d_16_source_6_source_pat_fsm_0[3:2] }), .Y(_09788_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33927_ ( .A(_stream_conv2d_16_source_6_source_pat_fsm_0[7:4]), .Y(_09789_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _33928_ ( .A({ _09791_, _09779_ }), .Y(_09790_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33929_ ( .A({ _09788_, _stream_conv2d_16_source_6_source_pat_fsm_0[0] }), .Y(_09791_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33930_ ( .A({ _09670_, _19447_, _09298_ }), .Y(_19479_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33931_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19012_, _19044_ }), .Y(_18980_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33932_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19006_, _19038_ }), .Y(_18974_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33933_ ( .A({ _09670_, _19652_, _09298_ }), .Y(_19684_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33934_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19005_, _19037_ }), .Y(_18973_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33935_ ( .A({ _09670_, _19651_, _09298_ }), .Y(_19683_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33936_ ( .A({ _19207_, _05987_, _09790_, _19239_ }), .Y(_19175_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33937_ ( .A({ _19191_, _05987_, _09790_, _19223_ }), .Y(_19159_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33938_ ( .A({ _19209_, _05987_, _09790_, _19241_ }), .Y(_19177_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33939_ ( .A({ _09670_, _19459_, _09298_ }), .Y(_19491_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _33940_ ( .A({ _09792_, _19271_, _09298_ }), .Y(_19303_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _33941_ ( .A({ _19367_, _05727_, _09303_, _19335_ }), .Y(_09792_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33942_ ( .A({ _09670_, _19443_, _09298_ }), .Y(_19475_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _33943_ ( .A({ _09793_, _19326_, _09303_ }), .Y(_19294_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _33944_ ( .A({ _19262_, _09298_, _19358_, _05727_ }), .Y(_09793_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33945_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[4], _05991_, _19466_, _09298_ }), .Y(_19498_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33946_ ( .A({ _09670_, _19833_, _09298_ }), .Y(_19865_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33947_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _18997_, _19029_ }), .Y(_18965_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33948_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19017_, _19049_ }), .Y(_18985_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33949_ ( .A({ _19202_, _05987_, _09790_, _19234_ }), .Y(_19170_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33950_ ( .A({ _19187_, _05987_, _09790_, _19219_ }), .Y(_19155_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _33951_ ( .A({ _19194_, _05987_, _09790_, _19226_ }), .Y(_19162_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _33952_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19108_, _19140_ }), .Y(_19076_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33953_ ( .A({ _09795_, _09803_, _stream_conv2d_16_source_8_source_pat_fsm_1[1] }), .Y(_09794_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33954_ ( .A({ _09802_, _09801_, _09796_ }), .Y(_09795_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33955_ ( .A({ _09800_, _09799_, _09798_, _09797_ }), .Y(_09796_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33956_ ( .A(_stream_conv2d_16_source_8_source_pat_fsm_1[23:20]), .Y(_09797_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33957_ ( .A(_stream_conv2d_16_source_8_source_pat_fsm_1[19:16]), .Y(_09798_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33958_ ( .A(_stream_conv2d_16_source_8_source_pat_fsm_1[31:28]), .Y(_09799_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33959_ ( .A(_stream_conv2d_16_source_8_source_pat_fsm_1[27:24]), .Y(_09800_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33960_ ( .A(_stream_conv2d_16_source_8_source_pat_fsm_1[15:12]), .Y(_09801_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33961_ ( .A(_stream_conv2d_16_source_8_source_pat_fsm_1[11:8]), .Y(_09802_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33962_ ( .A({ _09804_, _stream_conv2d_16_source_8_source_pat_fsm_1[3:2] }), .Y(_09803_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33963_ ( .A(_stream_conv2d_16_source_8_source_pat_fsm_1[7:4]), .Y(_09804_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33964_ ( .A({ _09670_, _19453_, _09298_ }), .Y(_19485_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33965_ ( .A({ _09670_, _19444_, _09298_ }), .Y(_19476_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _33966_ ( .A({ _09670_, _19469_, _09298_ }), .Y(_19501_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _33967_ ( .A({ _05965_, _09805_ }), .Y(_24057_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _33968_ ( .A({ _09806_, _09811_, _stream_conv2d_16_source_29_source_pat_fsm_12[0] }), .Y(_09805_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _33969_ ( .A({ _09810_, _09809_, _09807_ }), .Y(_09806_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _33970_ ( .A({ _09808_, _stream_conv2d_16_source_29_source_pat_fsm_12[3:2] }), .Y(_09807_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33971_ ( .A(_stream_conv2d_16_source_29_source_pat_fsm_12[7:4]), .Y(_09808_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33972_ ( .A(_stream_conv2d_16_source_29_source_pat_fsm_12[15:12]), .Y(_09809_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33973_ ( .A(_stream_conv2d_16_source_29_source_pat_fsm_12[11:8]), .Y(_09810_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _33974_ ( .A({ _09815_, _09814_, _09813_, _09812_ }), .Y(_09811_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33975_ ( .A(_stream_conv2d_16_source_29_source_pat_fsm_12[23:20]), .Y(_09812_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33976_ ( .A(_stream_conv2d_16_source_29_source_pat_fsm_12[19:16]), .Y(_09813_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33977_ ( .A(_stream_conv2d_16_source_29_source_pat_fsm_12[31:28]), .Y(_09814_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _33978_ ( .A(_stream_conv2d_16_source_29_source_pat_fsm_12[27:24]), .Y(_09815_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _33979_ ( .A({ _09806_, _stream_conv2d_16_source_29_source_pat_fsm_12[0], _09811_, _stream_conv2d_16_source_29_source_pat_fsm_12[1] }), .Y(_05965_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33980_ ( .A({ _18063_, _09816_, _18031_, _05965_ }), .Y(_17999_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _33981_ ( .A({ _09805_, _stream_conv2d_16_source_29_source_pat_fsm_12[1] }), .Y(_09816_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33982_ ( .A({ _18074_, _09816_, _18042_, _05965_ }), .Y(_18010_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33983_ ( .A({ _18085_, _09816_, _18053_, _05965_ }), .Y(_18021_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33984_ ( .A({ _18088_, _09816_, _18056_, _05965_ }), .Y(_18024_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33985_ ( .A({ _18089_, _09816_, _18057_, _05965_ }), .Y(_18025_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33986_ ( .A({ _18090_, _09816_, _18058_, _05965_ }), .Y(_18026_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33987_ ( .A({ _18091_, _09816_, _18059_, _05965_ }), .Y(_18027_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33988_ ( .A({ _18092_, _09816_, _18060_, _05965_ }), .Y(_18028_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33989_ ( .A({ _18093_, _09816_, _18061_, _05965_ }), .Y(_18029_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33990_ ( .A({ _18094_, _09816_, _18062_, _05965_ }), .Y(_18030_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33991_ ( .A({ _18064_, _09816_, _18032_, _05965_ }), .Y(_18000_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33992_ ( .A({ _18065_, _09816_, _18033_, _05965_ }), .Y(_18001_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33993_ ( .A({ _18066_, _09816_, _18034_, _05965_ }), .Y(_18002_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33994_ ( .A({ _18067_, _09816_, _18035_, _05965_ }), .Y(_18003_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33995_ ( .A({ _18068_, _09816_, _18036_, _05965_ }), .Y(_18004_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33996_ ( .A({ _18069_, _09816_, _18037_, _05965_ }), .Y(_18005_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33997_ ( .A({ _18070_, _09816_, _18038_, _05965_ }), .Y(_18006_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33998_ ( .A({ _18071_, _09816_, _18039_, _05965_ }), .Y(_18007_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _33999_ ( .A({ _18072_, _09816_, _18040_, _05965_ }), .Y(_18008_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34000_ ( .A({ _18073_, _09816_, _18041_, _05965_ }), .Y(_18009_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34001_ ( .A({ _18075_, _09816_, _18043_, _05965_ }), .Y(_18011_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34002_ ( .A({ _18076_, _09816_, _18044_, _05965_ }), .Y(_18012_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34003_ ( .A({ _18077_, _09816_, _18045_, _05965_ }), .Y(_18013_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34004_ ( .A({ _18078_, _09816_, _18046_, _05965_ }), .Y(_18014_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34005_ ( .A({ _18079_, _09816_, _18047_, _05965_ }), .Y(_18015_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34006_ ( .A({ _18080_, _09816_, _18048_, _05965_ }), .Y(_18016_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34007_ ( .A({ _18081_, _09816_, _18049_, _05965_ }), .Y(_18017_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34008_ ( .A({ _18082_, _09816_, _18050_, _05965_ }), .Y(_18018_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34009_ ( .A({ _18083_, _09816_, _18051_, _05965_ }), .Y(_18019_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34010_ ( .A({ _18084_, _09816_, _18052_, _05965_ }), .Y(_18020_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34011_ ( .A({ _18086_, _09816_, _18054_, _05965_ }), .Y(_18022_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34012_ ( .A({ _18087_, _09816_, _18055_, _05965_ }), .Y(_18023_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34013_ ( .A({ _05960_, _09817_ }), .Y(_24056_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34014_ ( .A({ _09826_, _09823_, _09818_ }), .Y(_09817_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34015_ ( .A({ _09822_, _09821_, _09820_, _09819_ }), .Y(_09818_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34016_ ( .A(_stream_conv2d_16_source_30_source_pat_fsm_13[23:20]), .Y(_09819_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34017_ ( .A(_stream_conv2d_16_source_30_source_pat_fsm_13[19:16]), .Y(_09820_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34018_ ( .A(_stream_conv2d_16_source_30_source_pat_fsm_13[31:28]), .Y(_09821_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34019_ ( .A(_stream_conv2d_16_source_30_source_pat_fsm_13[27:24]), .Y(_09822_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34020_ ( .A({ _09825_, _09824_ }), .Y(_09823_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34021_ ( .A(_stream_conv2d_16_source_30_source_pat_fsm_13[15:12]), .Y(_09824_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34022_ ( .A(_stream_conv2d_16_source_30_source_pat_fsm_13[11:8]), .Y(_09825_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34023_ ( .A({ _09827_, _stream_conv2d_16_source_30_source_pat_fsm_13[3:2], _stream_conv2d_16_source_30_source_pat_fsm_13[0] }), .Y(_09826_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34024_ ( .A(_stream_conv2d_16_source_30_source_pat_fsm_13[7:4]), .Y(_09827_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _34025_ ( .A({ _09828_, _09827_, _09823_, _09818_ }), .Y(_05960_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34026_ ( .A({ _stream_conv2d_16_source_30_source_pat_fsm_13[0], _stream_conv2d_16_source_30_source_pat_fsm_13[3:1] }), .Y(_09828_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34027_ ( .A({ _17967_, _09829_, _17935_, _05960_ }), .Y(_17903_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34028_ ( .A({ _09817_, _stream_conv2d_16_source_30_source_pat_fsm_13[1] }), .Y(_09829_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34029_ ( .A({ _17978_, _09829_, _17946_, _05960_ }), .Y(_17914_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34030_ ( .A({ _17989_, _09829_, _17957_, _05960_ }), .Y(_17925_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34031_ ( .A({ _17992_, _09829_, _17960_, _05960_ }), .Y(_17928_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34032_ ( .A({ _17993_, _09829_, _17961_, _05960_ }), .Y(_17929_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34033_ ( .A({ _17994_, _09829_, _17962_, _05960_ }), .Y(_17930_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34034_ ( .A({ _17995_, _09829_, _17963_, _05960_ }), .Y(_17931_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34035_ ( .A({ _17996_, _09829_, _17964_, _05960_ }), .Y(_17932_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34036_ ( .A({ _17997_, _09829_, _17965_, _05960_ }), .Y(_17933_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34037_ ( .A({ _17998_, _09829_, _17966_, _05960_ }), .Y(_17934_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34038_ ( .A({ _17968_, _09829_, _17936_, _05960_ }), .Y(_17904_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34039_ ( .A({ _17969_, _09829_, _17937_, _05960_ }), .Y(_17905_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34040_ ( .A({ _17970_, _09829_, _17938_, _05960_ }), .Y(_17906_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34041_ ( .A({ _17971_, _09829_, _17939_, _05960_ }), .Y(_17907_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34042_ ( .A({ _17972_, _09829_, _17940_, _05960_ }), .Y(_17908_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34043_ ( .A({ _17973_, _09829_, _17941_, _05960_ }), .Y(_17909_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34044_ ( .A({ _17974_, _09829_, _17942_, _05960_ }), .Y(_17910_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34045_ ( .A({ _17975_, _09829_, _17943_, _05960_ }), .Y(_17911_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34046_ ( .A({ _17976_, _09829_, _17944_, _05960_ }), .Y(_17912_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34047_ ( .A({ _17977_, _09829_, _17945_, _05960_ }), .Y(_17913_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34048_ ( .A({ _17979_, _09829_, _17947_, _05960_ }), .Y(_17915_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34049_ ( .A({ _17980_, _09829_, _17948_, _05960_ }), .Y(_17916_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34050_ ( .A({ _17981_, _09829_, _17949_, _05960_ }), .Y(_17917_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34051_ ( .A({ _17982_, _09829_, _17950_, _05960_ }), .Y(_17918_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34052_ ( .A({ _17983_, _09829_, _17951_, _05960_ }), .Y(_17919_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34053_ ( .A({ _17984_, _09829_, _17952_, _05960_ }), .Y(_17920_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34054_ ( .A({ _17985_, _09829_, _17953_, _05960_ }), .Y(_17921_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34055_ ( .A({ _17986_, _09829_, _17954_, _05960_ }), .Y(_17922_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34056_ ( .A({ _17987_, _09829_, _17955_, _05960_ }), .Y(_17923_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34057_ ( .A({ _17988_, _09829_, _17956_, _05960_ }), .Y(_17924_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34058_ ( .A({ _17990_, _09829_, _17958_, _05960_ }), .Y(_17926_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34059_ ( .A({ _17991_, _09829_, _17959_, _05960_ }), .Y(_17927_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34060_ ( .A({ _09835_, _09830_ }), .Y(matmul_29_dma_out_mask_0) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34061_ ( .A({ _09834_, _09833_, _09832_, _09831_ }), .Y(_09830_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34062_ ( .A(matmul_29_out_row_count[23:20]), .Y(_09831_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34063_ ( .A(matmul_29_out_row_count[19:16]), .Y(_09832_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34064_ ( .A(matmul_29_out_row_count[31:28]), .Y(_09833_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34065_ ( .A(matmul_29_out_row_count[27:24]), .Y(_09834_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34066_ ( .A({ _09839_, _09838_, _09837_, _09836_ }), .Y(_09835_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34067_ ( .A(matmul_29_out_row_count[7:4]), .Y(_09836_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34068_ ( .A(matmul_29_out_row_count[3:0]), .Y(_09837_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34069_ ( .A(matmul_29_out_row_count[15:12]), .Y(_09838_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34070_ ( .A(matmul_29_out_row_count[11:8]), .Y(_09839_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34071_ ( .A({ _09845_, _09840_ }), .Y(matmul_29_dma_pad_mask_0) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34072_ ( .A({ _09844_, _09843_, _09842_, _09841_ }), .Y(_09840_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34073_ ( .A(matmul_29_row_count[23:20]), .Y(_09841_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34074_ ( .A(matmul_29_row_count[19:16]), .Y(_09842_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34075_ ( .A(matmul_29_row_count[31:28]), .Y(_09843_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34076_ ( .A(matmul_29_row_count[27:24]), .Y(_09844_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34077_ ( .A({ _09849_, _09848_, _09847_, _09846_ }), .Y(_09845_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34078_ ( .A(matmul_29_row_count[7:4]), .Y(_09846_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34079_ ( .A(matmul_29_row_count[3:0]), .Y(_09847_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34080_ ( .A(matmul_29_row_count[15:12]), .Y(_09848_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34081_ ( .A(matmul_29_row_count[11:8]), .Y(_09849_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34082_ ( .A({ _09396_, _09857_, _09850_ }), .Y(max_pool_serial_18_dma_pad_mask_0) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _34083_ ( .A({ _09854_, max_pool_serial_18_row_count[3], cparam_max_pool_serial_18_act_num_col[3], _09851_ }), .Y(_09850_) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _34084_ ( .A({ cparam_max_pool_serial_18_act_num_col[2], _09852_, _09853_, max_pool_serial_18_row_count[2] }), .Y(_09851_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _34085_ ( .A({ cparam_max_pool_serial_18_act_num_col[0], max_pool_serial_18_row_count[0], cparam_max_pool_serial_18_act_num_col[1], max_pool_serial_18_row_count[1] }), .Y(_09852_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34086_ ( .A({ max_pool_serial_18_row_count[1], cparam_max_pool_serial_18_act_num_col[1] }), .Y(_09853_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34087_ ( .A({ _09856_, _09855_, max_pool_serial_18_row_count[7:6] }), .Y(_09854_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _34088_ ( .A({ max_pool_serial_18_row_count[4], cparam_max_pool_serial_18_act_num_col[4], max_pool_serial_18_row_count[5], cparam_max_pool_serial_18_act_num_col[5] }), .Y(_09855_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _34089_ ( .A({ cparam_max_pool_serial_18_act_num_col[4], max_pool_serial_18_row_count[4], cparam_max_pool_serial_18_act_num_col[5], max_pool_serial_18_row_count[5] }), .Y(_09856_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _34090_ ( .A({ _09855_, max_pool_serial_18_row_count[5], cparam_max_pool_serial_18_act_num_col[5] }), .Y(_09857_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _34091_ ( .A({ _03905_, cparam_max_pool_serial_18_act_num_col[3], _09859_ }), .Y(_09858_) );
  \$lut  #( .LUT(16'hddd4), .WIDTH(4) ) _34092_ ( .A({ _09861_, _09860_, _03902_, cparam_max_pool_serial_18_act_num_col[2] }), .Y(_09859_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34093_ ( .A({ _03891_, cparam_max_pool_serial_18_act_num_col[1] }), .Y(_09860_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _34094_ ( .A({ cparam_max_pool_serial_18_act_num_col[0], _03880_, cparam_max_pool_serial_18_act_num_col[1], _03891_ }), .Y(_09861_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _34095_ ( .A({ _03909_, _03908_ }), .Y(_09862_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34096_ ( .A({ _09868_, _09867_, _09866_, _09864_ }), .Y(_09863_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34097_ ( .A({ _09865_, _09862_, _03882_, _03910_ }), .Y(_09864_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34098_ ( .A({ _03890_, _03887_, _03885_, _03884_ }), .Y(_09865_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34099_ ( .A({ _03904_, _03903_, _03901_, _03900_ }), .Y(_09866_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34100_ ( .A({ _03899_, _03896_, _03894_, _03893_ }), .Y(_09867_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34101_ ( .A({ _03898_, _03897_, _03895_, _03892_ }), .Y(_09868_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34102_ ( .A({ _03889_, _03888_, _03886_, _03883_ }), .Y(_09869_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34103_ ( .A({ _09878_, _09877_, _09876_, _09871_ }), .Y(_09870_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34104_ ( .A({ _09875_, _09874_, _09873_, _09872_ }), .Y(_09871_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34105_ ( .A(conv2d_16_out_row_count[11:8]), .Y(_09872_) );
  \$lut  #( .LUT(16'h000b), .WIDTH(4) ) _34106_ ( .A({ conv2d_16_out_row_count[6], conv2d_16_out_row_count[7], conv2d_16_out_row_count[5], cparam_conv2d_16_act_num_row[5] }), .Y(_09873_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34107_ ( .A(conv2d_16_out_row_count[19:16]), .Y(_09874_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34108_ ( .A(conv2d_16_out_row_count[15:12]), .Y(_09875_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34109_ ( .A(conv2d_16_out_row_count[31:28]), .Y(_09876_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34110_ ( .A(conv2d_16_out_row_count[27:24]), .Y(_09877_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34111_ ( .A(conv2d_16_out_row_count[23:20]), .Y(_09878_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _34112_ ( .A({ cparam_conv2d_16_act_num_row[3], conv2d_16_out_row_count[3], cparam_conv2d_16_act_num_row[2], conv2d_16_out_row_count[2] }), .Y(_09879_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _34113_ ( .A({ conv2d_16_out_row_count[0], cparam_conv2d_16_act_num_row[0], cparam_conv2d_16_act_num_row[1], conv2d_16_out_row_count[1] }), .Y(_09880_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _34114_ ( .A({ cparam_conv2d_16_act_num_row[2], cparam_conv2d_16_act_num_row[3], conv2d_16_out_row_count[2], conv2d_16_out_row_count[3] }), .Y(_09881_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _34115_ ( .A({ cparam_conv2d_16_act_num_row[1], conv2d_16_out_row_count[1], cparam_conv2d_16_act_num_row[0], conv2d_16_out_row_count[0] }), .Y(_09882_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34116_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18725_, _18757_ }), .Y(_18693_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34117_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18424_, _18456_ }), .Y(_18392_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34118_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18714_, _18746_ }), .Y(_18682_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34119_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18919_, _18951_ }), .Y(_18887_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34120_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18703_, _18735_ }), .Y(_18671_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34121_ ( .A({ _09670_, _19461_, _09298_ }), .Y(_19493_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34122_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18914_, _18946_ }), .Y(_18882_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34123_ ( .A({ _09670_, _19458_, _09298_ }), .Y(_19490_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34124_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18913_, _18945_ }), .Y(_18881_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34125_ ( .A({ _20440_, _06930_, _07066_, _20472_ }), .Y(_05647_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34126_ ( .A({ _09670_, _19454_, _09298_ }), .Y(_19486_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34127_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18909_, _18941_ }), .Y(_18877_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34128_ ( .A({ _20438_, _06930_, _07066_, _20470_ }), .Y(_05648_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34129_ ( .A({ _09670_, _19452_, _09298_ }), .Y(_19484_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34130_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18908_, _18940_ }), .Y(_18876_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34131_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18535_, _18567_ }), .Y(_18503_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34132_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18423_, _18455_ }), .Y(_18391_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34133_ ( .A({ _20434_, _06930_, _07066_, _20466_ }), .Y(_05649_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34134_ ( .A({ _09670_, _19446_, _09298_ }), .Y(_19478_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34135_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18905_, _18937_ }), .Y(_18873_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34136_ ( .A({ _05976_, _07793_ }), .Y(_24064_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _34137_ ( .A({ _stream_conv2d_16_source_22_source_pat_fsm_5[1], _07794_, _07802_, _stream_conv2d_16_source_22_source_pat_fsm_5[0] }), .Y(_05976_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34138_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18534_, _18566_ }), .Y(_18502_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34139_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18422_, _18454_ }), .Y(_18390_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34140_ ( .A({ _20427_, _06930_, _07066_, _20459_ }), .Y(_05650_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34141_ ( .A({ _20426_, _06930_, _07066_, _20458_ }), .Y(_05651_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34142_ ( .A({ _20423_, _06930_, _07066_, _20455_ }), .Y(_05652_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34143_ ( .A({ _20421_, _06930_, _07066_, _20453_ }), .Y(_05653_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34144_ ( .A({ _20420_, _06930_, _07066_, _20452_ }), .Y(_05654_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34145_ ( .A({ _09670_, _19468_, _09298_ }), .Y(_19500_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34146_ ( .A({ _09883_, _19327_, _09303_ }), .Y(_19295_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34147_ ( .A({ _19263_, _09298_, _19359_, _05727_ }), .Y(_09883_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34148_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18900_, _18932_ }), .Y(_18868_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34149_ ( .A({ _20447_, _06930_, _07066_, _20479_ }), .Y(_05655_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34150_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[1], _05991_, _19451_, _09298_ }), .Y(_19483_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34151_ ( .A({ _09884_, _19321_, _09303_ }), .Y(_19289_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34152_ ( .A({ _19257_, _09298_, _19353_, _05727_ }), .Y(_09884_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34153_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18899_, _18931_ }), .Y(_18867_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34154_ ( .A({ _20446_, _06930_, _07066_, _20478_ }), .Y(_05656_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34155_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[0], _05991_, _19440_, _09298_ }), .Y(_19472_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34156_ ( .A({ _09885_, _19256_, _09298_ }), .Y(_19288_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34157_ ( .A({ _19352_, _05727_, _09303_, _19320_ }), .Y(_09885_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34158_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18897_, _18929_ }), .Y(_18865_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34159_ ( .A({ _20442_, _06930_, _07066_, _20474_ }), .Y(_05657_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34160_ ( .A({ _09886_, _19316_, _09303_ }), .Y(_19284_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34161_ ( .A({ _19252_, _09298_, _19348_, _05727_ }), .Y(_09886_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34162_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18926_, _18958_ }), .Y(_18894_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34163_ ( .A({ _09887_, _19312_, _09303_ }), .Y(_19280_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34164_ ( .A({ _19248_, _09298_, _19344_, _05727_ }), .Y(_09887_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34165_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18922_, _18954_ }), .Y(_18890_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34166_ ( .A({ _09888_, _19278_, _09298_ }), .Y(_19310_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34167_ ( .A({ _19374_, _05727_, _09303_, _19342_ }), .Y(_09888_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34168_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18921_, _18953_ }), .Y(_18889_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34169_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18532_, _18564_ }), .Y(_18500_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34170_ ( .A({ _09889_, _19274_, _09298_ }), .Y(_19306_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34171_ ( .A({ _19370_, _05727_, _09303_, _19338_ }), .Y(_09889_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34172_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18920_, _18952_ }), .Y(_18888_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34173_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18531_, _18563_ }), .Y(_18499_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34174_ ( .A({ _09890_, _05989_, _09305_ }), .Y(_19301_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _34175_ ( .A({ _09891_, _05727_, _19365_ }), .Y(_09890_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34176_ ( .A({ _19269_, _09298_, _09303_, _19333_ }), .Y(_09891_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34177_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18917_, _18949_ }), .Y(_18885_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34178_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18536_, _18568_ }), .Y(_18504_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34179_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19015_, _19047_ }), .Y(_18983_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34180_ ( .A({ _09371_, _stream_conv2d_16_source_23_source_pat_fsm_6[0], _18607_, _18639_ }), .Y(_18575_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34181_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18533_, _18565_ }), .Y(_18501_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34182_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19014_, _19046_ }), .Y(_18982_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34183_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18522_, _18554_ }), .Y(_18490_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34184_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19011_, _19043_ }), .Y(_18979_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34185_ ( .A({ _09252_, _stream_conv2d_16_source_24_source_pat_fsm_7[0], _18511_, _18543_ }), .Y(_18479_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34186_ ( .A({ _05970_, _09241_ }), .Y(_24061_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _34187_ ( .A({ _stream_conv2d_16_source_25_source_pat_fsm_8[1], _09242_, _09250_, _stream_conv2d_16_source_25_source_pat_fsm_8[0] }), .Y(_05970_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34188_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18439_, _18471_ }), .Y(_18407_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34189_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19010_, _19042_ }), .Y(_18978_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34190_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18823_, _18855_ }), .Y(_18791_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34191_ ( .A({ _09670_, _19658_, _09298_ }), .Y(_19690_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34192_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19009_, _19041_ }), .Y(_18977_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34193_ ( .A({ _09670_, _19657_, _09298_ }), .Y(_19689_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34194_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19008_, _19040_ }), .Y(_18976_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34195_ ( .A({ _09670_, _19655_, _09298_ }), .Y(_19687_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34196_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19007_, _19039_ }), .Y(_18975_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34197_ ( .A({ _09670_, _19654_, _09298_ }), .Y(_19686_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34198_ ( .A({ _09670_, _19653_, _09298_ }), .Y(_19685_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34199_ ( .A({ _09892_, _20369_, _09893_ }), .Y(_20305_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34200_ ( .A({ _20401_, _09285_, maxi_rready, _20337_ }), .Y(_09892_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34201_ ( .A({ _maxi_read_fsm[1], _09286_, _09275_, _maxi_read_fsm[0] }), .Y(_09893_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34202_ ( .A({ _09894_, _20368_, _09893_ }), .Y(_20304_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34203_ ( .A({ _20400_, _09285_, maxi_rready, _20336_ }), .Y(_09894_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34204_ ( .A({ _09895_, _20366_, _09893_ }), .Y(_20302_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34205_ ( .A({ _20398_, _09285_, maxi_rready, _20334_ }), .Y(_09895_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34206_ ( .A({ _09896_, _20365_, _09893_ }), .Y(_20301_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34207_ ( .A({ _20397_, _09285_, maxi_rready, _20333_ }), .Y(_09896_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34208_ ( .A({ _09897_, _20364_, _09893_ }), .Y(_20300_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34209_ ( .A({ _20396_, _09285_, maxi_rready, _20332_ }), .Y(_09897_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34210_ ( .A({ _09898_, _20395_, _09285_ }), .Y(_20299_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34211_ ( .A({ _20331_, maxi_rready, _09893_, _20363_ }), .Y(_09898_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34212_ ( .A({ _09899_, _20394_, _09285_ }), .Y(_20298_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34213_ ( .A({ _20330_, maxi_rready, _09893_, _20362_ }), .Y(_09899_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34214_ ( .A({ _09900_, _20361_, _09893_ }), .Y(_20297_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34215_ ( .A({ _20393_, _09285_, maxi_rready, _20329_ }), .Y(_09900_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34216_ ( .A({ _09901_, _20360_, _09893_ }), .Y(_20296_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34217_ ( .A({ _20392_, _09285_, maxi_rready, _20328_ }), .Y(_09901_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34218_ ( .A({ _09902_, _20359_, _09893_ }), .Y(_20295_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34219_ ( .A({ _20391_, _09285_, maxi_rready, _20327_ }), .Y(_09902_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34220_ ( .A({ _09903_, _20358_, _09893_ }), .Y(_20294_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34221_ ( .A({ _20390_, _09285_, maxi_rready, _20326_ }), .Y(_09903_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34222_ ( .A({ _09904_, _20357_, _09893_ }), .Y(_20293_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34223_ ( .A({ _20389_, _09285_, maxi_rready, _20325_ }), .Y(_09904_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34224_ ( .A({ _09905_, _20355_, _09893_ }), .Y(_20291_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34225_ ( .A({ _20387_, _09285_, maxi_rready, _20323_ }), .Y(_09905_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34226_ ( .A({ _09906_, _20354_, _09893_ }), .Y(_20290_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34227_ ( .A({ _20386_, _09285_, maxi_rready, _20322_ }), .Y(_09906_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34228_ ( .A({ _09907_, _20385_, _09285_ }), .Y(_20289_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34229_ ( .A({ _20321_, maxi_rready, _09893_, _20353_ }), .Y(_09907_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34230_ ( .A({ _09908_, _20384_, _09285_ }), .Y(_20288_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34231_ ( .A({ _20320_, maxi_rready, _09893_, _20352_ }), .Y(_09908_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34232_ ( .A({ _09909_, _20351_, _09893_ }), .Y(_20287_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34233_ ( .A({ _20383_, _09285_, maxi_rready, _20319_ }), .Y(_09909_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34234_ ( .A({ _09910_, _20350_, _09893_ }), .Y(_20286_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34235_ ( .A({ _20382_, _09285_, maxi_rready, _20318_ }), .Y(_09910_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34236_ ( .A({ _09911_, _20349_, _09893_ }), .Y(_20285_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34237_ ( .A({ _20381_, _09285_, maxi_rready, _20317_ }), .Y(_09911_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34238_ ( .A({ _09912_, _20348_, _09893_ }), .Y(_20284_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34239_ ( .A({ _20380_, _09285_, maxi_rready, _20316_ }), .Y(_09912_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34240_ ( .A({ _09913_, _20347_, _09893_ }), .Y(_20283_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34241_ ( .A({ _20379_, _09285_, maxi_rready, _20315_ }), .Y(_09913_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34242_ ( .A({ _09914_, _20346_, _09893_ }), .Y(_20282_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34243_ ( .A({ _20378_, _09285_, maxi_rready, _20314_ }), .Y(_09914_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34244_ ( .A({ _09915_, _20376_, _09893_ }), .Y(_20312_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34245_ ( .A({ _20408_, _09285_, maxi_rready, _20344_ }), .Y(_09915_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34246_ ( .A({ _09916_, _20407_, _09285_ }), .Y(_20311_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34247_ ( .A({ _20343_, maxi_rready, _09893_, _20375_ }), .Y(_09916_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34248_ ( .A({ _09917_, _20374_, _09893_ }), .Y(_20310_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34249_ ( .A({ _20406_, _09285_, maxi_rready, _20342_ }), .Y(_09917_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34250_ ( .A({ _09918_, _20373_, _09893_ }), .Y(_20309_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34251_ ( .A({ _20405_, _09285_, maxi_rready, _20341_ }), .Y(_09918_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34252_ ( .A({ _09919_, _20372_, _09893_ }), .Y(_20308_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34253_ ( .A({ _20404_, _09285_, maxi_rready, _20340_ }), .Y(_09919_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34254_ ( .A({ _09920_, _20371_, _09893_ }), .Y(_20307_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34255_ ( .A({ _20403_, _09285_, maxi_rready, _20339_ }), .Y(_09920_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34256_ ( .A({ _09921_, _20370_, _09893_ }), .Y(_20306_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34257_ ( .A({ _20402_, _09285_, maxi_rready, _20338_ }), .Y(_09921_) );
  \$lut  #( .LUT(16'hf8ff), .WIDTH(4) ) _34258_ ( .A({ _09922_, _09925_, _09285_, _20399_ }), .Y(_20303_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _34259_ ( .A({ _05994_, maxi_rready, _20335_ }), .Y(_09922_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34260_ ( .A({ _09923_, _maxi_read_fsm[0] }), .Y(_05994_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34261_ ( .A({ _09924_, _09274_ }), .Y(_09923_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34262_ ( .A({ _maxi_read_fsm[2], _09284_, _maxi_read_fsm[1], _maxi_read_fsm[3] }), .Y(_09924_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34263_ ( .A({ _20367_, _09893_ }), .Y(_09925_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34264_ ( .A({ _09926_, _20388_, _09285_ }), .Y(_20292_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _34265_ ( .A({ _09927_, _09893_, _20356_ }), .Y(_09926_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _34266_ ( .A({ _05996_, maxi_rready, _20324_ }), .Y(_09927_) );
  \$lut  #( .LUT(16'hf8ff), .WIDTH(4) ) _34267_ ( .A({ _09928_, _09929_, _09285_, _20377_ }), .Y(_20281_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _34268_ ( .A({ _05994_, maxi_rready, _20313_ }), .Y(_09928_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34269_ ( .A({ _20345_, _09893_ }), .Y(_09929_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34270_ ( .A({ _05996_, _09285_ }), .Y(_05658_) );
  \$lut  #( .LUT(16'hfeff), .WIDTH(4) ) _34271_ ( .A({ _05996_, _09923_, _09893_, _24072_ }), .Y(_24073_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34272_ ( .A({ _09670_, _19650_, _09298_ }), .Y(_19682_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34273_ ( .A({ _09670_, _19649_, _09298_ }), .Y(_19681_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34274_ ( .A({ _09670_, _19648_, _09298_ }), .Y(_19680_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34275_ ( .A({ _09670_, _19647_, _09298_ }), .Y(_19679_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34276_ ( .A({ _09670_, _19646_, _09298_ }), .Y(_19678_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34277_ ( .A({ _09670_, _19644_, _09298_ }), .Y(_19676_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34278_ ( .A({ _09670_, _19643_, _09298_ }), .Y(_19675_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34279_ ( .A({ _09670_, _19642_, _09298_ }), .Y(_19674_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34280_ ( .A({ _09670_, _19641_, _09298_ }), .Y(_19673_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34281_ ( .A({ _09670_, _19640_, _09298_ }), .Y(_19672_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34282_ ( .A({ _09670_, _19639_, _09298_ }), .Y(_19671_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34283_ ( .A({ _09670_, _19638_, _09298_ }), .Y(_19670_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34284_ ( .A({ _09670_, _19637_, _09298_ }), .Y(_19669_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34285_ ( .A({ _09670_, _19636_, _09298_ }), .Y(_19668_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34286_ ( .A({ _09670_, _19635_, _09298_ }), .Y(_19667_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34287_ ( .A({ _09670_, _19665_, _09298_ }), .Y(_19697_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34288_ ( .A({ _09670_, _19664_, _09298_ }), .Y(_19696_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34289_ ( .A({ _09670_, _19663_, _09298_ }), .Y(_19695_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34290_ ( .A({ _09670_, _19662_, _09298_ }), .Y(_19694_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34291_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[5], _05991_, _09298_, _19661_ }), .Y(_19693_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34292_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[4], _05991_, _09298_, _19660_ }), .Y(_19692_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34293_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[3], _05991_, _19659_, _09298_ }), .Y(_19691_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34294_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[2], _05991_, _09298_, _19656_ }), .Y(_19688_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34295_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[1], _05991_, _19645_, _09298_ }), .Y(_19677_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34296_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[0], _05991_, _09298_, _19634_ }), .Y(_19666_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34297_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19004_, _19036_ }), .Y(_18972_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34298_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18822_, _18854_ }), .Y(_18790_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34299_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19003_, _19035_ }), .Y(_18971_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34300_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18820_, _18852_ }), .Y(_18788_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34301_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18438_, _18470_ }), .Y(_18406_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34302_ ( .A({ _05969_, _08878_ }), .Y(_24060_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _34303_ ( .A({ _stream_conv2d_16_source_26_source_pat_fsm_9[1], _08879_, _08887_, _stream_conv2d_16_source_26_source_pat_fsm_9[0] }), .Y(_05969_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34304_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18344_, _18376_ }), .Y(_18312_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34305_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18321_, _18353_ }), .Y(_18289_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34306_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19001_, _19033_ }), .Y(_18969_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34307_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19000_, _19032_ }), .Y(_18968_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34308_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _18999_, _19031_ }), .Y(_18967_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34309_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _18998_, _19030_ }), .Y(_18966_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34310_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _18996_, _19028_ }), .Y(_18964_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34311_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _18995_, _19027_ }), .Y(_18963_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34312_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _18994_, _19026_ }), .Y(_18962_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34313_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _18993_, _19025_ }), .Y(_18961_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34314_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _18992_, _19024_ }), .Y(_18960_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34315_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19022_, _19054_ }), .Y(_18990_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34316_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19021_, _19053_ }), .Y(_18989_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34317_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19020_, _19052_ }), .Y(_18988_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34318_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19019_, _19051_ }), .Y(_18987_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34319_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19018_, _19050_ }), .Y(_18986_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34320_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19016_, _19048_ }), .Y(_18984_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34321_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _19002_, _19034_ }), .Y(_18970_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34322_ ( .A({ _09768_, _stream_conv2d_16_source_19_source_pat_fsm_2[0], _18991_, _19023_ }), .Y(_18959_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34323_ ( .A({ _05984_, _09768_ }), .Y(_24067_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _34324_ ( .A({ _09769_, _stream_conv2d_16_source_19_source_pat_fsm_2[1], _09777_, _stream_conv2d_16_source_19_source_pat_fsm_2[0] }), .Y(_05984_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34325_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18819_, _18851_ }), .Y(_18787_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34326_ ( .A({ _05975_, _09371_ }), .Y(_24063_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _34327_ ( .A({ _stream_conv2d_16_source_23_source_pat_fsm_6[1], _09372_, _09380_, _stream_conv2d_16_source_23_source_pat_fsm_6[0] }), .Y(_05975_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34328_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18818_, _18850_ }), .Y(_18786_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34329_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18817_, _18849_ }), .Y(_18785_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34330_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18816_, _18848_ }), .Y(_18784_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34331_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18815_, _18847_ }), .Y(_18783_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34332_ ( .A({ _06021_, _20409_, _06930_ }), .Y(_20410_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34333_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18814_, _18846_ }), .Y(_18782_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34334_ ( .A({ _19206_, _05987_, _09790_, _19238_ }), .Y(_19174_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34335_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18813_, _18845_ }), .Y(_18781_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34336_ ( .A({ _19204_, _05987_, _09790_, _19236_ }), .Y(_19172_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34337_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18812_, _18844_ }), .Y(_18780_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34338_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18727_, _18759_ }), .Y(_18695_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34339_ ( .A({ _19203_, _05987_, _09790_, _19235_ }), .Y(_19171_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34340_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18811_, _18843_ }), .Y(_18779_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34341_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18726_, _18758_ }), .Y(_18694_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34342_ ( .A({ _19201_, _05987_, _09790_, _19233_ }), .Y(_19169_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34343_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18809_, _18841_ }), .Y(_18777_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34344_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18724_, _18756_ }), .Y(_18692_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34345_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18436_, _18468_ }), .Y(_18404_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34346_ ( .A({ _19200_, _05987_, _09790_, _19232_ }), .Y(_19168_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34347_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18808_, _18840_ }), .Y(_18776_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34348_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18723_, _18755_ }), .Y(_18691_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34349_ ( .A({ _05973_, _09252_ }), .Y(_24062_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _34350_ ( .A({ _09253_, _stream_conv2d_16_source_24_source_pat_fsm_7[1], _09261_, _stream_conv2d_16_source_24_source_pat_fsm_7[0] }), .Y(_05973_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34351_ ( .A({ _19198_, _05987_, _09790_, _19230_ }), .Y(_19166_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34352_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18807_, _18839_ }), .Y(_18775_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34353_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18722_, _18754_ }), .Y(_18690_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34354_ ( .A({ _19197_, _05987_, _09790_, _19229_ }), .Y(_19165_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34355_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18806_, _18838_ }), .Y(_18774_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34356_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18721_, _18753_ }), .Y(_18689_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34357_ ( .A({ _19196_, _05987_, _09790_, _19228_ }), .Y(_19164_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34358_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18805_, _18837_ }), .Y(_18773_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34359_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18720_, _18752_ }), .Y(_18688_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34360_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18435_, _18467_ }), .Y(_18403_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34361_ ( .A({ _19195_, _05987_, _09790_, _19227_ }), .Y(_19163_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34362_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18804_, _18836_ }), .Y(_18772_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34363_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18719_, _18751_ }), .Y(_18687_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34364_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18434_, _18466_ }), .Y(_18402_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34365_ ( .A({ _19193_, _05987_, _09790_, _19225_ }), .Y(_19161_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34366_ ( .A({ _19192_, _05987_, _09790_, _19224_ }), .Y(_19160_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34367_ ( .A({ _19190_, _05987_, _09790_, _19222_ }), .Y(_19158_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34368_ ( .A({ _19189_, _05987_, _09790_, _19221_ }), .Y(_19157_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34369_ ( .A({ _19188_, _05987_, _09790_, _19220_ }), .Y(_19156_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34370_ ( .A({ _19186_, _05987_, _09790_, _19218_ }), .Y(_19154_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34371_ ( .A({ _19185_, _05987_, _09790_, _19217_ }), .Y(_19153_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34372_ ( .A({ _19184_, _05987_, _09790_, _19216_ }), .Y(_19152_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34373_ ( .A({ _19214_, _05987_, _09790_, _19246_ }), .Y(_19182_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34374_ ( .A({ _19213_, _05987_, _09790_, _19245_ }), .Y(_19181_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34375_ ( .A({ _19212_, _05987_, _09790_, _19244_ }), .Y(_19180_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34376_ ( .A({ _19211_, _05987_, _09790_, _19243_ }), .Y(_19179_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34377_ ( .A({ _19210_, _05987_, _09790_, _19242_ }), .Y(_19178_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34378_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19111_, _19143_ }), .Y(_19079_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34379_ ( .A({ _19208_, _05987_, _09790_, _19240_ }), .Y(_19176_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34380_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19110_, _19142_ }), .Y(_19078_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34381_ ( .A({ _19205_, _05987_, _09790_, _19237_ }), .Y(_19173_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34382_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19107_, _19139_ }), .Y(_19075_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34383_ ( .A({ _19183_, _05987_, _09790_, _19215_ }), .Y(_19151_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34384_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19106_, _19138_ }), .Y(_19074_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34385_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19105_, _19137_ }), .Y(_19073_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34386_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19104_, _19136_ }), .Y(_19072_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34387_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19103_, _19135_ }), .Y(_19071_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34388_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19102_, _19134_ }), .Y(_19070_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34389_ ( .A({ _05988_, _05987_, _09790_ }), .Y(_24069_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34390_ ( .A({ _stream_conv2d_16_source_6_source_pat_fsm_0[1], _09791_, _09780_ }), .Y(_05988_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34391_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19101_, _19133_ }), .Y(_19069_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34392_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19100_, _19132_ }), .Y(_19068_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34393_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19099_, _19131_ }), .Y(_19067_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34394_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19097_, _19129_ }), .Y(_19065_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34395_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19096_, _19128_ }), .Y(_19064_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34396_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19095_, _19127_ }), .Y(_19063_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34397_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19094_, _19126_ }), .Y(_19062_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34398_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19093_, _19125_ }), .Y(_19061_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34399_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18803_, _18835_ }), .Y(_18771_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34400_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18718_, _18750_ }), .Y(_18686_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34401_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19092_, _19124_ }), .Y(_19060_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34402_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18802_, _18834_ }), .Y(_18770_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34403_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18717_, _18749_ }), .Y(_18685_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34404_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19091_, _19123_ }), .Y(_19059_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34405_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18801_, _18833_ }), .Y(_18769_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34406_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18716_, _18748_ }), .Y(_18684_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34407_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19090_, _19122_ }), .Y(_19058_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34408_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18800_, _18832_ }), .Y(_18768_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34409_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18715_, _18747_ }), .Y(_18683_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34410_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19089_, _19121_ }), .Y(_19057_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34411_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18830_, _18862_ }), .Y(_18798_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34412_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18713_, _18745_ }), .Y(_18681_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34413_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19088_, _19120_ }), .Y(_19056_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34414_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18829_, _18861_ }), .Y(_18797_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34415_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18712_, _18744_ }), .Y(_18680_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34416_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19118_, _19150_ }), .Y(_19086_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34417_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18828_, _18860_ }), .Y(_18796_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34418_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18711_, _18743_ }), .Y(_18679_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34419_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19117_, _19149_ }), .Y(_19085_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34420_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18827_, _18859_ }), .Y(_18795_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34421_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18710_, _18742_ }), .Y(_18678_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34422_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19116_, _19148_ }), .Y(_19084_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34423_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18826_, _18858_ }), .Y(_18794_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34424_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18709_, _18741_ }), .Y(_18677_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34425_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19115_, _19147_ }), .Y(_19083_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34426_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18825_, _18857_ }), .Y(_18793_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34427_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18708_, _18740_ }), .Y(_18676_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34428_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19114_, _19146_ }), .Y(_19082_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34429_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18824_, _18856_ }), .Y(_18792_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34430_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18707_, _18739_ }), .Y(_18675_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34431_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19113_, _19145_ }), .Y(_19081_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34432_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18821_, _18853_ }), .Y(_18789_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34433_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18706_, _18738_ }), .Y(_18674_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34434_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19112_, _19144_ }), .Y(_19080_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34435_ ( .A({ _07879_, _stream_conv2d_16_source_21_source_pat_fsm_4[0], _18810_, _18842_ }), .Y(_18778_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34436_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18704_, _18736_ }), .Y(_18672_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34437_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19109_, _19141_ }), .Y(_19077_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34438_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18734_, _18766_ }), .Y(_18702_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34439_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18432_, _18464_ }), .Y(_18400_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34440_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19098_, _19130_ }), .Y(_19066_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34441_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18733_, _18765_ }), .Y(_18701_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34442_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18431_, _18463_ }), .Y(_18399_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34443_ ( .A({ _09794_, _stream_conv2d_16_source_8_source_pat_fsm_1[0], _19087_, _19119_ }), .Y(_19055_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34444_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18732_, _18764_ }), .Y(_18700_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34445_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18430_, _18462_ }), .Y(_18398_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34446_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18731_, _18763_ }), .Y(_18699_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34447_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18429_, _18461_ }), .Y(_18397_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34448_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18341_, _18373_ }), .Y(_18309_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34449_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18320_, _18352_ }), .Y(_18288_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34450_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18328_, _18360_ }), .Y(_18296_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34451_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18730_, _18762_ }), .Y(_18698_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34452_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18428_, _18460_ }), .Y(_18396_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34453_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18330_, _18362_ }), .Y(_18298_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34454_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18350_, _18382_ }), .Y(_18318_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34455_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18327_, _18359_ }), .Y(_18295_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34456_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18729_, _18761_ }), .Y(_18697_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34457_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18427_, _18459_ }), .Y(_18395_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34458_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18319_, _18351_ }), .Y(_18287_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34459_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18349_, _18381_ }), .Y(_18317_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34460_ ( .A({ _08878_, _stream_conv2d_16_source_26_source_pat_fsm_9[0], _18326_, _18358_ }), .Y(_18294_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34461_ ( .A({ _07793_, _stream_conv2d_16_source_22_source_pat_fsm_5[0], _18728_, _18760_ }), .Y(_18696_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34462_ ( .A({ _09241_, _stream_conv2d_16_source_25_source_pat_fsm_8[0], _18425_, _18457_ }), .Y(_18393_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34463_ ( .A({ _05985_, _09794_ }), .Y(_24068_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _34464_ ( .A({ _stream_conv2d_16_source_8_source_pat_fsm_1[1], _09795_, _09803_, _stream_conv2d_16_source_8_source_pat_fsm_1[0] }), .Y(_05985_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34465_ ( .A({ _09670_, _19464_, _09298_ }), .Y(_19496_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34466_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18918_, _18950_ }), .Y(_18886_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34467_ ( .A({ _09670_, _19463_, _09298_ }), .Y(_19495_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34468_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18916_, _18948_ }), .Y(_18884_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34469_ ( .A({ _09670_, _19460_, _09298_ }), .Y(_19492_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34470_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18915_, _18947_ }), .Y(_18883_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34471_ ( .A({ _09670_, _19457_, _09298_ }), .Y(_19489_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34472_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18912_, _18944_ }), .Y(_18880_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34473_ ( .A({ _09670_, _19456_, _09298_ }), .Y(_19488_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34474_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18911_, _18943_ }), .Y(_18879_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34475_ ( .A({ _20441_, _06930_, _07066_, _20473_ }), .Y(_05659_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34476_ ( .A({ _09670_, _19455_, _09298_ }), .Y(_19487_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34477_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18910_, _18942_ }), .Y(_18878_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34478_ ( .A({ _20437_, _06930_, _07066_, _20469_ }), .Y(_05660_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34479_ ( .A({ _09670_, _19450_, _09298_ }), .Y(_19482_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34480_ ( .A({ _20436_, _06930_, _07066_, _20468_ }), .Y(_05661_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34481_ ( .A({ _09670_, _19449_, _09298_ }), .Y(_19481_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34482_ ( .A({ _20435_, _06930_, _07066_, _20467_ }), .Y(_05662_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34483_ ( .A({ _09670_, _19448_, _09298_ }), .Y(_19480_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34484_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18907_, _18939_ }), .Y(_18875_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34485_ ( .A({ _20432_, _06930_, _07066_, _20464_ }), .Y(_05663_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34486_ ( .A({ _09670_, _19445_, _09298_ }), .Y(_19477_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34487_ ( .A({ _09930_, _19270_, _09298_ }), .Y(_19302_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34488_ ( .A({ _19366_, _05727_, _09303_, _19334_ }), .Y(_09930_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34489_ ( .A({ _20431_, _06930_, _07066_, _20463_ }), .Y(_05664_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34490_ ( .A({ _09670_, _19442_, _09298_ }), .Y(_19474_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34491_ ( .A({ _09931_, _19332_, _09303_ }), .Y(_19300_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34492_ ( .A({ _19268_, _09298_, _19364_, _05727_ }), .Y(_09931_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34493_ ( .A({ _20430_, _06930_, _07066_, _20462_ }), .Y(_05665_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34494_ ( .A({ _09670_, _19441_, _09298_ }), .Y(_19473_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34495_ ( .A({ _09932_, _19267_, _09298_ }), .Y(_19299_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34496_ ( .A({ _19363_, _05727_, _09303_, _19331_ }), .Y(_09932_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34497_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18904_, _18936_ }), .Y(_18872_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34498_ ( .A({ _05962_, _09933_ }), .Y(_24055_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _34499_ ( .A({ _09934_, _09939_, _stream_conv2d_16_source_31_source_pat_fsm_14[0] }), .Y(_09933_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34500_ ( .A({ _09938_, _09937_, _09935_ }), .Y(_09934_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34501_ ( .A({ _09936_, _stream_conv2d_16_source_31_source_pat_fsm_14[3:2] }), .Y(_09935_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34502_ ( .A(_stream_conv2d_16_source_31_source_pat_fsm_14[7:4]), .Y(_09936_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34503_ ( .A(_stream_conv2d_16_source_31_source_pat_fsm_14[15:12]), .Y(_09937_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34504_ ( .A(_stream_conv2d_16_source_31_source_pat_fsm_14[11:8]), .Y(_09938_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34505_ ( .A({ _09943_, _09942_, _09941_, _09940_ }), .Y(_09939_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34506_ ( .A(_stream_conv2d_16_source_31_source_pat_fsm_14[23:20]), .Y(_09940_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34507_ ( .A(_stream_conv2d_16_source_31_source_pat_fsm_14[19:16]), .Y(_09941_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34508_ ( .A(_stream_conv2d_16_source_31_source_pat_fsm_14[31:28]), .Y(_09942_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34509_ ( .A(_stream_conv2d_16_source_31_source_pat_fsm_14[27:24]), .Y(_09943_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _34510_ ( .A({ _09934_, _stream_conv2d_16_source_31_source_pat_fsm_14[0], _09939_, _stream_conv2d_16_source_31_source_pat_fsm_14[1] }), .Y(_05962_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34511_ ( .A({ _20425_, _06930_, _07066_, _20457_ }), .Y(_05666_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34512_ ( .A({ _09670_, _19471_, _09298_ }), .Y(_19503_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34513_ ( .A({ _09944_, _19266_, _09298_ }), .Y(_19298_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34514_ ( .A({ _19362_, _05727_, _09303_, _19330_ }), .Y(_09944_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34515_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18903_, _18935_ }), .Y(_18871_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34516_ ( .A({ _20424_, _06930_, _07066_, _20456_ }), .Y(_05667_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34517_ ( .A({ _09670_, _19470_, _09298_ }), .Y(_19502_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34518_ ( .A({ _09945_, _19329_, _09303_ }), .Y(_19297_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34519_ ( .A({ _19265_, _09298_, _19361_, _05727_ }), .Y(_09945_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34520_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18902_, _18934_ }), .Y(_18870_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34521_ ( .A({ _20422_, _06930_, _07066_, _20454_ }), .Y(_05668_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34522_ ( .A({ _09946_, _19328_, _09303_ }), .Y(_19296_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34523_ ( .A({ _19264_, _09298_, _19360_, _05727_ }), .Y(_09946_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34524_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18901_, _18933_ }), .Y(_18869_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34525_ ( .A({ _20419_, _06930_, _07066_, _20451_ }), .Y(_05669_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34526_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[5], _05991_, _19467_, _09298_ }), .Y(_19499_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34527_ ( .A({ _09947_, _19261_, _09298_ }), .Y(_19293_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34528_ ( .A({ _19357_, _05727_, _09303_, _19325_ }), .Y(_09947_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34529_ ( .A({ _20418_, _06930_, _07066_, _20450_ }), .Y(_05670_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34530_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[3], _05991_, _19465_, _09298_ }), .Y(_19497_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34531_ ( .A({ _09948_, _19324_, _09303_ }), .Y(_19292_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34532_ ( .A({ _19260_, _09298_, _19356_, _05727_ }), .Y(_09948_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34533_ ( .A({ _20448_, _06930_, _07066_, _20480_ }), .Y(_05671_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34534_ ( .A({ cparam_conv2d_16_stream_act_local_large_offset[2], _05991_, _19462_, _09298_ }), .Y(_19494_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34535_ ( .A({ _09949_, _19259_, _09298_ }), .Y(_19291_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34536_ ( .A({ _19355_, _05727_, _09303_, _19323_ }), .Y(_09949_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34537_ ( .A({ _20445_, _06930_, _07066_, _20477_ }), .Y(_05672_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34538_ ( .A({ _09950_, _19319_, _09303_ }), .Y(_19287_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34539_ ( .A({ _19255_, _09298_, _19351_, _05727_ }), .Y(_09950_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34540_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18898_, _18930_ }), .Y(_18866_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34541_ ( .A({ _20444_, _06930_, _07066_, _20476_ }), .Y(_05673_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34542_ ( .A({ _09951_, _19254_, _09298_ }), .Y(_19286_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34543_ ( .A({ _19350_, _05727_, _09303_, _19318_ }), .Y(_09951_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34544_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18896_, _18928_ }), .Y(_18864_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34545_ ( .A({ _20443_, _06930_, _07066_, _20475_ }), .Y(_05674_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34546_ ( .A({ _09952_, _19253_, _09298_ }), .Y(_19285_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34547_ ( .A({ _19349_, _05727_, _09303_, _19317_ }), .Y(_09952_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34548_ ( .A({ _20439_, _06930_, _07066_, _20471_ }), .Y(_05675_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34549_ ( .A({ _09953_, _19251_, _09298_ }), .Y(_19283_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34550_ ( .A({ _19347_, _05727_, _09303_, _19315_ }), .Y(_09953_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34551_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18925_, _18957_ }), .Y(_18893_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34552_ ( .A({ _20428_, _06930_, _07066_, _20460_ }), .Y(_05676_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34553_ ( .A({ _09954_, _19250_, _09298_ }), .Y(_19282_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34554_ ( .A({ _19346_, _05727_, _09303_, _19314_ }), .Y(_09954_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34555_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18924_, _18956_ }), .Y(_18892_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34556_ ( .A({ _20417_, _06930_, _07066_, _20449_ }), .Y(_05677_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34557_ ( .A({ _09955_, _19313_, _09303_ }), .Y(_19281_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34558_ ( .A({ _19249_, _09298_, _19345_, _05727_ }), .Y(_09955_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34559_ ( .A({ _09263_, _stream_conv2d_16_source_20_source_pat_fsm_3[0], _18923_, _18955_ }), .Y(_18891_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34560_ ( .A({ _17871_, _09956_, _17839_, _05962_ }), .Y(_17807_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34561_ ( .A({ _09933_, _stream_conv2d_16_source_31_source_pat_fsm_14[1] }), .Y(_09956_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34562_ ( .A({ _17882_, _09956_, _17850_, _05962_ }), .Y(_17818_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34563_ ( .A({ _17893_, _09956_, _17861_, _05962_ }), .Y(_17829_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34564_ ( .A({ _09957_, _19341_, _09303_ }), .Y(_19309_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34565_ ( .A({ _19277_, _09298_, _19373_, _05727_ }), .Y(_09957_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34566_ ( .A({ _09958_, _19340_, _09303_ }), .Y(_19308_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34567_ ( .A({ _19276_, _09298_, _19372_, _05727_ }), .Y(_09958_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34568_ ( .A({ _09959_, _19275_, _09298_ }), .Y(_19307_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34569_ ( .A({ _19371_, _05727_, _09303_, _19339_ }), .Y(_09959_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34570_ ( .A({ _17896_, _09956_, _17864_, _05962_ }), .Y(_17832_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34571_ ( .A({ _17897_, _09956_, _17865_, _05962_ }), .Y(_17833_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34572_ ( .A({ _17898_, _09956_, _17866_, _05962_ }), .Y(_17834_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34573_ ( .A({ _17899_, _09956_, _17867_, _05962_ }), .Y(_17835_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34574_ ( .A({ _17900_, _09956_, _17868_, _05962_ }), .Y(_17836_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34575_ ( .A({ _17901_, _09956_, _17869_, _05962_ }), .Y(_17837_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34576_ ( .A({ _09960_, _19273_, _09298_ }), .Y(_19305_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34577_ ( .A({ _19369_, _05727_, _09303_, _19337_ }), .Y(_09960_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34578_ ( .A({ _09961_, _19336_, _09303_ }), .Y(_19304_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34579_ ( .A({ _19272_, _09298_, _19368_, _05727_ }), .Y(_09961_) );
  \$lut  #( .LUT(16'h8fff), .WIDTH(4) ) _34580_ ( .A({ _09962_, _09304_, _09303_, _19322_ }), .Y(_19290_) );
  \$lut  #( .LUT(16'h0bbb), .WIDTH(4) ) _34581_ ( .A({ _19258_, _09298_, _19354_, _05727_ }), .Y(_09962_) );
  \$lut  #( .LUT(16'h8fff), .WIDTH(4) ) _34582_ ( .A({ _09963_, _05990_, _09298_, _19247_ }), .Y(_19279_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _34583_ ( .A({ _19343_, _05727_, _09303_, _19311_ }), .Y(_09963_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34584_ ( .A({ _17902_, _09956_, _17870_, _05962_ }), .Y(_17838_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34585_ ( .A({ _17872_, _09956_, _17840_, _05962_ }), .Y(_17808_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34586_ ( .A({ _17873_, _09956_, _17841_, _05962_ }), .Y(_17809_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34587_ ( .A({ _17874_, _09956_, _17842_, _05962_ }), .Y(_17810_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34588_ ( .A({ _17875_, _09956_, _17843_, _05962_ }), .Y(_17811_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34589_ ( .A({ _17876_, _09956_, _17844_, _05962_ }), .Y(_17812_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34590_ ( .A({ _17877_, _09956_, _17845_, _05962_ }), .Y(_17813_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34591_ ( .A({ _17878_, _09956_, _17846_, _05962_ }), .Y(_17814_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34592_ ( .A({ _17879_, _09956_, _17847_, _05962_ }), .Y(_17815_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34593_ ( .A({ _17880_, _09956_, _17848_, _05962_ }), .Y(_17816_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34594_ ( .A({ _17881_, _09956_, _17849_, _05962_ }), .Y(_17817_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34595_ ( .A({ _17883_, _09956_, _17851_, _05962_ }), .Y(_17819_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34596_ ( .A({ _17884_, _09956_, _17852_, _05962_ }), .Y(_17820_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34597_ ( .A({ _17885_, _09956_, _17853_, _05962_ }), .Y(_17821_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34598_ ( .A({ _17886_, _09956_, _17854_, _05962_ }), .Y(_17822_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34599_ ( .A({ _17887_, _09956_, _17855_, _05962_ }), .Y(_17823_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34600_ ( .A({ _17888_, _09956_, _17856_, _05962_ }), .Y(_17824_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34601_ ( .A({ _17889_, _09956_, _17857_, _05962_ }), .Y(_17825_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34602_ ( .A({ _17890_, _09956_, _17858_, _05962_ }), .Y(_17826_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34603_ ( .A({ _17891_, _09956_, _17859_, _05962_ }), .Y(_17827_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34604_ ( .A({ _17892_, _09956_, _17860_, _05962_ }), .Y(_17828_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34605_ ( .A({ _17894_, _09956_, _17862_, _05962_ }), .Y(_17830_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _34606_ ( .A({ _17895_, _09956_, _17863_, _05962_ }), .Y(_17831_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34607_ ( .A({ _20111_, _05996_, _09285_, _20177_ }), .Y(_20144_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34608_ ( .A({ _20110_, _05996_, _09285_, _20176_ }), .Y(_20143_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34609_ ( .A({ _20109_, _05996_, _09285_, _20175_ }), .Y(_20142_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34610_ ( .A({ _20107_, _05996_, _09285_, _20173_ }), .Y(_20140_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34611_ ( .A({ _20106_, _05996_, _09285_, _20172_ }), .Y(_20139_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34612_ ( .A({ _20433_, _06930_, _07066_, _20465_ }), .Y(_05678_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _34613_ ( .A({ _20429_, _06930_, _07066_, _20461_ }), .Y(_05679_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _34614_ ( .A({ _07066_, _05514_ }), .Y(_24074_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34615_ ( .A({ _09964_, _04442_, _08509_ }), .Y(_22879_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34616_ ( .A({ _04570_, _08507_, _04666_, _08508_ }), .Y(_09964_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34617_ ( .A({ _09965_, _04667_, _08508_ }), .Y(_22880_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34618_ ( .A({ _04571_, _08507_, _08509_, _04443_ }), .Y(_09965_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34619_ ( .A({ _09966_, _04480_, _08473_ }), .Y(_22853_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34620_ ( .A({ _04704_, _08474_, _08472_, _04608_ }), .Y(_09966_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34621_ ( .A({ _09967_, _04703_, _08474_ }), .Y(_22852_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _34622_ ( .A({ _04607_, _08472_, _08473_, _04479_ }), .Y(_09967_) );
  \$lut  #( .LUT(16'hfff8), .WIDTH(4) ) _34623_ ( .A({ _05681_, _05680_, _06901_, _06907_ }), .Y(_24090_) );
  \$lut  #( .LUT(16'hfff8), .WIDTH(4) ) _34624_ ( .A({ _05646_, _05682_, _06908_, _06917_ }), .Y(_24091_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34625_ ( .A({ _09142_, _05683_ }), .Y(_24092_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34626_ ( .A({ _09973_, _09968_ }), .Y(_tmp_1281) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34627_ ( .A({ _stream_matmul_29_fsm[1], _09972_, _09969_ }), .Y(_09968_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34628_ ( .A({ _09971_, _09970_, _stream_matmul_29_fsm[3:2] }), .Y(_09969_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34629_ ( .A(_stream_matmul_29_fsm[15:12]), .Y(_09970_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34630_ ( .A(_stream_matmul_29_fsm[11:8]), .Y(_09971_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34631_ ( .A(_stream_matmul_29_fsm[7:4]), .Y(_09972_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34632_ ( .A({ _stream_matmul_29_fsm[0], _09974_ }), .Y(_09973_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34633_ ( .A({ _09978_, _09977_, _09976_, _09975_ }), .Y(_09974_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34634_ ( .A(_stream_matmul_29_fsm[23:20]), .Y(_09975_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34635_ ( .A(_stream_matmul_29_fsm[19:16]), .Y(_09976_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34636_ ( .A(_stream_matmul_29_fsm[31:28]), .Y(_09977_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34637_ ( .A(_stream_matmul_29_fsm[27:24]), .Y(_09978_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34638_ ( .A({ _05685_, _tmp_1281 }), .Y(_24093_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34639_ ( .A({ _09980_, _09979_ }), .Y(_05685_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34640_ ( .A({ _09974_, _stream_matmul_29_fsm[0] }), .Y(_09979_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _34641_ ( .A({ _09969_, _09972_, _stream_matmul_29_fsm[1] }), .Y(_09980_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34642_ ( .A({ _23623_, _05685_, _23591_, _09981_ }), .Y(_23559_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34643_ ( .A({ _09979_, _09968_ }), .Y(_09981_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34644_ ( .A({ _23622_, _05685_, _23590_, _09981_ }), .Y(_23558_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34645_ ( .A({ _23620_, _05685_, _23588_, _09981_ }), .Y(_23556_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34646_ ( .A({ _23619_, _05685_, _23587_, _09981_ }), .Y(_23555_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34647_ ( .A({ _23618_, _05685_, _23586_, _09981_ }), .Y(_23554_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34648_ ( .A({ _23617_, _05685_, _23585_, _09981_ }), .Y(_23553_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34649_ ( .A({ _23616_, _05685_, _23584_, _09981_ }), .Y(_23552_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34650_ ( .A({ _23615_, _05685_, _23583_, _09981_ }), .Y(_23551_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34651_ ( .A({ _23614_, _05685_, _23582_, _09981_ }), .Y(_23550_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34652_ ( .A({ _23613_, _05685_, _23581_, _09981_ }), .Y(_23549_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34653_ ( .A({ _23612_, _05685_, _23580_, _09981_ }), .Y(_23548_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34654_ ( .A({ _23611_, _05685_, _23579_, _09981_ }), .Y(_23547_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34655_ ( .A({ _23609_, _05685_, _23577_, _09981_ }), .Y(_23545_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34656_ ( .A({ _23608_, _05685_, _23576_, _09981_ }), .Y(_23544_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34657_ ( .A({ _23607_, _05685_, _23575_, _09981_ }), .Y(_23543_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34658_ ( .A({ _23606_, _05685_, _23574_, _09981_ }), .Y(_23542_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34659_ ( .A({ _23605_, _05685_, _23573_, _09981_ }), .Y(_23541_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34660_ ( .A({ _23604_, _05685_, _23572_, _09981_ }), .Y(_23540_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34661_ ( .A({ _23603_, _05685_, _23571_, _09981_ }), .Y(_23539_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34662_ ( .A({ _23602_, _05685_, _23570_, _09981_ }), .Y(_23538_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34663_ ( .A({ _23601_, _05685_, _23569_, _09981_ }), .Y(_23537_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34664_ ( .A({ _23600_, _05685_, _23568_, _09981_ }), .Y(_23536_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34665_ ( .A({ _23630_, _05685_, _23598_, _09981_ }), .Y(_23566_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34666_ ( .A({ _23629_, _05685_, _23597_, _09981_ }), .Y(_23565_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34667_ ( .A({ _23628_, _05685_, _23596_, _09981_ }), .Y(_23564_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34668_ ( .A({ _23627_, _05685_, _23595_, _09981_ }), .Y(_23563_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34669_ ( .A({ _23626_, _05685_, _23594_, _09981_ }), .Y(_23562_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34670_ ( .A({ _23625_, _05685_, _23593_, _09981_ }), .Y(_23561_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34671_ ( .A({ _23624_, _05685_, _23592_, _09981_ }), .Y(_23560_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34672_ ( .A({ _23621_, _05685_, _23589_, _09981_ }), .Y(_23557_) );
  \$lut  #( .LUT(8'h8f), .WIDTH(3) ) _34673_ ( .A({ _09982_, _23578_, _09981_ }), .Y(_23546_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _34674_ ( .A({ _09983_, _05685_, _23610_ }), .Y(_09982_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34675_ ( .A({ _09980_, _09973_ }), .Y(_09983_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34676_ ( .A({ _23599_, _05685_, _23567_, _09981_ }), .Y(_23535_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _34677_ ( .A({ _09983_, _09981_, _24093_ }), .Y(_24094_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34678_ ( .A({ _stream_max_pool_serial_18_fsm[0], _09989_, _09984_ }), .Y(_tmp_1056) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34679_ ( .A({ _stream_max_pool_serial_18_fsm[1], _09988_, _09985_ }), .Y(_09984_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34680_ ( .A({ _09987_, _09986_, _stream_max_pool_serial_18_fsm[3:2] }), .Y(_09985_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34681_ ( .A(_stream_max_pool_serial_18_fsm[15:12]), .Y(_09986_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34682_ ( .A(_stream_max_pool_serial_18_fsm[11:8]), .Y(_09987_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34683_ ( .A(_stream_max_pool_serial_18_fsm[7:4]), .Y(_09988_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34684_ ( .A({ _09993_, _09992_, _09991_, _09990_ }), .Y(_09989_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34685_ ( .A(_stream_max_pool_serial_18_fsm[23:20]), .Y(_09990_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34686_ ( .A(_stream_max_pool_serial_18_fsm[19:16]), .Y(_09991_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34687_ ( .A(_stream_max_pool_serial_18_fsm[31:28]), .Y(_09992_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34688_ ( .A(_stream_max_pool_serial_18_fsm[27:24]), .Y(_09993_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34689_ ( .A({ _05686_, _tmp_1056 }), .Y(_24095_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34690_ ( .A({ _09995_, _09994_ }), .Y(_05686_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34691_ ( .A({ _09989_, _stream_max_pool_serial_18_fsm[0] }), .Y(_09994_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _34692_ ( .A({ _09985_, _09988_, _stream_max_pool_serial_18_fsm[1] }), .Y(_09995_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34693_ ( .A({ _23721_, _05686_, _23689_, _09996_ }), .Y(_23657_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34694_ ( .A({ _09994_, _09984_ }), .Y(_09996_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34695_ ( .A({ _23720_, _05686_, _23688_, _09996_ }), .Y(_23656_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34696_ ( .A({ _23718_, _05686_, _23686_, _09996_ }), .Y(_23654_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34697_ ( .A({ _23717_, _05686_, _23685_, _09996_ }), .Y(_23653_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34698_ ( .A({ _23716_, _05686_, _23684_, _09996_ }), .Y(_23652_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34699_ ( .A({ _23715_, _05686_, _23683_, _09996_ }), .Y(_23651_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34700_ ( .A({ _23714_, _05686_, _23682_, _09996_ }), .Y(_23650_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34701_ ( .A({ _23713_, _05686_, _23681_, _09996_ }), .Y(_23649_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34702_ ( .A({ _23712_, _05686_, _23680_, _09996_ }), .Y(_23648_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34703_ ( .A({ _23711_, _05686_, _23679_, _09996_ }), .Y(_23647_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34704_ ( .A({ _23710_, _05686_, _23678_, _09996_ }), .Y(_23646_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34705_ ( .A({ _23709_, _05686_, _23677_, _09996_ }), .Y(_23645_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34706_ ( .A({ _23707_, _05686_, _23675_, _09996_ }), .Y(_23643_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34707_ ( .A({ _23706_, _05686_, _23674_, _09996_ }), .Y(_23642_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34708_ ( .A({ _23705_, _05686_, _23673_, _09996_ }), .Y(_23641_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34709_ ( .A({ _23704_, _05686_, _23672_, _09996_ }), .Y(_23640_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34710_ ( .A({ _23703_, _05686_, _23671_, _09996_ }), .Y(_23639_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34711_ ( .A({ _23702_, _05686_, _23670_, _09996_ }), .Y(_23638_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34712_ ( .A({ _23701_, _05686_, _23669_, _09996_ }), .Y(_23637_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34713_ ( .A({ _23700_, _05686_, _23668_, _09996_ }), .Y(_23636_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34714_ ( .A({ _23699_, _05686_, _23667_, _09996_ }), .Y(_23635_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34715_ ( .A({ _23698_, _05686_, _23666_, _09996_ }), .Y(_23634_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34716_ ( .A({ _23728_, _05686_, _23696_, _09996_ }), .Y(_23664_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34717_ ( .A({ _23727_, _05686_, _23695_, _09996_ }), .Y(_23663_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34718_ ( .A({ _23726_, _05686_, _23694_, _09996_ }), .Y(_23662_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34719_ ( .A({ _23725_, _05686_, _23693_, _09996_ }), .Y(_23661_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34720_ ( .A({ _23724_, _05686_, _23692_, _09996_ }), .Y(_23660_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34721_ ( .A({ _23723_, _05686_, _23691_, _09996_ }), .Y(_23659_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34722_ ( .A({ _23722_, _05686_, _23690_, _09996_ }), .Y(_23658_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34723_ ( .A({ _23719_, _05686_, _23687_, _09996_ }), .Y(_23655_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34724_ ( .A({ _09997_, _23676_, _09996_ }), .Y(_23644_) );
  \$lut  #( .LUT(16'he000), .WIDTH(4) ) _34725_ ( .A({ _09989_, _09995_, _stream_max_pool_serial_18_fsm[0], _23708_ }), .Y(_09997_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34726_ ( .A({ _23697_, _05686_, _23665_, _09996_ }), .Y(_23633_) );
  \$lut  #( .LUT(8'he0), .WIDTH(3) ) _34727_ ( .A({ _09989_, _09984_, _09995_ }), .Y(_24096_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34728_ ( .A({ _stream_conv2d_16_fsm[0], _10003_, _09998_ }), .Y(_tmp_943) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34729_ ( .A({ _stream_conv2d_16_fsm[1], _10002_, _09999_ }), .Y(_09998_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34730_ ( .A({ _10001_, _10000_, _stream_conv2d_16_fsm[3:2] }), .Y(_09999_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34731_ ( .A(_stream_conv2d_16_fsm[15:12]), .Y(_10000_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34732_ ( .A(_stream_conv2d_16_fsm[11:8]), .Y(_10001_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34733_ ( .A(_stream_conv2d_16_fsm[7:4]), .Y(_10002_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34734_ ( .A({ _10007_, _10006_, _10005_, _10004_ }), .Y(_10003_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34735_ ( .A(_stream_conv2d_16_fsm[23:20]), .Y(_10004_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34736_ ( .A(_stream_conv2d_16_fsm[19:16]), .Y(_10005_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34737_ ( .A(_stream_conv2d_16_fsm[31:28]), .Y(_10006_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34738_ ( .A(_stream_conv2d_16_fsm[27:24]), .Y(_10007_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34739_ ( .A({ _05687_, _tmp_943 }), .Y(_24097_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34740_ ( .A({ _10009_, _10008_ }), .Y(_05687_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34741_ ( .A({ _10003_, _stream_conv2d_16_fsm[0] }), .Y(_10008_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _34742_ ( .A({ _09999_, _10002_, _stream_conv2d_16_fsm[1] }), .Y(_10009_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34743_ ( .A({ _23819_, _05687_, _23787_, _10010_ }), .Y(_23755_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _34744_ ( .A({ _10008_, _09998_ }), .Y(_10010_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34745_ ( .A({ _23818_, _05687_, _23786_, _10010_ }), .Y(_23754_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34746_ ( .A({ _23816_, _05687_, _23784_, _10010_ }), .Y(_23752_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34747_ ( .A({ _23815_, _05687_, _23783_, _10010_ }), .Y(_23751_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34748_ ( .A({ _23814_, _05687_, _23782_, _10010_ }), .Y(_23750_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34749_ ( .A({ _23813_, _05687_, _23781_, _10010_ }), .Y(_23749_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34750_ ( .A({ _23812_, _05687_, _23780_, _10010_ }), .Y(_23748_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34751_ ( .A({ _23811_, _05687_, _23779_, _10010_ }), .Y(_23747_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34752_ ( .A({ _23810_, _05687_, _23778_, _10010_ }), .Y(_23746_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34753_ ( .A({ _23809_, _05687_, _23777_, _10010_ }), .Y(_23745_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34754_ ( .A({ _23808_, _05687_, _23776_, _10010_ }), .Y(_23744_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34755_ ( .A({ _23807_, _05687_, _23775_, _10010_ }), .Y(_23743_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34756_ ( .A({ _23805_, _05687_, _23773_, _10010_ }), .Y(_23741_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34757_ ( .A({ _23804_, _05687_, _23772_, _10010_ }), .Y(_23740_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34758_ ( .A({ _23803_, _05687_, _23771_, _10010_ }), .Y(_23739_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34759_ ( .A({ _23802_, _05687_, _23770_, _10010_ }), .Y(_23738_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34760_ ( .A({ _23801_, _05687_, _23769_, _10010_ }), .Y(_23737_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34761_ ( .A({ _23800_, _05687_, _23768_, _10010_ }), .Y(_23736_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34762_ ( .A({ _23799_, _05687_, _23767_, _10010_ }), .Y(_23735_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34763_ ( .A({ _23798_, _05687_, _23766_, _10010_ }), .Y(_23734_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34764_ ( .A({ _23797_, _05687_, _23765_, _10010_ }), .Y(_23733_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34765_ ( .A({ _23796_, _05687_, _23764_, _10010_ }), .Y(_23732_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34766_ ( .A({ _23826_, _05687_, _23794_, _10010_ }), .Y(_23762_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34767_ ( .A({ _23825_, _05687_, _23793_, _10010_ }), .Y(_23761_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34768_ ( .A({ _23824_, _05687_, _23792_, _10010_ }), .Y(_23760_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34769_ ( .A({ _23823_, _05687_, _23791_, _10010_ }), .Y(_23759_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34770_ ( .A({ _23822_, _05687_, _23790_, _10010_ }), .Y(_23758_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34771_ ( .A({ _23821_, _05687_, _23789_, _10010_ }), .Y(_23757_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34772_ ( .A({ _23820_, _05687_, _23788_, _10010_ }), .Y(_23756_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34773_ ( .A({ _23817_, _05687_, _23785_, _10010_ }), .Y(_23753_) );
  \$lut  #( .LUT(8'hf8), .WIDTH(3) ) _34774_ ( .A({ _10011_, _23774_, _10010_ }), .Y(_23742_) );
  \$lut  #( .LUT(16'he000), .WIDTH(4) ) _34775_ ( .A({ _10003_, _10009_, _stream_conv2d_16_fsm[0], _23806_ }), .Y(_10011_) );
  \$lut  #( .LUT(16'h8f88), .WIDTH(4) ) _34776_ ( .A({ _23795_, _05687_, _23763_, _10010_ }), .Y(_23731_) );
  \$lut  #( .LUT(8'he0), .WIDTH(3) ) _34777_ ( .A({ _10003_, _09998_, _10009_ }), .Y(_24098_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34778_ ( .A({ _10012_, _saxi_register_fsm[0], _23883_, _23915_ }), .Y(_23851_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _34779_ ( .A({ _10013_, _10021_, _saxi_register_fsm[1] }), .Y(_10012_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _34780_ ( .A({ _10020_, _10019_, _10014_ }), .Y(_10013_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34781_ ( .A({ _10018_, _10017_, _10016_, _10015_ }), .Y(_10014_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34782_ ( .A(_saxi_register_fsm[23:20]), .Y(_10015_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34783_ ( .A(_saxi_register_fsm[19:16]), .Y(_10016_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34784_ ( .A(_saxi_register_fsm[31:28]), .Y(_10017_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34785_ ( .A(_saxi_register_fsm[27:24]), .Y(_10018_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34786_ ( .A(_saxi_register_fsm[15:12]), .Y(_10019_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34787_ ( .A(_saxi_register_fsm[11:8]), .Y(_10020_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _34788_ ( .A({ _10022_, _saxi_register_fsm[3:2] }), .Y(_10021_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34789_ ( .A(_saxi_register_fsm[7:4]), .Y(_10022_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34790_ ( .A({ _10012_, _saxi_register_fsm[0], _23882_, _23914_ }), .Y(_23850_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34791_ ( .A({ _10012_, _saxi_register_fsm[0], _23880_, _23912_ }), .Y(_23848_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34792_ ( .A({ _10012_, _saxi_register_fsm[0], _23879_, _23911_ }), .Y(_23847_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34793_ ( .A({ _10012_, _saxi_register_fsm[0], _23878_, _23910_ }), .Y(_23846_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34794_ ( .A({ _10012_, _saxi_register_fsm[0], _23877_, _23909_ }), .Y(_23845_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34795_ ( .A({ _10012_, _saxi_register_fsm[0], _23876_, _23908_ }), .Y(_23844_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34796_ ( .A({ _10012_, _saxi_register_fsm[0], _23875_, _23907_ }), .Y(_23843_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34797_ ( .A({ _10012_, _saxi_register_fsm[0], _23874_, _23906_ }), .Y(_23842_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34798_ ( .A({ _10012_, _saxi_register_fsm[0], _23873_, _23905_ }), .Y(_23841_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34799_ ( .A({ _10012_, _saxi_register_fsm[0], _23872_, _23904_ }), .Y(_23840_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34800_ ( .A({ _10012_, _saxi_register_fsm[0], _23871_, _23903_ }), .Y(_23839_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34801_ ( .A({ _10012_, _saxi_register_fsm[0], _23869_, _23901_ }), .Y(_23837_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34802_ ( .A({ _10012_, _saxi_register_fsm[0], _23868_, _23900_ }), .Y(_23836_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34803_ ( .A({ _10012_, _saxi_register_fsm[0], _23867_, _23899_ }), .Y(_23835_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34804_ ( .A({ _10012_, _saxi_register_fsm[0], _23866_, _23898_ }), .Y(_23834_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34805_ ( .A({ _10012_, _saxi_register_fsm[0], _23865_, _23897_ }), .Y(_23833_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34806_ ( .A({ _10012_, _saxi_register_fsm[0], _23864_, _23896_ }), .Y(_23832_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34807_ ( .A({ _10012_, _saxi_register_fsm[0], _23863_, _23895_ }), .Y(_23831_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34808_ ( .A({ _10012_, _saxi_register_fsm[0], _23862_, _23894_ }), .Y(_23830_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34809_ ( .A({ _10012_, _saxi_register_fsm[0], _23861_, _23893_ }), .Y(_23829_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34810_ ( .A({ _10012_, _saxi_register_fsm[0], _23860_, _23892_ }), .Y(_23828_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34811_ ( .A({ _10012_, _saxi_register_fsm[0], _23890_, _23922_ }), .Y(_23858_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34812_ ( .A({ _10012_, _saxi_register_fsm[0], _23889_, _23921_ }), .Y(_23857_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34813_ ( .A({ _10012_, _saxi_register_fsm[0], _23888_, _23920_ }), .Y(_23856_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34814_ ( .A({ _10012_, _saxi_register_fsm[0], _23887_, _23919_ }), .Y(_23855_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34815_ ( .A({ _10012_, _saxi_register_fsm[0], _23886_, _23918_ }), .Y(_23854_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34816_ ( .A({ _10012_, _saxi_register_fsm[0], _23885_, _23917_ }), .Y(_23853_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34817_ ( .A({ _10012_, _saxi_register_fsm[0], _23884_, _23916_ }), .Y(_23852_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34818_ ( .A({ _10012_, _saxi_register_fsm[0], _23881_, _23913_ }), .Y(_23849_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34819_ ( .A({ _10012_, _saxi_register_fsm[0], _23870_, _23902_ }), .Y(_23838_) );
  \$lut  #( .LUT(16'hca00), .WIDTH(4) ) _34820_ ( .A({ _10012_, _saxi_register_fsm[0], _23859_, _23891_ }), .Y(_23827_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34821_ ( .A({ _10013_, _saxi_register_fsm[1], _10021_, _saxi_register_fsm[0] }), .Y(saxi_wready) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _34822_ ( .A({ saxi_wready, _10012_ }), .Y(_24099_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34823_ ( .A({ _05929_, _13755_ }), .Y(_05515_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34824_ ( .A({ conv2d_16_control_param_index[0], conv2d_16_control_param_index[1] }), .Y(_05744_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34825_ ( .A({ max_pool_serial_18_control_param_index[0], max_pool_serial_18_control_param_index[1] }), .Y(_05745_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34826_ ( .A({ matmul_29_control_param_index[0], matmul_29_control_param_index[1] }), .Y(_05746_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34827_ ( .A({ conv2d_16_prev_row_select[0], conv2d_16_prev_row_select[1] }), .Y(_05747_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34828_ ( .A(conv2d_16_prev_row_select), .Y(_05748_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34829_ ( .A({ __tmp_464_2[0], __tmp_464_2[1] }), .Y(_05749_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34830_ ( .A(__tmp_464_2), .Y(_05750_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34831_ ( .A({ __tmp_464_2[0], __tmp_464_2[1] }), .Y(_05751_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34832_ ( .A({ __tmp_475_2[0], __tmp_475_2[1] }), .Y(_05752_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34833_ ( .A(__tmp_475_2), .Y(_05753_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34834_ ( .A({ __tmp_475_2[0], __tmp_475_2[1] }), .Y(_05754_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34835_ ( .A({ __tmp_495_2[0], __tmp_495_2[1] }), .Y(_05755_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34836_ ( .A(__tmp_495_2), .Y(_05756_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34837_ ( .A({ __tmp_495_2[0], __tmp_495_2[1] }), .Y(_05757_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34838_ ( .A({ __tmp_505_2[0], __tmp_505_2[1] }), .Y(_05758_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34839_ ( .A(__tmp_505_2), .Y(_05759_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34840_ ( .A({ __tmp_505_2[0], __tmp_505_2[1] }), .Y(_05760_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34841_ ( .A({ __tmp_515_2[0], __tmp_515_2[1] }), .Y(_05761_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34842_ ( .A(__tmp_515_2), .Y(_05762_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34843_ ( .A({ __tmp_515_2[0], __tmp_515_2[1] }), .Y(_05763_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34844_ ( .A({ __tmp_525_2[0], __tmp_525_2[1] }), .Y(_05764_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34845_ ( .A(__tmp_525_2), .Y(_05765_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34846_ ( .A({ __tmp_525_2[0], __tmp_525_2[1] }), .Y(_05766_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34847_ ( .A({ __tmp_535_2[0], __tmp_535_2[1] }), .Y(_05767_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34848_ ( .A(__tmp_535_2), .Y(_05768_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34849_ ( .A({ __tmp_535_2[0], __tmp_535_2[1] }), .Y(_05769_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34850_ ( .A({ __tmp_545_2[0], __tmp_545_2[1] }), .Y(_05770_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34851_ ( .A(__tmp_545_2), .Y(_05771_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34852_ ( .A({ __tmp_545_2[0], __tmp_545_2[1] }), .Y(_05772_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34853_ ( .A({ __tmp_555_2[0], __tmp_555_2[1] }), .Y(_05773_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34854_ ( .A(__tmp_555_2), .Y(_05774_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34855_ ( .A({ __tmp_555_2[0], __tmp_555_2[1] }), .Y(_05775_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34856_ ( .A({ __tmp_565_2[0], __tmp_565_2[1] }), .Y(_05776_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34857_ ( .A(__tmp_565_2), .Y(_05777_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34858_ ( .A({ __tmp_565_2[0], __tmp_565_2[1] }), .Y(_05778_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34859_ ( .A({ __tmp_575_2[0], __tmp_575_2[1] }), .Y(_05779_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34860_ ( .A(__tmp_575_2), .Y(_05780_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34861_ ( .A({ __tmp_575_2[0], __tmp_575_2[1] }), .Y(_05781_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34862_ ( .A({ __tmp_585_2[0], __tmp_585_2[1], __tmp_585_2[2] }), .Y(_05782_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34863_ ( .A({ __tmp_585_2[1:0], __tmp_585_2[2] }), .Y(_05783_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34864_ ( .A({ __tmp_585_2[1:0], __tmp_585_2[2] }), .Y(_05784_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34865_ ( .A(__tmp_585_2), .Y(_05785_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34866_ ( .A({ __tmp_585_2[2], __tmp_585_2[0], __tmp_585_2[1] }), .Y(_05786_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34867_ ( .A({ __tmp_585_2[1], __tmp_585_2[2], __tmp_585_2[0] }), .Y(_05787_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34868_ ( .A({ __tmp_585_2[1:0], __tmp_585_2[2] }), .Y(_05788_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34869_ ( .A({ __tmp_599_2[0], __tmp_599_2[1], __tmp_599_2[2] }), .Y(_05789_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34870_ ( .A({ __tmp_599_2[1:0], __tmp_599_2[2] }), .Y(_05790_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34871_ ( .A({ __tmp_599_2[1:0], __tmp_599_2[2] }), .Y(_05791_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34872_ ( .A(__tmp_599_2), .Y(_05792_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34873_ ( .A({ __tmp_599_2[2], __tmp_599_2[0], __tmp_599_2[1] }), .Y(_05793_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34874_ ( .A({ __tmp_599_2[1], __tmp_599_2[2], __tmp_599_2[0] }), .Y(_05794_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34875_ ( .A({ __tmp_599_2[1:0], __tmp_599_2[2] }), .Y(_05795_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34876_ ( .A({ __tmp_613_2[0], __tmp_613_2[1], __tmp_613_2[2] }), .Y(_05796_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34877_ ( .A({ __tmp_613_2[1:0], __tmp_613_2[2] }), .Y(_05797_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34878_ ( .A({ __tmp_613_2[1:0], __tmp_613_2[2] }), .Y(_05798_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34879_ ( .A(__tmp_613_2), .Y(_05799_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34880_ ( .A({ __tmp_613_2[2], __tmp_613_2[0], __tmp_613_2[1] }), .Y(_05800_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34881_ ( .A({ __tmp_613_2[1], __tmp_613_2[2], __tmp_613_2[0] }), .Y(_05801_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34882_ ( .A({ __tmp_613_2[1:0], __tmp_613_2[2] }), .Y(_05802_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34883_ ( .A({ __tmp_627_2[0], __tmp_627_2[1], __tmp_627_2[2] }), .Y(_05803_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34884_ ( .A({ __tmp_627_2[1:0], __tmp_627_2[2] }), .Y(_05804_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34885_ ( .A({ __tmp_627_2[1:0], __tmp_627_2[2] }), .Y(_05805_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34886_ ( .A(__tmp_627_2), .Y(_05806_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34887_ ( .A({ __tmp_627_2[2], __tmp_627_2[0], __tmp_627_2[1] }), .Y(_05807_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34888_ ( .A({ __tmp_627_2[1], __tmp_627_2[2], __tmp_627_2[0] }), .Y(_05808_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34889_ ( .A({ __tmp_627_2[1:0], __tmp_627_2[2] }), .Y(_05809_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34890_ ( .A({ __tmp_641_2[0], __tmp_641_2[1], __tmp_641_2[2] }), .Y(_05810_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34891_ ( .A({ __tmp_641_2[1:0], __tmp_641_2[2] }), .Y(_05811_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34892_ ( .A({ __tmp_641_2[1:0], __tmp_641_2[2] }), .Y(_05812_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34893_ ( .A(__tmp_641_2), .Y(_05813_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34894_ ( .A({ __tmp_641_2[2], __tmp_641_2[0], __tmp_641_2[1] }), .Y(_05814_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34895_ ( .A({ __tmp_641_2[1], __tmp_641_2[2], __tmp_641_2[0] }), .Y(_05815_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34896_ ( .A({ __tmp_641_2[1:0], __tmp_641_2[2] }), .Y(_05816_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34897_ ( .A({ __tmp_655_2[0], __tmp_655_2[1], __tmp_655_2[2] }), .Y(_05817_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34898_ ( .A({ __tmp_655_2[1:0], __tmp_655_2[2] }), .Y(_05818_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34899_ ( .A({ __tmp_655_2[1:0], __tmp_655_2[2] }), .Y(_05819_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34900_ ( .A(__tmp_655_2), .Y(_05820_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34901_ ( .A({ __tmp_655_2[2], __tmp_655_2[0], __tmp_655_2[1] }), .Y(_05821_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34902_ ( .A({ __tmp_655_2[1], __tmp_655_2[2], __tmp_655_2[0] }), .Y(_05822_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34903_ ( .A({ __tmp_655_2[1:0], __tmp_655_2[2] }), .Y(_05823_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34904_ ( .A({ __tmp_669_2[0], __tmp_669_2[1], __tmp_669_2[2] }), .Y(_05824_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34905_ ( .A({ __tmp_669_2[1:0], __tmp_669_2[2] }), .Y(_05825_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34906_ ( .A({ __tmp_669_2[1:0], __tmp_669_2[2] }), .Y(_05826_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34907_ ( .A(__tmp_669_2), .Y(_05827_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34908_ ( .A({ __tmp_669_2[2], __tmp_669_2[0], __tmp_669_2[1] }), .Y(_05828_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34909_ ( .A({ __tmp_669_2[1], __tmp_669_2[2], __tmp_669_2[0] }), .Y(_05829_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34910_ ( .A({ __tmp_669_2[1:0], __tmp_669_2[2] }), .Y(_05830_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34911_ ( .A({ __tmp_683_2[0], __tmp_683_2[1], __tmp_683_2[2] }), .Y(_05831_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34912_ ( .A({ __tmp_683_2[1:0], __tmp_683_2[2] }), .Y(_05832_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34913_ ( .A({ __tmp_683_2[1:0], __tmp_683_2[2] }), .Y(_05833_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34914_ ( .A(__tmp_683_2), .Y(_05834_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34915_ ( .A({ __tmp_683_2[2], __tmp_683_2[0], __tmp_683_2[1] }), .Y(_05835_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34916_ ( .A({ __tmp_683_2[1], __tmp_683_2[2], __tmp_683_2[0] }), .Y(_05836_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34917_ ( .A({ __tmp_683_2[1:0], __tmp_683_2[2] }), .Y(_05837_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34918_ ( .A({ __tmp_697_2[0], __tmp_697_2[1], __tmp_697_2[2] }), .Y(_05838_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34919_ ( .A({ __tmp_697_2[1:0], __tmp_697_2[2] }), .Y(_05839_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34920_ ( .A({ __tmp_697_2[1:0], __tmp_697_2[2] }), .Y(_05840_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34921_ ( .A(__tmp_697_2), .Y(_05841_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34922_ ( .A({ __tmp_697_2[2], __tmp_697_2[0], __tmp_697_2[1] }), .Y(_05842_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34923_ ( .A({ __tmp_697_2[1], __tmp_697_2[2], __tmp_697_2[0] }), .Y(_05843_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34924_ ( .A({ __tmp_697_2[1:0], __tmp_697_2[2] }), .Y(_05844_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34925_ ( .A({ conv2d_16_row_select[0], conv2d_16_row_select[1] }), .Y(_05845_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34926_ ( .A(conv2d_16_row_select), .Y(_05846_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34927_ ( .A({ __tmp_1027_2[0], __tmp_1027_2[1] }), .Y(_05847_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34928_ ( .A(__tmp_1027_2), .Y(_05848_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34929_ ( .A({ __tmp_1027_2[0], __tmp_1027_2[1] }), .Y(_05849_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34930_ ( .A({ __tmp_1170_2[0], __tmp_1170_2[1] }), .Y(_05850_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34931_ ( .A(__tmp_1170_2), .Y(_05851_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34932_ ( .A({ __tmp_1170_2[0], __tmp_1170_2[1] }), .Y(_05852_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34933_ ( .A({ __tmp_1181_2[0], __tmp_1181_2[1] }), .Y(_05853_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34934_ ( .A(__tmp_1181_2), .Y(_05854_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34935_ ( .A({ __tmp_1181_2[0], __tmp_1181_2[1] }), .Y(_05855_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34936_ ( .A({ __tmp_1201_2[0], __tmp_1201_2[1] }), .Y(_05856_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _34937_ ( .A(__tmp_1201_2), .Y(_05857_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34938_ ( .A({ __tmp_1201_2[0], __tmp_1201_2[1] }), .Y(_05858_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34939_ ( .A({ __tmp_1211_2[0], __tmp_1211_2[1], __tmp_1211_2[2] }), .Y(_05859_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34940_ ( .A({ __tmp_1211_2[1:0], __tmp_1211_2[2] }), .Y(_05860_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34941_ ( .A({ __tmp_1211_2[1:0], __tmp_1211_2[2] }), .Y(_05861_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34942_ ( .A(__tmp_1211_2), .Y(_05862_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34943_ ( .A({ __tmp_1211_2[2], __tmp_1211_2[0], __tmp_1211_2[1] }), .Y(_05863_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34944_ ( .A({ __tmp_1211_2[1], __tmp_1211_2[2], __tmp_1211_2[0] }), .Y(_05864_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34945_ ( .A({ __tmp_1211_2[1:0], __tmp_1211_2[2] }), .Y(_05865_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34946_ ( .A({ _10023_, _tmp_5[0], _tmp_5[1] }), .Y(_05866_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _34947_ ( .A(_tmp_5[3:2]), .Y(_10023_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34948_ ( .A({ _tmp_5[1], _10023_, _tmp_5[0] }), .Y(_05867_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34949_ ( .A({ _tmp_5[1:0], _10023_ }), .Y(_05868_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34950_ ( .A({ _10024_, _tmp_5[1:0] }), .Y(_05869_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34951_ ( .A({ _tmp_5[2], _tmp_5[3] }), .Y(_10024_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34952_ ( .A({ _10024_, _tmp_5[0], _tmp_5[1] }), .Y(_05870_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34953_ ( .A({ _tmp_5[1], _10024_, _tmp_5[0] }), .Y(_05871_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34954_ ( .A({ _tmp_5[1:0], _10024_ }), .Y(_05872_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _34955_ ( .A({ _10025_, _tmp_5[1:0] }), .Y(_05873_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _34956_ ( .A(_tmp_5[3:2]), .Y(_10025_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34957_ ( .A({ _10025_, _tmp_5[0], _tmp_5[1] }), .Y(_05874_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _34958_ ( .A({ _tmp_5[1], _10025_, _tmp_5[0] }), .Y(_05875_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _34959_ ( .A({ _tmp_5[1:0], _10025_ }), .Y(_05876_) );
  \$lut  #( .LUT(16'hefff), .WIDTH(4) ) _34960_ ( .A(_tmp_5), .Y(_05877_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _34961_ ( .A({ _tmp_5[2], _tmp_5[0], _tmp_5[3], _tmp_5[1] }), .Y(_05878_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34962_ ( .A({ _10027_, _10026_ }), .Y(_05879_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34963_ ( .A({ _stream_conv2d_16_source_28_source_ram_sel[3:2], _stream_conv2d_16_source_28_source_ram_sel[7:6] }), .Y(_10026_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34964_ ( .A({ _stream_conv2d_16_source_28_source_ram_sel[5:4], _stream_conv2d_16_source_28_source_ram_sel[1:0] }), .Y(_10027_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34965_ ( .A({ _10029_, _10028_ }), .Y(_05880_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34966_ ( .A({ _stream_matmul_29_source_20_source_ram_sel[2], _stream_matmul_29_source_20_source_ram_sel[7:5] }), .Y(_10028_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34967_ ( .A({ _stream_matmul_29_source_20_source_ram_sel[4:3], _stream_matmul_29_source_20_source_ram_sel[1:0] }), .Y(_10029_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34968_ ( .A({ _10031_, _10030_ }), .Y(_05881_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34969_ ( .A({ _stream_conv2d_16_source_29_source_ram_sel[3:2], _stream_conv2d_16_source_29_source_ram_sel[0], _stream_conv2d_16_source_29_source_ram_sel[7] }), .Y(_10030_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34970_ ( .A({ _stream_conv2d_16_source_29_source_ram_sel[6:4], _stream_conv2d_16_source_29_source_ram_sel[1] }), .Y(_10031_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34971_ ( .A({ _10033_, _10032_ }), .Y(_05882_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34972_ ( .A({ _stream_conv2d_16_source_30_source_ram_sel[3:1], _stream_conv2d_16_source_30_source_ram_sel[7] }), .Y(_10032_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34973_ ( .A({ _stream_conv2d_16_source_30_source_ram_sel[6:4], _stream_conv2d_16_source_30_source_ram_sel[0] }), .Y(_10033_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34974_ ( .A({ _10035_, _10034_ }), .Y(_05883_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _34975_ ( .A(_stream_conv2d_16_source_31_source_ram_sel[3:0]), .Y(_10034_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34976_ ( .A(_stream_conv2d_16_source_31_source_ram_sel[7:4]), .Y(_10035_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34977_ ( .A({ _10037_, _10036_ }), .Y(_05884_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34978_ ( .A({ _stream_conv2d_16_source_32_source_ram_sel[4], _stream_conv2d_16_source_32_source_ram_sel[7:5] }), .Y(_10036_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34979_ ( .A(_stream_conv2d_16_source_32_source_ram_sel[3:0]), .Y(_10037_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34980_ ( .A({ _10039_, _10038_ }), .Y(_05885_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34981_ ( .A({ _stream_conv2d_16_source_33_source_ram_sel[4], _stream_conv2d_16_source_33_source_ram_sel[0], _stream_conv2d_16_source_33_source_ram_sel[7:6] }), .Y(_10038_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34982_ ( .A({ _stream_conv2d_16_source_33_source_ram_sel[5], _stream_conv2d_16_source_33_source_ram_sel[3:1] }), .Y(_10039_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34983_ ( .A({ _10041_, _10040_ }), .Y(_05886_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34984_ ( .A({ _stream_conv2d_16_source_34_source_ram_sel[4], _stream_conv2d_16_source_34_source_ram_sel[1], _stream_conv2d_16_source_34_source_ram_sel[7:6] }), .Y(_10040_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34985_ ( .A({ _stream_conv2d_16_source_34_source_ram_sel[5], _stream_conv2d_16_source_34_source_ram_sel[3:2], _stream_conv2d_16_source_34_source_ram_sel[0] }), .Y(_10041_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34986_ ( .A({ _10043_, _10042_ }), .Y(_05887_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _34987_ ( .A({ _stream_conv2d_16_source_35_source_ram_sel[4], _stream_conv2d_16_source_35_source_ram_sel[1:0], _stream_conv2d_16_source_35_source_ram_sel[7] }), .Y(_10042_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34988_ ( .A({ _stream_conv2d_16_source_35_source_ram_sel[6:5], _stream_conv2d_16_source_35_source_ram_sel[3:2] }), .Y(_10043_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34989_ ( .A({ _10045_, _10044_ }), .Y(_05888_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _34990_ ( .A({ _stream_conv2d_16_source_36_source_ram_sel[4], _stream_conv2d_16_source_36_source_ram_sel[2], _stream_conv2d_16_source_36_source_ram_sel[7:6] }), .Y(_10044_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34991_ ( .A({ _stream_conv2d_16_source_36_source_ram_sel[5], _stream_conv2d_16_source_36_source_ram_sel[3], _stream_conv2d_16_source_36_source_ram_sel[1:0] }), .Y(_10045_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34992_ ( .A({ _10047_, _10046_ }), .Y(_05889_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34993_ ( .A({ _stream_conv2d_16_source_8_source_ram_sel[1], _stream_conv2d_16_source_8_source_ram_sel[7:5] }), .Y(_10046_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34994_ ( .A({ _stream_conv2d_16_source_8_source_ram_sel[4:2], _stream_conv2d_16_source_8_source_ram_sel[0] }), .Y(_10047_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34995_ ( .A({ _10049_, _10048_ }), .Y(_05890_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34996_ ( .A({ _stream_matmul_29_source_8_source_ram_sel[1], _stream_matmul_29_source_8_source_ram_sel[7:5] }), .Y(_10048_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _34997_ ( .A({ _stream_matmul_29_source_8_source_ram_sel[4:2], _stream_matmul_29_source_8_source_ram_sel[0] }), .Y(_10049_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _34998_ ( .A({ _10051_, _10050_ }), .Y(_05891_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _34999_ ( .A({ _stream_conv2d_16_source_6_source_ram_sel[0], _stream_conv2d_16_source_6_source_ram_sel[7:5] }), .Y(_10050_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35000_ ( .A(_stream_conv2d_16_source_6_source_ram_sel[4:1]), .Y(_10051_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35001_ ( .A({ _10053_, _10052_ }), .Y(_05892_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35002_ ( .A({ _stream_max_pool_serial_18_source_1_source_ram_sel[0], _stream_max_pool_serial_18_source_1_source_ram_sel[7:5] }), .Y(_10052_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35003_ ( .A(_stream_max_pool_serial_18_source_1_source_ram_sel[4:1]), .Y(_10053_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35004_ ( .A({ _10055_, _10054_ }), .Y(_05893_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35005_ ( .A({ _stream_conv2d_16_source_19_source_ram_sel[1:0], _stream_conv2d_16_source_19_source_ram_sel[7:6] }), .Y(_10054_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35006_ ( .A(_stream_conv2d_16_source_19_source_ram_sel[5:2]), .Y(_10055_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35007_ ( .A({ _10057_, _10056_ }), .Y(_05894_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35008_ ( .A({ _stream_matmul_29_source_6_source_ram_sel[0], _stream_matmul_29_source_6_source_ram_sel[7:5] }), .Y(_10056_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35009_ ( .A(_stream_matmul_29_source_6_source_ram_sel[4:1]), .Y(_10057_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35010_ ( .A({ _10059_, _10058_ }), .Y(_05895_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35011_ ( .A({ _stream_conv2d_16_source_20_source_ram_sel[2], _stream_conv2d_16_source_20_source_ram_sel[7:5] }), .Y(_10058_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35012_ ( .A({ _stream_conv2d_16_source_20_source_ram_sel[4:3], _stream_conv2d_16_source_20_source_ram_sel[1:0] }), .Y(_10059_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35013_ ( .A({ _10061_, _10060_ }), .Y(_05896_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35014_ ( .A({ _stream_matmul_29_source_19_source_ram_sel[1:0], _stream_matmul_29_source_19_source_ram_sel[7:6] }), .Y(_10060_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35015_ ( .A(_stream_matmul_29_source_19_source_ram_sel[5:2]), .Y(_10061_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35016_ ( .A({ _10063_, _10062_ }), .Y(_05897_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35017_ ( .A({ _stream_conv2d_16_source_21_source_ram_sel[2], _stream_conv2d_16_source_21_source_ram_sel[0], _stream_conv2d_16_source_21_source_ram_sel[7:6] }), .Y(_10062_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35018_ ( .A({ _stream_conv2d_16_source_21_source_ram_sel[5:3], _stream_conv2d_16_source_21_source_ram_sel[1] }), .Y(_10063_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35019_ ( .A({ _10065_, _10064_ }), .Y(_05898_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35020_ ( .A({ _stream_conv2d_16_source_22_source_ram_sel[2:1], _stream_conv2d_16_source_22_source_ram_sel[7:6] }), .Y(_10064_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35021_ ( .A({ _stream_conv2d_16_source_22_source_ram_sel[5:3], _stream_conv2d_16_source_22_source_ram_sel[0] }), .Y(_10065_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35022_ ( .A({ _10067_, _10066_ }), .Y(_05899_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35023_ ( .A({ _stream_conv2d_16_source_23_source_ram_sel[2:0], _stream_conv2d_16_source_23_source_ram_sel[7] }), .Y(_10066_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35024_ ( .A(_stream_conv2d_16_source_23_source_ram_sel[6:3]), .Y(_10067_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35025_ ( .A({ _10069_, _10068_ }), .Y(_05900_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35026_ ( .A({ _stream_conv2d_16_source_24_source_ram_sel[3], _stream_conv2d_16_source_24_source_ram_sel[7:5] }), .Y(_10068_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35027_ ( .A({ _stream_conv2d_16_source_24_source_ram_sel[4], _stream_conv2d_16_source_24_source_ram_sel[2:0] }), .Y(_10069_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35028_ ( .A({ _10071_, _10070_ }), .Y(_05901_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35029_ ( .A({ _stream_conv2d_16_source_25_source_ram_sel[3], _stream_conv2d_16_source_25_source_ram_sel[0], _stream_conv2d_16_source_25_source_ram_sel[7:6] }), .Y(_10070_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35030_ ( .A({ _stream_conv2d_16_source_25_source_ram_sel[5:4], _stream_conv2d_16_source_25_source_ram_sel[2:1] }), .Y(_10071_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35031_ ( .A({ _10073_, _10072_ }), .Y(_05902_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35032_ ( .A({ _stream_conv2d_16_source_26_source_ram_sel[3], _stream_conv2d_16_source_26_source_ram_sel[1], _stream_conv2d_16_source_26_source_ram_sel[7:6] }), .Y(_10072_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35033_ ( .A({ _stream_conv2d_16_source_26_source_ram_sel[5:4], _stream_conv2d_16_source_26_source_ram_sel[2], _stream_conv2d_16_source_26_source_ram_sel[0] }), .Y(_10073_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35034_ ( .A({ _10075_, _10074_ }), .Y(_05903_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35035_ ( .A({ _stream_conv2d_16_source_27_source_ram_sel[3], _stream_conv2d_16_source_27_source_ram_sel[1:0], _stream_conv2d_16_source_27_source_ram_sel[7] }), .Y(_10074_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35036_ ( .A({ _stream_conv2d_16_source_27_source_ram_sel[6:4], _stream_conv2d_16_source_27_source_ram_sel[2] }), .Y(_10075_) );
  \$lut  #( .LUT(16'hefff), .WIDTH(4) ) _35037_ ( .A({ cparam_conv2d_16_bias_num[0], _10076_, cparam_conv2d_16_bias_num[6:5] }), .Y(_05904_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35038_ ( .A(cparam_conv2d_16_bias_num[4:1]), .Y(_10076_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _35039_ ( .A({ _10077_, cparam_matmul_29_bias_num[5:4] }), .Y(_05905_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35040_ ( .A({ cparam_matmul_29_bias_num[0], _10078_, cparam_matmul_29_bias_num[8:7] }), .Y(_10077_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35041_ ( .A({ cparam_matmul_29_bias_num[6], cparam_matmul_29_bias_num[3:1] }), .Y(_10078_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35042_ ( .A({ _10084_, _10079_ }), .Y(_06885_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35043_ ( .A({ _10083_, _10082_, _10081_, _10080_ }), .Y(_10079_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35044_ ( .A(_saxi_register_4[23:20]), .Y(_10080_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35045_ ( .A(_saxi_register_4[19:16]), .Y(_10081_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35046_ ( .A(_saxi_register_4[31:28]), .Y(_10082_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35047_ ( .A(_saxi_register_4[27:24]), .Y(_10083_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35048_ ( .A({ _10088_, _10087_, _10086_, _10085_ }), .Y(_10084_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35049_ ( .A(_saxi_register_4[7:4]), .Y(_10085_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35050_ ( .A(_saxi_register_4[3:0]), .Y(_10086_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35051_ ( .A(_saxi_register_4[15:12]), .Y(_10087_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35052_ ( .A(_saxi_register_4[11:8]), .Y(_10088_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35053_ ( .A({ _10094_, _10089_ }), .Y(_19569_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35054_ ( .A({ _10093_, _10092_, _10091_, _10090_ }), .Y(_10089_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35055_ ( .A({ _24115_, _24114_, _24113_, _24112_ }), .Y(_10090_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35056_ ( .A({ _24110_, _24109_, _24108_, _24107_ }), .Y(_10091_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35057_ ( .A({ _24124_, _24123_, _24121_, _24120_ }), .Y(_10092_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35058_ ( .A({ _24119_, _24118_, _24117_, _24116_ }), .Y(_10093_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35059_ ( .A({ _10098_, _10097_, _10096_, _10095_ }), .Y(_10094_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35060_ ( .A({ _24129_, _24128_, _24127_, _24126_ }), .Y(_10095_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35061_ ( .A({ _24125_, _24122_, _24111_, _24100_ }), .Y(_10096_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35062_ ( .A({ _24106_, _24105_, _24104_, _24103_ }), .Y(_10097_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35063_ ( .A({ _24102_, _24101_, _24131_, _24130_ }), .Y(_10098_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35064_ ( .A({ _10104_, _10099_ }), .Y(_19504_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35065_ ( .A({ _10103_, _10102_, _10101_, _10100_ }), .Y(_10099_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35066_ ( .A({ _24147_, _24146_, _24145_, _24144_ }), .Y(_10100_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35067_ ( .A({ _24142_, _24141_, _24140_, _24139_ }), .Y(_10101_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35068_ ( .A({ _24156_, _24155_, _24153_, _24152_ }), .Y(_10102_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35069_ ( .A({ _24151_, _24150_, _24149_, _24148_ }), .Y(_10103_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35070_ ( .A({ _10108_, _10107_, _10106_, _10105_ }), .Y(_10104_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35071_ ( .A({ _24161_, _24160_, _24159_, _24158_ }), .Y(_10105_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35072_ ( .A({ _24157_, _24154_, _24143_, _24132_ }), .Y(_10106_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35073_ ( .A({ _24138_, _24137_, _24136_, _24135_ }), .Y(_10107_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35074_ ( .A({ _24134_, _24133_, _24163_, _24162_ }), .Y(_10108_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _35075_ ( .A({ conv2d_16_col_select[0], conv2d_16_col_select[1] }), .Y(_05906_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _35076_ ( .A(conv2d_16_col_select), .Y(_05907_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35077_ ( .A({ _10114_, _10109_ }), .Y(_19439_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35078_ ( .A({ _10113_, _10112_, _10111_, _10110_ }), .Y(_10109_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35079_ ( .A({ _24179_, _24178_, _24177_, _24176_ }), .Y(_10110_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35080_ ( .A({ _24174_, _24173_, _24172_, _24171_ }), .Y(_10111_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35081_ ( .A({ _24188_, _24187_, _24185_, _24184_ }), .Y(_10112_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35082_ ( .A({ _24183_, _24182_, _24181_, _24180_ }), .Y(_10113_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35083_ ( .A({ _10118_, _10117_, _10116_, _10115_ }), .Y(_10114_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35084_ ( .A({ _24193_, _24192_, _24191_, _24190_ }), .Y(_10115_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35085_ ( .A({ _24189_, _24186_, _24175_, _24164_ }), .Y(_10116_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35086_ ( .A({ _24170_, _24169_, _24168_, _24167_ }), .Y(_10117_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35087_ ( .A({ _24166_, _24165_, _24195_, _24194_ }), .Y(_10118_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35088_ ( .A({ _stream_matmul_29_source_20_source_pat_fsm_3[0], _09209_ }), .Y(_05909_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35089_ ( .A({ _stream_matmul_29_source_19_source_pat_fsm_2[1], _09220_ }), .Y(_05910_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35090_ ( .A({ _stream_matmul_29_source_8_source_pat_fsm_1[1], _09185_ }), .Y(_05914_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35091_ ( .A({ _stream_matmul_29_source_6_source_pat_fsm_0[1], _09172_ }), .Y(_05915_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _35092_ ( .A({ _10128_, _10127_, _10124_, _10119_ }), .Y(_05918_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35093_ ( .A({ _10123_, _10122_, _10121_, _10120_ }), .Y(_10119_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35094_ ( .A(_d1_control_matmul_29[23:20]), .Y(_10120_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35095_ ( .A(_d1_control_matmul_29[19:16]), .Y(_10121_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35096_ ( .A(_d1_control_matmul_29[31:28]), .Y(_10122_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35097_ ( .A(_d1_control_matmul_29[27:24]), .Y(_10123_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35098_ ( .A({ _10126_, _10125_ }), .Y(_10124_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35099_ ( .A(_d1_control_matmul_29[15:12]), .Y(_10125_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35100_ ( .A(_d1_control_matmul_29[11:8]), .Y(_10126_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35101_ ( .A({ _d1_control_matmul_29[5], _d1_control_matmul_29[1:0], _d1_control_matmul_29[4] }), .Y(_10127_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35102_ ( .A({ _d1_control_matmul_29[7:6], _d1_control_matmul_29[2], _d1_control_matmul_29[3] }), .Y(_10128_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _35103_ ( .A({ _10130_, _10119_, _10129_ }), .Y(_05919_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35104_ ( .A({ _d1_control_matmul_29[2:1], _10124_, _d1_control_matmul_29[0] }), .Y(_10129_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _35105_ ( .A({ _10131_, _d1_control_matmul_29[4:3] }), .Y(_10130_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _35106_ ( .A(_d1_control_matmul_29[7:5]), .Y(_10131_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35107_ ( .A({ _10132_, _10129_ }), .Y(_05921_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35108_ ( .A({ _d1_control_matmul_29[3], _10133_, _10119_ }), .Y(_10132_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35109_ ( .A({ _10131_, _d1_control_matmul_29[4] }), .Y(_10133_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35110_ ( .A({ _10134_, _10132_ }), .Y(_05922_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35111_ ( .A({ _10124_, _d1_control_matmul_29[2:0] }), .Y(_10134_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _35112_ ( .A({ _10135_, _10133_, _10124_, _10119_ }), .Y(_05923_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35113_ ( .A({ _d1_control_matmul_29[0], _d1_control_matmul_29[1], _d1_control_matmul_29[2], _d1_control_matmul_29[3] }), .Y(_10135_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _35114_ ( .A({ _08038_, _08090_, control_matmul_29[1] }), .Y(_05925_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35115_ ( .A({ control_matmul_29[1], _08081_ }), .Y(_05927_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _35116_ ( .A({ _08081_, control_matmul_29[1] }), .Y(_05930_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _35117_ ( .A({ _10145_, _10140_, _10136_ }), .Y(_05938_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35118_ ( .A({ _d1_control_max_pool_serial_18[0], _d1_control_max_pool_serial_18[1], _10137_, _d1_control_max_pool_serial_18[2] }), .Y(_10136_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35119_ ( .A({ _10139_, _10138_ }), .Y(_10137_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35120_ ( .A(_d1_control_max_pool_serial_18[15:12]), .Y(_10138_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35121_ ( .A(_d1_control_max_pool_serial_18[11:8]), .Y(_10139_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35122_ ( .A({ _10144_, _10143_, _10142_, _10141_ }), .Y(_10140_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35123_ ( .A(_d1_control_max_pool_serial_18[23:20]), .Y(_10141_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35124_ ( .A(_d1_control_max_pool_serial_18[19:16]), .Y(_10142_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35125_ ( .A(_d1_control_max_pool_serial_18[31:28]), .Y(_10143_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35126_ ( .A(_d1_control_max_pool_serial_18[27:24]), .Y(_10144_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _35127_ ( .A({ _10146_, _d1_control_max_pool_serial_18[7:6] }), .Y(_10145_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _35128_ ( .A({ _d1_control_max_pool_serial_18[4], _d1_control_max_pool_serial_18[5], _d1_control_max_pool_serial_18[3] }), .Y(_10146_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _35129_ ( .A({ _d1_control_max_pool_serial_18[3], _10147_, _10140_, _10136_ }), .Y(_05939_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35130_ ( .A({ _d1_control_max_pool_serial_18[7:6], _d1_control_max_pool_serial_18[4], _d1_control_max_pool_serial_18[5] }), .Y(_10147_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _35131_ ( .A({ _10148_, _10147_, _10137_, _10140_ }), .Y(_05940_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35132_ ( .A({ _d1_control_max_pool_serial_18[0], _d1_control_max_pool_serial_18[2:1], _d1_control_max_pool_serial_18[3] }), .Y(_10148_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _35133_ ( .A({ _07082_, _07080_, _07070_ }), .Y(_05941_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35134_ ( .A({ _07080_, _07095_ }), .Y(_05943_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35135_ ( .A({ _07091_, _07092_ }), .Y(_05944_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35136_ ( .A({ _10154_, _10149_ }), .Y(_05946_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35137_ ( .A({ _10153_, _10152_, _10151_, _10150_ }), .Y(_10149_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35138_ ( .A(_d1__maxi_write_fsm[24:21]), .Y(_10150_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35139_ ( .A(_d1__maxi_write_fsm[20:17]), .Y(_10151_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35140_ ( .A({ _d1__maxi_write_fsm[2], _d1__maxi_write_fsm[31:29] }), .Y(_10152_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35141_ ( .A(_d1__maxi_write_fsm[28:25]), .Y(_10153_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35142_ ( .A({ _10158_, _10157_, _10156_, _10155_ }), .Y(_10154_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35143_ ( .A(_d1__maxi_write_fsm[8:5]), .Y(_10155_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35144_ ( .A({ _d1__maxi_write_fsm[4:3], _d1__maxi_write_fsm[1:0] }), .Y(_10156_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35145_ ( .A(_d1__maxi_write_fsm[16:13]), .Y(_10157_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35146_ ( .A(_d1__maxi_write_fsm[12:9]), .Y(_10158_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35147_ ( .A({ _stream_conv2d_16_source_36_source_pat_fsm_19[1], _06970_ }), .Y(_05950_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35148_ ( .A({ _stream_conv2d_16_source_35_source_pat_fsm_18[1], _06983_ }), .Y(_05951_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35149_ ( .A({ _stream_conv2d_16_source_34_source_pat_fsm_17[1], _06958_ }), .Y(_05953_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35150_ ( .A({ _stream_conv2d_16_source_33_source_pat_fsm_16[1], _06946_ }), .Y(_05955_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35151_ ( .A({ _stream_conv2d_16_source_32_source_pat_fsm_15[1], _06934_ }), .Y(_05957_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35152_ ( .A({ _stream_conv2d_16_source_31_source_pat_fsm_14[1], _09933_ }), .Y(_05958_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35153_ ( .A({ _stream_conv2d_16_source_30_source_pat_fsm_13[1], _09817_ }), .Y(_05961_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35154_ ( .A({ _stream_conv2d_16_source_29_source_pat_fsm_12[1], _09805_ }), .Y(_05963_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35155_ ( .A({ _stream_conv2d_16_source_28_source_pat_fsm_11[1], _09475_ }), .Y(_05964_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35156_ ( .A({ _stream_conv2d_16_source_27_source_pat_fsm_10[0], _06995_ }), .Y(_05968_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35157_ ( .A({ _stream_conv2d_16_source_26_source_pat_fsm_9[0], _08878_ }), .Y(_05971_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35158_ ( .A({ _stream_conv2d_16_source_24_source_pat_fsm_7[0], _09252_ }), .Y(_05972_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35159_ ( .A({ _stream_conv2d_16_source_25_source_pat_fsm_8[0], _09241_ }), .Y(_05974_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35160_ ( .A({ _stream_conv2d_16_source_23_source_pat_fsm_6[0], _09371_ }), .Y(_05977_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35161_ ( .A({ _stream_conv2d_16_source_22_source_pat_fsm_5[0], _07793_ }), .Y(_05979_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35162_ ( .A({ _stream_conv2d_16_source_21_source_pat_fsm_4[0], _07879_ }), .Y(_05981_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35163_ ( .A({ _stream_conv2d_16_source_20_source_pat_fsm_3[0], _09263_ }), .Y(_05982_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35164_ ( .A({ _stream_conv2d_16_source_19_source_pat_fsm_2[0], _09768_ }), .Y(_05983_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35165_ ( .A({ _stream_conv2d_16_source_8_source_pat_fsm_1[0], _09794_ }), .Y(_05986_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35166_ ( .A({ _10167_, _10159_ }), .Y(_05992_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35167_ ( .A({ _10160_, _10166_, _10165_, _d1__maxi_read_fsm[3] }), .Y(_10159_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35168_ ( .A({ _10164_, _10163_, _10162_, _10161_ }), .Y(_10160_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35169_ ( .A({ _d1__maxi_read_fsm[22:21], _d1__maxi_read_fsm[19], _d1__maxi_read_fsm[16] }), .Y(_10161_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35170_ ( .A({ _d1__maxi_read_fsm[31], _d1__maxi_read_fsm[28], _d1__maxi_read_fsm[26:25] }), .Y(_10162_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35171_ ( .A({ _d1__maxi_read_fsm[23], _d1__maxi_read_fsm[20], _d1__maxi_read_fsm[18:17] }), .Y(_10163_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35172_ ( .A({ _d1__maxi_read_fsm[30:29], _d1__maxi_read_fsm[27], _d1__maxi_read_fsm[24] }), .Y(_10164_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35173_ ( .A({ _d1__maxi_read_fsm[15], _d1__maxi_read_fsm[13], _d1__maxi_read_fsm[11], _d1__maxi_read_fsm[9] }), .Y(_10165_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35174_ ( .A({ _d1__maxi_read_fsm[14], _d1__maxi_read_fsm[12], _d1__maxi_read_fsm[10], _d1__maxi_read_fsm[8] }), .Y(_10166_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35175_ ( .A({ _d1__maxi_read_fsm[2], _10168_, _d1__maxi_read_fsm[1:0] }), .Y(_10167_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35176_ ( .A(_d1__maxi_read_fsm[7:4]), .Y(_10168_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35177_ ( .A({ _10169_, _10159_ }), .Y(_05993_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35178_ ( .A({ _10168_, _d1__maxi_read_fsm[1:0], _d1__maxi_read_fsm[2] }), .Y(_10169_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _35179_ ( .A({ _d1_control_conv2d_16[5], _10179_, _10170_ }), .Y(_05997_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35180_ ( .A({ _d1_control_conv2d_16[4], _10176_, _10171_ }), .Y(_10170_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35181_ ( .A({ _10175_, _10174_, _10173_, _10172_ }), .Y(_10171_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35182_ ( .A(_d1_control_conv2d_16[23:20]), .Y(_10172_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35183_ ( .A(_d1_control_conv2d_16[19:16]), .Y(_10173_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35184_ ( .A(_d1_control_conv2d_16[31:28]), .Y(_10174_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35185_ ( .A(_d1_control_conv2d_16[27:24]), .Y(_10175_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35186_ ( .A({ _10178_, _10177_, _d1_control_conv2d_16[7:6] }), .Y(_10176_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35187_ ( .A(_d1_control_conv2d_16[15:12]), .Y(_10177_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35188_ ( .A(_d1_control_conv2d_16[11:8]), .Y(_10178_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _35189_ ( .A({ _10180_, _d1_control_conv2d_16[2], _d1_control_conv2d_16[3] }), .Y(_10179_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35190_ ( .A({ _d1_control_conv2d_16[0], _d1_control_conv2d_16[1] }), .Y(_10180_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _35191_ ( .A({ _10181_, _d1_control_conv2d_16[1:0] }), .Y(_05998_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35192_ ( .A({ _10183_, _10182_ }), .Y(_10181_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35193_ ( .A({ _10176_, _d1_control_conv2d_16[4] }), .Y(_10182_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35194_ ( .A({ _d1_control_conv2d_16[2], _d1_control_conv2d_16[5], _10171_, _d1_control_conv2d_16[3] }), .Y(_10183_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _35195_ ( .A({ _d1_control_conv2d_16[0], _10181_, _d1_control_conv2d_16[1] }), .Y(_05999_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _35196_ ( .A({ _d1_control_conv2d_16[2], _d1_control_conv2d_16[3], _10185_, _10184_ }), .Y(_06000_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35197_ ( .A({ _10170_, _d1_control_conv2d_16[5] }), .Y(_10184_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35198_ ( .A({ _d1_control_conv2d_16[0], _d1_control_conv2d_16[1] }), .Y(_10185_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35199_ ( .A({ _10186_, _10184_ }), .Y(_06001_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35200_ ( .A({ _d1_control_conv2d_16[2:1], _d1_control_conv2d_16[3], _d1_control_conv2d_16[0] }), .Y(_10186_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _35201_ ( .A({ _10184_, _d1_control_conv2d_16[3], _10180_, _d1_control_conv2d_16[2] }), .Y(_06002_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _35202_ ( .A({ _d1_control_conv2d_16[2], _10184_, _10185_, _d1_control_conv2d_16[3] }), .Y(_06003_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _35203_ ( .A({ _d1_control_conv2d_16[2], _d1_control_conv2d_16[3], _10185_, _10187_ }), .Y(_06004_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _35204_ ( .A({ _10182_, _10171_, _d1_control_conv2d_16[5] }), .Y(_10187_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35205_ ( .A({ _10186_, _10187_ }), .Y(_06005_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _35206_ ( .A({ _10187_, _d1_control_conv2d_16[3], _10180_, _d1_control_conv2d_16[2] }), .Y(_06006_) );
  \$lut  #( .LUT(16'hefff), .WIDTH(4) ) _35207_ ( .A({ _10185_, _10187_, _d1_control_conv2d_16[2], _d1_control_conv2d_16[3] }), .Y(_06007_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35208_ ( .A({ _07486_, _07918_ }), .Y(_06009_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35209_ ( .A({ _07464_, _07905_ }), .Y(_06010_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35210_ ( .A({ _06933_, _07905_ }), .Y(_06011_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35211_ ( .A({ _07466_, _07930_ }), .Y(_06018_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35212_ ( .A({ _07908_, _07930_ }), .Y(_06019_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35213_ ( .A({ _07461_, _07930_ }), .Y(_06020_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35214_ ( .A({ _08682_, _09039_ }), .Y(_06022_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35215_ ( .A({ _06900_, _09039_ }), .Y(_06023_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35216_ ( .A({ _06902_, _09039_ }), .Y(_06024_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35217_ ( .A({ _06904_, _06886_ }), .Y(_06025_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35218_ ( .A({ _08576_, _06886_ }), .Y(_06026_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _35219_ ( .A({ _10012_, _saxi_register_fsm[0] }), .Y(_05688_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35220_ ( .A({ conv2d_16_control_param_index[0], conv2d_16_control_param_index[1] }), .Y(_05689_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35221_ ( .A({ max_pool_serial_18_control_param_index[0], max_pool_serial_18_control_param_index[1] }), .Y(_05690_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35222_ ( .A({ matmul_29_control_param_index[0], matmul_29_control_param_index[1] }), .Y(_05691_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35223_ ( .A({ conv2d_16_prev_row_select[0], conv2d_16_prev_row_select[1] }), .Y(_05692_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35224_ ( .A({ __tmp_464_2[0], __tmp_464_2[1] }), .Y(_05693_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35225_ ( .A({ __tmp_475_2[0], __tmp_475_2[1] }), .Y(_05694_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35226_ ( .A({ __tmp_495_2[0], __tmp_495_2[1] }), .Y(_05695_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35227_ ( .A({ __tmp_505_2[0], __tmp_505_2[1] }), .Y(_05696_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35228_ ( .A({ __tmp_515_2[0], __tmp_515_2[1] }), .Y(_05697_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35229_ ( .A({ __tmp_525_2[0], __tmp_525_2[1] }), .Y(_05698_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35230_ ( .A({ __tmp_535_2[0], __tmp_535_2[1] }), .Y(_05699_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35231_ ( .A({ __tmp_545_2[0], __tmp_545_2[1] }), .Y(_05700_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35232_ ( .A({ __tmp_555_2[0], __tmp_555_2[1] }), .Y(_05701_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35233_ ( .A({ __tmp_565_2[0], __tmp_565_2[1] }), .Y(_05702_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35234_ ( .A({ __tmp_575_2[0], __tmp_575_2[1] }), .Y(_05703_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _35235_ ( .A({ __tmp_585_2[1:0], __tmp_585_2[2] }), .Y(_05704_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _35236_ ( .A({ __tmp_599_2[1:0], __tmp_599_2[2] }), .Y(_05705_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _35237_ ( .A({ __tmp_613_2[1:0], __tmp_613_2[2] }), .Y(_05706_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _35238_ ( .A({ __tmp_627_2[1:0], __tmp_627_2[2] }), .Y(_05707_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _35239_ ( .A({ __tmp_641_2[1:0], __tmp_641_2[2] }), .Y(_05708_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _35240_ ( .A({ __tmp_655_2[1:0], __tmp_655_2[2] }), .Y(_05709_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _35241_ ( .A({ __tmp_669_2[1:0], __tmp_669_2[2] }), .Y(_05710_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _35242_ ( .A({ __tmp_683_2[1:0], __tmp_683_2[2] }), .Y(_05711_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _35243_ ( .A({ __tmp_697_2[1:0], __tmp_697_2[2] }), .Y(_05712_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35244_ ( .A({ conv2d_16_row_select[0], conv2d_16_row_select[1] }), .Y(_05713_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35245_ ( .A({ __tmp_1027_2[0], __tmp_1027_2[1] }), .Y(_05714_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35246_ ( .A({ __tmp_1170_2[0], __tmp_1170_2[1] }), .Y(_05715_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35247_ ( .A({ __tmp_1181_2[0], __tmp_1181_2[1] }), .Y(_05716_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35248_ ( .A({ __tmp_1201_2[0], __tmp_1201_2[1] }), .Y(_05717_) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _35249_ ( .A({ __tmp_1211_2[1:0], __tmp_1211_2[2] }), .Y(_05718_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _35250_ ( .A({ _10023_, _tmp_5[1:0] }), .Y(_05719_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _35251_ ( .A({ _10194_, _10192_, _10188_ }), .Y(_05720_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35252_ ( .A({ _10191_, _10190_, _10189_ }), .Y(_10188_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _35253_ ( .A(_reduceadd_count_17[32:30]), .Y(_10189_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35254_ ( .A(_reduceadd_count_17[29:26]), .Y(_10190_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35255_ ( .A(_reduceadd_count_17[25:22]), .Y(_10191_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _35256_ ( .A({ _10193_, _reduceadd_count_17[1:0] }), .Y(_10192_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35257_ ( .A(_reduceadd_count_17[5:2]), .Y(_10193_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35258_ ( .A({ _10198_, _10197_, _10196_, _10195_ }), .Y(_10194_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35259_ ( .A(_reduceadd_count_17[13:10]), .Y(_10195_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35260_ ( .A(_reduceadd_count_17[9:6]), .Y(_10196_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35261_ ( .A(_reduceadd_count_17[21:18]), .Y(_10197_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35262_ ( .A(_reduceadd_count_17[17:14]), .Y(_10198_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _35263_ ( .A({ _10199_, _reducemax_count_211[4:3] }), .Y(_05721_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35264_ ( .A({ _10200_, _reducemax_count_211[8:6] }), .Y(_10199_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35265_ ( .A({ _reducemax_count_211[5], _reducemax_count_211[2:0] }), .Y(_10200_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35266_ ( .A({ _10206_, _10201_ }), .Y(_05722_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35267_ ( .A({ _10205_, _10204_, _10203_, _10202_ }), .Y(_10201_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35268_ ( .A(conv2d_16_out_ram_select[23:20]), .Y(_10202_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35269_ ( .A(conv2d_16_out_ram_select[19:16]), .Y(_10203_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35270_ ( .A(conv2d_16_out_ram_select[31:28]), .Y(_10204_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35271_ ( .A(conv2d_16_out_ram_select[27:24]), .Y(_10205_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35272_ ( .A({ _10210_, _10209_, _10208_, _10207_ }), .Y(_10206_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35273_ ( .A(conv2d_16_out_ram_select[7:4]), .Y(_10207_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35274_ ( .A(conv2d_16_out_ram_select[3:0]), .Y(_10208_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35275_ ( .A(conv2d_16_out_ram_select[15:12]), .Y(_10209_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35276_ ( .A(conv2d_16_out_ram_select[11:8]), .Y(_10210_) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35277_ ( .A({ conv2d_16_col_select[0], conv2d_16_col_select[1] }), .Y(_05723_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35278_ ( .A({ _10216_, _10211_ }), .Y(_05724_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35279_ ( .A({ _10215_, _10214_, _10213_, _10212_ }), .Y(_10211_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35280_ ( .A(matmul_29_out_ram_select[23:20]), .Y(_10212_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35281_ ( .A(matmul_29_out_ram_select[19:16]), .Y(_10213_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35282_ ( .A(matmul_29_out_ram_select[31:28]), .Y(_10214_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35283_ ( .A(matmul_29_out_ram_select[27:24]), .Y(_10215_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35284_ ( .A({ _10220_, _10219_, _10218_, _10217_ }), .Y(_10216_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35285_ ( .A(matmul_29_out_ram_select[7:4]), .Y(_10217_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35286_ ( .A(matmul_29_out_ram_select[3:0]), .Y(_10218_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35287_ ( .A(matmul_29_out_ram_select[15:12]), .Y(_10219_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35288_ ( .A(matmul_29_out_ram_select[11:8]), .Y(_10220_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35289_ ( .A({ _tmp_68[0], _tmp_68[1], _tmp_68[3:2] }), .Y(_06028_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35290_ ( .A({ _tmp_99[0], _tmp_99[1], _tmp_99[3:2] }), .Y(_06037_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35291_ ( .A({ _tmp_130[0], _tmp_130[1], _tmp_130[3:2] }), .Y(_06046_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35292_ ( .A({ _tmp_161[0], _tmp_161[1], _tmp_161[3:2] }), .Y(_06055_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35293_ ( .A({ _tmp_192[0], _tmp_192[1], _tmp_192[3:2] }), .Y(_06064_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35294_ ( .A({ _tmp_223[0], _tmp_223[1], _tmp_223[3:2] }), .Y(_06073_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35295_ ( .A({ _tmp_254[0], _tmp_254[1], _tmp_254[3:2] }), .Y(_06082_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35296_ ( .A({ _tmp_285[0], _tmp_285[1], _tmp_285[3:2] }), .Y(_06091_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35297_ ( .A({ _tmp_68[0], _tmp_68[1], _tmp_68[3:2] }), .Y(_06029_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35298_ ( .A({ _tmp_99[0], _tmp_99[1], _tmp_99[3:2] }), .Y(_06038_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35299_ ( .A({ _tmp_130[0], _tmp_130[1], _tmp_130[3:2] }), .Y(_06047_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35300_ ( .A({ _tmp_161[0], _tmp_161[1], _tmp_161[3:2] }), .Y(_06056_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35301_ ( .A({ _tmp_192[0], _tmp_192[1], _tmp_192[3:2] }), .Y(_06065_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35302_ ( .A({ _tmp_223[0], _tmp_223[1], _tmp_223[3:2] }), .Y(_06074_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35303_ ( .A({ _tmp_254[0], _tmp_254[1], _tmp_254[3:2] }), .Y(_06083_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35304_ ( .A({ _tmp_285[0], _tmp_285[1], _tmp_285[3:2] }), .Y(_06092_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35305_ ( .A({ _tmp_68[1:0], _tmp_68[3:2] }), .Y(_06030_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35306_ ( .A({ _tmp_99[1:0], _tmp_99[3:2] }), .Y(_06039_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35307_ ( .A({ _tmp_130[1:0], _tmp_130[3:2] }), .Y(_06048_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35308_ ( .A({ _tmp_161[1:0], _tmp_161[3:2] }), .Y(_06057_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35309_ ( .A({ _tmp_192[1:0], _tmp_192[3:2] }), .Y(_06066_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35310_ ( .A({ _tmp_223[1:0], _tmp_223[3:2] }), .Y(_06075_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35311_ ( .A({ _tmp_254[1:0], _tmp_254[3:2] }), .Y(_06084_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35312_ ( .A({ _tmp_285[1:0], _tmp_285[3:2] }), .Y(_06093_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35313_ ( .A({ _tmp_68[0], _tmp_68[1], _tmp_68[3:2] }), .Y(_06031_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35314_ ( .A({ _tmp_99[0], _tmp_99[1], _tmp_99[3:2] }), .Y(_06040_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35315_ ( .A({ _tmp_130[0], _tmp_130[1], _tmp_130[3:2] }), .Y(_06049_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35316_ ( .A({ _tmp_161[0], _tmp_161[1], _tmp_161[3:2] }), .Y(_06058_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35317_ ( .A({ _tmp_192[0], _tmp_192[1], _tmp_192[3:2] }), .Y(_06067_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35318_ ( .A({ _tmp_223[0], _tmp_223[1], _tmp_223[3:2] }), .Y(_06076_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35319_ ( .A({ _tmp_254[0], _tmp_254[1], _tmp_254[3:2] }), .Y(_06085_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35320_ ( .A({ _tmp_285[0], _tmp_285[1], _tmp_285[3:2] }), .Y(_06094_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35321_ ( .A({ _tmp_68[2], _tmp_68[0], _tmp_68[1], _tmp_68[3] }), .Y(_06032_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35322_ ( .A({ _tmp_99[2], _tmp_99[0], _tmp_99[1], _tmp_99[3] }), .Y(_06041_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35323_ ( .A({ _tmp_130[2], _tmp_130[0], _tmp_130[1], _tmp_130[3] }), .Y(_06050_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35324_ ( .A({ _tmp_161[2], _tmp_161[0], _tmp_161[1], _tmp_161[3] }), .Y(_06059_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35325_ ( .A({ _tmp_192[2], _tmp_192[0], _tmp_192[1], _tmp_192[3] }), .Y(_06068_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35326_ ( .A({ _tmp_223[2], _tmp_223[0], _tmp_223[1], _tmp_223[3] }), .Y(_06077_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35327_ ( .A({ _tmp_254[2], _tmp_254[0], _tmp_254[1], _tmp_254[3] }), .Y(_06086_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35328_ ( .A({ _tmp_285[2], _tmp_285[0], _tmp_285[1], _tmp_285[3] }), .Y(_06095_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35329_ ( .A({ _tmp_68[0], _tmp_68[2:1], _tmp_68[3] }), .Y(_06033_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35330_ ( .A({ _tmp_99[0], _tmp_99[2:1], _tmp_99[3] }), .Y(_06042_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35331_ ( .A({ _tmp_130[0], _tmp_130[2:1], _tmp_130[3] }), .Y(_06051_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35332_ ( .A({ _tmp_161[0], _tmp_161[2:1], _tmp_161[3] }), .Y(_06060_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35333_ ( .A({ _tmp_192[0], _tmp_192[2:1], _tmp_192[3] }), .Y(_06069_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35334_ ( .A({ _tmp_223[0], _tmp_223[2:1], _tmp_223[3] }), .Y(_06078_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35335_ ( .A({ _tmp_254[0], _tmp_254[2:1], _tmp_254[3] }), .Y(_06087_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35336_ ( .A({ _tmp_285[0], _tmp_285[2:1], _tmp_285[3] }), .Y(_06096_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35337_ ( .A({ _tmp_68[2:0], _tmp_68[3] }), .Y(_06034_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35338_ ( .A({ _tmp_99[2:0], _tmp_99[3] }), .Y(_06043_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35339_ ( .A({ _tmp_130[2:0], _tmp_130[3] }), .Y(_06052_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35340_ ( .A({ _tmp_161[2:0], _tmp_161[3] }), .Y(_06061_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35341_ ( .A({ _tmp_192[2:0], _tmp_192[3] }), .Y(_06070_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35342_ ( .A({ _tmp_223[2:0], _tmp_223[3] }), .Y(_06079_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35343_ ( .A({ _tmp_254[2:0], _tmp_254[3] }), .Y(_06088_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35344_ ( .A({ _tmp_285[2:0], _tmp_285[3] }), .Y(_06097_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35345_ ( .A({ _tmp_68[0], _tmp_68[1], _tmp_68[2], _tmp_68[3] }), .Y(_06035_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35346_ ( .A({ _tmp_99[0], _tmp_99[1], _tmp_99[2], _tmp_99[3] }), .Y(_06044_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35347_ ( .A({ _tmp_130[0], _tmp_130[1], _tmp_130[2], _tmp_130[3] }), .Y(_06053_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35348_ ( .A({ _tmp_161[0], _tmp_161[1], _tmp_161[2], _tmp_161[3] }), .Y(_06062_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35349_ ( .A({ _tmp_192[0], _tmp_192[1], _tmp_192[2], _tmp_192[3] }), .Y(_06071_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35350_ ( .A({ _tmp_223[0], _tmp_223[1], _tmp_223[2], _tmp_223[3] }), .Y(_06080_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35351_ ( .A({ _tmp_254[0], _tmp_254[1], _tmp_254[2], _tmp_254[3] }), .Y(_06089_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35352_ ( .A({ _tmp_285[0], _tmp_285[1], _tmp_285[2], _tmp_285[3] }), .Y(_06098_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35353_ ( .A({ _tmp_68[3], _tmp_68[0], _tmp_68[1], _tmp_68[2] }), .Y(_06027_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35354_ ( .A({ _tmp_99[3], _tmp_99[0], _tmp_99[1], _tmp_99[2] }), .Y(_06036_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35355_ ( .A({ _tmp_130[3], _tmp_130[0], _tmp_130[1], _tmp_130[2] }), .Y(_06045_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35356_ ( .A({ _tmp_161[3], _tmp_161[0], _tmp_161[1], _tmp_161[2] }), .Y(_06054_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35357_ ( .A({ _tmp_192[3], _tmp_192[0], _tmp_192[1], _tmp_192[2] }), .Y(_06063_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35358_ ( .A({ _tmp_223[3], _tmp_223[0], _tmp_223[1], _tmp_223[2] }), .Y(_06072_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35359_ ( .A({ _tmp_254[3], _tmp_254[0], _tmp_254[1], _tmp_254[2] }), .Y(_06081_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35360_ ( .A({ _tmp_285[3], _tmp_285[0], _tmp_285[1], _tmp_285[2] }), .Y(_06090_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35361_ ( .A({ _tmp_303[0], _tmp_303[1] }), .Y(_06101_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35362_ ( .A({ _tmp_316[0], _tmp_316[1] }), .Y(_06104_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35363_ ( .A({ _tmp_329[0], _tmp_329[1] }), .Y(_06107_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35364_ ( .A({ _tmp_342[0], _tmp_342[1] }), .Y(_06110_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35365_ ( .A({ _tmp_303[0], _tmp_303[1] }), .Y(_06102_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35366_ ( .A({ _tmp_316[0], _tmp_316[1] }), .Y(_06105_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35367_ ( .A({ _tmp_329[0], _tmp_329[1] }), .Y(_06108_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35368_ ( .A({ _tmp_342[0], _tmp_342[1] }), .Y(_06111_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35369_ ( .A(_tmp_303), .Y(_06100_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35370_ ( .A(_tmp_316), .Y(_06103_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35371_ ( .A(_tmp_329), .Y(_06106_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35372_ ( .A(_tmp_342), .Y(_06109_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35373_ ( .A({ _tmp_360[0], _tmp_360[1] }), .Y(_06113_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35374_ ( .A({ _tmp_373[0], _tmp_373[1] }), .Y(_06116_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35375_ ( .A({ _tmp_386[0], _tmp_386[1] }), .Y(_06119_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35376_ ( .A({ _tmp_399[0], _tmp_399[1] }), .Y(_06122_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35377_ ( .A({ _tmp_360[0], _tmp_360[1] }), .Y(_06114_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35378_ ( .A({ _tmp_373[0], _tmp_373[1] }), .Y(_06117_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35379_ ( .A({ _tmp_386[0], _tmp_386[1] }), .Y(_06120_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35380_ ( .A({ _tmp_399[0], _tmp_399[1] }), .Y(_06123_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35381_ ( .A(_tmp_360), .Y(_06112_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35382_ ( .A(_tmp_373), .Y(_06115_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35383_ ( .A(_tmp_386), .Y(_06118_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35384_ ( .A(_tmp_399), .Y(_06121_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35385_ ( .A({ _tmp_417[0], _tmp_417[1] }), .Y(_06125_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35386_ ( .A({ _tmp_430[0], _tmp_430[1] }), .Y(_06128_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35387_ ( .A({ _tmp_443[0], _tmp_443[1] }), .Y(_06131_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35388_ ( .A({ _tmp_456[0], _tmp_456[1] }), .Y(_06134_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35389_ ( .A({ _tmp_417[0], _tmp_417[1] }), .Y(_06126_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35390_ ( .A({ _tmp_430[0], _tmp_430[1] }), .Y(_06129_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35391_ ( .A({ _tmp_443[0], _tmp_443[1] }), .Y(_06132_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35392_ ( .A({ _tmp_456[0], _tmp_456[1] }), .Y(_06135_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35393_ ( .A(_tmp_417), .Y(_06124_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35394_ ( .A(_tmp_430), .Y(_06127_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35395_ ( .A(_tmp_443), .Y(_06130_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35396_ ( .A(_tmp_456), .Y(_06133_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35397_ ( .A({ _10230_, _10228_, _10221_ }), .Y(_06099_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35398_ ( .A({ _10227_, _10222_, _maxi_write_size[2:1] }), .Y(_10221_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35399_ ( .A({ _10226_, _10225_, _10224_, _10223_ }), .Y(_10222_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35400_ ( .A(_maxi_write_size[14:11]), .Y(_10223_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35401_ ( .A(_maxi_write_size[10:7]), .Y(_10224_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35402_ ( .A(_maxi_write_size[22:19]), .Y(_10225_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35403_ ( .A(_maxi_write_size[18:15]), .Y(_10226_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35404_ ( .A(_maxi_write_size[6:3]), .Y(_10227_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35405_ ( .A({ _maxi_write_size[0], _10229_, _maxi_write_size[32:31] }), .Y(_10228_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35406_ ( .A({ _maxi_write_size[29:28], _maxi_write_size[26], _maxi_write_size[23] }), .Y(_10229_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35407_ ( .A({ _maxi_write_size[30], _maxi_write_size[27], _maxi_write_size[25:24] }), .Y(_10230_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35408_ ( .A(__variable_wdata_215), .Y(_06136_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35409_ ( .A({ __variable_wdata_215[0], __variable_wdata_215[1] }), .Y(_06137_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35410_ ( .A(__variable_wdata_215), .Y(_06138_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35411_ ( .A(__variable_wdata_216), .Y(_06139_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35412_ ( .A({ __variable_wdata_216[0], __variable_wdata_216[1] }), .Y(_06140_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35413_ ( .A(__variable_wdata_216), .Y(_06141_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35414_ ( .A({ __variable_wdata_849[0], __variable_wdata_849[1] }), .Y(_06144_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35415_ ( .A({ __variable_wdata_849[0], __variable_wdata_849[1] }), .Y(_06145_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35416_ ( .A({ _tmp_3, saxi_bvalid, _06878_, _05688_ }), .Y(saxi_awready) );
  \$lut  #( .LUT(4'he), .WIDTH(2) ) _35417_ ( .A({ _tmp_1, _tmp_2 }), .Y(_06878_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _35418_ ( .A({ _tmp_4, _06878_, _05688_ }), .Y(saxi_arready) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _35419_ ( .A({ conv2d_16_row_count[5], _10232_, _10237_, _05317_ }), .Y(_10231_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35420_ ( .A({ _10236_, _10235_, _10234_, _10233_ }), .Y(_10232_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35421_ ( .A({ conv2d_16_row_count[2], _05312_ }), .Y(_10233_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _35422_ ( .A({ _05290_, conv2d_16_row_count[0], conv2d_16_row_count[1], _05301_ }), .Y(_10234_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35423_ ( .A({ _05312_, conv2d_16_row_count[2], _05315_, conv2d_16_row_count[3] }), .Y(_10235_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35424_ ( .A({ conv2d_16_row_count[3], _05315_, conv2d_16_row_count[4], _05316_ }), .Y(_10236_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35425_ ( .A({ _05316_, conv2d_16_row_count[4] }), .Y(_10237_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35426_ ( .A({ _05292_, conv2d_16_row_count[11:10], _05291_ }), .Y(_10238_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35427_ ( .A({ _05318_, conv2d_16_row_count[6] }), .Y(_10239_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35428_ ( .A({ conv2d_16_row_count[7], _05319_, conv2d_16_row_count[6], _05318_ }), .Y(_10240_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35429_ ( .A({ _10243_, _10238_, _10242_ }), .Y(_10241_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35430_ ( .A({ conv2d_16_row_count[8], _05320_, _05321_, conv2d_16_row_count[9] }), .Y(_10242_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35431_ ( .A({ conv2d_16_row_count[10], conv2d_16_row_count[11], _05291_, _05292_ }), .Y(_10243_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35432_ ( .A({ _05296_, conv2d_16_row_count[15:14], _05295_ }), .Y(_10244_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _35433_ ( .A({ _10246_, _10253_, _10248_, _10254_ }), .Y(_10245_) );
  \$lut  #( .LUT(16'h0bff), .WIDTH(4) ) _35434_ ( .A({ _10247_, _10252_, _10250_, _10251_ }), .Y(_10246_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35435_ ( .A({ _10249_, _10248_ }), .Y(_10247_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35436_ ( .A({ _05305_, conv2d_16_row_count[23:22], _05304_ }), .Y(_10248_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35437_ ( .A({ conv2d_16_row_count[20], _05302_, _05303_, conv2d_16_row_count[21] }), .Y(_10249_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35438_ ( .A({ _05300_, conv2d_16_row_count[19:18], _05299_ }), .Y(_10250_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35439_ ( .A({ conv2d_16_row_count[16], _05297_, _05298_, conv2d_16_row_count[17] }), .Y(_10251_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35440_ ( .A({ conv2d_16_row_count[18], conv2d_16_row_count[19], _05299_, _05300_ }), .Y(_10252_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35441_ ( .A({ conv2d_16_row_count[22], conv2d_16_row_count[23], _05304_, _05305_ }), .Y(_10253_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _35442_ ( .A({ conv2d_16_row_count[20], _05302_, _05303_, conv2d_16_row_count[21] }), .Y(_10254_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35443_ ( .A({ _10256_, _10250_, _10247_ }), .Y(_10255_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35444_ ( .A({ conv2d_16_row_count[17], _05298_, conv2d_16_row_count[16], _05297_ }), .Y(_10256_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35445_ ( .A({ _10259_, _10244_, _10258_ }), .Y(_10257_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35446_ ( .A({ conv2d_16_row_count[12], _05293_, _05294_, conv2d_16_row_count[13] }), .Y(_10258_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35447_ ( .A({ conv2d_16_row_count[14], conv2d_16_row_count[15], _05295_, _05296_ }), .Y(_10259_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35448_ ( .A({ _10264_, _10261_ }), .Y(_10260_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35449_ ( .A({ _10263_, _10262_ }), .Y(_10261_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35450_ ( .A({ conv2d_16_row_count[30], _05313_, conv2d_16_row_count[31], _05314_ }), .Y(_10262_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35451_ ( .A({ conv2d_16_row_count[29], _05311_, conv2d_16_row_count[28], _05310_ }), .Y(_10263_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35452_ ( .A({ _05309_, conv2d_16_row_count[27], _05308_, conv2d_16_row_count[26] }), .Y(_10264_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _35453_ ( .A({ conv2d_16_row_count[28], _05310_, _05311_, conv2d_16_row_count[29] }), .Y(_10265_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35454_ ( .A({ conv2d_16_row_count[26], _05308_, _05309_, conv2d_16_row_count[27] }), .Y(_10266_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35455_ ( .A({ conv2d_16_row_count[30], conv2d_16_row_count[31], _05313_, _05314_ }), .Y(_10267_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35456_ ( .A({ conv2d_16_row_count[24], conv2d_16_row_count[25], _05306_, _05307_ }), .Y(_10268_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35457_ ( .A({ conv2d_16_row_count[4], conv2d_16_row_count[2], conv2d_16_row_count[3], conv2d_16_row_count[1] }), .Y(_10269_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35458_ ( .A({ _05306_, conv2d_16_row_count[24], conv2d_16_row_count[25], _05307_ }), .Y(_10270_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35459_ ( .A({ _05315_, _05347_ }), .Y(_10271_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35460_ ( .A({ _05290_, _05322_, _05333_, _05301_ }), .Y(_10272_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35461_ ( .A({ _05347_, _05315_, _05348_, _05316_ }), .Y(_10273_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35462_ ( .A({ _05349_, _05317_ }), .Y(_10274_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35463_ ( .A({ _05316_, _05348_, _05317_, _05349_ }), .Y(_10275_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35464_ ( .A({ _10278_, _10277_, _05319_, _05351_ }), .Y(_10276_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35465_ ( .A({ _05324_, _05292_, _05323_, _05291_ }), .Y(_10277_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35466_ ( .A({ _05353_, _05321_, _05352_, _05320_ }), .Y(_10278_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35467_ ( .A({ _05318_, _05350_ }), .Y(_10279_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35468_ ( .A({ _05351_, _05319_, _05350_, _05318_ }), .Y(_10280_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _35469_ ( .A({ _10282_, _10277_, _10283_ }), .Y(_10281_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35470_ ( .A({ _05323_, _05324_, _05291_, _05292_ }), .Y(_10282_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35471_ ( .A({ _05352_, _05353_, _05320_, _05321_ }), .Y(_10283_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35472_ ( .A({ _05328_, _05296_, _05327_, _05295_ }), .Y(_10284_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35473_ ( .A({ _05326_, _05294_, _05325_, _05293_ }), .Y(_10285_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35474_ ( .A({ _05327_, _05328_, _05295_, _05296_ }), .Y(_10286_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35475_ ( .A({ _05325_, _05326_, _05293_, _05294_ }), .Y(_10287_) );
  \$lut  #( .LUT(16'h000b), .WIDTH(4) ) _35476_ ( .A({ _10297_, _10289_, _10291_, _10293_ }), .Y(_10288_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _35477_ ( .A({ _10290_, _10295_, _10296_, _10294_ }), .Y(_10289_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35478_ ( .A({ _10293_, _10291_, _05302_, _05334_ }), .Y(_10290_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35479_ ( .A({ _10292_, _05303_, _05335_ }), .Y(_10291_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35480_ ( .A({ _05337_, _05305_, _05336_, _05304_ }), .Y(_10292_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35481_ ( .A({ _05334_, _05302_, _05335_, _05303_ }), .Y(_10293_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35482_ ( .A({ _05332_, _05300_, _05331_, _05299_ }), .Y(_10294_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35483_ ( .A({ _05331_, _05332_, _05299_, _05300_ }), .Y(_10295_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35484_ ( .A({ _05329_, _05330_, _05297_, _05298_ }), .Y(_10296_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35485_ ( .A({ _05336_, _05337_, _05304_, _05305_ }), .Y(_10297_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35486_ ( .A({ _10299_, _05306_, _05338_ }), .Y(_10298_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35487_ ( .A({ _10304_, _10300_, _05307_, _05339_ }), .Y(_10299_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35488_ ( .A({ _10303_, _10301_, _05310_, _05342_ }), .Y(_10300_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35489_ ( .A({ _10302_, _05346_, _05314_ }), .Y(_10301_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35490_ ( .A({ _05313_, _05345_, _05311_, _05343_ }), .Y(_10302_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35491_ ( .A({ _05342_, _05310_, _05343_, _05311_ }), .Y(_10303_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35492_ ( .A({ _05341_, _05309_, _05340_, _05308_ }), .Y(_10304_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35493_ ( .A({ _10306_, _10294_, _10290_ }), .Y(_10305_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35494_ ( .A({ _05330_, _05298_, _05329_, _05297_ }), .Y(_10306_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35495_ ( .A({ _05340_, _05341_, _05308_, _05309_ }), .Y(_10307_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35496_ ( .A({ _05345_, _05346_, _05313_, _05314_ }), .Y(_10308_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35497_ ( .A({ _10313_, _10312_, _10311_, _10310_ }), .Y(_10309_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35498_ ( .A({ _05337_, _05336_, _05335_, _05334_ }), .Y(_10310_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35499_ ( .A({ _05332_, _05331_, _05330_, _05329_ }), .Y(_10311_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35500_ ( .A({ _05346_, _05345_, _05343_, _05342_ }), .Y(_10312_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35501_ ( .A({ _05341_, _05340_, _05339_, _05338_ }), .Y(_10313_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35502_ ( .A({ _10318_, _10317_, _10316_, _10315_ }), .Y(_10314_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35503_ ( .A({ _05351_, _05350_, _05349_, _05348_ }), .Y(_10315_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35504_ ( .A({ _05347_, _05344_, _05333_, _05322_ }), .Y(_10316_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35505_ ( .A({ _05324_, _05323_, _05353_, _05352_ }), .Y(_10317_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35506_ ( .A({ _05328_, _05327_, _05326_, _05325_ }), .Y(_10318_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _35507_ ( .A({ _10329_, _10320_, _10332_ }), .Y(_10319_) );
  \$lut  #( .LUT(16'h00f4), .WIDTH(4) ) _35508_ ( .A({ _10326_, _10327_, _10328_, _10321_ }), .Y(_10320_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _35509_ ( .A({ _10325_, _10324_, _10322_, _10323_ }), .Y(_10321_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35510_ ( .A({ _05376_, _05312_ }), .Y(_10322_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35511_ ( .A({ _05290_, _05354_, _05365_, _05301_ }), .Y(_10323_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35512_ ( .A({ _05312_, _05376_, _05315_, _05379_ }), .Y(_10324_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35513_ ( .A({ _05379_, _05315_, _05380_, _05316_ }), .Y(_10325_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35514_ ( .A({ _05318_, _05382_ }), .Y(_10326_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35515_ ( .A({ _05381_, _05317_ }), .Y(_10327_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35516_ ( .A({ _05316_, _05380_, _05317_, _05381_ }), .Y(_10328_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35517_ ( .A({ _10331_, _10330_, _05319_, _05383_ }), .Y(_10329_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35518_ ( .A({ _05356_, _05292_, _05355_, _05291_ }), .Y(_10330_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35519_ ( .A({ _05385_, _05321_, _05384_, _05320_ }), .Y(_10331_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35520_ ( .A({ _05383_, _05319_, _05382_, _05318_ }), .Y(_10332_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35521_ ( .A({ _10336_, _10334_ }), .Y(_10333_) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _35522_ ( .A({ _10330_, _05385_, _05321_, _10335_ }), .Y(_10334_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35523_ ( .A({ _05384_, _05320_ }), .Y(_10335_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35524_ ( .A({ _05355_, _05356_, _05291_, _05292_ }), .Y(_10336_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35525_ ( .A({ _05360_, _05296_, _05359_, _05295_ }), .Y(_10337_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35526_ ( .A({ _05294_, _05358_, _05357_, _05293_ }), .Y(_10338_) );
  \$lut  #( .LUT(16'h9000), .WIDTH(4) ) _35527_ ( .A({ _10344_, _10340_, _05298_, _05362_ }), .Y(_10339_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35528_ ( .A({ _10341_, _05361_, _05297_ }), .Y(_10340_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35529_ ( .A({ _10343_, _10342_ }), .Y(_10341_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35530_ ( .A({ _05369_, _05305_, _05368_, _05304_ }), .Y(_10342_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35531_ ( .A({ _05303_, _05367_, _05366_, _05302_ }), .Y(_10343_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35532_ ( .A({ _05364_, _05300_, _05363_, _05299_ }), .Y(_10344_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _35533_ ( .A({ _05357_, _05293_, _05294_, _05358_ }), .Y(_10345_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35534_ ( .A({ _05359_, _05360_, _05295_, _05296_ }), .Y(_10346_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35535_ ( .A({ _10348_, _10364_, _10365_ }), .Y(_10347_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _35536_ ( .A({ _10363_, _10349_, _10360_, _10362_ }), .Y(_10348_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35537_ ( .A({ _10359_, _10358_, _10355_, _10350_ }), .Y(_10349_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35538_ ( .A({ _10354_, _10353_, _10352_, _10351_ }), .Y(_10350_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35539_ ( .A({ _05378_, _05377_, _05375_, _05374_ }), .Y(_10351_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35540_ ( .A({ _05373_, _05372_, _05371_, _05370_ }), .Y(_10352_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35541_ ( .A({ _05369_, _05368_, _05367_, _05366_ }), .Y(_10353_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35542_ ( .A({ _05364_, _05363_, _05362_, _05361_ }), .Y(_10354_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35543_ ( .A({ _10357_, _10356_ }), .Y(_10355_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35544_ ( .A({ _05360_, _05359_, _05358_, _05357_ }), .Y(_10356_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35545_ ( .A({ _05356_, _05355_, _05385_, _05384_ }), .Y(_10357_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35546_ ( .A({ _05383_, _05382_, _05381_, _05380_ }), .Y(_10358_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35547_ ( .A({ _05379_, _05376_, _05365_, _05354_ }), .Y(_10359_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35548_ ( .A({ _10361_, _05378_, _05314_ }), .Y(_10360_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35549_ ( .A({ _05313_, _05377_, _05311_, _05375_ }), .Y(_10361_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35550_ ( .A({ _05374_, _05310_, _05375_, _05311_ }), .Y(_10362_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35551_ ( .A({ _05377_, _05378_, _05313_, _05314_ }), .Y(_10363_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35552_ ( .A({ _10362_, _10360_, _05310_, _05374_ }), .Y(_10364_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _35553_ ( .A({ _10368_, _10366_, _10367_ }), .Y(_10365_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35554_ ( .A({ _05309_, _05373_, _05308_, _05372_ }), .Y(_10366_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35555_ ( .A({ _05370_, _05371_, _05306_, _05307_ }), .Y(_10367_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35556_ ( .A({ _05372_, _05308_, _05309_, _05373_ }), .Y(_10368_) );
  \$lut  #( .LUT(16'hf4ff), .WIDTH(4) ) _35557_ ( .A({ _10373_, _10370_, _10342_, _10374_ }), .Y(_10369_) );
  \$lut  #( .LUT(16'hf400), .WIDTH(4) ) _35558_ ( .A({ _10341_, _10372_, _10344_, _10371_ }), .Y(_10370_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35559_ ( .A({ _05361_, _05297_, _05298_, _05362_ }), .Y(_10371_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35560_ ( .A({ _05363_, _05364_, _05299_, _05300_ }), .Y(_10372_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35561_ ( .A({ _05368_, _05369_, _05304_, _05305_ }), .Y(_10373_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35562_ ( .A({ _05366_, _05302_, _05303_, _05367_ }), .Y(_10374_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35563_ ( .A({ _10376_, _10366_, _10364_ }), .Y(_10375_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35564_ ( .A({ _05306_, _05370_, _05371_, _05307_ }), .Y(_10376_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35565_ ( .A({ _10428_, _10377_ }), .Y(conv2d_16_stream_pad_mask_0_0) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35566_ ( .A({ _10426_, _10424_, _10416_, _13120_ }), .Y(_10377_) );
  \$lut  #( .LUT(16'h00f4), .WIDTH(4) ) _35567_ ( .A({ _10384_, _10385_, _10386_, _10379_ }), .Y(_10378_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _35568_ ( .A({ _10380_, _10383_, _10382_, _10381_ }), .Y(_10379_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35569_ ( .A({ conv2d_16_col_count[3], _05315_, conv2d_16_col_count[4], _05316_ }), .Y(_10380_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35570_ ( .A({ conv2d_16_col_count[2], _05312_ }), .Y(_10381_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35571_ ( .A({ _05290_, conv2d_16_col_count[0], conv2d_16_col_count[1], _05301_ }), .Y(_10382_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35572_ ( .A({ _05312_, conv2d_16_col_count[2], _05315_, conv2d_16_col_count[3] }), .Y(_10383_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35573_ ( .A({ _05318_, conv2d_16_col_count[6] }), .Y(_10384_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35574_ ( .A({ conv2d_16_col_count[5], _05317_ }), .Y(_10385_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35575_ ( .A({ _05316_, conv2d_16_col_count[4], _05317_, conv2d_16_col_count[5] }), .Y(_10386_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35576_ ( .A({ conv2d_16_col_count[11], _05292_, conv2d_16_col_count[10], _05291_ }), .Y(_10387_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _35577_ ( .A({ _10389_, _10390_, _10387_ }), .Y(_10388_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35578_ ( .A({ conv2d_16_col_count[10], conv2d_16_col_count[11], _05291_, _05292_ }), .Y(_10389_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35579_ ( .A({ conv2d_16_col_count[8], _05320_, _05321_, conv2d_16_col_count[9] }), .Y(_10390_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35580_ ( .A({ conv2d_16_col_count[7], _05319_, conv2d_16_col_count[6], _05318_ }), .Y(_10391_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35581_ ( .A({ _10407_, _10402_, _10397_, _10393_ }), .Y(_10392_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35582_ ( .A({ _10396_, _10394_, _05310_, conv2d_16_col_count[28] }), .Y(_10393_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _35583_ ( .A({ _10395_, conv2d_16_col_count[29], _05311_ }), .Y(_10394_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35584_ ( .A({ _05313_, conv2d_16_col_count[30], conv2d_16_col_count[31], _05314_ }), .Y(_10395_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35585_ ( .A({ conv2d_16_col_count[28], _05310_, conv2d_16_col_count[29], _05311_ }), .Y(_10396_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _35586_ ( .A({ _10398_, _10400_, _10401_ }), .Y(_10397_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35587_ ( .A({ _10399_, _05309_, conv2d_16_col_count[27] }), .Y(_10398_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35588_ ( .A({ _05308_, conv2d_16_col_count[26], _05307_, conv2d_16_col_count[25] }), .Y(_10399_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35589_ ( .A({ conv2d_16_col_count[25], _05307_, conv2d_16_col_count[24], _05306_ }), .Y(_10400_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35590_ ( .A({ _05306_, conv2d_16_col_count[24] }), .Y(_10401_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _35591_ ( .A({ _10403_, _10405_, _10406_ }), .Y(_10402_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35592_ ( .A({ _10404_, conv2d_16_col_count[23], _05305_ }), .Y(_10403_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35593_ ( .A({ conv2d_16_col_count[22], _05304_, _05303_, conv2d_16_col_count[21] }), .Y(_10404_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35594_ ( .A({ conv2d_16_col_count[20], _05302_, conv2d_16_col_count[21], _05303_ }), .Y(_10405_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35595_ ( .A({ _05302_, conv2d_16_col_count[20] }), .Y(_10406_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35596_ ( .A({ _10409_, _10408_ }), .Y(_10407_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35597_ ( .A({ conv2d_16_col_count[19], _05300_, conv2d_16_col_count[18], _05299_ }), .Y(_10408_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35598_ ( .A({ _05298_, conv2d_16_col_count[17:16], _05297_ }), .Y(_10409_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35599_ ( .A({ _10412_, _10411_ }), .Y(_10410_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35600_ ( .A({ conv2d_16_col_count[15], _05296_, conv2d_16_col_count[14], _05295_ }), .Y(_10411_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35601_ ( .A({ conv2d_16_col_count[12], _05293_, _05294_, conv2d_16_col_count[13] }), .Y(_10412_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35602_ ( .A({ _10415_, _10411_, _10414_ }), .Y(_10413_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35603_ ( .A({ conv2d_16_col_count[12], _05293_, _05294_, conv2d_16_col_count[13] }), .Y(_10414_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35604_ ( .A({ conv2d_16_col_count[14], conv2d_16_col_count[15], _05295_, _05296_ }), .Y(_10415_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _35605_ ( .A({ _10393_, _10417_, _10423_ }), .Y(_10416_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _35606_ ( .A({ _10398_, _10400_, _10401_, _10418_ }), .Y(_10417_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35607_ ( .A({ _10422_, _10403_, _10405_, _10419_ }), .Y(_10418_) );
  \$lut  #( .LUT(16'h004f), .WIDTH(4) ) _35608_ ( .A({ _10406_, _10421_, _10408_, _10420_ }), .Y(_10419_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35609_ ( .A({ conv2d_16_col_count[16], _05297_, _05298_, conv2d_16_col_count[17] }), .Y(_10420_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35610_ ( .A({ conv2d_16_col_count[18], conv2d_16_col_count[19], _05299_, _05300_ }), .Y(_10421_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35611_ ( .A({ conv2d_16_col_count[22], conv2d_16_col_count[23], _05304_, _05305_ }), .Y(_10422_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35612_ ( .A({ conv2d_16_col_count[26], _05308_, _05309_, conv2d_16_col_count[27] }), .Y(_10423_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _35613_ ( .A({ _10425_, conv2d_16_col_count[4], conv2d_16_col_count[2] }), .Y(_10424_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35614_ ( .A({ _09491_, conv2d_16_col_count[3], conv2d_16_col_count[1:0] }), .Y(_10425_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35615_ ( .A({ _10427_, _10394_, _10396_ }), .Y(_10426_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35616_ ( .A({ conv2d_16_col_count[30], conv2d_16_col_count[31], _05313_, _05314_ }), .Y(_10427_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35617_ ( .A({ _10456_, _10484_, _10478_, _10429_ }), .Y(_10428_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35618_ ( .A({ _10444_, _10453_, _10450_, _13123_ }), .Y(_10429_) );
  \$lut  #( .LUT(16'h00f4), .WIDTH(4) ) _35619_ ( .A({ _10436_, _10437_, _10438_, _10431_ }), .Y(_10430_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _35620_ ( .A({ _10435_, _10434_, _10432_, _10433_ }), .Y(_10431_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35621_ ( .A({ _05290_, conv2d_16_row_count_buf[0], conv2d_16_row_count_buf[1], _05301_ }), .Y(_10432_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35622_ ( .A({ conv2d_16_row_count_buf[2], _05312_, _05315_, conv2d_16_row_count_buf[3] }), .Y(_10433_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _35623_ ( .A({ conv2d_16_row_count_buf[2], _05312_, _05315_, conv2d_16_row_count_buf[3] }), .Y(_10434_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35624_ ( .A({ conv2d_16_row_count_buf[3], _05315_, conv2d_16_row_count_buf[4], _05316_ }), .Y(_10435_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35625_ ( .A({ _05318_, conv2d_16_row_count_buf[6] }), .Y(_10436_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35626_ ( .A({ conv2d_16_row_count_buf[5], _05317_ }), .Y(_10437_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35627_ ( .A({ _05316_, conv2d_16_row_count_buf[4], _05317_, conv2d_16_row_count_buf[5] }), .Y(_10438_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35628_ ( .A({ conv2d_16_row_count_buf[11], _05292_, conv2d_16_row_count_buf[10], _05291_ }), .Y(_10439_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35629_ ( .A({ conv2d_16_row_count_buf[10], conv2d_16_row_count_buf[11], _05291_, _05292_ }), .Y(_10440_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35630_ ( .A({ _10442_, _10439_, _05319_, conv2d_16_row_count_buf[7] }), .Y(_10441_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35631_ ( .A({ conv2d_16_row_count_buf[9], _05321_, conv2d_16_row_count_buf[8], _05320_ }), .Y(_10442_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35632_ ( .A({ conv2d_16_row_count_buf[7], _05319_, conv2d_16_row_count_buf[6], _05318_ }), .Y(_10443_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35633_ ( .A({ _10449_, _10448_, _10445_ }), .Y(_10444_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35634_ ( .A({ _10447_, _10446_ }), .Y(_10445_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35635_ ( .A({ conv2d_16_row_count_buf[23], _05305_, conv2d_16_row_count_buf[22], _05304_ }), .Y(_10446_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35636_ ( .A({ _05303_, conv2d_16_row_count_buf[21:20], _05302_ }), .Y(_10447_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35637_ ( .A({ conv2d_16_row_count_buf[19], _05300_, conv2d_16_row_count_buf[18], _05299_ }), .Y(_10448_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35638_ ( .A({ _05298_, conv2d_16_row_count_buf[17:16], _05297_ }), .Y(_10449_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35639_ ( .A({ _10452_, _10451_ }), .Y(_10450_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35640_ ( .A({ conv2d_16_row_count_buf[15], _05296_, conv2d_16_row_count_buf[14], _05295_ }), .Y(_10451_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35641_ ( .A({ _05294_, conv2d_16_row_count_buf[13:12], _05293_ }), .Y(_10452_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _35642_ ( .A({ _10455_, _10451_, _10454_ }), .Y(_10453_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _35643_ ( .A({ conv2d_16_row_count_buf[12], _05293_, _05294_, conv2d_16_row_count_buf[13] }), .Y(_10454_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35644_ ( .A({ conv2d_16_row_count_buf[14], conv2d_16_row_count_buf[15], _05295_, _05296_ }), .Y(_10455_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _35645_ ( .A({ _10477_, _10457_, _10467_, _10472_ }), .Y(_10456_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _35646_ ( .A({ _10463_, _10465_, _10466_, _10458_ }), .Y(_10457_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35647_ ( .A({ _10462_, _10459_, _10461_ }), .Y(_10458_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35648_ ( .A({ _10460_, _05309_, conv2d_16_row_count_buf[27] }), .Y(_10459_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35649_ ( .A({ _05308_, conv2d_16_row_count_buf[26], _05307_, conv2d_16_row_count_buf[25] }), .Y(_10460_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35650_ ( .A({ conv2d_16_row_count_buf[25], _05307_, conv2d_16_row_count_buf[24], _05306_ }), .Y(_10461_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35651_ ( .A({ conv2d_16_row_count_buf[26], _05308_, _05309_, conv2d_16_row_count_buf[27] }), .Y(_10462_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35652_ ( .A({ _10464_, conv2d_16_row_count_buf[31], _05314_ }), .Y(_10463_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35653_ ( .A({ _05313_, conv2d_16_row_count_buf[30], _05311_, conv2d_16_row_count_buf[29] }), .Y(_10464_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35654_ ( .A({ conv2d_16_row_count_buf[28], _05310_, conv2d_16_row_count_buf[29], _05311_ }), .Y(_10465_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35655_ ( .A({ _05310_, conv2d_16_row_count_buf[28] }), .Y(_10466_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35656_ ( .A({ _10471_, _10470_, _10469_, _10468_ }), .Y(_10467_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35657_ ( .A(conv2d_16_row_count_buf[23:20]), .Y(_10468_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35658_ ( .A(conv2d_16_row_count_buf[19:16]), .Y(_10469_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35659_ ( .A(conv2d_16_row_count_buf[31:28]), .Y(_10470_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35660_ ( .A(conv2d_16_row_count_buf[27:24]), .Y(_10471_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35661_ ( .A({ _10476_, _10475_, _10474_, _10473_ }), .Y(_10472_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35662_ ( .A(conv2d_16_row_count_buf[7:4]), .Y(_10473_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35663_ ( .A(conv2d_16_row_count_buf[3:0]), .Y(_10474_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35664_ ( .A(conv2d_16_row_count_buf[15:12]), .Y(_10475_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35665_ ( .A(conv2d_16_row_count_buf[11:8]), .Y(_10476_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35666_ ( .A({ conv2d_16_row_count_buf[30], conv2d_16_row_count_buf[31], _05313_, _05314_ }), .Y(_10477_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _35667_ ( .A({ _10483_, _10479_, _10446_, _10482_ }), .Y(_10478_) );
  \$lut  #( .LUT(16'h8f00), .WIDTH(4) ) _35668_ ( .A({ _10445_, _10481_, _10480_, _10448_ }), .Y(_10479_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _35669_ ( .A({ conv2d_16_row_count_buf[16], _05297_, _05298_, conv2d_16_row_count_buf[17] }), .Y(_10480_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35670_ ( .A({ conv2d_16_row_count_buf[18], conv2d_16_row_count_buf[19], _05299_, _05300_ }), .Y(_10481_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35671_ ( .A({ conv2d_16_row_count_buf[20], _05302_, _05303_, conv2d_16_row_count_buf[21] }), .Y(_10482_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35672_ ( .A({ conv2d_16_row_count_buf[22], conv2d_16_row_count_buf[23], _05304_, _05305_ }), .Y(_10483_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35673_ ( .A({ _10461_, _10485_, _10463_, _10459_ }), .Y(_10484_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _35674_ ( .A({ _10465_, _10466_, conv2d_16_row_count_buf[24], _05306_ }), .Y(_10485_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35675_ ( .A({ _10486_, _10428_ }), .Y(conv2d_16_stream_pad_mask_0_1) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _35676_ ( .A({ _10533_, _10523_, _10487_ }), .Y(_10486_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35677_ ( .A({ _13126_, _10520_, _10517_, _10488_ }), .Y(_10487_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35678_ ( .A({ _10501_, _10498_, _10504_, _10489_ }), .Y(_10488_) );
  \$lut  #( .LUT(16'hf100), .WIDTH(4) ) _35679_ ( .A({ _10497_, _10495_, _10496_, _10490_ }), .Y(_10489_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35680_ ( .A({ _10494_, _10493_, _10492_, _10491_ }), .Y(_10490_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35681_ ( .A({ _05408_, _05312_ }), .Y(_10491_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _35682_ ( .A({ _05290_, _05386_, _05397_, _05301_ }), .Y(_10492_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35683_ ( .A({ _05312_, _05408_, _05315_, _05411_ }), .Y(_10493_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35684_ ( .A({ _05411_, _05315_, _05412_, _05316_ }), .Y(_10494_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35685_ ( .A({ _05413_, _05317_ }), .Y(_10495_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35686_ ( .A({ _05316_, _05412_ }), .Y(_10496_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35687_ ( .A({ _05317_, _05413_, _05318_, _05414_ }), .Y(_10497_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35688_ ( .A({ _10500_, _10499_, _05319_, _05415_ }), .Y(_10498_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35689_ ( .A({ _05388_, _05292_, _05387_, _05291_ }), .Y(_10499_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35690_ ( .A({ _05321_, _05417_, _05416_, _05320_ }), .Y(_10500_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35691_ ( .A({ _10503_, _10499_, _10502_ }), .Y(_10501_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35692_ ( .A({ _05416_, _05320_, _05321_, _05417_ }), .Y(_10502_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35693_ ( .A({ _05387_, _05388_, _05291_, _05292_ }), .Y(_10503_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35694_ ( .A({ _05415_, _05319_, _05414_, _05318_ }), .Y(_10504_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35695_ ( .A({ _10508_, _10506_, _05310_, _05406_ }), .Y(_10505_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35696_ ( .A({ _10507_, _05410_, _05314_ }), .Y(_10506_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35697_ ( .A({ _05313_, _05409_, _05311_, _05407_ }), .Y(_10507_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35698_ ( .A({ _05406_, _05310_, _05407_, _05311_ }), .Y(_10508_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _35699_ ( .A({ _10512_, _10510_, _05398_, _05302_ }), .Y(_10509_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _35700_ ( .A({ _10511_, _05399_, _05303_ }), .Y(_10510_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35701_ ( .A({ _05401_, _05305_, _05400_, _05304_ }), .Y(_10511_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35702_ ( .A({ _05398_, _05302_, _05399_, _05303_ }), .Y(_10512_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35703_ ( .A({ _10515_, _10514_ }), .Y(_10513_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35704_ ( .A({ _05309_, _05405_, _05308_, _05404_ }), .Y(_10514_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35705_ ( .A({ _05306_, _05402_, _05403_, _05307_ }), .Y(_10515_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35706_ ( .A({ _05396_, _05300_, _05395_, _05299_ }), .Y(_10516_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35707_ ( .A({ _10519_, _10518_ }), .Y(_10517_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35708_ ( .A({ _05392_, _05296_, _05391_, _05295_ }), .Y(_10518_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35709_ ( .A({ _05294_, _05390_, _05293_, _05389_ }), .Y(_10519_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35710_ ( .A({ _10522_, _10518_, _10521_ }), .Y(_10520_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35711_ ( .A({ _05389_, _05293_, _05294_, _05390_ }), .Y(_10521_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35712_ ( .A({ _05391_, _05392_, _05295_, _05296_ }), .Y(_10522_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _35713_ ( .A({ _10505_, _10524_, _10530_ }), .Y(_10523_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35714_ ( .A({ _10513_, _10528_, _10509_, _10525_ }), .Y(_10524_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _35715_ ( .A({ _05300_, _05396_, _10526_ }), .Y(_10525_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _35716_ ( .A({ _05299_, _05395_, _10527_ }), .Y(_10526_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35717_ ( .A({ _05393_, _05297_, _05298_, _05394_ }), .Y(_10527_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35718_ ( .A({ _10529_, _10510_, _10512_ }), .Y(_10528_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35719_ ( .A({ _05400_, _05401_, _05304_, _05305_ }), .Y(_10529_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _35720_ ( .A({ _10531_, _10514_, _10532_ }), .Y(_10530_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _35721_ ( .A({ _05404_, _05308_, _05309_, _05405_ }), .Y(_10531_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35722_ ( .A({ _05402_, _05403_, _05306_, _05307_ }), .Y(_10532_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _35723_ ( .A({ _10545_, _10534_, _10506_, _10508_ }), .Y(_10533_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35724_ ( .A({ _10544_, _10543_, _10540_, _10535_ }), .Y(_10534_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35725_ ( .A({ _10539_, _10538_, _10537_, _10536_ }), .Y(_10535_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35726_ ( .A({ _05410_, _05409_, _05407_, _05406_ }), .Y(_10536_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35727_ ( .A({ _05405_, _05404_, _05403_, _05402_ }), .Y(_10537_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35728_ ( .A({ _05401_, _05400_, _05399_, _05398_ }), .Y(_10538_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35729_ ( .A({ _05396_, _05395_, _05394_, _05393_ }), .Y(_10539_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35730_ ( .A({ _10542_, _10541_ }), .Y(_10540_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35731_ ( .A({ _05392_, _05391_, _05390_, _05389_ }), .Y(_10541_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35732_ ( .A({ _05388_, _05387_, _05417_, _05416_ }), .Y(_10542_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35733_ ( .A({ _05415_, _05414_, _05413_, _05412_ }), .Y(_10543_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35734_ ( .A({ _05411_, _05408_, _05397_, _05386_ }), .Y(_10544_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35735_ ( .A({ _05409_, _05410_, _05313_, _05314_ }), .Y(_10545_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35736_ ( .A({ _10546_, _10428_ }), .Y(conv2d_16_stream_pad_mask_0_2) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35737_ ( .A({ _10583_, _10605_, _10578_, _10547_ }), .Y(_10546_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35738_ ( .A({ _10565_, _10575_, _10572_, _10548_ }), .Y(_10547_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35739_ ( .A({ _10561_, _10558_, _10564_, _10549_ }), .Y(_10548_) );
  \$lut  #( .LUT(16'h00f4), .WIDTH(4) ) _35740_ ( .A({ _10555_, _10556_, _10557_, _10550_ }), .Y(_10549_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _35741_ ( .A({ _10554_, _10553_, _10551_, _10552_ }), .Y(_10550_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35742_ ( .A({ _05440_, _05312_ }), .Y(_10551_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35743_ ( .A({ _05290_, _05418_, _05429_, _05301_ }), .Y(_10552_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35744_ ( .A({ _05312_, _05440_, _05315_, _05443_ }), .Y(_10553_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35745_ ( .A({ _05443_, _05315_, _05444_, _05316_ }), .Y(_10554_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35746_ ( .A({ _05318_, _05446_ }), .Y(_10555_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35747_ ( .A({ _05445_, _05317_ }), .Y(_10556_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35748_ ( .A({ _05316_, _05444_, _05317_, _05445_ }), .Y(_10557_) );
  \$lut  #( .LUT(16'h9000), .WIDTH(4) ) _35749_ ( .A({ _10560_, _10559_, _05321_, _05449_ }), .Y(_10558_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35750_ ( .A({ _05420_, _05292_, _05419_, _05291_ }), .Y(_10559_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35751_ ( .A({ _05448_, _05320_, _05319_, _05447_ }), .Y(_10560_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35752_ ( .A({ _10563_, _10559_, _10562_ }), .Y(_10561_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35753_ ( .A({ _05448_, _05320_, _05321_, _05449_ }), .Y(_10562_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35754_ ( .A({ _05419_, _05420_, _05291_, _05292_ }), .Y(_10563_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35755_ ( .A({ _05447_, _05319_, _05446_, _05318_ }), .Y(_10564_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35756_ ( .A({ _10571_, _10570_, _10566_ }), .Y(_10565_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _35757_ ( .A({ _10569_, _10567_, _05430_, _05302_ }), .Y(_10566_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35758_ ( .A({ _10568_, _05433_, _05305_ }), .Y(_10567_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35759_ ( .A({ _05432_, _05304_, _05303_, _05431_ }), .Y(_10568_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35760_ ( .A({ _05430_, _05302_, _05431_, _05303_ }), .Y(_10569_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35761_ ( .A({ _05428_, _05300_, _05427_, _05299_ }), .Y(_10570_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35762_ ( .A({ _05298_, _05426_, _05425_, _05297_ }), .Y(_10571_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35763_ ( .A({ _10574_, _10573_ }), .Y(_10572_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35764_ ( .A({ _05424_, _05296_, _05423_, _05295_ }), .Y(_10573_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35765_ ( .A({ _05294_, _05422_, _05293_, _05421_ }), .Y(_10574_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35766_ ( .A({ _10577_, _10573_, _10576_ }), .Y(_10575_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35767_ ( .A({ _05421_, _05293_, _05294_, _05422_ }), .Y(_10576_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35768_ ( .A({ _05423_, _05424_, _05295_, _05296_ }), .Y(_10577_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _35769_ ( .A({ _10582_, _10579_, _10567_, _10569_ }), .Y(_10578_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _35770_ ( .A({ _10566_, _10580_, _10581_, _10570_ }), .Y(_10579_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35771_ ( .A({ _05427_, _05428_, _05299_, _05300_ }), .Y(_10580_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _35772_ ( .A({ _05425_, _05297_, _05298_, _05426_ }), .Y(_10581_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35773_ ( .A({ _05432_, _05433_, _05304_, _05305_ }), .Y(_10582_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _35774_ ( .A({ _10604_, _10591_, _10584_, _10602_ }), .Y(_10583_) );
  \$lut  #( .LUT(16'hf400), .WIDTH(4) ) _35775_ ( .A({ _10590_, _10585_, _05310_, _05438_ }), .Y(_10584_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35776_ ( .A({ _10589_, _10586_, _10588_ }), .Y(_10585_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35777_ ( .A({ _10587_, _05308_, _05436_ }), .Y(_10586_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35778_ ( .A({ _05309_, _05437_, _05307_, _05435_ }), .Y(_10587_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35779_ ( .A({ _05435_, _05307_, _05434_, _05306_ }), .Y(_10588_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35780_ ( .A({ _05436_, _05308_, _05309_, _05437_ }), .Y(_10589_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35781_ ( .A({ _05438_, _05310_, _05439_, _05311_ }), .Y(_10590_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _35782_ ( .A({ _10592_, _10597_, _10595_, _05443_ }), .Y(_10591_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35783_ ( .A({ _10594_, _10593_ }), .Y(_10592_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35784_ ( .A({ _05433_, _05432_, _05431_, _05430_ }), .Y(_10593_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35785_ ( .A({ _05428_, _05427_, _05426_, _05425_ }), .Y(_10594_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35786_ ( .A({ _10596_, _05440_, _05429_, _05418_ }), .Y(_10595_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35787_ ( .A({ _05447_, _05446_, _05445_, _05444_ }), .Y(_10596_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35788_ ( .A({ _10601_, _10600_, _10599_, _10598_ }), .Y(_10597_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35789_ ( .A({ _05442_, _05441_, _05439_, _05438_ }), .Y(_10598_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35790_ ( .A({ _05437_, _05436_, _05435_, _05434_ }), .Y(_10599_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35791_ ( .A({ _05424_, _05423_, _05422_, _05421_ }), .Y(_10600_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35792_ ( .A({ _05420_, _05419_, _05449_, _05448_ }), .Y(_10601_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35793_ ( .A({ _10603_, _05442_, _05314_ }), .Y(_10602_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35794_ ( .A({ _05313_, _05441_, _05311_, _05439_ }), .Y(_10603_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35795_ ( .A({ _05441_, _05442_, _05313_, _05314_ }), .Y(_10604_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35796_ ( .A({ _10602_, _10606_ }), .Y(_10605_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35797_ ( .A({ _10607_, _10590_, _10588_, _10586_ }), .Y(_10606_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35798_ ( .A({ _05310_, _05438_, _05306_, _05434_ }), .Y(_10607_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35799_ ( .A({ _10608_, _10377_ }), .Y(conv2d_16_stream_pad_mask_1_0) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35800_ ( .A({ _10645_, _10667_, _10640_, _10609_ }), .Y(_10608_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35801_ ( .A({ _10627_, _10637_, _10634_, _10610_ }), .Y(_10609_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35802_ ( .A({ _10623_, _10620_, _10626_, _10611_ }), .Y(_10610_) );
  \$lut  #( .LUT(16'hf100), .WIDTH(4) ) _35803_ ( .A({ _10619_, _10617_, _10618_, _10612_ }), .Y(_10611_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _35804_ ( .A({ _10616_, _10615_, _10613_, _10614_ }), .Y(_10612_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35805_ ( .A({ _05290_, _05450_, _05461_, _05301_ }), .Y(_10613_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35806_ ( .A({ _05472_, _05312_, _05315_, _05475_ }), .Y(_10614_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35807_ ( .A({ _05476_, _05316_ }), .Y(_10615_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35808_ ( .A({ _05472_, _05475_, _05312_, _05315_ }), .Y(_10616_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35809_ ( .A({ _05477_, _05317_ }), .Y(_10617_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35810_ ( .A({ _05316_, _05476_ }), .Y(_10618_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35811_ ( .A({ _05317_, _05477_, _05318_, _05478_ }), .Y(_10619_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35812_ ( .A({ _10622_, _10621_, _05319_, _05479_ }), .Y(_10620_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35813_ ( .A({ _05452_, _05292_, _05451_, _05291_ }), .Y(_10621_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35814_ ( .A({ _05321_, _05481_, _05480_, _05320_ }), .Y(_10622_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35815_ ( .A({ _10625_, _10621_, _10624_ }), .Y(_10623_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35816_ ( .A({ _05480_, _05320_, _05321_, _05481_ }), .Y(_10624_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35817_ ( .A({ _05451_, _05452_, _05291_, _05292_ }), .Y(_10625_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35818_ ( .A({ _05479_, _05319_, _05478_, _05318_ }), .Y(_10626_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35819_ ( .A({ _10633_, _10632_, _10628_ }), .Y(_10627_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _35820_ ( .A({ _10631_, _10629_, _05462_, _05302_ }), .Y(_10628_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35821_ ( .A({ _10630_, _05465_, _05305_ }), .Y(_10629_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35822_ ( .A({ _05464_, _05304_, _05303_, _05463_ }), .Y(_10630_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35823_ ( .A({ _05462_, _05302_, _05463_, _05303_ }), .Y(_10631_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35824_ ( .A({ _05460_, _05300_, _05459_, _05299_ }), .Y(_10632_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35825_ ( .A({ _05298_, _05458_, _05457_, _05297_ }), .Y(_10633_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35826_ ( .A({ _10635_, _05294_, _05454_ }), .Y(_10634_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35827_ ( .A({ _10636_, _05293_, _05453_ }), .Y(_10635_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35828_ ( .A({ _05456_, _05296_, _05455_, _05295_ }), .Y(_10636_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _35829_ ( .A({ _10639_, _10636_, _10638_ }), .Y(_10637_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35830_ ( .A({ _05453_, _05293_, _05294_, _05454_ }), .Y(_10638_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35831_ ( .A({ _05455_, _05456_, _05295_, _05296_ }), .Y(_10639_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _35832_ ( .A({ _10644_, _10641_, _10629_, _10631_ }), .Y(_10640_) );
  \$lut  #( .LUT(16'hf400), .WIDTH(4) ) _35833_ ( .A({ _10628_, _10643_, _10632_, _10642_ }), .Y(_10641_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35834_ ( .A({ _05457_, _05297_, _05298_, _05458_ }), .Y(_10642_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35835_ ( .A({ _05459_, _05460_, _05299_, _05300_ }), .Y(_10643_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35836_ ( .A({ _05464_, _05465_, _05304_, _05305_ }), .Y(_10644_) );
  \$lut  #( .LUT(16'h0d00), .WIDTH(4) ) _35837_ ( .A({ _10666_, _10653_, _10646_, _10664_ }), .Y(_10645_) );
  \$lut  #( .LUT(16'hf400), .WIDTH(4) ) _35838_ ( .A({ _10652_, _10647_, _05310_, _05470_ }), .Y(_10646_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35839_ ( .A({ _10651_, _10648_, _10650_ }), .Y(_10647_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35840_ ( .A({ _10649_, _05309_, _05469_ }), .Y(_10648_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35841_ ( .A({ _05308_, _05468_, _05307_, _05467_ }), .Y(_10649_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35842_ ( .A({ _05467_, _05307_, _05466_, _05306_ }), .Y(_10650_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35843_ ( .A({ _05468_, _05308_, _05309_, _05469_ }), .Y(_10651_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35844_ ( .A({ _05470_, _05310_, _05471_, _05311_ }), .Y(_10652_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35845_ ( .A({ _10663_, _10662_, _10657_, _10654_ }), .Y(_10653_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35846_ ( .A({ _10656_, _10655_ }), .Y(_10654_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35847_ ( .A({ _05465_, _05464_, _05463_, _05462_ }), .Y(_10655_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35848_ ( .A({ _05460_, _05459_, _05458_, _05457_ }), .Y(_10656_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35849_ ( .A({ _10661_, _10660_, _10659_, _10658_ }), .Y(_10657_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35850_ ( .A({ _05452_, _05451_, _05481_, _05480_ }), .Y(_10658_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35851_ ( .A({ _05456_, _05455_, _05454_, _05453_ }), .Y(_10659_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35852_ ( .A({ _05479_, _05478_, _05477_, _05476_ }), .Y(_10660_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35853_ ( .A({ _05475_, _05472_, _05461_, _05450_ }), .Y(_10661_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35854_ ( .A({ _05474_, _05473_, _05471_, _05470_ }), .Y(_10662_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35855_ ( .A({ _05469_, _05468_, _05467_, _05466_ }), .Y(_10663_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35856_ ( .A({ _10665_, _05474_, _05314_ }), .Y(_10664_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35857_ ( .A({ _05313_, _05473_, _05311_, _05471_ }), .Y(_10665_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35858_ ( .A({ _05473_, _05474_, _05313_, _05314_ }), .Y(_10666_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35859_ ( .A({ _10648_, _10668_ }), .Y(_10667_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35860_ ( .A({ _10669_, _10650_, _10652_, _10664_ }), .Y(_10668_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35861_ ( .A({ _05310_, _05470_, _05306_, _05466_ }), .Y(_10669_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35862_ ( .A({ _10608_, _10486_ }), .Y(conv2d_16_stream_pad_mask_1_1) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35863_ ( .A({ _10608_, _10546_ }), .Y(conv2d_16_stream_pad_mask_1_2) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35864_ ( .A({ _10670_, _10377_ }), .Y(conv2d_16_stream_pad_mask_2_0) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35865_ ( .A({ _10707_, _10729_, _10702_, _10671_ }), .Y(_10670_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35866_ ( .A({ _10689_, _10699_, _10696_, _10672_ }), .Y(_10671_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _35867_ ( .A({ _10685_, _10682_, _10688_, _10673_ }), .Y(_10672_) );
  \$lut  #( .LUT(16'h00f4), .WIDTH(4) ) _35868_ ( .A({ _10679_, _10680_, _10681_, _10674_ }), .Y(_10673_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _35869_ ( .A({ _10678_, _10677_, _10675_, _10676_ }), .Y(_10674_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35870_ ( .A({ _05290_, _05482_, _05493_, _05301_ }), .Y(_10675_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35871_ ( .A({ _05504_, _05312_, _05315_, _05507_ }), .Y(_10676_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35872_ ( .A({ _05508_, _05316_ }), .Y(_10677_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35873_ ( .A({ _05504_, _05507_, _05312_, _05315_ }), .Y(_10678_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35874_ ( .A({ _05318_, _05510_ }), .Y(_10679_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35875_ ( .A({ _05509_, _05317_ }), .Y(_10680_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35876_ ( .A({ _05316_, _05508_, _05317_, _05509_ }), .Y(_10681_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35877_ ( .A({ _10684_, _10683_, _05319_, _05511_ }), .Y(_10682_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35878_ ( .A({ _05484_, _05292_, _05483_, _05291_ }), .Y(_10683_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35879_ ( .A({ _05321_, _05513_, _05512_, _05320_ }), .Y(_10684_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35880_ ( .A({ _10687_, _10683_, _10686_ }), .Y(_10685_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35881_ ( .A({ _05512_, _05320_, _05321_, _05513_ }), .Y(_10686_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35882_ ( .A({ _05483_, _05484_, _05291_, _05292_ }), .Y(_10687_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35883_ ( .A({ _05511_, _05319_, _05510_, _05318_ }), .Y(_10688_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35884_ ( .A({ _10695_, _10694_, _10690_ }), .Y(_10689_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _35885_ ( .A({ _10693_, _10691_, _05494_, _05302_ }), .Y(_10690_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35886_ ( .A({ _10692_, _05497_, _05305_ }), .Y(_10691_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35887_ ( .A({ _05496_, _05304_, _05303_, _05495_ }), .Y(_10692_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35888_ ( .A({ _05494_, _05302_, _05495_, _05303_ }), .Y(_10693_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35889_ ( .A({ _05492_, _05300_, _05491_, _05299_ }), .Y(_10694_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35890_ ( .A({ _05298_, _05490_, _05489_, _05297_ }), .Y(_10695_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35891_ ( .A({ _10698_, _10697_ }), .Y(_10696_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35892_ ( .A({ _05488_, _05296_, _05487_, _05295_ }), .Y(_10697_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35893_ ( .A({ _05294_, _05486_, _05293_, _05485_ }), .Y(_10698_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _35894_ ( .A({ _10701_, _10697_, _10700_ }), .Y(_10699_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _35895_ ( .A({ _05485_, _05293_, _05294_, _05486_ }), .Y(_10700_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35896_ ( .A({ _05487_, _05488_, _05295_, _05296_ }), .Y(_10701_) );
  \$lut  #( .LUT(16'h0b00), .WIDTH(4) ) _35897_ ( .A({ _10706_, _10703_, _10691_, _10693_ }), .Y(_10702_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _35898_ ( .A({ _10690_, _10704_, _10705_, _10694_ }), .Y(_10703_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35899_ ( .A({ _05491_, _05492_, _05299_, _05300_ }), .Y(_10704_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _35900_ ( .A({ _05489_, _05297_, _05298_, _05490_ }), .Y(_10705_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35901_ ( .A({ _05496_, _05497_, _05304_, _05305_ }), .Y(_10706_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _35902_ ( .A({ _10728_, _10717_, _10716_, _10708_ }), .Y(_10707_) );
  \$lut  #( .LUT(16'hf800), .WIDTH(4) ) _35903_ ( .A({ _10709_, _10714_, _10715_, _10713_ }), .Y(_10708_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _35904_ ( .A({ _10712_, _10710_, _05310_, _05502_ }), .Y(_10709_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _35905_ ( .A({ _10711_, _05506_, _05314_ }), .Y(_10710_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _35906_ ( .A({ _05313_, _05505_, _05311_, _05503_ }), .Y(_10711_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35907_ ( .A({ _05502_, _05310_, _05503_, _05311_ }), .Y(_10712_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35908_ ( .A({ _05309_, _05501_, _05308_, _05500_ }), .Y(_10713_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _35909_ ( .A({ _05500_, _05308_, _05309_, _05501_ }), .Y(_10714_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _35910_ ( .A({ _05498_, _05499_, _05306_, _05307_ }), .Y(_10715_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35911_ ( .A({ _10710_, _10712_ }), .Y(_10716_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35912_ ( .A({ _10727_, _10726_, _10721_, _10718_ }), .Y(_10717_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35913_ ( .A({ _10720_, _10719_ }), .Y(_10718_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35914_ ( .A({ _05497_, _05496_, _05495_, _05494_ }), .Y(_10719_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35915_ ( .A({ _05492_, _05491_, _05490_, _05489_ }), .Y(_10720_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35916_ ( .A({ _10725_, _10724_, _10723_, _10722_ }), .Y(_10721_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35917_ ( .A({ _05511_, _05510_, _05509_, _05508_ }), .Y(_10722_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35918_ ( .A({ _05507_, _05504_, _05493_, _05482_ }), .Y(_10723_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35919_ ( .A({ _05488_, _05487_, _05486_, _05485_ }), .Y(_10724_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35920_ ( .A({ _05484_, _05483_, _05513_, _05512_ }), .Y(_10725_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35921_ ( .A({ _05506_, _05505_, _05503_, _05502_ }), .Y(_10726_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35922_ ( .A({ _05501_, _05500_, _05499_, _05498_ }), .Y(_10727_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _35923_ ( .A({ _05505_, _05506_, _05313_, _05314_ }), .Y(_10728_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35924_ ( .A({ _10730_, _10713_, _10709_ }), .Y(_10729_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _35925_ ( .A({ _05306_, _05498_, _05499_, _05307_ }), .Y(_10730_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35926_ ( .A({ _10670_, _10486_ }), .Y(conv2d_16_stream_pad_mask_2_1) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35927_ ( .A({ _10670_, _10546_ }), .Y(conv2d_16_stream_pad_mask_2_2) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35928_ ( .A({ _09303_, _stream_conv2d_16_source_busy }), .Y(_06874_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35929_ ( .A({ _10737_, _10736_, _10731_ }), .Y(_stream_conv2d_16_done) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _35930_ ( .A({ _10735_, _10734_, _10732_ }), .Y(_10731_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35931_ ( .A({ _stream_conv2d_16_source_8_idle, _stream_conv2d_16_source_6_idle, _stream_conv2d_16_source_36_idle, _10733_ }), .Y(_10732_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35932_ ( .A({ _stream_conv2d_16_source_35_idle, _stream_conv2d_16_source_34_idle, _stream_conv2d_16_source_33_idle, _stream_conv2d_16_source_32_idle }), .Y(_10733_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35933_ ( .A({ _stream_conv2d_16_source_31_idle, _stream_conv2d_16_source_30_idle, _stream_conv2d_16_source_29_idle, _stream_conv2d_16_source_28_idle }), .Y(_10734_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35934_ ( .A({ _stream_conv2d_16_source_27_idle, _stream_conv2d_16_source_26_idle, _stream_conv2d_16_source_25_idle, _stream_conv2d_16_source_24_idle }), .Y(_10735_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35935_ ( .A({ _stream_conv2d_16_source_23_idle, _stream_conv2d_16_source_22_idle, _stream_conv2d_16_source_21_idle, _stream_conv2d_16_source_20_idle }), .Y(_10736_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35936_ ( .A({ _stream_conv2d_16_source_19_idle, _stream_conv2d_16_source_14_idle, _stream_conv2d_16_source_12_idle, _stream_conv2d_16_source_10_idle }), .Y(_10737_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35937_ ( .A({ _13131_, _10738_ }), .Y(max_pool_serial_18_stream_pad_mask_0_0) );
  \$lut  #( .LUT(16'hb200), .WIDTH(4) ) _35938_ ( .A({ _10742_, cparam_max_pool_serial_18_act_num_col[5], max_pool_serial_18_col_count[5], _13128_ }), .Y(_10738_) );
  \$lut  #( .LUT(16'ha8fe), .WIDTH(4) ) _35939_ ( .A({ cparam_max_pool_serial_18_act_num_col[2], _10740_, _10741_, max_pool_serial_18_col_count[2] }), .Y(_10739_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35940_ ( .A({ cparam_max_pool_serial_18_act_num_col[1], max_pool_serial_18_col_count[1], cparam_max_pool_serial_18_act_num_col[0], max_pool_serial_18_col_count[0] }), .Y(_10740_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35941_ ( .A({ max_pool_serial_18_col_count[1], cparam_max_pool_serial_18_act_num_col[1] }), .Y(_10741_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _35942_ ( .A({ _09391_, _09387_ }), .Y(_10742_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _35943_ ( .A({ max_pool_serial_18_row_count_buf[3], cparam_max_pool_serial_18_act_num_col[3], _10744_ }), .Y(_10743_) );
  \$lut  #( .LUT(16'hddd4), .WIDTH(4) ) _35944_ ( .A({ _10746_, _10745_, max_pool_serial_18_row_count_buf[2], cparam_max_pool_serial_18_act_num_col[2] }), .Y(_10744_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35945_ ( .A({ max_pool_serial_18_row_count_buf[1], cparam_max_pool_serial_18_act_num_col[1] }), .Y(_10745_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35946_ ( .A({ cparam_max_pool_serial_18_act_num_col[0], max_pool_serial_18_row_count_buf[0], cparam_max_pool_serial_18_act_num_col[1], max_pool_serial_18_row_count_buf[1] }), .Y(_10746_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35947_ ( .A(max_pool_serial_18_row_count_buf[7:6]), .Y(_10747_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35948_ ( .A({ _10753_, _10752_, _10751_, _10749_ }), .Y(_10748_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35949_ ( .A({ _10750_, _10747_, max_pool_serial_18_row_count_buf[11], max_pool_serial_18_row_count_buf[8] }), .Y(_10749_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35950_ ( .A({ max_pool_serial_18_row_count_buf[19], max_pool_serial_18_row_count_buf[16], max_pool_serial_18_row_count_buf[14:13] }), .Y(_10750_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35951_ ( .A(max_pool_serial_18_row_count_buf[31:28]), .Y(_10751_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35952_ ( .A({ max_pool_serial_18_row_count_buf[27], max_pool_serial_18_row_count_buf[24], max_pool_serial_18_row_count_buf[22:21] }), .Y(_10752_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35953_ ( .A({ max_pool_serial_18_row_count_buf[26:25], max_pool_serial_18_row_count_buf[23], max_pool_serial_18_row_count_buf[20] }), .Y(_10753_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35954_ ( .A({ max_pool_serial_18_row_count_buf[18:17], max_pool_serial_18_row_count_buf[15], max_pool_serial_18_row_count_buf[12] }), .Y(_10754_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35955_ ( .A({ _13134_, _13131_ }), .Y(max_pool_serial_18_stream_pad_mask_0_1) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _35956_ ( .A({ _03937_, cparam_max_pool_serial_18_act_num_col[3], _10756_ }), .Y(_10755_) );
  \$lut  #( .LUT(16'hddd4), .WIDTH(4) ) _35957_ ( .A({ _10758_, _10757_, _03934_, cparam_max_pool_serial_18_act_num_col[2] }), .Y(_10756_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35958_ ( .A({ _03923_, cparam_max_pool_serial_18_act_num_col[1] }), .Y(_10757_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35959_ ( .A({ cparam_max_pool_serial_18_act_num_col[0], _03912_, cparam_max_pool_serial_18_act_num_col[1], _03923_ }), .Y(_10758_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35960_ ( .A({ _03941_, _03940_ }), .Y(_10759_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35961_ ( .A({ _10765_, _10764_, _10763_, _10761_ }), .Y(_10760_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35962_ ( .A({ _10762_, _10759_, _03914_, _03942_ }), .Y(_10761_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35963_ ( .A({ _03922_, _03919_, _03917_, _03916_ }), .Y(_10762_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35964_ ( .A({ _03936_, _03935_, _03933_, _03932_ }), .Y(_10763_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35965_ ( .A({ _03931_, _03928_, _03926_, _03925_ }), .Y(_10764_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35966_ ( .A({ _03930_, _03929_, _03927_, _03924_ }), .Y(_10765_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35967_ ( .A({ _03921_, _03920_, _03918_, _03915_ }), .Y(_10766_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35968_ ( .A({ _13136_, _10738_ }), .Y(max_pool_serial_18_stream_pad_mask_1_0) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _35969_ ( .A({ _03970_, cparam_max_pool_serial_18_act_num_col[4], _10768_ }), .Y(_10767_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _35970_ ( .A({ _03969_, cparam_max_pool_serial_18_act_num_col[3], _10769_ }), .Y(_10768_) );
  \$lut  #( .LUT(16'hddd4), .WIDTH(4) ) _35971_ ( .A({ _10771_, _10770_, _03966_, cparam_max_pool_serial_18_act_num_col[2] }), .Y(_10769_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _35972_ ( .A({ _03955_, cparam_max_pool_serial_18_act_num_col[1] }), .Y(_10770_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _35973_ ( .A({ cparam_max_pool_serial_18_act_num_col[0], _03944_, cparam_max_pool_serial_18_act_num_col[1], _03955_ }), .Y(_10771_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _35974_ ( .A({ _03973_, _03972_ }), .Y(_10772_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35975_ ( .A({ _10778_, _10777_, _10776_, _10774_ }), .Y(_10773_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _35976_ ( .A({ _10775_, _10772_, _03946_, _03974_ }), .Y(_10774_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35977_ ( .A({ _03954_, _03951_, _03949_, _03948_ }), .Y(_10775_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35978_ ( .A({ _03968_, _03967_, _03965_, _03964_ }), .Y(_10776_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35979_ ( .A({ _03963_, _03960_, _03958_, _03957_ }), .Y(_10777_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35980_ ( .A({ _03962_, _03961_, _03959_, _03956_ }), .Y(_10778_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35981_ ( .A({ _03953_, _03952_, _03950_, _03947_ }), .Y(_10779_) );
  \$lut  #( .LUT(4'h7), .WIDTH(2) ) _35982_ ( .A({ _13136_, _13134_ }), .Y(max_pool_serial_18_stream_pad_mask_1_1) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _35983_ ( .A({ _10795_, _10790_, _10785_, _10780_ }), .Y(matmul_29_stream_pad_mask_0_0) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35984_ ( .A({ _10784_, _10783_, _10782_, _10781_ }), .Y(_10780_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35985_ ( .A(matmul_29_row_count_buf[22:19]), .Y(_10781_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35986_ ( .A(matmul_29_row_count_buf[18:15]), .Y(_10782_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35987_ ( .A(matmul_29_row_count_buf[30:27]), .Y(_10783_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35988_ ( .A(matmul_29_row_count_buf[26:23]), .Y(_10784_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35989_ ( .A({ _10789_, _10788_, _10787_, _10786_ }), .Y(_10785_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35990_ ( .A(matmul_29_row_count_buf[6:3]), .Y(_10786_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35991_ ( .A({ matmul_29_row_count_buf[2:1], matmul_29_col_count[0], matmul_29_row_count_buf[0] }), .Y(_10787_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35992_ ( .A(matmul_29_row_count_buf[14:11]), .Y(_10788_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35993_ ( .A(matmul_29_row_count_buf[10:7]), .Y(_10789_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35994_ ( .A({ _10794_, _10793_, _10792_, _10791_ }), .Y(_10790_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35995_ ( .A(matmul_29_col_count[23:20]), .Y(_10791_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35996_ ( .A(matmul_29_col_count[19:16]), .Y(_10792_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35997_ ( .A(matmul_29_col_count[31:28]), .Y(_10793_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _35998_ ( .A(matmul_29_col_count[27:24]), .Y(_10794_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _35999_ ( .A({ _10799_, _10798_, _10797_, _10796_ }), .Y(_10795_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36000_ ( .A(matmul_29_col_count[7:4]), .Y(_10796_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36001_ ( .A({ matmul_29_col_count[3:1], matmul_29_row_count_buf[31] }), .Y(_10797_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36002_ ( .A(matmul_29_col_count[15:12]), .Y(_10798_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36003_ ( .A(matmul_29_col_count[11:8]), .Y(_10799_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36004_ ( .A({ _08872_, _stream_matmul_29_source_busy }), .Y(_06177_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36005_ ( .A({ _stream_matmul_29_source_8_idle, _stream_matmul_29_source_6_idle, _stream_matmul_29_source_20_idle, _10800_ }), .Y(_stream_matmul_29_done) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36006_ ( .A({ _stream_matmul_29_source_19_idle, _stream_matmul_29_source_14_idle, _stream_matmul_29_source_12_idle, _stream_matmul_29_source_10_idle }), .Y(_10800_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _36007_ ( .A({ _tmp_1357, maxi_wready, maxi_wvalid }), .Y(_06178_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _36008_ ( .A({ _tmp_1120, maxi_wready, maxi_wvalid }), .Y(_06179_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _36009_ ( .A({ _tmp_1020, maxi_wready, maxi_wvalid }), .Y(_06180_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36010_ ( .A({ maxi_arvalid, maxi_arready }), .Y(_06182_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36011_ ( .A({ _09893_, _10801_, _06182_ }), .Y(_06181_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36012_ ( .A({ _10802_, _tmp_20[4:3] }), .Y(_10801_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36013_ ( .A({ _10803_, _tmp_20[8:6] }), .Y(_10802_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36014_ ( .A({ _tmp_20[5], _tmp_20[2:0] }), .Y(_10803_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36015_ ( .A({ _10804_, _10801_ }), .Y(_06183_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36016_ ( .A({ maxi_rvalid, maxi_rready }), .Y(_10804_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36017_ ( .A({ _07033_, _10805_, _06186_ }), .Y(_06184_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36018_ ( .A({ _10806_, _tmp_1019[0] }), .Y(_10805_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36019_ ( .A({ _10808_, _10807_ }), .Y(_10806_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36020_ ( .A(_tmp_1019[8:5]), .Y(_10807_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36021_ ( .A(_tmp_1019[4:1]), .Y(_10808_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36022_ ( .A({ maxi_awvalid, maxi_awready }), .Y(_06186_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36023_ ( .A({ _10818_, _10816_, _10809_, _06184_ }), .Y(_06185_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36024_ ( .A({ _10815_, _10810_, _maxi_write_cur_size[1:0] }), .Y(_10809_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36025_ ( .A({ _10814_, _10813_, _10812_, _10811_ }), .Y(_10810_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36026_ ( .A(_maxi_write_cur_size[13:10]), .Y(_10811_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36027_ ( .A(_maxi_write_cur_size[9:6]), .Y(_10812_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36028_ ( .A(_maxi_write_cur_size[21:18]), .Y(_10813_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36029_ ( .A(_maxi_write_cur_size[17:14]), .Y(_10814_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36030_ ( .A(_maxi_write_cur_size[5:2]), .Y(_10815_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36031_ ( .A({ _10817_, _maxi_write_cur_size[32:30] }), .Y(_10816_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36032_ ( .A({ _maxi_write_cur_size[28:27], _maxi_write_cur_size[25], _maxi_write_cur_size[22] }), .Y(_10817_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36033_ ( .A({ _maxi_write_cur_size[29], _maxi_write_cur_size[26], _maxi_write_cur_size[24:23] }), .Y(_10818_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _36034_ ( .A({ _dataflow_cat_valid_98, _10820_, _10819_ }), .Y(_06187_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36035_ ( .A({ _07030_, _06189_, _10805_ }), .Y(_10819_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36036_ ( .A({ maxi_wvalid, maxi_wready }), .Y(_06189_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _36037_ ( .A({ _maxi_write_op_sel[0], _10821_, _10822_, _maxi_write_op_sel[1] }), .Y(_10820_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36038_ ( .A(_maxi_write_op_sel[7:4]), .Y(_10821_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36039_ ( .A(_maxi_write_op_sel[3:2]), .Y(_10822_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36040_ ( .A({ _10823_, _06187_ }), .Y(_06188_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36041_ ( .A({ _tmp_1019[0], _10806_ }), .Y(_10823_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _36042_ ( .A({ _dataflow_cat_valid_107, _10824_, _10819_ }), .Y(_06190_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _36043_ ( .A({ _10821_, _maxi_write_op_sel[1], _10822_, _maxi_write_op_sel[0] }), .Y(_10824_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36044_ ( .A({ _10823_, _06190_ }), .Y(_06191_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _36045_ ( .A({ _dataflow_cat_valid_167, _10825_, _10819_ }), .Y(_06192_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36046_ ( .A({ _maxi_write_op_sel[0], _maxi_write_op_sel[1], _10822_, _10821_ }), .Y(_10825_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36047_ ( .A({ _10823_, _06192_ }), .Y(_06193_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36048_ ( .A({ _dataflow_slice_valid_3, _10826_ }), .Y(_06194_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36049_ ( .A({ _tmp_13, _10827_ }), .Y(_10826_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36050_ ( .A({ _10828_, _tmp_12[0], _tmp_12[33:32] }), .Y(_10827_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36051_ ( .A({ _10837_, _10836_, _10834_, _10829_ }), .Y(_10828_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36052_ ( .A({ _10833_, _10832_, _10831_, _10830_ }), .Y(_10829_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36053_ ( .A({ _tmp_12[24], _tmp_12[21], _tmp_12[19:18] }), .Y(_10830_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36054_ ( .A({ _tmp_12[31], _tmp_12[29:28], _tmp_12[25] }), .Y(_10831_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36055_ ( .A({ _tmp_12[7:6], _tmp_12[4], _tmp_12[1] }), .Y(_10832_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36056_ ( .A({ _tmp_12[16], _tmp_12[13], _tmp_12[11:10] }), .Y(_10833_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36057_ ( .A({ _10835_, _tmp_12[30], _tmp_12[27:26] }), .Y(_10834_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36058_ ( .A({ _tmp_12[23:22], _tmp_12[20], _tmp_12[17] }), .Y(_10835_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36059_ ( .A({ _tmp_12[8], _tmp_12[5], _tmp_12[3:2] }), .Y(_10836_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36060_ ( .A({ _tmp_12[15:14], _tmp_12[12], _tmp_12[9] }), .Y(_10837_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36061_ ( .A({ _wvalid_11, _06194_ }), .Y(_06195_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36062_ ( .A({ _dataflow_slice_valid_6, _10838_ }), .Y(_06197_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36063_ ( .A({ _tmp_15, _10839_ }), .Y(_10838_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36064_ ( .A({ _10840_, _tmp_14[0], _tmp_14[33:32] }), .Y(_10839_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36065_ ( .A({ _10849_, _10848_, _10846_, _10841_ }), .Y(_10840_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36066_ ( .A({ _10845_, _10844_, _10843_, _10842_ }), .Y(_10841_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36067_ ( .A({ _tmp_14[24], _tmp_14[21], _tmp_14[19:18] }), .Y(_10842_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36068_ ( .A({ _tmp_14[31], _tmp_14[29:28], _tmp_14[25] }), .Y(_10843_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36069_ ( .A({ _tmp_14[7:6], _tmp_14[4], _tmp_14[1] }), .Y(_10844_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36070_ ( .A({ _tmp_14[16], _tmp_14[13], _tmp_14[11:10] }), .Y(_10845_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36071_ ( .A({ _10847_, _tmp_14[30], _tmp_14[27:26] }), .Y(_10846_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36072_ ( .A({ _tmp_14[23:22], _tmp_14[20], _tmp_14[17] }), .Y(_10847_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36073_ ( .A({ _tmp_14[8], _tmp_14[5], _tmp_14[3:2] }), .Y(_10848_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36074_ ( .A({ _tmp_14[15:14], _tmp_14[12], _tmp_14[9] }), .Y(_10849_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36075_ ( .A({ _wvalid_11, _06197_ }), .Y(_06198_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36076_ ( .A({ _dataflow_slice_valid_9, _10850_ }), .Y(_06200_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36077_ ( .A({ _tmp_17, _10851_ }), .Y(_10850_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36078_ ( .A({ _10852_, _tmp_16[0], _tmp_16[33:32] }), .Y(_10851_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36079_ ( .A({ _10861_, _10860_, _10858_, _10853_ }), .Y(_10852_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36080_ ( .A({ _10857_, _10856_, _10855_, _10854_ }), .Y(_10853_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36081_ ( .A({ _tmp_16[24], _tmp_16[21], _tmp_16[19:18] }), .Y(_10854_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36082_ ( .A({ _tmp_16[31], _tmp_16[29:28], _tmp_16[25] }), .Y(_10855_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36083_ ( .A({ _tmp_16[7:6], _tmp_16[4], _tmp_16[1] }), .Y(_10856_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36084_ ( .A({ _tmp_16[16], _tmp_16[13], _tmp_16[11:10] }), .Y(_10857_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36085_ ( .A({ _10859_, _tmp_16[30], _tmp_16[27:26] }), .Y(_10858_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36086_ ( .A({ _tmp_16[23:22], _tmp_16[20], _tmp_16[17] }), .Y(_10859_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36087_ ( .A({ _tmp_16[8], _tmp_16[5], _tmp_16[3:2] }), .Y(_10860_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36088_ ( .A({ _tmp_16[15:14], _tmp_16[12], _tmp_16[9] }), .Y(_10861_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36089_ ( .A({ _wvalid_11, _06200_ }), .Y(_06201_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36090_ ( .A({ _dataflow_slice_valid_12, _10862_ }), .Y(_06203_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36091_ ( .A({ _tmp_19, _10863_ }), .Y(_10862_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36092_ ( .A({ _10864_, _tmp_18[0], _tmp_18[33:32] }), .Y(_10863_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36093_ ( .A({ _10873_, _10872_, _10870_, _10865_ }), .Y(_10864_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36094_ ( .A({ _10869_, _10868_, _10867_, _10866_ }), .Y(_10865_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36095_ ( .A({ _tmp_18[24], _tmp_18[21], _tmp_18[19:18] }), .Y(_10866_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36096_ ( .A({ _tmp_18[31], _tmp_18[29:28], _tmp_18[25] }), .Y(_10867_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36097_ ( .A({ _tmp_18[7:6], _tmp_18[4], _tmp_18[1] }), .Y(_10868_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36098_ ( .A({ _tmp_18[16], _tmp_18[13], _tmp_18[11:10] }), .Y(_10869_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36099_ ( .A({ _10871_, _tmp_18[30], _tmp_18[27:26] }), .Y(_10870_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36100_ ( .A({ _tmp_18[23:22], _tmp_18[20], _tmp_18[17] }), .Y(_10871_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36101_ ( .A({ _tmp_18[8], _tmp_18[5], _tmp_18[3:2] }), .Y(_10872_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36102_ ( .A({ _tmp_18[15:14], _tmp_18[12], _tmp_18[9] }), .Y(_10873_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36103_ ( .A({ _wvalid_11, _06203_ }), .Y(_06204_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36104_ ( .A({ _dataflow_slice_valid_16, _10874_ }), .Y(_06206_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36105_ ( .A({ _tmp_26, _10875_ }), .Y(_10874_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36106_ ( .A({ _10876_, _tmp_25[0], _tmp_25[33:32] }), .Y(_10875_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36107_ ( .A({ _10885_, _10884_, _10882_, _10877_ }), .Y(_10876_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36108_ ( .A({ _10881_, _10880_, _10879_, _10878_ }), .Y(_10877_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36109_ ( .A({ _tmp_25[24], _tmp_25[21], _tmp_25[19:18] }), .Y(_10878_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36110_ ( .A({ _tmp_25[31], _tmp_25[29:28], _tmp_25[25] }), .Y(_10879_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36111_ ( .A({ _tmp_25[7:6], _tmp_25[4], _tmp_25[1] }), .Y(_10880_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36112_ ( .A({ _tmp_25[16], _tmp_25[13], _tmp_25[11:10] }), .Y(_10881_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36113_ ( .A({ _10883_, _tmp_25[30], _tmp_25[27:26] }), .Y(_10882_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36114_ ( .A({ _tmp_25[23:22], _tmp_25[20], _tmp_25[17] }), .Y(_10883_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36115_ ( .A({ _tmp_25[8], _tmp_25[5], _tmp_25[3:2] }), .Y(_10884_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36116_ ( .A({ _tmp_25[15:14], _tmp_25[12], _tmp_25[9] }), .Y(_10885_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36117_ ( .A({ _wvalid_24, _06206_ }), .Y(_06207_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36118_ ( .A({ _dataflow_slice_valid_19, _10886_ }), .Y(_06209_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36119_ ( .A({ _tmp_28, _10887_ }), .Y(_10886_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36120_ ( .A({ _10888_, _tmp_27[0], _tmp_27[33:32] }), .Y(_10887_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36121_ ( .A({ _10897_, _10896_, _10894_, _10889_ }), .Y(_10888_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36122_ ( .A({ _10893_, _10892_, _10891_, _10890_ }), .Y(_10889_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36123_ ( .A({ _tmp_27[24], _tmp_27[21], _tmp_27[19:18] }), .Y(_10890_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36124_ ( .A({ _tmp_27[31], _tmp_27[29:28], _tmp_27[25] }), .Y(_10891_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36125_ ( .A({ _tmp_27[7:6], _tmp_27[4], _tmp_27[1] }), .Y(_10892_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36126_ ( .A({ _tmp_27[16], _tmp_27[13], _tmp_27[11:10] }), .Y(_10893_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36127_ ( .A({ _10895_, _tmp_27[30], _tmp_27[27:26] }), .Y(_10894_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36128_ ( .A({ _tmp_27[23:22], _tmp_27[20], _tmp_27[17] }), .Y(_10895_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36129_ ( .A({ _tmp_27[8], _tmp_27[5], _tmp_27[3:2] }), .Y(_10896_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36130_ ( .A({ _tmp_27[15:14], _tmp_27[12], _tmp_27[9] }), .Y(_10897_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36131_ ( .A({ _wvalid_24, _06209_ }), .Y(_06210_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36132_ ( .A({ _dataflow_slice_valid_22, _10898_ }), .Y(_06212_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36133_ ( .A({ _tmp_30, _10899_ }), .Y(_10898_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36134_ ( .A({ _10900_, _tmp_29[0], _tmp_29[33:32] }), .Y(_10899_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36135_ ( .A({ _10909_, _10908_, _10906_, _10901_ }), .Y(_10900_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36136_ ( .A({ _10905_, _10904_, _10903_, _10902_ }), .Y(_10901_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36137_ ( .A({ _tmp_29[24], _tmp_29[21], _tmp_29[19:18] }), .Y(_10902_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36138_ ( .A({ _tmp_29[31], _tmp_29[29:28], _tmp_29[25] }), .Y(_10903_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36139_ ( .A({ _tmp_29[7:6], _tmp_29[4], _tmp_29[1] }), .Y(_10904_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36140_ ( .A({ _tmp_29[16], _tmp_29[13], _tmp_29[11:10] }), .Y(_10905_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36141_ ( .A({ _10907_, _tmp_29[30], _tmp_29[27:26] }), .Y(_10906_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36142_ ( .A({ _tmp_29[23:22], _tmp_29[20], _tmp_29[17] }), .Y(_10907_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36143_ ( .A({ _tmp_29[8], _tmp_29[5], _tmp_29[3:2] }), .Y(_10908_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36144_ ( .A({ _tmp_29[15:14], _tmp_29[12], _tmp_29[9] }), .Y(_10909_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36145_ ( .A({ _wvalid_24, _06212_ }), .Y(_06213_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36146_ ( .A({ _dataflow_slice_valid_25, _10910_ }), .Y(_06215_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36147_ ( .A({ _tmp_32, _10911_ }), .Y(_10910_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36148_ ( .A({ _10912_, _tmp_31[0], _tmp_31[33:32] }), .Y(_10911_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36149_ ( .A({ _10921_, _10920_, _10918_, _10913_ }), .Y(_10912_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36150_ ( .A({ _10917_, _10916_, _10915_, _10914_ }), .Y(_10913_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36151_ ( .A({ _tmp_31[24], _tmp_31[21], _tmp_31[19:18] }), .Y(_10914_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36152_ ( .A({ _tmp_31[31], _tmp_31[29:28], _tmp_31[25] }), .Y(_10915_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36153_ ( .A({ _tmp_31[7:6], _tmp_31[4], _tmp_31[1] }), .Y(_10916_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36154_ ( .A({ _tmp_31[16], _tmp_31[13], _tmp_31[11:10] }), .Y(_10917_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36155_ ( .A({ _10919_, _tmp_31[30], _tmp_31[27:26] }), .Y(_10918_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36156_ ( .A({ _tmp_31[23:22], _tmp_31[20], _tmp_31[17] }), .Y(_10919_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36157_ ( .A({ _tmp_31[8], _tmp_31[5], _tmp_31[3:2] }), .Y(_10920_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36158_ ( .A({ _tmp_31[15:14], _tmp_31[12], _tmp_31[9] }), .Y(_10921_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36159_ ( .A({ _wvalid_24, _06215_ }), .Y(_06216_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _36160_ ( .A({ _dataflow_slice_valid_29, _tmp_40, _10922_ }), .Y(_06218_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36161_ ( .A({ _10923_, _tmp_39[0], _tmp_39[33:32] }), .Y(_10922_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36162_ ( .A({ _10932_, _10931_, _10929_, _10924_ }), .Y(_10923_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36163_ ( .A({ _10928_, _10927_, _10926_, _10925_ }), .Y(_10924_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36164_ ( .A({ _tmp_39[24], _tmp_39[21], _tmp_39[19:18] }), .Y(_10925_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36165_ ( .A({ _tmp_39[31], _tmp_39[29:28], _tmp_39[25] }), .Y(_10926_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36166_ ( .A({ _tmp_39[7:6], _tmp_39[4], _tmp_39[1] }), .Y(_10927_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36167_ ( .A({ _tmp_39[16], _tmp_39[13], _tmp_39[11:10] }), .Y(_10928_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36168_ ( .A({ _10930_, _tmp_39[30], _tmp_39[27:26] }), .Y(_10929_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36169_ ( .A({ _tmp_39[23:22], _tmp_39[20], _tmp_39[17] }), .Y(_10930_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36170_ ( .A({ _tmp_39[8], _tmp_39[5], _tmp_39[3:2] }), .Y(_10931_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36171_ ( .A({ _tmp_39[15:14], _tmp_39[12], _tmp_39[9] }), .Y(_10932_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36172_ ( .A({ _wvalid_37, _06218_ }), .Y(_06219_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _36173_ ( .A({ _dataflow_slice_valid_32, _tmp_71, _10933_ }), .Y(_06221_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36174_ ( .A({ _10934_, _tmp_70[0], _tmp_70[33:32] }), .Y(_10933_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36175_ ( .A({ _10943_, _10942_, _10940_, _10935_ }), .Y(_10934_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36176_ ( .A({ _10939_, _10938_, _10937_, _10936_ }), .Y(_10935_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36177_ ( .A({ _tmp_70[24], _tmp_70[21], _tmp_70[19:18] }), .Y(_10936_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36178_ ( .A({ _tmp_70[31], _tmp_70[29:28], _tmp_70[25] }), .Y(_10937_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36179_ ( .A({ _tmp_70[7:6], _tmp_70[4], _tmp_70[1] }), .Y(_10938_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36180_ ( .A({ _tmp_70[16], _tmp_70[13], _tmp_70[11:10] }), .Y(_10939_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36181_ ( .A({ _10941_, _tmp_70[30], _tmp_70[27:26] }), .Y(_10940_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36182_ ( .A({ _tmp_70[23:22], _tmp_70[20], _tmp_70[17] }), .Y(_10941_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36183_ ( .A({ _tmp_70[8], _tmp_70[5], _tmp_70[3:2] }), .Y(_10942_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36184_ ( .A({ _tmp_70[15:14], _tmp_70[12], _tmp_70[9] }), .Y(_10943_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36185_ ( .A({ _wvalid_37, _06221_ }), .Y(_06222_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _36186_ ( .A({ _dataflow_slice_valid_35, _tmp_102, _10944_ }), .Y(_06224_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36187_ ( .A({ _10945_, _tmp_101[0], _tmp_101[33:32] }), .Y(_10944_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36188_ ( .A({ _10954_, _10953_, _10951_, _10946_ }), .Y(_10945_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36189_ ( .A({ _10950_, _10949_, _10948_, _10947_ }), .Y(_10946_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36190_ ( .A({ _tmp_101[24], _tmp_101[21], _tmp_101[19:18] }), .Y(_10947_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36191_ ( .A({ _tmp_101[31], _tmp_101[29:28], _tmp_101[25] }), .Y(_10948_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36192_ ( .A({ _tmp_101[7:6], _tmp_101[4], _tmp_101[1] }), .Y(_10949_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36193_ ( .A({ _tmp_101[16], _tmp_101[13], _tmp_101[11:10] }), .Y(_10950_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36194_ ( .A({ _10952_, _tmp_101[30], _tmp_101[27:26] }), .Y(_10951_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36195_ ( .A({ _tmp_101[23:22], _tmp_101[20], _tmp_101[17] }), .Y(_10952_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36196_ ( .A({ _tmp_101[8], _tmp_101[5], _tmp_101[3:2] }), .Y(_10953_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36197_ ( .A({ _tmp_101[15:14], _tmp_101[12], _tmp_101[9] }), .Y(_10954_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36198_ ( .A({ _wvalid_37, _06224_ }), .Y(_06225_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _36199_ ( .A({ _dataflow_slice_valid_38, _tmp_133, _10955_ }), .Y(_06227_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36200_ ( .A({ _10956_, _tmp_132[0], _tmp_132[33:32] }), .Y(_10955_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36201_ ( .A({ _10965_, _10964_, _10962_, _10957_ }), .Y(_10956_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36202_ ( .A({ _10961_, _10960_, _10959_, _10958_ }), .Y(_10957_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36203_ ( .A({ _tmp_132[24], _tmp_132[21], _tmp_132[19:18] }), .Y(_10958_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36204_ ( .A({ _tmp_132[31], _tmp_132[29:28], _tmp_132[25] }), .Y(_10959_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36205_ ( .A({ _tmp_132[7:6], _tmp_132[4], _tmp_132[1] }), .Y(_10960_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36206_ ( .A({ _tmp_132[16], _tmp_132[13], _tmp_132[11:10] }), .Y(_10961_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36207_ ( .A({ _10963_, _tmp_132[30], _tmp_132[27:26] }), .Y(_10962_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36208_ ( .A({ _tmp_132[23:22], _tmp_132[20], _tmp_132[17] }), .Y(_10963_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36209_ ( .A({ _tmp_132[8], _tmp_132[5], _tmp_132[3:2] }), .Y(_10964_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36210_ ( .A({ _tmp_132[15:14], _tmp_132[12], _tmp_132[9] }), .Y(_10965_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36211_ ( .A({ _wvalid_37, _06227_ }), .Y(_06228_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _36212_ ( .A({ _dataflow_slice_valid_41, _tmp_164, _10966_ }), .Y(_06230_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36213_ ( .A({ _10967_, _tmp_163[0], _tmp_163[33:32] }), .Y(_10966_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36214_ ( .A({ _10976_, _10975_, _10973_, _10968_ }), .Y(_10967_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36215_ ( .A({ _10972_, _10971_, _10970_, _10969_ }), .Y(_10968_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36216_ ( .A({ _tmp_163[24], _tmp_163[21], _tmp_163[19:18] }), .Y(_10969_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36217_ ( .A({ _tmp_163[31], _tmp_163[29:28], _tmp_163[25] }), .Y(_10970_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36218_ ( .A({ _tmp_163[7:6], _tmp_163[4], _tmp_163[1] }), .Y(_10971_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36219_ ( .A({ _tmp_163[16], _tmp_163[13], _tmp_163[11:10] }), .Y(_10972_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36220_ ( .A({ _10974_, _tmp_163[30], _tmp_163[27:26] }), .Y(_10973_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36221_ ( .A({ _tmp_163[23:22], _tmp_163[20], _tmp_163[17] }), .Y(_10974_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36222_ ( .A({ _tmp_163[8], _tmp_163[5], _tmp_163[3:2] }), .Y(_10975_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36223_ ( .A({ _tmp_163[15:14], _tmp_163[12], _tmp_163[9] }), .Y(_10976_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36224_ ( .A({ _wvalid_37, _06230_ }), .Y(_06231_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _36225_ ( .A({ _dataflow_slice_valid_44, _tmp_195, _10977_ }), .Y(_06233_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36226_ ( .A({ _10978_, _tmp_194[0], _tmp_194[33:32] }), .Y(_10977_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36227_ ( .A({ _10987_, _10986_, _10984_, _10979_ }), .Y(_10978_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36228_ ( .A({ _10983_, _10982_, _10981_, _10980_ }), .Y(_10979_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36229_ ( .A({ _tmp_194[24], _tmp_194[21], _tmp_194[19:18] }), .Y(_10980_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36230_ ( .A({ _tmp_194[31], _tmp_194[29:28], _tmp_194[25] }), .Y(_10981_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36231_ ( .A({ _tmp_194[7:6], _tmp_194[4], _tmp_194[1] }), .Y(_10982_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36232_ ( .A({ _tmp_194[16], _tmp_194[13], _tmp_194[11:10] }), .Y(_10983_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36233_ ( .A({ _10985_, _tmp_194[30], _tmp_194[27:26] }), .Y(_10984_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36234_ ( .A({ _tmp_194[23:22], _tmp_194[20], _tmp_194[17] }), .Y(_10985_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36235_ ( .A({ _tmp_194[8], _tmp_194[5], _tmp_194[3:2] }), .Y(_10986_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36236_ ( .A({ _tmp_194[15:14], _tmp_194[12], _tmp_194[9] }), .Y(_10987_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36237_ ( .A({ _wvalid_37, _06233_ }), .Y(_06234_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _36238_ ( .A({ _dataflow_slice_valid_47, _tmp_226, _10988_ }), .Y(_06236_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36239_ ( .A({ _10989_, _tmp_225[0], _tmp_225[33:32] }), .Y(_10988_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36240_ ( .A({ _10998_, _10997_, _10995_, _10990_ }), .Y(_10989_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36241_ ( .A({ _10994_, _10993_, _10992_, _10991_ }), .Y(_10990_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36242_ ( .A({ _tmp_225[24], _tmp_225[21], _tmp_225[19:18] }), .Y(_10991_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36243_ ( .A({ _tmp_225[31], _tmp_225[29:28], _tmp_225[25] }), .Y(_10992_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36244_ ( .A({ _tmp_225[7:6], _tmp_225[4], _tmp_225[1] }), .Y(_10993_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36245_ ( .A({ _tmp_225[16], _tmp_225[13], _tmp_225[11:10] }), .Y(_10994_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36246_ ( .A({ _10996_, _tmp_225[30], _tmp_225[27:26] }), .Y(_10995_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36247_ ( .A({ _tmp_225[23:22], _tmp_225[20], _tmp_225[17] }), .Y(_10996_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36248_ ( .A({ _tmp_225[8], _tmp_225[5], _tmp_225[3:2] }), .Y(_10997_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36249_ ( .A({ _tmp_225[15:14], _tmp_225[12], _tmp_225[9] }), .Y(_10998_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36250_ ( .A({ _wvalid_37, _06236_ }), .Y(_06237_) );
  \$lut  #( .LUT(8'h1f), .WIDTH(3) ) _36251_ ( .A({ _dataflow_slice_valid_50, _tmp_257, _10999_ }), .Y(_06239_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36252_ ( .A({ _11000_, _tmp_256[0], _tmp_256[33:32] }), .Y(_10999_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36253_ ( .A({ _11009_, _11008_, _11006_, _11001_ }), .Y(_11000_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36254_ ( .A({ _11005_, _11004_, _11003_, _11002_ }), .Y(_11001_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36255_ ( .A({ _tmp_256[24], _tmp_256[21], _tmp_256[19:18] }), .Y(_11002_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36256_ ( .A({ _tmp_256[31], _tmp_256[29:28], _tmp_256[25] }), .Y(_11003_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36257_ ( .A({ _tmp_256[7:6], _tmp_256[4], _tmp_256[1] }), .Y(_11004_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36258_ ( .A({ _tmp_256[16], _tmp_256[13], _tmp_256[11:10] }), .Y(_11005_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36259_ ( .A({ _11007_, _tmp_256[30], _tmp_256[27:26] }), .Y(_11006_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36260_ ( .A({ _tmp_256[23:22], _tmp_256[20], _tmp_256[17] }), .Y(_11007_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36261_ ( .A({ _tmp_256[8], _tmp_256[5], _tmp_256[3:2] }), .Y(_11008_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36262_ ( .A({ _tmp_256[15:14], _tmp_256[12], _tmp_256[9] }), .Y(_11009_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36263_ ( .A({ _wvalid_37, _06239_ }), .Y(_06240_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36264_ ( .A({ _dataflow_slice_valid_54, _11010_ }), .Y(_06242_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36265_ ( .A({ _tmp_293, _11011_ }), .Y(_11010_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36266_ ( .A({ _11012_, _tmp_292[0], _tmp_292[33:32] }), .Y(_11011_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36267_ ( .A({ _11021_, _11020_, _11018_, _11013_ }), .Y(_11012_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36268_ ( .A({ _11017_, _11016_, _11015_, _11014_ }), .Y(_11013_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36269_ ( .A({ _tmp_292[24], _tmp_292[21], _tmp_292[19:18] }), .Y(_11014_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36270_ ( .A({ _tmp_292[31], _tmp_292[29:28], _tmp_292[25] }), .Y(_11015_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36271_ ( .A({ _tmp_292[7:6], _tmp_292[4], _tmp_292[1] }), .Y(_11016_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36272_ ( .A({ _tmp_292[16], _tmp_292[13], _tmp_292[11:10] }), .Y(_11017_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36273_ ( .A({ _11019_, _tmp_292[30], _tmp_292[27:26] }), .Y(_11018_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36274_ ( .A({ _tmp_292[23:22], _tmp_292[20], _tmp_292[17] }), .Y(_11019_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36275_ ( .A({ _tmp_292[8], _tmp_292[5], _tmp_292[3:2] }), .Y(_11020_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36276_ ( .A({ _tmp_292[15:14], _tmp_292[12], _tmp_292[9] }), .Y(_11021_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36277_ ( .A({ _wvalid_290, _06242_ }), .Y(_06243_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36278_ ( .A({ _dataflow_slice_valid_57, _11022_ }), .Y(_06245_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36279_ ( .A({ _tmp_306, _11023_ }), .Y(_11022_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36280_ ( .A({ _11024_, _tmp_305[0], _tmp_305[33:32] }), .Y(_11023_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36281_ ( .A({ _11033_, _11032_, _11030_, _11025_ }), .Y(_11024_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36282_ ( .A({ _11029_, _11028_, _11027_, _11026_ }), .Y(_11025_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36283_ ( .A({ _tmp_305[24], _tmp_305[21], _tmp_305[19:18] }), .Y(_11026_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36284_ ( .A({ _tmp_305[31], _tmp_305[29:28], _tmp_305[25] }), .Y(_11027_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36285_ ( .A({ _tmp_305[7:6], _tmp_305[4], _tmp_305[1] }), .Y(_11028_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36286_ ( .A({ _tmp_305[16], _tmp_305[13], _tmp_305[11:10] }), .Y(_11029_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36287_ ( .A({ _11031_, _tmp_305[30], _tmp_305[27:26] }), .Y(_11030_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36288_ ( .A({ _tmp_305[23:22], _tmp_305[20], _tmp_305[17] }), .Y(_11031_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36289_ ( .A({ _tmp_305[8], _tmp_305[5], _tmp_305[3:2] }), .Y(_11032_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36290_ ( .A({ _tmp_305[15:14], _tmp_305[12], _tmp_305[9] }), .Y(_11033_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36291_ ( .A({ _wvalid_290, _06245_ }), .Y(_06246_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36292_ ( .A({ _dataflow_slice_valid_60, _11034_ }), .Y(_06248_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36293_ ( .A({ _tmp_319, _11035_ }), .Y(_11034_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36294_ ( .A({ _11036_, _tmp_318[0], _tmp_318[33:32] }), .Y(_11035_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36295_ ( .A({ _11045_, _11044_, _11042_, _11037_ }), .Y(_11036_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36296_ ( .A({ _11041_, _11040_, _11039_, _11038_ }), .Y(_11037_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36297_ ( .A({ _tmp_318[24], _tmp_318[21], _tmp_318[19:18] }), .Y(_11038_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36298_ ( .A({ _tmp_318[31], _tmp_318[29:28], _tmp_318[25] }), .Y(_11039_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36299_ ( .A({ _tmp_318[7:6], _tmp_318[4], _tmp_318[1] }), .Y(_11040_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36300_ ( .A({ _tmp_318[16], _tmp_318[13], _tmp_318[11:10] }), .Y(_11041_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36301_ ( .A({ _11043_, _tmp_318[30], _tmp_318[27:26] }), .Y(_11042_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36302_ ( .A({ _tmp_318[23:22], _tmp_318[20], _tmp_318[17] }), .Y(_11043_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36303_ ( .A({ _tmp_318[8], _tmp_318[5], _tmp_318[3:2] }), .Y(_11044_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36304_ ( .A({ _tmp_318[15:14], _tmp_318[12], _tmp_318[9] }), .Y(_11045_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36305_ ( .A({ _wvalid_290, _06248_ }), .Y(_06249_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36306_ ( .A({ _dataflow_slice_valid_63, _11046_ }), .Y(_06251_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36307_ ( .A({ _tmp_332, _11047_ }), .Y(_11046_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36308_ ( .A({ _11048_, _tmp_331[0], _tmp_331[33:32] }), .Y(_11047_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36309_ ( .A({ _11057_, _11056_, _11054_, _11049_ }), .Y(_11048_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36310_ ( .A({ _11053_, _11052_, _11051_, _11050_ }), .Y(_11049_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36311_ ( .A({ _tmp_331[24], _tmp_331[21], _tmp_331[19:18] }), .Y(_11050_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36312_ ( .A({ _tmp_331[31], _tmp_331[29:28], _tmp_331[25] }), .Y(_11051_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36313_ ( .A({ _tmp_331[7:6], _tmp_331[4], _tmp_331[1] }), .Y(_11052_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36314_ ( .A({ _tmp_331[16], _tmp_331[13], _tmp_331[11:10] }), .Y(_11053_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36315_ ( .A({ _11055_, _tmp_331[30], _tmp_331[27:26] }), .Y(_11054_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36316_ ( .A({ _tmp_331[23:22], _tmp_331[20], _tmp_331[17] }), .Y(_11055_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36317_ ( .A({ _tmp_331[8], _tmp_331[5], _tmp_331[3:2] }), .Y(_11056_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36318_ ( .A({ _tmp_331[15:14], _tmp_331[12], _tmp_331[9] }), .Y(_11057_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36319_ ( .A({ _wvalid_290, _06251_ }), .Y(_06252_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36320_ ( .A({ _dataflow_slice_valid_67, _11058_ }), .Y(_06254_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36321_ ( .A({ _tmp_350, _11059_ }), .Y(_11058_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36322_ ( .A({ _11060_, _tmp_349[0], _tmp_349[33:32] }), .Y(_11059_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36323_ ( .A({ _11069_, _11068_, _11066_, _11061_ }), .Y(_11060_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36324_ ( .A({ _11065_, _11064_, _11063_, _11062_ }), .Y(_11061_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36325_ ( .A({ _tmp_349[24], _tmp_349[21], _tmp_349[19:18] }), .Y(_11062_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36326_ ( .A({ _tmp_349[31], _tmp_349[29:28], _tmp_349[25] }), .Y(_11063_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36327_ ( .A({ _tmp_349[7:6], _tmp_349[4], _tmp_349[1] }), .Y(_11064_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36328_ ( .A({ _tmp_349[16], _tmp_349[13], _tmp_349[11:10] }), .Y(_11065_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36329_ ( .A({ _11067_, _tmp_349[30], _tmp_349[27:26] }), .Y(_11066_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36330_ ( .A({ _tmp_349[23:22], _tmp_349[20], _tmp_349[17] }), .Y(_11067_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36331_ ( .A({ _tmp_349[8], _tmp_349[5], _tmp_349[3:2] }), .Y(_11068_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36332_ ( .A({ _tmp_349[15:14], _tmp_349[12], _tmp_349[9] }), .Y(_11069_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36333_ ( .A({ _wvalid_347, _06254_ }), .Y(_06255_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36334_ ( .A({ _dataflow_slice_valid_70, _11070_ }), .Y(_06257_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36335_ ( .A({ _tmp_363, _11071_ }), .Y(_11070_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36336_ ( .A({ _11072_, _tmp_362[0], _tmp_362[33:32] }), .Y(_11071_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36337_ ( .A({ _11081_, _11080_, _11078_, _11073_ }), .Y(_11072_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36338_ ( .A({ _11077_, _11076_, _11075_, _11074_ }), .Y(_11073_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36339_ ( .A({ _tmp_362[24], _tmp_362[21], _tmp_362[19:18] }), .Y(_11074_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36340_ ( .A({ _tmp_362[31], _tmp_362[29:28], _tmp_362[25] }), .Y(_11075_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36341_ ( .A({ _tmp_362[7:6], _tmp_362[4], _tmp_362[1] }), .Y(_11076_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36342_ ( .A({ _tmp_362[16], _tmp_362[13], _tmp_362[11:10] }), .Y(_11077_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36343_ ( .A({ _11079_, _tmp_362[30], _tmp_362[27:26] }), .Y(_11078_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36344_ ( .A({ _tmp_362[23:22], _tmp_362[20], _tmp_362[17] }), .Y(_11079_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36345_ ( .A({ _tmp_362[8], _tmp_362[5], _tmp_362[3:2] }), .Y(_11080_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36346_ ( .A({ _tmp_362[15:14], _tmp_362[12], _tmp_362[9] }), .Y(_11081_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36347_ ( .A({ _wvalid_347, _06257_ }), .Y(_06258_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36348_ ( .A({ _dataflow_slice_valid_73, _11082_ }), .Y(_06260_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36349_ ( .A({ _tmp_376, _11083_ }), .Y(_11082_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36350_ ( .A({ _11084_, _tmp_375[0], _tmp_375[33:32] }), .Y(_11083_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36351_ ( .A({ _11093_, _11092_, _11090_, _11085_ }), .Y(_11084_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36352_ ( .A({ _11089_, _11088_, _11087_, _11086_ }), .Y(_11085_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36353_ ( .A({ _tmp_375[24], _tmp_375[21], _tmp_375[19:18] }), .Y(_11086_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36354_ ( .A({ _tmp_375[31], _tmp_375[29:28], _tmp_375[25] }), .Y(_11087_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36355_ ( .A({ _tmp_375[7:6], _tmp_375[4], _tmp_375[1] }), .Y(_11088_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36356_ ( .A({ _tmp_375[16], _tmp_375[13], _tmp_375[11:10] }), .Y(_11089_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36357_ ( .A({ _11091_, _tmp_375[30], _tmp_375[27:26] }), .Y(_11090_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36358_ ( .A({ _tmp_375[23:22], _tmp_375[20], _tmp_375[17] }), .Y(_11091_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36359_ ( .A({ _tmp_375[8], _tmp_375[5], _tmp_375[3:2] }), .Y(_11092_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36360_ ( .A({ _tmp_375[15:14], _tmp_375[12], _tmp_375[9] }), .Y(_11093_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36361_ ( .A({ _wvalid_347, _06260_ }), .Y(_06261_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36362_ ( .A({ _dataflow_slice_valid_76, _11094_ }), .Y(_06263_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36363_ ( .A({ _tmp_389, _11095_ }), .Y(_11094_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36364_ ( .A({ _11096_, _tmp_388[0], _tmp_388[33:32] }), .Y(_11095_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36365_ ( .A({ _11105_, _11104_, _11102_, _11097_ }), .Y(_11096_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36366_ ( .A({ _11101_, _11100_, _11099_, _11098_ }), .Y(_11097_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36367_ ( .A({ _tmp_388[24], _tmp_388[21], _tmp_388[19:18] }), .Y(_11098_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36368_ ( .A({ _tmp_388[31], _tmp_388[29:28], _tmp_388[25] }), .Y(_11099_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36369_ ( .A({ _tmp_388[7:6], _tmp_388[4], _tmp_388[1] }), .Y(_11100_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36370_ ( .A({ _tmp_388[16], _tmp_388[13], _tmp_388[11:10] }), .Y(_11101_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36371_ ( .A({ _11103_, _tmp_388[30], _tmp_388[27:26] }), .Y(_11102_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36372_ ( .A({ _tmp_388[23:22], _tmp_388[20], _tmp_388[17] }), .Y(_11103_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36373_ ( .A({ _tmp_388[8], _tmp_388[5], _tmp_388[3:2] }), .Y(_11104_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36374_ ( .A({ _tmp_388[15:14], _tmp_388[12], _tmp_388[9] }), .Y(_11105_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36375_ ( .A({ _wvalid_347, _06263_ }), .Y(_06264_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36376_ ( .A({ _dataflow_slice_valid_80, _11106_ }), .Y(_06266_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36377_ ( .A({ _tmp_407, _11107_ }), .Y(_11106_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36378_ ( .A({ _11108_, _tmp_406[0], _tmp_406[33:32] }), .Y(_11107_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36379_ ( .A({ _11117_, _11116_, _11114_, _11109_ }), .Y(_11108_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36380_ ( .A({ _11113_, _11112_, _11111_, _11110_ }), .Y(_11109_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36381_ ( .A({ _tmp_406[24], _tmp_406[21], _tmp_406[19:18] }), .Y(_11110_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36382_ ( .A({ _tmp_406[31], _tmp_406[29:28], _tmp_406[25] }), .Y(_11111_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36383_ ( .A({ _tmp_406[7:6], _tmp_406[4], _tmp_406[1] }), .Y(_11112_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36384_ ( .A({ _tmp_406[16], _tmp_406[13], _tmp_406[11:10] }), .Y(_11113_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36385_ ( .A({ _11115_, _tmp_406[30], _tmp_406[27:26] }), .Y(_11114_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36386_ ( .A({ _tmp_406[23:22], _tmp_406[20], _tmp_406[17] }), .Y(_11115_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36387_ ( .A({ _tmp_406[8], _tmp_406[5], _tmp_406[3:2] }), .Y(_11116_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36388_ ( .A({ _tmp_406[15:14], _tmp_406[12], _tmp_406[9] }), .Y(_11117_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36389_ ( .A({ _wvalid_404, _06266_ }), .Y(_06267_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36390_ ( .A({ _dataflow_slice_valid_83, _11118_ }), .Y(_06269_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36391_ ( .A({ _tmp_420, _11119_ }), .Y(_11118_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36392_ ( .A({ _11120_, _tmp_419[0], _tmp_419[33:32] }), .Y(_11119_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36393_ ( .A({ _11129_, _11128_, _11126_, _11121_ }), .Y(_11120_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36394_ ( .A({ _11125_, _11124_, _11123_, _11122_ }), .Y(_11121_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36395_ ( .A({ _tmp_419[24], _tmp_419[21], _tmp_419[19:18] }), .Y(_11122_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36396_ ( .A({ _tmp_419[31], _tmp_419[29:28], _tmp_419[25] }), .Y(_11123_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36397_ ( .A({ _tmp_419[7:6], _tmp_419[4], _tmp_419[1] }), .Y(_11124_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36398_ ( .A({ _tmp_419[16], _tmp_419[13], _tmp_419[11:10] }), .Y(_11125_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36399_ ( .A({ _11127_, _tmp_419[30], _tmp_419[27:26] }), .Y(_11126_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36400_ ( .A({ _tmp_419[23:22], _tmp_419[20], _tmp_419[17] }), .Y(_11127_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36401_ ( .A({ _tmp_419[8], _tmp_419[5], _tmp_419[3:2] }), .Y(_11128_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36402_ ( .A({ _tmp_419[15:14], _tmp_419[12], _tmp_419[9] }), .Y(_11129_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36403_ ( .A({ _wvalid_404, _06269_ }), .Y(_06270_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36404_ ( .A({ _dataflow_slice_valid_86, _11130_ }), .Y(_06272_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36405_ ( .A({ _tmp_433, _11131_ }), .Y(_11130_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36406_ ( .A({ _11132_, _tmp_432[0], _tmp_432[33:32] }), .Y(_11131_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36407_ ( .A({ _11141_, _11140_, _11138_, _11133_ }), .Y(_11132_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36408_ ( .A({ _11137_, _11136_, _11135_, _11134_ }), .Y(_11133_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36409_ ( .A({ _tmp_432[24], _tmp_432[21], _tmp_432[19:18] }), .Y(_11134_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36410_ ( .A({ _tmp_432[31], _tmp_432[29:28], _tmp_432[25] }), .Y(_11135_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36411_ ( .A({ _tmp_432[7:6], _tmp_432[4], _tmp_432[1] }), .Y(_11136_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36412_ ( .A({ _tmp_432[16], _tmp_432[13], _tmp_432[11:10] }), .Y(_11137_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36413_ ( .A({ _11139_, _tmp_432[30], _tmp_432[27:26] }), .Y(_11138_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36414_ ( .A({ _tmp_432[23:22], _tmp_432[20], _tmp_432[17] }), .Y(_11139_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36415_ ( .A({ _tmp_432[8], _tmp_432[5], _tmp_432[3:2] }), .Y(_11140_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36416_ ( .A({ _tmp_432[15:14], _tmp_432[12], _tmp_432[9] }), .Y(_11141_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36417_ ( .A({ _wvalid_404, _06272_ }), .Y(_06273_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36418_ ( .A({ _dataflow_slice_valid_89, _11142_ }), .Y(_06275_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36419_ ( .A({ _tmp_446, _11143_ }), .Y(_11142_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36420_ ( .A({ _11144_, _tmp_445[0], _tmp_445[33:32] }), .Y(_11143_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36421_ ( .A({ _11153_, _11152_, _11150_, _11145_ }), .Y(_11144_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36422_ ( .A({ _11149_, _11148_, _11147_, _11146_ }), .Y(_11145_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36423_ ( .A({ _tmp_445[24], _tmp_445[21], _tmp_445[19:18] }), .Y(_11146_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36424_ ( .A({ _tmp_445[31], _tmp_445[29:28], _tmp_445[25] }), .Y(_11147_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36425_ ( .A({ _tmp_445[7:6], _tmp_445[4], _tmp_445[1] }), .Y(_11148_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36426_ ( .A({ _tmp_445[16], _tmp_445[13], _tmp_445[11:10] }), .Y(_11149_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36427_ ( .A({ _11151_, _tmp_445[30], _tmp_445[27:26] }), .Y(_11150_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36428_ ( .A({ _tmp_445[23:22], _tmp_445[20], _tmp_445[17] }), .Y(_11151_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36429_ ( .A({ _tmp_445[8], _tmp_445[5], _tmp_445[3:2] }), .Y(_11152_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36430_ ( .A({ _tmp_445[15:14], _tmp_445[12], _tmp_445[9] }), .Y(_11153_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36431_ ( .A({ _wvalid_404, _06275_ }), .Y(_06276_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36432_ ( .A({ _dataflow_slice_valid_111, _11154_ }), .Y(_06278_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36433_ ( .A({ _tmp_1125, _11155_ }), .Y(_11154_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36434_ ( .A({ _11156_, _tmp_1124[0], _tmp_1124[33:32] }), .Y(_11155_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36435_ ( .A({ _11165_, _11164_, _11162_, _11157_ }), .Y(_11156_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36436_ ( .A({ _11161_, _11160_, _11159_, _11158_ }), .Y(_11157_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36437_ ( .A({ _tmp_1124[24], _tmp_1124[21], _tmp_1124[19:18] }), .Y(_11158_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36438_ ( .A({ _tmp_1124[31], _tmp_1124[29:28], _tmp_1124[25] }), .Y(_11159_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36439_ ( .A({ _tmp_1124[7:6], _tmp_1124[4], _tmp_1124[1] }), .Y(_11160_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36440_ ( .A({ _tmp_1124[16], _tmp_1124[13], _tmp_1124[11:10] }), .Y(_11161_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36441_ ( .A({ _11163_, _tmp_1124[30], _tmp_1124[27:26] }), .Y(_11162_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36442_ ( .A({ _tmp_1124[23:22], _tmp_1124[20], _tmp_1124[17] }), .Y(_11163_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36443_ ( .A({ _tmp_1124[8], _tmp_1124[5], _tmp_1124[3:2] }), .Y(_11164_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36444_ ( .A({ _tmp_1124[15:14], _tmp_1124[12], _tmp_1124[9] }), .Y(_11165_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36445_ ( .A({ _wvalid_1123, _06278_ }), .Y(_06279_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36446_ ( .A({ _dataflow_slice_valid_114, _11166_ }), .Y(_06281_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36447_ ( .A({ _tmp_1127, _11167_ }), .Y(_11166_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36448_ ( .A({ _11168_, _tmp_1126[0], _tmp_1126[33:32] }), .Y(_11167_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36449_ ( .A({ _11177_, _11176_, _11174_, _11169_ }), .Y(_11168_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36450_ ( .A({ _11173_, _11172_, _11171_, _11170_ }), .Y(_11169_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36451_ ( .A({ _tmp_1126[24], _tmp_1126[21], _tmp_1126[19:18] }), .Y(_11170_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36452_ ( .A({ _tmp_1126[31], _tmp_1126[29:28], _tmp_1126[25] }), .Y(_11171_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36453_ ( .A({ _tmp_1126[7:6], _tmp_1126[4], _tmp_1126[1] }), .Y(_11172_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36454_ ( .A({ _tmp_1126[16], _tmp_1126[13], _tmp_1126[11:10] }), .Y(_11173_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36455_ ( .A({ _11175_, _tmp_1126[30], _tmp_1126[27:26] }), .Y(_11174_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36456_ ( .A({ _tmp_1126[23:22], _tmp_1126[20], _tmp_1126[17] }), .Y(_11175_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36457_ ( .A({ _tmp_1126[8], _tmp_1126[5], _tmp_1126[3:2] }), .Y(_11176_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36458_ ( .A({ _tmp_1126[15:14], _tmp_1126[12], _tmp_1126[9] }), .Y(_11177_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36459_ ( .A({ _wvalid_1123, _06281_ }), .Y(_06282_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36460_ ( .A({ _dataflow_slice_valid_117, _11178_ }), .Y(_06284_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36461_ ( .A({ _tmp_1129, _11179_ }), .Y(_11178_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36462_ ( .A({ _11180_, _tmp_1128[0], _tmp_1128[33:32] }), .Y(_11179_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36463_ ( .A({ _11189_, _11188_, _11186_, _11181_ }), .Y(_11180_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36464_ ( .A({ _11185_, _11184_, _11183_, _11182_ }), .Y(_11181_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36465_ ( .A({ _tmp_1128[24], _tmp_1128[21], _tmp_1128[19:18] }), .Y(_11182_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36466_ ( .A({ _tmp_1128[31], _tmp_1128[29:28], _tmp_1128[25] }), .Y(_11183_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36467_ ( .A({ _tmp_1128[7:6], _tmp_1128[4], _tmp_1128[1] }), .Y(_11184_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36468_ ( .A({ _tmp_1128[16], _tmp_1128[13], _tmp_1128[11:10] }), .Y(_11185_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36469_ ( .A({ _11187_, _tmp_1128[30], _tmp_1128[27:26] }), .Y(_11186_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36470_ ( .A({ _tmp_1128[23:22], _tmp_1128[20], _tmp_1128[17] }), .Y(_11187_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36471_ ( .A({ _tmp_1128[8], _tmp_1128[5], _tmp_1128[3:2] }), .Y(_11188_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36472_ ( .A({ _tmp_1128[15:14], _tmp_1128[12], _tmp_1128[9] }), .Y(_11189_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36473_ ( .A({ _wvalid_1123, _06284_ }), .Y(_06285_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36474_ ( .A({ _dataflow_slice_valid_120, _11190_ }), .Y(_06287_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36475_ ( .A({ _tmp_1131, _11191_ }), .Y(_11190_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36476_ ( .A({ _11192_, _tmp_1130[0], _tmp_1130[33:32] }), .Y(_11191_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36477_ ( .A({ _11201_, _11200_, _11198_, _11193_ }), .Y(_11192_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36478_ ( .A({ _11197_, _11196_, _11195_, _11194_ }), .Y(_11193_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36479_ ( .A({ _tmp_1130[24], _tmp_1130[21], _tmp_1130[19:18] }), .Y(_11194_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36480_ ( .A({ _tmp_1130[31], _tmp_1130[29:28], _tmp_1130[25] }), .Y(_11195_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36481_ ( .A({ _tmp_1130[7:6], _tmp_1130[4], _tmp_1130[1] }), .Y(_11196_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36482_ ( .A({ _tmp_1130[16], _tmp_1130[13], _tmp_1130[11:10] }), .Y(_11197_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36483_ ( .A({ _11199_, _tmp_1130[30], _tmp_1130[27:26] }), .Y(_11198_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36484_ ( .A({ _tmp_1130[23:22], _tmp_1130[20], _tmp_1130[17] }), .Y(_11199_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36485_ ( .A({ _tmp_1130[8], _tmp_1130[5], _tmp_1130[3:2] }), .Y(_11200_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36486_ ( .A({ _tmp_1130[15:14], _tmp_1130[12], _tmp_1130[9] }), .Y(_11201_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36487_ ( .A({ _wvalid_1123, _06287_ }), .Y(_06288_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36488_ ( .A({ _dataflow_slice_valid_124, _11202_ }), .Y(_06290_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36489_ ( .A({ _tmp_1137, _11203_ }), .Y(_11202_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36490_ ( .A({ _11204_, _tmp_1136[0], _tmp_1136[33:32] }), .Y(_11203_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36491_ ( .A({ _11213_, _11212_, _11210_, _11205_ }), .Y(_11204_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36492_ ( .A({ _11209_, _11208_, _11207_, _11206_ }), .Y(_11205_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36493_ ( .A({ _tmp_1136[24], _tmp_1136[21], _tmp_1136[19:18] }), .Y(_11206_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36494_ ( .A({ _tmp_1136[31], _tmp_1136[29:28], _tmp_1136[25] }), .Y(_11207_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36495_ ( .A({ _tmp_1136[7:6], _tmp_1136[4], _tmp_1136[1] }), .Y(_11208_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36496_ ( .A({ _tmp_1136[16], _tmp_1136[13], _tmp_1136[11:10] }), .Y(_11209_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36497_ ( .A({ _11211_, _tmp_1136[30], _tmp_1136[27:26] }), .Y(_11210_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36498_ ( .A({ _tmp_1136[23:22], _tmp_1136[20], _tmp_1136[17] }), .Y(_11211_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36499_ ( .A({ _tmp_1136[8], _tmp_1136[5], _tmp_1136[3:2] }), .Y(_11212_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36500_ ( .A({ _tmp_1136[15:14], _tmp_1136[12], _tmp_1136[9] }), .Y(_11213_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36501_ ( .A({ _wvalid_1135, _06290_ }), .Y(_06291_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36502_ ( .A({ _dataflow_slice_valid_127, _11214_ }), .Y(_06293_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36503_ ( .A({ _tmp_1139, _11215_ }), .Y(_11214_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36504_ ( .A({ _11216_, _tmp_1138[0], _tmp_1138[33:32] }), .Y(_11215_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36505_ ( .A({ _11225_, _11224_, _11222_, _11217_ }), .Y(_11216_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36506_ ( .A({ _11221_, _11220_, _11219_, _11218_ }), .Y(_11217_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36507_ ( .A({ _tmp_1138[24], _tmp_1138[21], _tmp_1138[19:18] }), .Y(_11218_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36508_ ( .A({ _tmp_1138[31], _tmp_1138[29:28], _tmp_1138[25] }), .Y(_11219_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36509_ ( .A({ _tmp_1138[7:6], _tmp_1138[4], _tmp_1138[1] }), .Y(_11220_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36510_ ( .A({ _tmp_1138[16], _tmp_1138[13], _tmp_1138[11:10] }), .Y(_11221_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36511_ ( .A({ _11223_, _tmp_1138[30], _tmp_1138[27:26] }), .Y(_11222_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36512_ ( .A({ _tmp_1138[23:22], _tmp_1138[20], _tmp_1138[17] }), .Y(_11223_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36513_ ( .A({ _tmp_1138[8], _tmp_1138[5], _tmp_1138[3:2] }), .Y(_11224_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36514_ ( .A({ _tmp_1138[15:14], _tmp_1138[12], _tmp_1138[9] }), .Y(_11225_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36515_ ( .A({ _wvalid_1135, _06293_ }), .Y(_06294_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36516_ ( .A({ _dataflow_slice_valid_130, _11226_ }), .Y(_06296_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36517_ ( .A({ _tmp_1141, _11227_ }), .Y(_11226_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36518_ ( .A({ _11228_, _tmp_1140[0], _tmp_1140[33:32] }), .Y(_11227_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36519_ ( .A({ _11237_, _11236_, _11234_, _11229_ }), .Y(_11228_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36520_ ( .A({ _11233_, _11232_, _11231_, _11230_ }), .Y(_11229_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36521_ ( .A({ _tmp_1140[24], _tmp_1140[21], _tmp_1140[19:18] }), .Y(_11230_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36522_ ( .A({ _tmp_1140[31], _tmp_1140[29:28], _tmp_1140[25] }), .Y(_11231_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36523_ ( .A({ _tmp_1140[7:6], _tmp_1140[4], _tmp_1140[1] }), .Y(_11232_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36524_ ( .A({ _tmp_1140[16], _tmp_1140[13], _tmp_1140[11:10] }), .Y(_11233_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36525_ ( .A({ _11235_, _tmp_1140[30], _tmp_1140[27:26] }), .Y(_11234_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36526_ ( .A({ _tmp_1140[23:22], _tmp_1140[20], _tmp_1140[17] }), .Y(_11235_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36527_ ( .A({ _tmp_1140[8], _tmp_1140[5], _tmp_1140[3:2] }), .Y(_11236_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36528_ ( .A({ _tmp_1140[15:14], _tmp_1140[12], _tmp_1140[9] }), .Y(_11237_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36529_ ( .A({ _wvalid_1135, _06296_ }), .Y(_06297_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36530_ ( .A({ _dataflow_slice_valid_133, _11238_ }), .Y(_06299_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36531_ ( .A({ _tmp_1143, _11239_ }), .Y(_11238_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36532_ ( .A({ _11240_, _tmp_1142[0], _tmp_1142[33:32] }), .Y(_11239_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36533_ ( .A({ _11249_, _11248_, _11246_, _11241_ }), .Y(_11240_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36534_ ( .A({ _11245_, _11244_, _11243_, _11242_ }), .Y(_11241_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36535_ ( .A({ _tmp_1142[24], _tmp_1142[21], _tmp_1142[19:18] }), .Y(_11242_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36536_ ( .A({ _tmp_1142[31], _tmp_1142[29:28], _tmp_1142[25] }), .Y(_11243_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36537_ ( .A({ _tmp_1142[7:6], _tmp_1142[4], _tmp_1142[1] }), .Y(_11244_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36538_ ( .A({ _tmp_1142[16], _tmp_1142[13], _tmp_1142[11:10] }), .Y(_11245_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36539_ ( .A({ _11247_, _tmp_1142[30], _tmp_1142[27:26] }), .Y(_11246_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36540_ ( .A({ _tmp_1142[23:22], _tmp_1142[20], _tmp_1142[17] }), .Y(_11247_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36541_ ( .A({ _tmp_1142[8], _tmp_1142[5], _tmp_1142[3:2] }), .Y(_11248_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36542_ ( .A({ _tmp_1142[15:14], _tmp_1142[12], _tmp_1142[9] }), .Y(_11249_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36543_ ( .A({ _wvalid_1135, _06299_ }), .Y(_06300_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36544_ ( .A({ _dataflow_slice_valid_136, _11250_ }), .Y(_06302_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36545_ ( .A({ _tmp_1145, _11251_ }), .Y(_11250_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36546_ ( .A({ _11252_, _tmp_1144[0], _tmp_1144[33:32] }), .Y(_11251_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36547_ ( .A({ _11261_, _11260_, _11258_, _11253_ }), .Y(_11252_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36548_ ( .A({ _11257_, _11256_, _11255_, _11254_ }), .Y(_11253_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36549_ ( .A({ _tmp_1144[24], _tmp_1144[21], _tmp_1144[19:18] }), .Y(_11254_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36550_ ( .A({ _tmp_1144[31], _tmp_1144[29:28], _tmp_1144[25] }), .Y(_11255_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36551_ ( .A({ _tmp_1144[7:6], _tmp_1144[4], _tmp_1144[1] }), .Y(_11256_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36552_ ( .A({ _tmp_1144[16], _tmp_1144[13], _tmp_1144[11:10] }), .Y(_11257_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36553_ ( .A({ _11259_, _tmp_1144[30], _tmp_1144[27:26] }), .Y(_11258_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36554_ ( .A({ _tmp_1144[23:22], _tmp_1144[20], _tmp_1144[17] }), .Y(_11259_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36555_ ( .A({ _tmp_1144[8], _tmp_1144[5], _tmp_1144[3:2] }), .Y(_11260_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36556_ ( .A({ _tmp_1144[15:14], _tmp_1144[12], _tmp_1144[9] }), .Y(_11261_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36557_ ( .A({ _wvalid_1135, _06302_ }), .Y(_06303_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36558_ ( .A({ _dataflow_slice_valid_139, _11262_ }), .Y(_06305_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36559_ ( .A({ _tmp_1147, _11263_ }), .Y(_11262_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36560_ ( .A({ _11264_, _tmp_1146[0], _tmp_1146[33:32] }), .Y(_11263_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36561_ ( .A({ _11273_, _11272_, _11270_, _11265_ }), .Y(_11264_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36562_ ( .A({ _11269_, _11268_, _11267_, _11266_ }), .Y(_11265_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36563_ ( .A({ _tmp_1146[24], _tmp_1146[21], _tmp_1146[19:18] }), .Y(_11266_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36564_ ( .A({ _tmp_1146[31], _tmp_1146[29:28], _tmp_1146[25] }), .Y(_11267_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36565_ ( .A({ _tmp_1146[7:6], _tmp_1146[4], _tmp_1146[1] }), .Y(_11268_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36566_ ( .A({ _tmp_1146[16], _tmp_1146[13], _tmp_1146[11:10] }), .Y(_11269_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36567_ ( .A({ _11271_, _tmp_1146[30], _tmp_1146[27:26] }), .Y(_11270_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36568_ ( .A({ _tmp_1146[23:22], _tmp_1146[20], _tmp_1146[17] }), .Y(_11271_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36569_ ( .A({ _tmp_1146[8], _tmp_1146[5], _tmp_1146[3:2] }), .Y(_11272_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36570_ ( .A({ _tmp_1146[15:14], _tmp_1146[12], _tmp_1146[9] }), .Y(_11273_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36571_ ( .A({ _wvalid_1135, _06305_ }), .Y(_06306_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36572_ ( .A({ _dataflow_slice_valid_142, _11274_ }), .Y(_06308_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36573_ ( .A({ _tmp_1149, _11275_ }), .Y(_11274_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36574_ ( .A({ _11276_, _tmp_1148[0], _tmp_1148[33:32] }), .Y(_11275_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36575_ ( .A({ _11285_, _11284_, _11282_, _11277_ }), .Y(_11276_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36576_ ( .A({ _11281_, _11280_, _11279_, _11278_ }), .Y(_11277_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36577_ ( .A({ _tmp_1148[24], _tmp_1148[21], _tmp_1148[19:18] }), .Y(_11278_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36578_ ( .A({ _tmp_1148[31], _tmp_1148[29:28], _tmp_1148[25] }), .Y(_11279_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36579_ ( .A({ _tmp_1148[7:6], _tmp_1148[4], _tmp_1148[1] }), .Y(_11280_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36580_ ( .A({ _tmp_1148[16], _tmp_1148[13], _tmp_1148[11:10] }), .Y(_11281_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36581_ ( .A({ _11283_, _tmp_1148[30], _tmp_1148[27:26] }), .Y(_11282_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36582_ ( .A({ _tmp_1148[23:22], _tmp_1148[20], _tmp_1148[17] }), .Y(_11283_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36583_ ( .A({ _tmp_1148[8], _tmp_1148[5], _tmp_1148[3:2] }), .Y(_11284_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36584_ ( .A({ _tmp_1148[15:14], _tmp_1148[12], _tmp_1148[9] }), .Y(_11285_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36585_ ( .A({ _wvalid_1135, _06308_ }), .Y(_06309_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36586_ ( .A({ _dataflow_slice_valid_145, _11286_ }), .Y(_06311_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36587_ ( .A({ _tmp_1151, _11287_ }), .Y(_11286_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36588_ ( .A({ _11288_, _tmp_1150[0], _tmp_1150[33:32] }), .Y(_11287_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36589_ ( .A({ _11297_, _11296_, _11294_, _11289_ }), .Y(_11288_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36590_ ( .A({ _11293_, _11292_, _11291_, _11290_ }), .Y(_11289_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36591_ ( .A({ _tmp_1150[24], _tmp_1150[21], _tmp_1150[19:18] }), .Y(_11290_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36592_ ( .A({ _tmp_1150[31], _tmp_1150[29:28], _tmp_1150[25] }), .Y(_11291_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36593_ ( .A({ _tmp_1150[7:6], _tmp_1150[4], _tmp_1150[1] }), .Y(_11292_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36594_ ( .A({ _tmp_1150[16], _tmp_1150[13], _tmp_1150[11:10] }), .Y(_11293_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36595_ ( .A({ _11295_, _tmp_1150[30], _tmp_1150[27:26] }), .Y(_11294_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36596_ ( .A({ _tmp_1150[23:22], _tmp_1150[20], _tmp_1150[17] }), .Y(_11295_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36597_ ( .A({ _tmp_1150[8], _tmp_1150[5], _tmp_1150[3:2] }), .Y(_11296_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36598_ ( .A({ _tmp_1150[15:14], _tmp_1150[12], _tmp_1150[9] }), .Y(_11297_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36599_ ( .A({ _wvalid_1135, _06311_ }), .Y(_06312_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36600_ ( .A({ _dataflow_slice_valid_149, _11298_ }), .Y(_06314_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36601_ ( .A({ _tmp_1156, _11299_ }), .Y(_11298_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36602_ ( .A({ _11300_, _tmp_1155[0], _tmp_1155[33:32] }), .Y(_11299_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36603_ ( .A({ _11309_, _11308_, _11306_, _11301_ }), .Y(_11300_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36604_ ( .A({ _11305_, _11304_, _11303_, _11302_ }), .Y(_11301_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36605_ ( .A({ _tmp_1155[24], _tmp_1155[21], _tmp_1155[19:18] }), .Y(_11302_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36606_ ( .A({ _tmp_1155[31], _tmp_1155[29:28], _tmp_1155[25] }), .Y(_11303_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36607_ ( .A({ _tmp_1155[7:6], _tmp_1155[4], _tmp_1155[1] }), .Y(_11304_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36608_ ( .A({ _tmp_1155[16], _tmp_1155[13], _tmp_1155[11:10] }), .Y(_11305_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36609_ ( .A({ _11307_, _tmp_1155[30], _tmp_1155[27:26] }), .Y(_11306_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36610_ ( .A({ _tmp_1155[23:22], _tmp_1155[20], _tmp_1155[17] }), .Y(_11307_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36611_ ( .A({ _tmp_1155[8], _tmp_1155[5], _tmp_1155[3:2] }), .Y(_11308_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36612_ ( .A({ _tmp_1155[15:14], _tmp_1155[12], _tmp_1155[9] }), .Y(_11309_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36613_ ( .A({ _wvalid_1154, _06314_ }), .Y(_06315_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36614_ ( .A({ _dataflow_slice_valid_152, _11310_ }), .Y(_06317_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36615_ ( .A({ _tmp_1158, _11311_ }), .Y(_11310_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36616_ ( .A({ _11312_, _tmp_1157[0], _tmp_1157[33:32] }), .Y(_11311_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36617_ ( .A({ _11321_, _11320_, _11318_, _11313_ }), .Y(_11312_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36618_ ( .A({ _11317_, _11316_, _11315_, _11314_ }), .Y(_11313_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36619_ ( .A({ _tmp_1157[24], _tmp_1157[21], _tmp_1157[19:18] }), .Y(_11314_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36620_ ( .A({ _tmp_1157[31], _tmp_1157[29:28], _tmp_1157[25] }), .Y(_11315_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36621_ ( .A({ _tmp_1157[7:6], _tmp_1157[4], _tmp_1157[1] }), .Y(_11316_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36622_ ( .A({ _tmp_1157[16], _tmp_1157[13], _tmp_1157[11:10] }), .Y(_11317_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36623_ ( .A({ _11319_, _tmp_1157[30], _tmp_1157[27:26] }), .Y(_11318_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36624_ ( .A({ _tmp_1157[23:22], _tmp_1157[20], _tmp_1157[17] }), .Y(_11319_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36625_ ( .A({ _tmp_1157[8], _tmp_1157[5], _tmp_1157[3:2] }), .Y(_11320_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36626_ ( .A({ _tmp_1157[15:14], _tmp_1157[12], _tmp_1157[9] }), .Y(_11321_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36627_ ( .A({ _wvalid_1154, _06317_ }), .Y(_06318_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36628_ ( .A({ _dataflow_slice_valid_155, _11322_ }), .Y(_06320_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36629_ ( .A({ _tmp_1160, _11323_ }), .Y(_11322_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36630_ ( .A({ _11324_, _tmp_1159[0], _tmp_1159[33:32] }), .Y(_11323_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36631_ ( .A({ _11333_, _11332_, _11330_, _11325_ }), .Y(_11324_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36632_ ( .A({ _11329_, _11328_, _11327_, _11326_ }), .Y(_11325_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36633_ ( .A({ _tmp_1159[24], _tmp_1159[21], _tmp_1159[19:18] }), .Y(_11326_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36634_ ( .A({ _tmp_1159[31], _tmp_1159[29:28], _tmp_1159[25] }), .Y(_11327_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36635_ ( .A({ _tmp_1159[7:6], _tmp_1159[4], _tmp_1159[1] }), .Y(_11328_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36636_ ( .A({ _tmp_1159[16], _tmp_1159[13], _tmp_1159[11:10] }), .Y(_11329_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36637_ ( .A({ _11331_, _tmp_1159[30], _tmp_1159[27:26] }), .Y(_11330_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36638_ ( .A({ _tmp_1159[23:22], _tmp_1159[20], _tmp_1159[17] }), .Y(_11331_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36639_ ( .A({ _tmp_1159[8], _tmp_1159[5], _tmp_1159[3:2] }), .Y(_11332_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36640_ ( .A({ _tmp_1159[15:14], _tmp_1159[12], _tmp_1159[9] }), .Y(_11333_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36641_ ( .A({ _wvalid_1154, _06320_ }), .Y(_06321_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36642_ ( .A({ _dataflow_slice_valid_158, _11334_ }), .Y(_06323_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _36643_ ( .A({ _tmp_1162, _11335_ }), .Y(_11334_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36644_ ( .A({ _11336_, _tmp_1161[0], _tmp_1161[33:32] }), .Y(_11335_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36645_ ( .A({ _11345_, _11344_, _11342_, _11337_ }), .Y(_11336_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36646_ ( .A({ _11341_, _11340_, _11339_, _11338_ }), .Y(_11337_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36647_ ( .A({ _tmp_1161[24], _tmp_1161[21], _tmp_1161[19:18] }), .Y(_11338_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36648_ ( .A({ _tmp_1161[31], _tmp_1161[29:28], _tmp_1161[25] }), .Y(_11339_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36649_ ( .A({ _tmp_1161[7:6], _tmp_1161[4], _tmp_1161[1] }), .Y(_11340_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36650_ ( .A({ _tmp_1161[16], _tmp_1161[13], _tmp_1161[11:10] }), .Y(_11341_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36651_ ( .A({ _11343_, _tmp_1161[30], _tmp_1161[27:26] }), .Y(_11342_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36652_ ( .A({ _tmp_1161[23:22], _tmp_1161[20], _tmp_1161[17] }), .Y(_11343_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36653_ ( .A({ _tmp_1161[8], _tmp_1161[5], _tmp_1161[3:2] }), .Y(_11344_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36654_ ( .A({ _tmp_1161[15:14], _tmp_1161[12], _tmp_1161[9] }), .Y(_11345_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36655_ ( .A({ _wvalid_1154, _06323_ }), .Y(_06324_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36656_ ( .A({ saxi_bready, saxi_bvalid }), .Y(_06326_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36657_ ( .A({ saxi_awvalid, saxi_awready }), .Y(_06328_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36658_ ( .A({ saxi_arvalid, saxi_arready }), .Y(_06329_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36659_ ( .A({ saxi_rvalid, saxi_rready }), .Y(_06331_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36660_ ( .A({ _tmp_7, _06330_, _05719_ }), .Y(_06332_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36661_ ( .A({ _saxi_register_fsm[0], _10012_, _06331_ }), .Y(_06330_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36662_ ( .A({ _tmp_7, _06330_, _05866_ }), .Y(_06333_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36663_ ( .A({ _tmp_7, _06330_, _05867_ }), .Y(_06334_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36664_ ( .A({ _tmp_7, _06330_, _05868_ }), .Y(_06335_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36665_ ( .A({ _tmp_7, _06330_, _05869_ }), .Y(_06336_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36666_ ( .A({ _tmp_7, _06330_, _05870_ }), .Y(_06337_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36667_ ( .A({ _tmp_7, _06330_, _05871_ }), .Y(_06338_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36668_ ( .A({ _tmp_7, _06330_, _05872_ }), .Y(_06339_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36669_ ( .A({ _tmp_7, _06330_, _05873_ }), .Y(_06340_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36670_ ( .A({ _tmp_7, _06330_, _05874_ }), .Y(_06341_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36671_ ( .A({ _tmp_7, _06330_, _05875_ }), .Y(_06342_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36672_ ( .A({ _tmp_7, _06330_, _05876_ }), .Y(_06343_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36673_ ( .A({ _tmp_7, _06330_, _05877_ }), .Y(_06344_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36674_ ( .A({ _tmp_7, _06330_, _05878_ }), .Y(_06345_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36675_ ( .A({ _06327_, _05719_ }), .Y(_06346_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36676_ ( .A({ saxi_wvalid, saxi_wready }), .Y(_06327_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36677_ ( .A({ _06327_, _05866_ }), .Y(_06347_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36678_ ( .A({ _06327_, _05867_ }), .Y(_06348_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36679_ ( .A({ _06327_, _05868_ }), .Y(_06349_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36680_ ( .A({ _06327_, _05869_ }), .Y(_06350_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36681_ ( .A({ _06327_, _05870_ }), .Y(_06351_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36682_ ( .A({ _06327_, _05871_ }), .Y(_06352_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36683_ ( .A({ _06327_, _05872_ }), .Y(_06353_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36684_ ( .A({ _06327_, _05873_ }), .Y(_06354_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36685_ ( .A({ _06327_, _05874_ }), .Y(_06355_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36686_ ( .A({ _06327_, _05875_ }), .Y(_06356_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36687_ ( .A({ _06327_, _05876_ }), .Y(_06357_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36688_ ( .A({ _06327_, _05877_ }), .Y(_06358_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36689_ ( .A({ _06327_, _05878_ }), .Y(_06359_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36690_ ( .A({ _maxi_read_start, _maxi_read_op_sel[1:0], _11346_ }), .Y(_06360_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36691_ ( .A({ _11347_, _maxi_read_op_sel[3:2] }), .Y(_11346_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36692_ ( .A(_maxi_read_op_sel[7:4]), .Y(_11347_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36693_ ( .A({ _06360_, _10922_ }), .Y(_06361_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36694_ ( .A({ _dataflow_slice_valid_29, _tmp_40, _10922_ }), .Y(_06220_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36695_ ( .A({ _11350_, _11349_, _11348_, _06220_ }), .Y(_06362_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _36696_ ( .A(_tmp_38[10:8]), .Y(_11348_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36697_ ( .A(_tmp_38[7:4]), .Y(_11349_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36698_ ( .A(_tmp_38[3:0]), .Y(_11350_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36699_ ( .A({ _06027_, _06362_ }), .Y(_06363_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36700_ ( .A({ _06028_, _06220_ }), .Y(_06364_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36701_ ( .A({ _06029_, _06220_ }), .Y(_06365_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36702_ ( .A({ _06030_, _06220_ }), .Y(_06366_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36703_ ( .A({ _06031_, _06220_ }), .Y(_06367_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36704_ ( .A({ _06032_, _06220_ }), .Y(_06368_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36705_ ( .A({ _06033_, _06220_ }), .Y(_06369_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36706_ ( .A({ _06034_, _06220_ }), .Y(_06370_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36707_ ( .A({ _06035_, _06220_ }), .Y(_06371_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36708_ ( .A({ _06027_, _06220_ }), .Y(_06372_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36709_ ( .A({ _11351_, _06220_ }), .Y(_06373_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36710_ ( .A({ _10923_, _tmp_39[33:32] }), .Y(_11351_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36711_ ( .A({ _maxi_read_start, _11352_, _maxi_read_op_sel[1:0] }), .Y(_06374_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36712_ ( .A({ _maxi_read_op_sel[3], _11347_, _maxi_read_op_sel[2] }), .Y(_11352_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36713_ ( .A({ _06374_, _11203_ }), .Y(_06375_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36714_ ( .A({ _dataflow_slice_valid_124, _11202_ }), .Y(_06292_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36715_ ( .A({ _11353_, _06292_ }), .Y(_06376_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36716_ ( .A({ _tmp_1136[0], _11204_, _tmp_1136[33:32] }), .Y(_11353_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36717_ ( .A({ _06360_, _10933_ }), .Y(_06377_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36718_ ( .A({ _dataflow_slice_valid_32, _tmp_71, _10933_ }), .Y(_06223_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36719_ ( .A({ _11356_, _11355_, _11354_, _06223_ }), .Y(_06378_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _36720_ ( .A(_tmp_69[10:8]), .Y(_11354_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36721_ ( .A(_tmp_69[7:4]), .Y(_11355_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36722_ ( .A(_tmp_69[3:0]), .Y(_11356_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36723_ ( .A({ _06036_, _06378_ }), .Y(_06379_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36724_ ( .A({ _06037_, _06223_ }), .Y(_06380_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36725_ ( .A({ _06038_, _06223_ }), .Y(_06381_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36726_ ( .A({ _06039_, _06223_ }), .Y(_06382_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36727_ ( .A({ _06040_, _06223_ }), .Y(_06383_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36728_ ( .A({ _06041_, _06223_ }), .Y(_06384_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36729_ ( .A({ _06042_, _06223_ }), .Y(_06385_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36730_ ( .A({ _06043_, _06223_ }), .Y(_06386_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36731_ ( .A({ _06044_, _06223_ }), .Y(_06387_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36732_ ( .A({ _06036_, _06223_ }), .Y(_06388_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36733_ ( .A({ _11357_, _06223_ }), .Y(_06389_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36734_ ( .A({ _10934_, _tmp_70[33:32] }), .Y(_11357_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36735_ ( .A({ _06374_, _11215_ }), .Y(_06390_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36736_ ( .A({ _dataflow_slice_valid_127, _11214_ }), .Y(_06295_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36737_ ( .A({ _11358_, _06295_ }), .Y(_06391_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36738_ ( .A({ _tmp_1138[0], _11216_, _tmp_1138[33:32] }), .Y(_11358_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36739_ ( .A({ _06360_, _10944_ }), .Y(_06392_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36740_ ( .A({ _dataflow_slice_valid_35, _tmp_102, _10944_ }), .Y(_06226_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36741_ ( .A({ _11361_, _11360_, _11359_, _06226_ }), .Y(_06393_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _36742_ ( .A(_tmp_100[10:8]), .Y(_11359_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36743_ ( .A(_tmp_100[7:4]), .Y(_11360_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36744_ ( .A(_tmp_100[3:0]), .Y(_11361_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36745_ ( .A({ _06045_, _06393_ }), .Y(_06394_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36746_ ( .A({ _06046_, _06226_ }), .Y(_06395_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36747_ ( .A({ _06047_, _06226_ }), .Y(_06396_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36748_ ( .A({ _06048_, _06226_ }), .Y(_06397_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36749_ ( .A({ _06049_, _06226_ }), .Y(_06398_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36750_ ( .A({ _06050_, _06226_ }), .Y(_06399_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36751_ ( .A({ _06051_, _06226_ }), .Y(_06400_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36752_ ( .A({ _06052_, _06226_ }), .Y(_06401_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36753_ ( .A({ _06053_, _06226_ }), .Y(_06402_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36754_ ( .A({ _06045_, _06226_ }), .Y(_06403_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36755_ ( .A({ _11362_, _06226_ }), .Y(_06404_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36756_ ( .A({ _10945_, _tmp_101[33:32] }), .Y(_11362_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36757_ ( .A({ _06374_, _11227_ }), .Y(_06405_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36758_ ( .A({ _dataflow_slice_valid_130, _11226_ }), .Y(_06298_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36759_ ( .A({ _11363_, _06298_ }), .Y(_06406_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36760_ ( .A({ _tmp_1140[0], _11228_, _tmp_1140[33:32] }), .Y(_11363_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36761_ ( .A({ _06360_, _10955_ }), .Y(_06407_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36762_ ( .A({ _dataflow_slice_valid_38, _tmp_133, _10955_ }), .Y(_06229_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36763_ ( .A({ _11366_, _11365_, _11364_, _06229_ }), .Y(_06408_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _36764_ ( .A(_tmp_131[10:8]), .Y(_11364_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36765_ ( .A(_tmp_131[7:4]), .Y(_11365_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36766_ ( .A(_tmp_131[3:0]), .Y(_11366_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36767_ ( .A({ _06054_, _06408_ }), .Y(_06409_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36768_ ( .A({ _06055_, _06229_ }), .Y(_06410_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36769_ ( .A({ _06056_, _06229_ }), .Y(_06411_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36770_ ( .A({ _06057_, _06229_ }), .Y(_06412_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36771_ ( .A({ _06058_, _06229_ }), .Y(_06413_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36772_ ( .A({ _06059_, _06229_ }), .Y(_06414_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36773_ ( .A({ _06060_, _06229_ }), .Y(_06415_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36774_ ( .A({ _06061_, _06229_ }), .Y(_06416_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36775_ ( .A({ _06062_, _06229_ }), .Y(_06417_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36776_ ( .A({ _06054_, _06229_ }), .Y(_06418_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36777_ ( .A({ _11367_, _06229_ }), .Y(_06419_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36778_ ( .A({ _10956_, _tmp_132[33:32] }), .Y(_11367_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36779_ ( .A({ _06374_, _11239_ }), .Y(_06420_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36780_ ( .A({ _dataflow_slice_valid_133, _11238_ }), .Y(_06301_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36781_ ( .A({ _11368_, _06301_ }), .Y(_06421_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36782_ ( .A({ _tmp_1142[0], _11240_, _tmp_1142[33:32] }), .Y(_11368_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36783_ ( .A({ _06360_, _10966_ }), .Y(_06422_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36784_ ( .A({ _dataflow_slice_valid_41, _tmp_164, _10966_ }), .Y(_06232_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36785_ ( .A({ _11371_, _11370_, _11369_, _06232_ }), .Y(_06423_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _36786_ ( .A(_tmp_162[10:8]), .Y(_11369_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36787_ ( .A(_tmp_162[7:4]), .Y(_11370_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36788_ ( .A(_tmp_162[3:0]), .Y(_11371_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36789_ ( .A({ _06063_, _06423_ }), .Y(_06424_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36790_ ( .A({ _06064_, _06232_ }), .Y(_06425_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36791_ ( .A({ _06065_, _06232_ }), .Y(_06426_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36792_ ( .A({ _06066_, _06232_ }), .Y(_06427_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36793_ ( .A({ _06067_, _06232_ }), .Y(_06428_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36794_ ( .A({ _06068_, _06232_ }), .Y(_06429_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36795_ ( .A({ _06069_, _06232_ }), .Y(_06430_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36796_ ( .A({ _06070_, _06232_ }), .Y(_06431_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36797_ ( .A({ _06071_, _06232_ }), .Y(_06432_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36798_ ( .A({ _06063_, _06232_ }), .Y(_06433_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36799_ ( .A({ _11372_, _06232_ }), .Y(_06434_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36800_ ( .A({ _10967_, _tmp_163[33:32] }), .Y(_11372_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36801_ ( .A({ _06374_, _11251_ }), .Y(_06435_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36802_ ( .A({ _dataflow_slice_valid_136, _11250_ }), .Y(_06304_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36803_ ( .A({ _11373_, _06304_ }), .Y(_06436_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36804_ ( .A({ _tmp_1144[0], _11252_, _tmp_1144[33:32] }), .Y(_11373_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36805_ ( .A({ _06360_, _10977_ }), .Y(_06437_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36806_ ( .A({ _dataflow_slice_valid_44, _tmp_195, _10977_ }), .Y(_06235_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36807_ ( .A({ _11376_, _11375_, _11374_, _06235_ }), .Y(_06438_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _36808_ ( .A(_tmp_193[10:8]), .Y(_11374_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36809_ ( .A(_tmp_193[7:4]), .Y(_11375_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36810_ ( .A(_tmp_193[3:0]), .Y(_11376_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36811_ ( .A({ _06072_, _06438_ }), .Y(_06439_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36812_ ( .A({ _06073_, _06235_ }), .Y(_06440_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36813_ ( .A({ _06074_, _06235_ }), .Y(_06441_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36814_ ( .A({ _06075_, _06235_ }), .Y(_06442_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36815_ ( .A({ _06076_, _06235_ }), .Y(_06443_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36816_ ( .A({ _06077_, _06235_ }), .Y(_06444_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36817_ ( .A({ _06078_, _06235_ }), .Y(_06445_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36818_ ( .A({ _06079_, _06235_ }), .Y(_06446_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36819_ ( .A({ _06080_, _06235_ }), .Y(_06447_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36820_ ( .A({ _06072_, _06235_ }), .Y(_06448_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36821_ ( .A({ _11377_, _06235_ }), .Y(_06449_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36822_ ( .A({ _10978_, _tmp_194[33:32] }), .Y(_11377_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36823_ ( .A({ _06374_, _11263_ }), .Y(_06450_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36824_ ( .A({ _dataflow_slice_valid_139, _11262_ }), .Y(_06307_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36825_ ( .A({ _11378_, _06307_ }), .Y(_06451_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36826_ ( .A({ _tmp_1146[0], _11264_, _tmp_1146[33:32] }), .Y(_11378_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36827_ ( .A({ _06360_, _10988_ }), .Y(_06452_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36828_ ( .A({ _dataflow_slice_valid_47, _tmp_226, _10988_ }), .Y(_06238_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36829_ ( .A({ _11381_, _11380_, _11379_, _06238_ }), .Y(_06453_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _36830_ ( .A(_tmp_224[10:8]), .Y(_11379_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36831_ ( .A(_tmp_224[7:4]), .Y(_11380_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36832_ ( .A(_tmp_224[3:0]), .Y(_11381_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36833_ ( .A({ _06081_, _06453_ }), .Y(_06454_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36834_ ( .A({ _06082_, _06238_ }), .Y(_06455_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36835_ ( .A({ _06083_, _06238_ }), .Y(_06456_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36836_ ( .A({ _06084_, _06238_ }), .Y(_06457_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36837_ ( .A({ _06085_, _06238_ }), .Y(_06458_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36838_ ( .A({ _06086_, _06238_ }), .Y(_06459_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36839_ ( .A({ _06087_, _06238_ }), .Y(_06460_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36840_ ( .A({ _06088_, _06238_ }), .Y(_06461_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36841_ ( .A({ _06089_, _06238_ }), .Y(_06462_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36842_ ( .A({ _06081_, _06238_ }), .Y(_06463_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36843_ ( .A({ _11382_, _06238_ }), .Y(_06464_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36844_ ( .A({ _10989_, _tmp_225[33:32] }), .Y(_11382_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36845_ ( .A({ _06374_, _11275_ }), .Y(_06465_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36846_ ( .A({ _dataflow_slice_valid_142, _11274_ }), .Y(_06310_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36847_ ( .A({ _11383_, _06310_ }), .Y(_06466_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36848_ ( .A({ _tmp_1148[0], _11276_, _tmp_1148[33:32] }), .Y(_11383_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36849_ ( .A({ _06360_, _10999_ }), .Y(_06467_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36850_ ( .A({ _dataflow_slice_valid_50, _tmp_257, _10999_ }), .Y(_06241_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36851_ ( .A({ _11386_, _11385_, _11384_, _06241_ }), .Y(_06468_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _36852_ ( .A(_tmp_255[10:8]), .Y(_11384_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36853_ ( .A(_tmp_255[7:4]), .Y(_11385_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36854_ ( .A(_tmp_255[3:0]), .Y(_11386_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36855_ ( .A({ _06090_, _06468_ }), .Y(_06469_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36856_ ( .A({ _06091_, _06241_ }), .Y(_06470_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36857_ ( .A({ _06092_, _06241_ }), .Y(_06471_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36858_ ( .A({ _06093_, _06241_ }), .Y(_06472_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36859_ ( .A({ _06094_, _06241_ }), .Y(_06473_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36860_ ( .A({ _06095_, _06241_ }), .Y(_06474_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36861_ ( .A({ _06096_, _06241_ }), .Y(_06475_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36862_ ( .A({ _06097_, _06241_ }), .Y(_06476_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36863_ ( .A({ _06098_, _06241_ }), .Y(_06477_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36864_ ( .A({ _06090_, _06241_ }), .Y(_06478_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36865_ ( .A({ _11387_, _06241_ }), .Y(_06479_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36866_ ( .A({ _11000_, _tmp_256[33:32] }), .Y(_11387_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36867_ ( .A({ _stream_conv2d_16_source_28_source_ram_renable, _05879_ }), .Y(_tmp_597) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36868_ ( .A({ _06374_, _11287_ }), .Y(_06480_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36869_ ( .A({ _dataflow_slice_valid_145, _11286_ }), .Y(_06313_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36870_ ( .A({ _11388_, _06313_ }), .Y(_06481_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36871_ ( .A({ _tmp_1150[0], _11288_, _tmp_1150[33:32] }), .Y(_11388_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36872_ ( .A({ _stream_matmul_29_source_20_source_ram_renable, _05880_ }), .Y(_tmp_1223) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36873_ ( .A({ _stream_conv2d_16_source_29_source_ram_renable, _05881_ }), .Y(_tmp_611) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36874_ ( .A({ _stream_conv2d_16_source_30_source_ram_renable, _05882_ }), .Y(_tmp_625) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36875_ ( .A({ _stream_conv2d_16_source_31_source_ram_renable, _05883_ }), .Y(_tmp_639) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36876_ ( .A({ _stream_conv2d_16_source_32_source_ram_renable, _05884_ }), .Y(_tmp_653) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36877_ ( .A({ _stream_conv2d_16_source_33_source_ram_renable, _05885_ }), .Y(_tmp_667) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36878_ ( .A({ _stream_conv2d_16_source_34_source_ram_renable, _05886_ }), .Y(_tmp_681) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36879_ ( .A({ _stream_conv2d_16_source_35_source_ram_renable, _05887_ }), .Y(_tmp_695) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36880_ ( .A({ _stream_conv2d_16_source_36_source_ram_renable, _05888_ }), .Y(_tmp_709) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _36881_ ( .A({ _maxi_read_start, _maxi_read_op_sel[1], _11346_, _maxi_read_op_sel[0] }), .Y(_06482_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36882_ ( .A({ _06482_, _10875_ }), .Y(_06483_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36883_ ( .A({ _dataflow_slice_valid_16, _10874_ }), .Y(_06208_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36884_ ( .A({ _11389_, _06208_ }), .Y(_06484_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36885_ ( .A({ _tmp_25[0], _10876_, _tmp_25[33:32] }), .Y(_11389_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36886_ ( .A({ _11390_, _stream_max_pool_serial_18_sink_3_sink_waddr[1] }), .Y(_06485_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36887_ ( .A({ _11391_, _stream_max_pool_serial_18_sink_3_sink_waddr[0] }), .Y(_11390_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36888_ ( .A({ _11393_, _11392_, _stream_max_pool_serial_18_sink_3_sink_ram_sel[2], _stream_max_pool_serial_18_sink_3_sink_ram_sel[0] }), .Y(_11391_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _36889_ ( .A({ _stream_max_pool_serial_18_sink_3_sink_ram_sel[1], _stream_max_pool_serial_18_sink_3_sink_wenable, _stream_max_pool_serial_18_sink_3_sink_ram_sel[7] }), .Y(_11392_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36890_ ( .A(_stream_max_pool_serial_18_sink_3_sink_ram_sel[6:3]), .Y(_11393_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36891_ ( .A({ _tmp_1072, _06493_ }), .Y(_tmp_1077) );
  \$lut  #( .LUT(16'h8f00), .WIDTH(4) ) _36892_ ( .A({ _06492_, _dataflow_cat_valid_107, _10819_, _10824_ }), .Y(_06493_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36893_ ( .A({ _tmp_1108, _tmp_1096, _tmp_1084, _tmp_1072 }), .Y(_06492_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _36894_ ( .A({ _tmp_1080, _06493_, _tmp_1072 }), .Y(_06486_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _36895_ ( .A({ _tmp_1079, _06493_, _tmp_1072 }), .Y(_06487_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36896_ ( .A({ _maxi_write_start, _10824_ }), .Y(_06488_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36897_ ( .A({ _06488_, _11394_, _tmp_1082, _tmp_1081 }), .Y(_06489_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36898_ ( .A({ _11395_, _tmp_1083[0] }), .Y(_11394_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36899_ ( .A({ _11405_, _11400_, _11398_, _11396_ }), .Y(_11395_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36900_ ( .A({ _11397_, _tmp_1083[33:31] }), .Y(_11396_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36901_ ( .A({ _tmp_1083[29:28], _tmp_1083[26], _tmp_1083[23] }), .Y(_11397_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36902_ ( .A({ _11399_, _tmp_1083[2:1] }), .Y(_11398_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36903_ ( .A(_tmp_1083[6:3]), .Y(_11399_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36904_ ( .A({ _11404_, _11403_, _11402_, _11401_ }), .Y(_11400_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36905_ ( .A(_tmp_1083[14:11]), .Y(_11401_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36906_ ( .A(_tmp_1083[10:7]), .Y(_11402_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36907_ ( .A(_tmp_1083[22:19]), .Y(_11403_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36908_ ( .A(_tmp_1083[18:15]), .Y(_11404_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36909_ ( .A({ _tmp_1083[30], _tmp_1083[27], _tmp_1083[25:24] }), .Y(_11405_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _36910_ ( .A({ _11394_, _06493_, _tmp_1072 }), .Y(_06490_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _36911_ ( .A({ _11395_, _tmp_1083[0], _06493_, _tmp_1072 }), .Y(_06491_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36912_ ( .A({ _06482_, _10887_ }), .Y(_06494_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36913_ ( .A({ _dataflow_slice_valid_19, _10886_ }), .Y(_06211_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36914_ ( .A({ _11406_, _06211_ }), .Y(_06495_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36915_ ( .A({ _tmp_27[0], _10888_, _tmp_27[33:32] }), .Y(_11406_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36916_ ( .A({ _11407_, _stream_max_pool_serial_18_sink_3_sink_waddr[1] }), .Y(_06496_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36917_ ( .A({ _stream_max_pool_serial_18_sink_3_sink_waddr[0], _11391_ }), .Y(_11407_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36918_ ( .A({ _tmp_1084, _06493_ }), .Y(_tmp_1089) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _36919_ ( .A({ _tmp_1092, _06493_, _tmp_1084 }), .Y(_06497_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _36920_ ( .A({ _tmp_1091, _06493_, _tmp_1084 }), .Y(_06498_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36921_ ( .A({ _06488_, _11408_, _tmp_1094, _tmp_1093 }), .Y(_06499_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36922_ ( .A({ _11409_, _tmp_1095[0] }), .Y(_11408_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36923_ ( .A({ _11419_, _11414_, _11412_, _11410_ }), .Y(_11409_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36924_ ( .A({ _11411_, _tmp_1095[33:31] }), .Y(_11410_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36925_ ( .A({ _tmp_1095[29:28], _tmp_1095[26], _tmp_1095[23] }), .Y(_11411_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36926_ ( .A({ _11413_, _tmp_1095[2:1] }), .Y(_11412_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36927_ ( .A(_tmp_1095[6:3]), .Y(_11413_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36928_ ( .A({ _11418_, _11417_, _11416_, _11415_ }), .Y(_11414_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36929_ ( .A(_tmp_1095[14:11]), .Y(_11415_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36930_ ( .A(_tmp_1095[10:7]), .Y(_11416_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36931_ ( .A(_tmp_1095[22:19]), .Y(_11417_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36932_ ( .A(_tmp_1095[18:15]), .Y(_11418_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36933_ ( .A({ _tmp_1095[30], _tmp_1095[27], _tmp_1095[25:24] }), .Y(_11419_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _36934_ ( .A({ _11408_, _06493_, _tmp_1084 }), .Y(_06500_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _36935_ ( .A({ _11409_, _tmp_1095[0], _06493_, _tmp_1084 }), .Y(_06501_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36936_ ( .A({ _06482_, _10899_ }), .Y(_06502_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36937_ ( .A({ _dataflow_slice_valid_22, _10898_ }), .Y(_06214_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36938_ ( .A({ _11420_, _06214_ }), .Y(_06503_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36939_ ( .A({ _tmp_29[0], _10900_, _tmp_29[33:32] }), .Y(_11420_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36940_ ( .A({ _stream_max_pool_serial_18_sink_3_sink_waddr[1], _11390_ }), .Y(_06504_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36941_ ( .A({ _tmp_1096, _06493_ }), .Y(_tmp_1101) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _36942_ ( .A({ _tmp_1104, _06493_, _tmp_1096 }), .Y(_06505_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _36943_ ( .A({ _tmp_1103, _06493_, _tmp_1096 }), .Y(_06506_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36944_ ( .A({ _06488_, _11421_, _tmp_1106, _tmp_1105 }), .Y(_06507_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36945_ ( .A({ _11422_, _tmp_1107[0] }), .Y(_11421_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36946_ ( .A({ _11432_, _11427_, _11425_, _11423_ }), .Y(_11422_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36947_ ( .A({ _11424_, _tmp_1107[33:31] }), .Y(_11423_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36948_ ( .A({ _tmp_1107[29:28], _tmp_1107[26], _tmp_1107[23] }), .Y(_11424_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36949_ ( .A({ _11426_, _tmp_1107[2:1] }), .Y(_11425_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36950_ ( .A(_tmp_1107[6:3]), .Y(_11426_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36951_ ( .A({ _11431_, _11430_, _11429_, _11428_ }), .Y(_11427_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36952_ ( .A(_tmp_1107[14:11]), .Y(_11428_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36953_ ( .A(_tmp_1107[10:7]), .Y(_11429_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36954_ ( .A(_tmp_1107[22:19]), .Y(_11430_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36955_ ( .A(_tmp_1107[18:15]), .Y(_11431_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36956_ ( .A({ _tmp_1107[30], _tmp_1107[27], _tmp_1107[25:24] }), .Y(_11432_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _36957_ ( .A({ _11421_, _06493_, _tmp_1096 }), .Y(_06508_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _36958_ ( .A({ _11422_, _tmp_1107[0], _06493_, _tmp_1096 }), .Y(_06509_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36959_ ( .A({ _06482_, _10911_ }), .Y(_06510_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36960_ ( .A({ _dataflow_slice_valid_25, _10910_ }), .Y(_06217_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36961_ ( .A({ _11433_, _06217_ }), .Y(_06511_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36962_ ( .A({ _tmp_31[0], _10912_, _tmp_31[33:32] }), .Y(_11433_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36963_ ( .A({ _stream_conv2d_16_source_8_source_ram_renable, _05889_ }), .Y(_tmp_483) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36964_ ( .A({ _stream_max_pool_serial_18_sink_3_sink_waddr[1], _11407_ }), .Y(_06512_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36965_ ( .A({ _tmp_1108, _06493_ }), .Y(_tmp_1113) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _36966_ ( .A({ _tmp_1116, _06493_, _tmp_1108 }), .Y(_06513_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _36967_ ( .A({ _tmp_1115, _06493_, _tmp_1108 }), .Y(_06514_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36968_ ( .A({ _06488_, _11434_, _tmp_1118, _tmp_1117 }), .Y(_06515_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36969_ ( .A({ _11435_, _tmp_1119[0] }), .Y(_11434_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36970_ ( .A({ _11445_, _11440_, _11438_, _11436_ }), .Y(_11435_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _36971_ ( .A({ _11437_, _tmp_1119[33:31] }), .Y(_11436_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36972_ ( .A({ _tmp_1119[29:28], _tmp_1119[26], _tmp_1119[23] }), .Y(_11437_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _36973_ ( .A({ _11439_, _tmp_1119[2:1] }), .Y(_11438_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36974_ ( .A(_tmp_1119[6:3]), .Y(_11439_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36975_ ( .A({ _11444_, _11443_, _11442_, _11441_ }), .Y(_11440_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36976_ ( .A(_tmp_1119[14:11]), .Y(_11441_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36977_ ( .A(_tmp_1119[10:7]), .Y(_11442_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36978_ ( .A(_tmp_1119[22:19]), .Y(_11443_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36979_ ( .A(_tmp_1119[18:15]), .Y(_11444_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36980_ ( .A({ _tmp_1119[30], _tmp_1119[27], _tmp_1119[25:24] }), .Y(_11445_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _36981_ ( .A({ _11434_, _06493_, _tmp_1108 }), .Y(_06516_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _36982_ ( .A({ _11435_, _tmp_1119[0], _06493_, _tmp_1108 }), .Y(_06517_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36983_ ( .A({ _stream_matmul_29_source_8_source_ram_renable, _05890_ }), .Y(_tmp_1189) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _36984_ ( .A({ _maxi_read_start, _11346_, _maxi_read_op_sel[0], _maxi_read_op_sel[1] }), .Y(_06518_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36985_ ( .A({ _06518_, _10827_ }), .Y(_06519_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36986_ ( .A({ _dataflow_slice_valid_3, _10826_ }), .Y(_06196_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36987_ ( .A({ _11446_, _06196_ }), .Y(_06520_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36988_ ( .A({ _tmp_12[0], _10828_, _tmp_12[33:32] }), .Y(_11446_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36989_ ( .A({ _11447_, _stream_matmul_29_sink_21_sink_waddr[1] }), .Y(_06521_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _36990_ ( .A({ _11448_, _stream_matmul_29_sink_21_sink_waddr[0] }), .Y(_11447_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _36991_ ( .A({ _11450_, _11449_, _stream_matmul_29_sink_21_sink_ram_sel[3], _stream_matmul_29_sink_21_sink_ram_sel[1] }), .Y(_11448_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _36992_ ( .A({ _stream_matmul_29_sink_21_sink_ram_sel[2], _stream_matmul_29_sink_21_sink_ram_sel[0], _stream_matmul_29_sink_21_sink_wenable }), .Y(_11449_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _36993_ ( .A(_stream_matmul_29_sink_21_sink_ram_sel[7:4]), .Y(_11450_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _36994_ ( .A({ _tmp_1309, _06529_ }), .Y(_tmp_1314) );
  \$lut  #( .LUT(16'h8f00), .WIDTH(4) ) _36995_ ( .A({ _06528_, _dataflow_cat_valid_167, _10819_, _10825_ }), .Y(_06529_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _36996_ ( .A({ _tmp_1345, _tmp_1333, _tmp_1321, _tmp_1309 }), .Y(_06528_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _36997_ ( .A({ _tmp_1317, _06529_, _tmp_1309 }), .Y(_06522_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _36998_ ( .A({ _tmp_1316, _06529_, _tmp_1309 }), .Y(_06523_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _36999_ ( .A({ _maxi_write_start, _10825_ }), .Y(_06524_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37000_ ( .A({ _06524_, _11451_, _tmp_1319, _tmp_1318 }), .Y(_06525_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37001_ ( .A({ _11452_, _tmp_1320[0] }), .Y(_11451_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37002_ ( .A({ _11462_, _11457_, _11455_, _11453_ }), .Y(_11452_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37003_ ( .A({ _11454_, _tmp_1320[33:31] }), .Y(_11453_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37004_ ( .A({ _tmp_1320[29:28], _tmp_1320[26], _tmp_1320[23] }), .Y(_11454_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37005_ ( .A({ _11456_, _tmp_1320[2:1] }), .Y(_11455_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37006_ ( .A(_tmp_1320[6:3]), .Y(_11456_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37007_ ( .A({ _11461_, _11460_, _11459_, _11458_ }), .Y(_11457_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37008_ ( .A(_tmp_1320[14:11]), .Y(_11458_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37009_ ( .A(_tmp_1320[10:7]), .Y(_11459_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37010_ ( .A(_tmp_1320[22:19]), .Y(_11460_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37011_ ( .A(_tmp_1320[18:15]), .Y(_11461_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37012_ ( .A({ _tmp_1320[30], _tmp_1320[27], _tmp_1320[25:24] }), .Y(_11462_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _37013_ ( .A({ _11451_, _06529_, _tmp_1309 }), .Y(_06526_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _37014_ ( .A({ _11452_, _tmp_1320[0], _06529_, _tmp_1309 }), .Y(_06527_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37015_ ( .A({ _06518_, _10839_ }), .Y(_06530_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37016_ ( .A({ _dataflow_slice_valid_6, _10838_ }), .Y(_06199_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37017_ ( .A({ _11463_, _06199_ }), .Y(_06531_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37018_ ( .A({ _tmp_14[0], _10840_, _tmp_14[33:32] }), .Y(_11463_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37019_ ( .A({ _11464_, _stream_matmul_29_sink_21_sink_waddr[1] }), .Y(_06532_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37020_ ( .A({ _stream_matmul_29_sink_21_sink_waddr[0], _11448_ }), .Y(_11464_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _37021_ ( .A({ _tmp_1321, _06529_ }), .Y(_tmp_1326) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37022_ ( .A({ _tmp_1329, _06529_, _tmp_1321 }), .Y(_06533_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37023_ ( .A({ _tmp_1328, _06529_, _tmp_1321 }), .Y(_06534_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37024_ ( .A({ _06524_, _11465_, _tmp_1331, _tmp_1330 }), .Y(_06535_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37025_ ( .A({ _11466_, _tmp_1332[0] }), .Y(_11465_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37026_ ( .A({ _11476_, _11471_, _11469_, _11467_ }), .Y(_11466_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37027_ ( .A({ _11468_, _tmp_1332[33:31] }), .Y(_11467_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37028_ ( .A({ _tmp_1332[29:28], _tmp_1332[26], _tmp_1332[23] }), .Y(_11468_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37029_ ( .A({ _11470_, _tmp_1332[2:1] }), .Y(_11469_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37030_ ( .A(_tmp_1332[6:3]), .Y(_11470_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37031_ ( .A({ _11475_, _11474_, _11473_, _11472_ }), .Y(_11471_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37032_ ( .A(_tmp_1332[14:11]), .Y(_11472_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37033_ ( .A(_tmp_1332[10:7]), .Y(_11473_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37034_ ( .A(_tmp_1332[22:19]), .Y(_11474_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37035_ ( .A(_tmp_1332[18:15]), .Y(_11475_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37036_ ( .A({ _tmp_1332[30], _tmp_1332[27], _tmp_1332[25:24] }), .Y(_11476_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _37037_ ( .A({ _11465_, _06529_, _tmp_1321 }), .Y(_06536_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _37038_ ( .A({ _11466_, _tmp_1332[0], _06529_, _tmp_1321 }), .Y(_06537_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37039_ ( .A({ _06518_, _10851_ }), .Y(_06538_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37040_ ( .A({ _dataflow_slice_valid_9, _10850_ }), .Y(_06202_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37041_ ( .A({ _11477_, _06202_ }), .Y(_06539_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37042_ ( .A({ _tmp_16[0], _10852_, _tmp_16[33:32] }), .Y(_11477_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37043_ ( .A({ _stream_matmul_29_sink_21_sink_waddr[1], _11447_ }), .Y(_06540_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _37044_ ( .A({ _tmp_1333, _06529_ }), .Y(_tmp_1338) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37045_ ( .A({ _tmp_1341, _06529_, _tmp_1333 }), .Y(_06541_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37046_ ( .A({ _tmp_1340, _06529_, _tmp_1333 }), .Y(_06542_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37047_ ( .A({ _06524_, _11478_, _tmp_1343, _tmp_1342 }), .Y(_06543_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37048_ ( .A({ _11479_, _tmp_1344[0] }), .Y(_11478_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37049_ ( .A({ _11489_, _11484_, _11482_, _11480_ }), .Y(_11479_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37050_ ( .A({ _11481_, _tmp_1344[33:31] }), .Y(_11480_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37051_ ( .A({ _tmp_1344[29:28], _tmp_1344[26], _tmp_1344[23] }), .Y(_11481_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37052_ ( .A({ _11483_, _tmp_1344[2:1] }), .Y(_11482_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37053_ ( .A(_tmp_1344[6:3]), .Y(_11483_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37054_ ( .A({ _11488_, _11487_, _11486_, _11485_ }), .Y(_11484_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37055_ ( .A(_tmp_1344[14:11]), .Y(_11485_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37056_ ( .A(_tmp_1344[10:7]), .Y(_11486_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37057_ ( .A(_tmp_1344[22:19]), .Y(_11487_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37058_ ( .A(_tmp_1344[18:15]), .Y(_11488_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37059_ ( .A({ _tmp_1344[30], _tmp_1344[27], _tmp_1344[25:24] }), .Y(_11489_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _37060_ ( .A({ _11478_, _06529_, _tmp_1333 }), .Y(_06544_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _37061_ ( .A({ _11479_, _tmp_1344[0], _06529_, _tmp_1333 }), .Y(_06545_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37062_ ( .A({ _06518_, _10863_ }), .Y(_06546_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37063_ ( .A({ _dataflow_slice_valid_12, _10862_ }), .Y(_06205_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37064_ ( .A({ _11490_, _06205_ }), .Y(_06547_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37065_ ( .A({ _tmp_18[0], _10864_, _tmp_18[33:32] }), .Y(_11490_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37066_ ( .A({ _stream_conv2d_16_source_6_source_ram_renable, _05891_ }), .Y(_tmp_472) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37067_ ( .A({ _stream_max_pool_serial_18_source_1_source_ram_renable, _05892_ }), .Y(_tmp_1035) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37068_ ( .A({ _stream_matmul_29_sink_21_sink_waddr[1], _11464_ }), .Y(_06548_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _37069_ ( .A({ _tmp_1345, _06529_ }), .Y(_tmp_1350) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37070_ ( .A({ _tmp_1353, _06529_, _tmp_1345 }), .Y(_06549_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37071_ ( .A({ _tmp_1352, _06529_, _tmp_1345 }), .Y(_06550_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37072_ ( .A({ _06524_, _11491_, _tmp_1355, _tmp_1354 }), .Y(_06551_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37073_ ( .A({ _11492_, _tmp_1356[0] }), .Y(_11491_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37074_ ( .A({ _11502_, _11497_, _11495_, _11493_ }), .Y(_11492_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37075_ ( .A({ _11494_, _tmp_1356[33:31] }), .Y(_11493_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37076_ ( .A({ _tmp_1356[29:28], _tmp_1356[26], _tmp_1356[23] }), .Y(_11494_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37077_ ( .A({ _11496_, _tmp_1356[2:1] }), .Y(_11495_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37078_ ( .A(_tmp_1356[6:3]), .Y(_11496_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37079_ ( .A({ _11501_, _11500_, _11499_, _11498_ }), .Y(_11497_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37080_ ( .A(_tmp_1356[14:11]), .Y(_11498_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37081_ ( .A(_tmp_1356[10:7]), .Y(_11499_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37082_ ( .A(_tmp_1356[22:19]), .Y(_11500_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37083_ ( .A(_tmp_1356[18:15]), .Y(_11501_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37084_ ( .A({ _tmp_1356[30], _tmp_1356[27], _tmp_1356[25:24] }), .Y(_11502_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _37085_ ( .A({ _11491_, _06529_, _tmp_1345 }), .Y(_06552_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _37086_ ( .A({ _11492_, _tmp_1356[0], _06529_, _tmp_1345 }), .Y(_06553_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37087_ ( .A({ _maxi_read_start, _11503_, _maxi_read_op_sel[1:0] }), .Y(_06554_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _37088_ ( .A({ _11347_, _maxi_read_op_sel[2], _maxi_read_op_sel[3] }), .Y(_11503_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37089_ ( .A({ _06554_, _11011_ }), .Y(_06555_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37090_ ( .A({ _dataflow_slice_valid_54, _11010_ }), .Y(_06244_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37091_ ( .A({ _dataflow_slice_valid_54, _11504_, _11010_ }), .Y(_06556_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37092_ ( .A({ _11506_, _11505_, _tmp_291[1:0] }), .Y(_11504_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37093_ ( .A(_tmp_291[9:6]), .Y(_11505_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37094_ ( .A(_tmp_291[5:2]), .Y(_11506_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37095_ ( .A({ _06100_, _06556_ }), .Y(_06557_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37096_ ( .A({ _06101_, _06244_ }), .Y(_06558_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37097_ ( .A({ _06102_, _06244_ }), .Y(_06559_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37098_ ( .A({ _06100_, _06244_ }), .Y(_06560_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37099_ ( .A({ _11507_, _06244_ }), .Y(_06561_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37100_ ( .A({ _tmp_292[0], _11012_, _tmp_292[33:32] }), .Y(_11507_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37101_ ( .A({ _maxi_read_start, _maxi_read_op_sel[1:0], _11503_ }), .Y(_06562_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37102_ ( .A({ _06562_, _11155_ }), .Y(_06563_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37103_ ( .A({ _dataflow_slice_valid_111, _11154_ }), .Y(_06280_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37104_ ( .A({ _11508_, _06280_ }), .Y(_06564_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37105_ ( .A({ _tmp_1124[0], _11156_, _tmp_1124[33:32] }), .Y(_11508_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37106_ ( .A({ _06554_, _11023_ }), .Y(_06565_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37107_ ( .A({ _dataflow_slice_valid_57, _11022_ }), .Y(_06247_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37108_ ( .A({ _dataflow_slice_valid_57, _11509_, _11022_ }), .Y(_06566_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37109_ ( .A({ _11511_, _11510_, _tmp_304[1:0] }), .Y(_11509_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37110_ ( .A(_tmp_304[9:6]), .Y(_11510_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37111_ ( .A(_tmp_304[5:2]), .Y(_11511_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37112_ ( .A({ _06103_, _06566_ }), .Y(_06567_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37113_ ( .A({ _06104_, _06247_ }), .Y(_06568_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37114_ ( .A({ _06105_, _06247_ }), .Y(_06569_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37115_ ( .A({ _06103_, _06247_ }), .Y(_06570_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37116_ ( .A({ _11512_, _06247_ }), .Y(_06571_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37117_ ( .A({ _tmp_305[0], _11024_, _tmp_305[33:32] }), .Y(_11512_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37118_ ( .A({ _06562_, _11167_ }), .Y(_06572_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37119_ ( .A({ _dataflow_slice_valid_114, _11166_ }), .Y(_06283_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37120_ ( .A({ _11513_, _06283_ }), .Y(_06573_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37121_ ( .A({ _tmp_1126[0], _11168_, _tmp_1126[33:32] }), .Y(_11513_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37122_ ( .A({ _06554_, _11035_ }), .Y(_06574_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37123_ ( .A({ _dataflow_slice_valid_60, _11034_ }), .Y(_06250_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37124_ ( .A({ _dataflow_slice_valid_60, _11514_, _11034_ }), .Y(_06575_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37125_ ( .A({ _11516_, _11515_, _tmp_317[1:0] }), .Y(_11514_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37126_ ( .A(_tmp_317[9:6]), .Y(_11515_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37127_ ( .A(_tmp_317[5:2]), .Y(_11516_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37128_ ( .A({ _06106_, _06575_ }), .Y(_06576_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37129_ ( .A({ _06107_, _06250_ }), .Y(_06577_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37130_ ( .A({ _06108_, _06250_ }), .Y(_06578_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37131_ ( .A({ _06106_, _06250_ }), .Y(_06579_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37132_ ( .A({ _11517_, _06250_ }), .Y(_06580_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37133_ ( .A({ _tmp_318[0], _11036_, _tmp_318[33:32] }), .Y(_11517_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37134_ ( .A({ _06562_, _11179_ }), .Y(_06581_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37135_ ( .A({ _dataflow_slice_valid_117, _11178_ }), .Y(_06286_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37136_ ( .A({ _11518_, _06286_ }), .Y(_06582_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37137_ ( .A({ _tmp_1128[0], _11180_, _tmp_1128[33:32] }), .Y(_11518_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37138_ ( .A({ _06554_, _11047_ }), .Y(_06583_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37139_ ( .A({ _dataflow_slice_valid_63, _11046_ }), .Y(_06253_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37140_ ( .A({ _dataflow_slice_valid_63, _11519_, _11046_ }), .Y(_06584_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37141_ ( .A({ _11521_, _11520_, _tmp_330[1:0] }), .Y(_11519_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37142_ ( .A(_tmp_330[9:6]), .Y(_11520_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37143_ ( .A(_tmp_330[5:2]), .Y(_11521_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37144_ ( .A({ _06109_, _06584_ }), .Y(_06585_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37145_ ( .A({ _06110_, _06253_ }), .Y(_06586_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37146_ ( .A({ _06111_, _06253_ }), .Y(_06587_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37147_ ( .A({ _06109_, _06253_ }), .Y(_06588_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37148_ ( .A({ _11522_, _06253_ }), .Y(_06589_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37149_ ( .A({ _tmp_331[0], _11048_, _tmp_331[33:32] }), .Y(_11522_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37150_ ( .A({ _stream_conv2d_16_source_19_source_ram_renable, _05893_ }), .Y(_tmp_503) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37151_ ( .A({ _06562_, _11191_ }), .Y(_06590_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37152_ ( .A({ _dataflow_slice_valid_120, _11190_ }), .Y(_06289_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37153_ ( .A({ _11523_, _06289_ }), .Y(_06591_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37154_ ( .A({ _tmp_1130[0], _11192_, _tmp_1130[33:32] }), .Y(_11523_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37155_ ( .A({ _stream_matmul_29_source_6_source_ram_renable, _05894_ }), .Y(_tmp_1178) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _37156_ ( .A({ _maxi_read_start, _11352_, _maxi_read_op_sel[0], _maxi_read_op_sel[1] }), .Y(_06592_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37157_ ( .A({ _06592_, _11299_ }), .Y(_06593_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37158_ ( .A({ _dataflow_slice_valid_149, _11298_ }), .Y(_06316_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37159_ ( .A({ _11524_, _06316_ }), .Y(_06594_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37160_ ( .A({ _tmp_1155[0], _11300_, _tmp_1155[33:32] }), .Y(_11524_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37161_ ( .A({ _06592_, _11311_ }), .Y(_06595_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37162_ ( .A({ _dataflow_slice_valid_152, _11310_ }), .Y(_06319_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37163_ ( .A({ _11525_, _06319_ }), .Y(_06596_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37164_ ( .A({ _tmp_1157[0], _11312_, _tmp_1157[33:32] }), .Y(_11525_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37165_ ( .A({ _06592_, _11323_ }), .Y(_06597_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37166_ ( .A({ _dataflow_slice_valid_155, _11322_ }), .Y(_06322_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37167_ ( .A({ _11526_, _06322_ }), .Y(_06598_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37168_ ( .A({ _tmp_1159[0], _11324_, _tmp_1159[33:32] }), .Y(_11526_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37169_ ( .A({ _stream_conv2d_16_source_20_source_ram_renable, _05895_ }), .Y(_tmp_513) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37170_ ( .A({ _06592_, _11335_ }), .Y(_06599_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37171_ ( .A({ _dataflow_slice_valid_158, _11334_ }), .Y(_06325_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37172_ ( .A({ _11527_, _06325_ }), .Y(_06600_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37173_ ( .A({ _tmp_1161[0], _11336_, _tmp_1161[33:32] }), .Y(_11527_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37174_ ( .A({ _stream_matmul_29_source_19_source_ram_renable, _05896_ }), .Y(_tmp_1209) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37175_ ( .A({ _stream_conv2d_16_source_21_source_ram_renable, _05897_ }), .Y(_tmp_523) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _37176_ ( .A({ _maxi_read_start, _11503_, _maxi_read_op_sel[0], _maxi_read_op_sel[1] }), .Y(_06601_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37177_ ( .A({ _06601_, _11059_ }), .Y(_06602_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37178_ ( .A({ _dataflow_slice_valid_67, _11058_ }), .Y(_06256_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37179_ ( .A({ _dataflow_slice_valid_67, _11528_, _11058_ }), .Y(_06603_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37180_ ( .A({ _11530_, _11529_, _tmp_348[1:0] }), .Y(_11528_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37181_ ( .A(_tmp_348[9:6]), .Y(_11529_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37182_ ( .A(_tmp_348[5:2]), .Y(_11530_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37183_ ( .A({ _06112_, _06603_ }), .Y(_06604_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37184_ ( .A({ _06113_, _06256_ }), .Y(_06605_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37185_ ( .A({ _06114_, _06256_ }), .Y(_06606_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37186_ ( .A({ _06112_, _06256_ }), .Y(_06607_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37187_ ( .A({ _11531_, _06256_ }), .Y(_06608_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37188_ ( .A({ _tmp_349[0], _11060_, _tmp_349[33:32] }), .Y(_11531_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37189_ ( .A({ _06601_, _11071_ }), .Y(_06609_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37190_ ( .A({ _dataflow_slice_valid_70, _11070_ }), .Y(_06259_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37191_ ( .A({ _dataflow_slice_valid_70, _11532_, _11070_ }), .Y(_06610_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37192_ ( .A({ _11534_, _11533_, _tmp_361[1:0] }), .Y(_11532_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37193_ ( .A(_tmp_361[9:6]), .Y(_11533_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37194_ ( .A(_tmp_361[5:2]), .Y(_11534_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37195_ ( .A({ _06115_, _06610_ }), .Y(_06611_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37196_ ( .A({ _06116_, _06259_ }), .Y(_06612_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37197_ ( .A({ _06117_, _06259_ }), .Y(_06613_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37198_ ( .A({ _06115_, _06259_ }), .Y(_06614_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37199_ ( .A({ _11535_, _06259_ }), .Y(_06615_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37200_ ( .A({ _tmp_362[0], _11072_, _tmp_362[33:32] }), .Y(_11535_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37201_ ( .A({ _06601_, _11083_ }), .Y(_06616_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37202_ ( .A({ _dataflow_slice_valid_73, _11082_ }), .Y(_06262_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37203_ ( .A({ _dataflow_slice_valid_73, _11536_, _11082_ }), .Y(_06617_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37204_ ( .A({ _11538_, _11537_, _tmp_374[1:0] }), .Y(_11536_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37205_ ( .A(_tmp_374[9:6]), .Y(_11537_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37206_ ( .A(_tmp_374[5:2]), .Y(_11538_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37207_ ( .A({ _06118_, _06617_ }), .Y(_06618_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37208_ ( .A({ _06119_, _06262_ }), .Y(_06619_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37209_ ( .A({ _06120_, _06262_ }), .Y(_06620_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37210_ ( .A({ _06118_, _06262_ }), .Y(_06621_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37211_ ( .A({ _11539_, _06262_ }), .Y(_06622_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37212_ ( .A({ _tmp_375[0], _11084_, _tmp_375[33:32] }), .Y(_11539_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37213_ ( .A({ _06601_, _11095_ }), .Y(_06623_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37214_ ( .A({ _dataflow_slice_valid_76, _11094_ }), .Y(_06265_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37215_ ( .A({ _dataflow_slice_valid_76, _11540_, _11094_ }), .Y(_06624_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37216_ ( .A({ _11542_, _11541_, _tmp_387[1:0] }), .Y(_11540_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37217_ ( .A(_tmp_387[9:6]), .Y(_11541_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37218_ ( .A(_tmp_387[5:2]), .Y(_11542_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37219_ ( .A({ _06121_, _06624_ }), .Y(_06625_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37220_ ( .A({ _06122_, _06265_ }), .Y(_06626_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37221_ ( .A({ _06123_, _06265_ }), .Y(_06627_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37222_ ( .A({ _06121_, _06265_ }), .Y(_06628_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37223_ ( .A({ _11543_, _06265_ }), .Y(_06629_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37224_ ( .A({ _tmp_388[0], _11096_, _tmp_388[33:32] }), .Y(_11543_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37225_ ( .A({ _stream_conv2d_16_source_22_source_ram_renable, _05898_ }), .Y(_tmp_533) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37226_ ( .A({ _stream_conv2d_16_source_23_source_ram_renable, _05899_ }), .Y(_tmp_543) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37227_ ( .A({ _stream_conv2d_16_source_24_source_ram_renable, _05900_ }), .Y(_tmp_553) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _37228_ ( .A({ _maxi_read_start, _maxi_read_op_sel[1], _11503_, _maxi_read_op_sel[0] }), .Y(_06630_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37229_ ( .A({ _06630_, _11107_ }), .Y(_06631_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37230_ ( .A({ _dataflow_slice_valid_80, _11106_ }), .Y(_06268_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37231_ ( .A({ _dataflow_slice_valid_80, _11544_, _11106_ }), .Y(_06632_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37232_ ( .A({ _11546_, _11545_, _tmp_405[1:0] }), .Y(_11544_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37233_ ( .A(_tmp_405[9:6]), .Y(_11545_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37234_ ( .A(_tmp_405[5:2]), .Y(_11546_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37235_ ( .A({ _06124_, _06632_ }), .Y(_06633_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37236_ ( .A({ _06125_, _06268_ }), .Y(_06634_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37237_ ( .A({ _06126_, _06268_ }), .Y(_06635_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37238_ ( .A({ _06124_, _06268_ }), .Y(_06636_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37239_ ( .A({ _11547_, _06268_ }), .Y(_06637_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37240_ ( .A({ _tmp_406[0], _11108_, _tmp_406[33:32] }), .Y(_11547_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37241_ ( .A({ _06630_, _11119_ }), .Y(_06638_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37242_ ( .A({ _dataflow_slice_valid_83, _11118_ }), .Y(_06271_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37243_ ( .A({ _dataflow_slice_valid_83, _11548_, _11118_ }), .Y(_06639_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37244_ ( .A({ _11550_, _11549_, _tmp_418[1:0] }), .Y(_11548_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37245_ ( .A(_tmp_418[9:6]), .Y(_11549_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37246_ ( .A(_tmp_418[5:2]), .Y(_11550_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37247_ ( .A({ _06127_, _06639_ }), .Y(_06640_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37248_ ( .A({ _06128_, _06271_ }), .Y(_06641_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37249_ ( .A({ _06129_, _06271_ }), .Y(_06642_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37250_ ( .A({ _06127_, _06271_ }), .Y(_06643_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37251_ ( .A({ _11551_, _06271_ }), .Y(_06644_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37252_ ( .A({ _tmp_419[0], _11120_, _tmp_419[33:32] }), .Y(_11551_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37253_ ( .A({ _06630_, _11131_ }), .Y(_06645_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37254_ ( .A({ _dataflow_slice_valid_86, _11130_ }), .Y(_06274_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37255_ ( .A({ _dataflow_slice_valid_86, _11552_, _11130_ }), .Y(_06646_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37256_ ( .A({ _11554_, _11553_, _tmp_431[1:0] }), .Y(_11552_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37257_ ( .A(_tmp_431[9:6]), .Y(_11553_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37258_ ( .A(_tmp_431[5:2]), .Y(_11554_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37259_ ( .A({ _06130_, _06646_ }), .Y(_06647_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37260_ ( .A({ _06131_, _06274_ }), .Y(_06648_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37261_ ( .A({ _06132_, _06274_ }), .Y(_06649_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37262_ ( .A({ _06130_, _06274_ }), .Y(_06650_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37263_ ( .A({ _11555_, _06274_ }), .Y(_06651_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37264_ ( .A({ _tmp_432[0], _11132_, _tmp_432[33:32] }), .Y(_11555_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37265_ ( .A({ _06630_, _11143_ }), .Y(_06652_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37266_ ( .A({ _dataflow_slice_valid_89, _11142_ }), .Y(_06277_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37267_ ( .A({ _dataflow_slice_valid_89, _11556_, _11142_ }), .Y(_06653_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37268_ ( .A({ _11558_, _11557_, _tmp_444[1:0] }), .Y(_11556_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37269_ ( .A(_tmp_444[9:6]), .Y(_11557_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37270_ ( .A(_tmp_444[5:2]), .Y(_11558_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37271_ ( .A({ _06133_, _06653_ }), .Y(_06654_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37272_ ( .A({ _06134_, _06277_ }), .Y(_06655_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37273_ ( .A({ _06135_, _06277_ }), .Y(_06656_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37274_ ( .A({ _06133_, _06277_ }), .Y(_06657_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37275_ ( .A({ _11559_, _06277_ }), .Y(_06658_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37276_ ( .A({ _tmp_445[0], _11144_, _tmp_445[33:32] }), .Y(_11559_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37277_ ( .A({ _stream_conv2d_16_source_25_source_ram_renable, _05901_ }), .Y(_tmp_563) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37278_ ( .A({ _stream_conv2d_16_source_26_source_ram_renable, _05902_ }), .Y(_tmp_573) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37279_ ( .A({ _stream_conv2d_16_source_27_source_ram_renable, _05903_ }), .Y(_tmp_583) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37280_ ( .A({ _11560_, _stream_conv2d_16_sink_37_sink_waddr[1] }), .Y(_06659_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37281_ ( .A({ _11561_, _stream_conv2d_16_sink_37_sink_waddr[0] }), .Y(_11560_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37282_ ( .A({ _11562_, _stream_conv2d_16_sink_37_sink_ram_sel[7:6] }), .Y(_11561_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37283_ ( .A({ _stream_conv2d_16_sink_37_sink_ram_sel[4], _stream_conv2d_16_sink_37_sink_ram_sel[2], _stream_conv2d_16_sink_37_sink_ram_sel[0], _11563_ }), .Y(_11562_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37284_ ( .A({ _stream_conv2d_16_sink_37_sink_wenable, _stream_conv2d_16_sink_37_sink_ram_sel[5], _stream_conv2d_16_sink_37_sink_ram_sel[3], _stream_conv2d_16_sink_37_sink_ram_sel[1] }), .Y(_11563_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _37285_ ( .A({ _tmp_971, _06667_ }), .Y(_tmp_976) );
  \$lut  #( .LUT(16'h8f00), .WIDTH(4) ) _37286_ ( .A({ _06666_, _dataflow_cat_valid_98, _10819_, _10820_ }), .Y(_06667_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37287_ ( .A({ _tmp_1007, _tmp_995, _tmp_983, _tmp_971 }), .Y(_06666_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37288_ ( .A({ _tmp_979, _06667_, _tmp_971 }), .Y(_06660_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37289_ ( .A({ _tmp_978, _06667_, _tmp_971 }), .Y(_06661_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37290_ ( .A({ _maxi_write_start, _10820_ }), .Y(_06662_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37291_ ( .A({ _06662_, _11564_, _tmp_981, _tmp_980 }), .Y(_06663_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37292_ ( .A({ _11565_, _tmp_982[0] }), .Y(_11564_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37293_ ( .A({ _11575_, _11570_, _11568_, _11566_ }), .Y(_11565_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37294_ ( .A({ _11567_, _tmp_982[33:31] }), .Y(_11566_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37295_ ( .A({ _tmp_982[29:28], _tmp_982[26], _tmp_982[23] }), .Y(_11567_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37296_ ( .A({ _11569_, _tmp_982[2:1] }), .Y(_11568_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37297_ ( .A(_tmp_982[6:3]), .Y(_11569_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37298_ ( .A({ _11574_, _11573_, _11572_, _11571_ }), .Y(_11570_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37299_ ( .A(_tmp_982[14:11]), .Y(_11571_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37300_ ( .A(_tmp_982[10:7]), .Y(_11572_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37301_ ( .A(_tmp_982[22:19]), .Y(_11573_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37302_ ( .A(_tmp_982[18:15]), .Y(_11574_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37303_ ( .A({ _tmp_982[30], _tmp_982[27], _tmp_982[25:24] }), .Y(_11575_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _37304_ ( .A({ _11564_, _06667_, _tmp_971 }), .Y(_06664_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _37305_ ( .A({ _11565_, _tmp_982[0], _06667_, _tmp_971 }), .Y(_06665_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37306_ ( .A({ _11576_, _stream_conv2d_16_sink_37_sink_waddr[1] }), .Y(_06668_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37307_ ( .A({ _stream_conv2d_16_sink_37_sink_waddr[0], _11561_ }), .Y(_11576_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _37308_ ( .A({ _tmp_983, _06667_ }), .Y(_tmp_988) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37309_ ( .A({ _tmp_991, _06667_, _tmp_983 }), .Y(_06669_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37310_ ( .A({ _tmp_990, _06667_, _tmp_983 }), .Y(_06670_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37311_ ( .A({ _06662_, _11577_, _tmp_993, _tmp_992 }), .Y(_06671_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37312_ ( .A({ _11578_, _tmp_994[0] }), .Y(_11577_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37313_ ( .A({ _11588_, _11583_, _11581_, _11579_ }), .Y(_11578_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37314_ ( .A({ _11580_, _tmp_994[33:31] }), .Y(_11579_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37315_ ( .A({ _tmp_994[29:28], _tmp_994[26], _tmp_994[23] }), .Y(_11580_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37316_ ( .A({ _11582_, _tmp_994[2:1] }), .Y(_11581_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37317_ ( .A(_tmp_994[6:3]), .Y(_11582_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37318_ ( .A({ _11587_, _11586_, _11585_, _11584_ }), .Y(_11583_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37319_ ( .A(_tmp_994[14:11]), .Y(_11584_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37320_ ( .A(_tmp_994[10:7]), .Y(_11585_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37321_ ( .A(_tmp_994[22:19]), .Y(_11586_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37322_ ( .A(_tmp_994[18:15]), .Y(_11587_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37323_ ( .A({ _tmp_994[30], _tmp_994[27], _tmp_994[25:24] }), .Y(_11588_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _37324_ ( .A({ _11577_, _06667_, _tmp_983 }), .Y(_06672_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _37325_ ( .A({ _11578_, _tmp_994[0], _06667_, _tmp_983 }), .Y(_06673_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37326_ ( .A({ _stream_conv2d_16_sink_37_sink_waddr[1], _11560_ }), .Y(_06674_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _37327_ ( .A({ _tmp_995, _06667_ }), .Y(_tmp_1000) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37328_ ( .A({ _tmp_1003, _06667_, _tmp_995 }), .Y(_06675_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37329_ ( .A({ _tmp_1002, _06667_, _tmp_995 }), .Y(_06676_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37330_ ( .A({ _06662_, _11589_, _tmp_1005, _tmp_1004 }), .Y(_06677_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37331_ ( .A({ _11590_, _tmp_1006[0] }), .Y(_11589_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37332_ ( .A({ _11600_, _11595_, _11593_, _11591_ }), .Y(_11590_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37333_ ( .A({ _11592_, _tmp_1006[33:31] }), .Y(_11591_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37334_ ( .A({ _tmp_1006[29:28], _tmp_1006[26], _tmp_1006[23] }), .Y(_11592_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37335_ ( .A({ _11594_, _tmp_1006[2:1] }), .Y(_11593_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37336_ ( .A(_tmp_1006[6:3]), .Y(_11594_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37337_ ( .A({ _11599_, _11598_, _11597_, _11596_ }), .Y(_11595_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37338_ ( .A(_tmp_1006[14:11]), .Y(_11596_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37339_ ( .A(_tmp_1006[10:7]), .Y(_11597_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37340_ ( .A(_tmp_1006[22:19]), .Y(_11598_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37341_ ( .A(_tmp_1006[18:15]), .Y(_11599_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37342_ ( .A({ _tmp_1006[30], _tmp_1006[27], _tmp_1006[25:24] }), .Y(_11600_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _37343_ ( .A({ _11589_, _06667_, _tmp_995 }), .Y(_06678_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _37344_ ( .A({ _11590_, _tmp_1006[0], _06667_, _tmp_995 }), .Y(_06679_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37345_ ( .A({ _stream_conv2d_16_sink_37_sink_waddr[1], _11576_ }), .Y(_06680_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _37346_ ( .A({ _tmp_1007, _06667_ }), .Y(_tmp_1012) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37347_ ( .A({ _tmp_1015, _06667_, _tmp_1007 }), .Y(_06681_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _37348_ ( .A({ _tmp_1014, _06667_, _tmp_1007 }), .Y(_06682_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37349_ ( .A({ _06662_, _11601_, _tmp_1017, _tmp_1016 }), .Y(_06683_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37350_ ( .A({ _11602_, _tmp_1018[0] }), .Y(_11601_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37351_ ( .A({ _11612_, _11607_, _11605_, _11603_ }), .Y(_11602_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37352_ ( .A({ _11604_, _tmp_1018[33:31] }), .Y(_11603_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37353_ ( .A({ _tmp_1018[29:28], _tmp_1018[26], _tmp_1018[23] }), .Y(_11604_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37354_ ( .A({ _11606_, _tmp_1018[2:1] }), .Y(_11605_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37355_ ( .A(_tmp_1018[6:3]), .Y(_11606_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37356_ ( .A({ _11611_, _11610_, _11609_, _11608_ }), .Y(_11607_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37357_ ( .A(_tmp_1018[14:11]), .Y(_11608_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37358_ ( .A(_tmp_1018[10:7]), .Y(_11609_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37359_ ( .A(_tmp_1018[22:19]), .Y(_11610_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37360_ ( .A(_tmp_1018[18:15]), .Y(_11611_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37361_ ( .A({ _tmp_1018[30], _tmp_1018[27], _tmp_1018[25:24] }), .Y(_11612_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _37362_ ( .A({ _11601_, _06667_, _tmp_1007 }), .Y(_06684_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _37363_ ( .A({ _11602_, _tmp_1018[0], _06667_, _tmp_1007 }), .Y(_06685_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37364_ ( .A({ _11613_, _05987_ }), .Y(_06687_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37365_ ( .A({ _11623_, _11622_, _11621_, _11614_ }), .Y(_11613_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37366_ ( .A({ _11620_, _11615_, _source_stream_conv2d_16_source_6_pat_count_0[1:0] }), .Y(_11614_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37367_ ( .A({ _11619_, _11618_, _11617_, _11616_ }), .Y(_11615_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37368_ ( .A(_source_stream_conv2d_16_source_6_pat_count_0[13:10]), .Y(_11616_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37369_ ( .A(_source_stream_conv2d_16_source_6_pat_count_0[9:6]), .Y(_11617_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37370_ ( .A(_source_stream_conv2d_16_source_6_pat_count_0[21:18]), .Y(_11618_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37371_ ( .A(_source_stream_conv2d_16_source_6_pat_count_0[17:14]), .Y(_11619_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37372_ ( .A(_source_stream_conv2d_16_source_6_pat_count_0[5:2]), .Y(_11620_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _37373_ ( .A(_source_stream_conv2d_16_source_6_pat_count_0[32:30]), .Y(_11621_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37374_ ( .A(_source_stream_conv2d_16_source_6_pat_count_0[29:26]), .Y(_11622_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37375_ ( .A(_source_stream_conv2d_16_source_6_pat_count_0[25:22]), .Y(_11623_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37376_ ( .A({ _11624_, _06687_ }), .Y(_06688_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37377_ ( .A({ _11634_, _11632_, _11625_ }), .Y(_11624_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37378_ ( .A({ _11631_, _11626_, _source_stream_conv2d_16_source_6_pat_count_1[1:0] }), .Y(_11625_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37379_ ( .A({ _11630_, _11629_, _11628_, _11627_ }), .Y(_11626_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37380_ ( .A(_source_stream_conv2d_16_source_6_pat_count_1[13:10]), .Y(_11627_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37381_ ( .A(_source_stream_conv2d_16_source_6_pat_count_1[9:6]), .Y(_11628_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37382_ ( .A(_source_stream_conv2d_16_source_6_pat_count_1[21:18]), .Y(_11629_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37383_ ( .A(_source_stream_conv2d_16_source_6_pat_count_1[17:14]), .Y(_11630_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37384_ ( .A(_source_stream_conv2d_16_source_6_pat_count_1[5:2]), .Y(_11631_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37385_ ( .A({ _11633_, _source_stream_conv2d_16_source_6_pat_count_1[32:30] }), .Y(_11632_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37386_ ( .A({ _source_stream_conv2d_16_source_6_pat_count_1[28:27], _source_stream_conv2d_16_source_6_pat_count_1[25], _source_stream_conv2d_16_source_6_pat_count_1[22] }), .Y(_11633_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37387_ ( .A({ _source_stream_conv2d_16_source_6_pat_count_1[29], _source_stream_conv2d_16_source_6_pat_count_1[26], _source_stream_conv2d_16_source_6_pat_count_1[24:23] }), .Y(_11634_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37388_ ( .A({ _11635_, _11624_, _06687_ }), .Y(_06689_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37389_ ( .A({ _11645_, _11640_, _11638_, _11636_ }), .Y(_11635_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37390_ ( .A({ _11637_, _source_stream_conv2d_16_source_6_pat_count_2[32:30] }), .Y(_11636_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37391_ ( .A({ _source_stream_conv2d_16_source_6_pat_count_2[28:27], _source_stream_conv2d_16_source_6_pat_count_2[25], _source_stream_conv2d_16_source_6_pat_count_2[22] }), .Y(_11637_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37392_ ( .A({ _11639_, _source_stream_conv2d_16_source_6_pat_count_2[1:0] }), .Y(_11638_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37393_ ( .A(_source_stream_conv2d_16_source_6_pat_count_2[5:2]), .Y(_11639_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37394_ ( .A({ _11644_, _11643_, _11642_, _11641_ }), .Y(_11640_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37395_ ( .A(_source_stream_conv2d_16_source_6_pat_count_2[13:10]), .Y(_11641_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37396_ ( .A(_source_stream_conv2d_16_source_6_pat_count_2[9:6]), .Y(_11642_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37397_ ( .A(_source_stream_conv2d_16_source_6_pat_count_2[21:18]), .Y(_11643_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37398_ ( .A(_source_stream_conv2d_16_source_6_pat_count_2[17:14]), .Y(_11644_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37399_ ( .A({ _source_stream_conv2d_16_source_6_pat_count_2[29], _source_stream_conv2d_16_source_6_pat_count_2[26], _source_stream_conv2d_16_source_6_pat_count_2[24:23] }), .Y(_11645_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37400_ ( .A({ _06837_, _05987_ }), .Y(_06690_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37401_ ( .A({ _11646_, _11624_, _11613_ }), .Y(_06837_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37402_ ( .A({ _11656_, _11654_, _11647_, _11635_ }), .Y(_11646_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37403_ ( .A({ _11653_, _11648_, _source_stream_conv2d_16_source_6_pat_count_3[1:0] }), .Y(_11647_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37404_ ( .A({ _11652_, _11651_, _11650_, _11649_ }), .Y(_11648_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37405_ ( .A(_source_stream_conv2d_16_source_6_pat_count_3[13:10]), .Y(_11649_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37406_ ( .A(_source_stream_conv2d_16_source_6_pat_count_3[9:6]), .Y(_11650_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37407_ ( .A(_source_stream_conv2d_16_source_6_pat_count_3[21:18]), .Y(_11651_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37408_ ( .A(_source_stream_conv2d_16_source_6_pat_count_3[17:14]), .Y(_11652_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37409_ ( .A(_source_stream_conv2d_16_source_6_pat_count_3[5:2]), .Y(_11653_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37410_ ( .A({ _11655_, _source_stream_conv2d_16_source_6_pat_count_3[32:30] }), .Y(_11654_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37411_ ( .A({ _source_stream_conv2d_16_source_6_pat_count_3[28:27], _source_stream_conv2d_16_source_6_pat_count_3[25], _source_stream_conv2d_16_source_6_pat_count_3[22] }), .Y(_11655_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37412_ ( .A({ _source_stream_conv2d_16_source_6_pat_count_3[29], _source_stream_conv2d_16_source_6_pat_count_3[26], _source_stream_conv2d_16_source_6_pat_count_3[24:23] }), .Y(_11656_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37413_ ( .A({ _11657_, _05986_ }), .Y(_06692_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37414_ ( .A({ _11667_, _11662_, _11660_, _11658_ }), .Y(_11657_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37415_ ( .A({ _11659_, _source_stream_conv2d_16_source_8_pat_count_0[32:30] }), .Y(_11658_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37416_ ( .A({ _source_stream_conv2d_16_source_8_pat_count_0[28:27], _source_stream_conv2d_16_source_8_pat_count_0[25], _source_stream_conv2d_16_source_8_pat_count_0[22] }), .Y(_11659_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37417_ ( .A({ _11661_, _source_stream_conv2d_16_source_8_pat_count_0[1:0] }), .Y(_11660_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37418_ ( .A(_source_stream_conv2d_16_source_8_pat_count_0[5:2]), .Y(_11661_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37419_ ( .A({ _11666_, _11665_, _11664_, _11663_ }), .Y(_11662_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37420_ ( .A(_source_stream_conv2d_16_source_8_pat_count_0[13:10]), .Y(_11663_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37421_ ( .A(_source_stream_conv2d_16_source_8_pat_count_0[9:6]), .Y(_11664_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37422_ ( .A(_source_stream_conv2d_16_source_8_pat_count_0[21:18]), .Y(_11665_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37423_ ( .A(_source_stream_conv2d_16_source_8_pat_count_0[17:14]), .Y(_11666_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37424_ ( .A({ _source_stream_conv2d_16_source_8_pat_count_0[29], _source_stream_conv2d_16_source_8_pat_count_0[26], _source_stream_conv2d_16_source_8_pat_count_0[24:23] }), .Y(_11667_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37425_ ( .A({ _11668_, _06692_ }), .Y(_06693_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37426_ ( .A({ _11678_, _11676_, _11669_ }), .Y(_11668_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37427_ ( .A({ _11675_, _11670_, _source_stream_conv2d_16_source_8_pat_count_1[1:0] }), .Y(_11669_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37428_ ( .A({ _11674_, _11673_, _11672_, _11671_ }), .Y(_11670_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37429_ ( .A(_source_stream_conv2d_16_source_8_pat_count_1[13:10]), .Y(_11671_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37430_ ( .A(_source_stream_conv2d_16_source_8_pat_count_1[9:6]), .Y(_11672_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37431_ ( .A(_source_stream_conv2d_16_source_8_pat_count_1[21:18]), .Y(_11673_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37432_ ( .A(_source_stream_conv2d_16_source_8_pat_count_1[17:14]), .Y(_11674_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37433_ ( .A(_source_stream_conv2d_16_source_8_pat_count_1[5:2]), .Y(_11675_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37434_ ( .A({ _11677_, _source_stream_conv2d_16_source_8_pat_count_1[32:30] }), .Y(_11676_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37435_ ( .A({ _source_stream_conv2d_16_source_8_pat_count_1[28:27], _source_stream_conv2d_16_source_8_pat_count_1[25], _source_stream_conv2d_16_source_8_pat_count_1[22] }), .Y(_11677_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37436_ ( .A({ _source_stream_conv2d_16_source_8_pat_count_1[29], _source_stream_conv2d_16_source_8_pat_count_1[26], _source_stream_conv2d_16_source_8_pat_count_1[24:23] }), .Y(_11678_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37437_ ( .A({ _11679_, _11668_, _06692_ }), .Y(_06694_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37438_ ( .A({ _11689_, _11684_, _11682_, _11680_ }), .Y(_11679_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37439_ ( .A({ _11681_, _source_stream_conv2d_16_source_8_pat_count_2[32:30] }), .Y(_11680_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37440_ ( .A({ _source_stream_conv2d_16_source_8_pat_count_2[28:27], _source_stream_conv2d_16_source_8_pat_count_2[25], _source_stream_conv2d_16_source_8_pat_count_2[22] }), .Y(_11681_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37441_ ( .A({ _11683_, _source_stream_conv2d_16_source_8_pat_count_2[1:0] }), .Y(_11682_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37442_ ( .A(_source_stream_conv2d_16_source_8_pat_count_2[5:2]), .Y(_11683_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37443_ ( .A({ _11688_, _11687_, _11686_, _11685_ }), .Y(_11684_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37444_ ( .A(_source_stream_conv2d_16_source_8_pat_count_2[13:10]), .Y(_11685_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37445_ ( .A(_source_stream_conv2d_16_source_8_pat_count_2[9:6]), .Y(_11686_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37446_ ( .A(_source_stream_conv2d_16_source_8_pat_count_2[21:18]), .Y(_11687_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37447_ ( .A(_source_stream_conv2d_16_source_8_pat_count_2[17:14]), .Y(_11688_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37448_ ( .A({ _source_stream_conv2d_16_source_8_pat_count_2[29], _source_stream_conv2d_16_source_8_pat_count_2[26], _source_stream_conv2d_16_source_8_pat_count_2[24:23] }), .Y(_11689_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37449_ ( .A({ _06838_, _05986_ }), .Y(_06695_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37450_ ( .A({ _11690_, _11679_, _11657_, _11668_ }), .Y(_06838_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37451_ ( .A({ _11700_, _11695_, _11693_, _11691_ }), .Y(_11690_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37452_ ( .A({ _11692_, _source_stream_conv2d_16_source_8_pat_count_3[32:30] }), .Y(_11691_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37453_ ( .A({ _source_stream_conv2d_16_source_8_pat_count_3[28:27], _source_stream_conv2d_16_source_8_pat_count_3[25], _source_stream_conv2d_16_source_8_pat_count_3[22] }), .Y(_11692_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37454_ ( .A({ _11694_, _source_stream_conv2d_16_source_8_pat_count_3[1:0] }), .Y(_11693_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37455_ ( .A(_source_stream_conv2d_16_source_8_pat_count_3[5:2]), .Y(_11694_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37456_ ( .A({ _11699_, _11698_, _11697_, _11696_ }), .Y(_11695_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37457_ ( .A(_source_stream_conv2d_16_source_8_pat_count_3[13:10]), .Y(_11696_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37458_ ( .A(_source_stream_conv2d_16_source_8_pat_count_3[9:6]), .Y(_11697_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37459_ ( .A(_source_stream_conv2d_16_source_8_pat_count_3[21:18]), .Y(_11698_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37460_ ( .A(_source_stream_conv2d_16_source_8_pat_count_3[17:14]), .Y(_11699_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37461_ ( .A({ _source_stream_conv2d_16_source_8_pat_count_3[29], _source_stream_conv2d_16_source_8_pat_count_3[26], _source_stream_conv2d_16_source_8_pat_count_3[24:23] }), .Y(_11700_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37462_ ( .A({ _11701_, _05983_ }), .Y(_06697_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37463_ ( .A({ _11711_, _11710_, _11709_, _11702_ }), .Y(_11701_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37464_ ( .A({ _11708_, _11703_, _source_stream_conv2d_16_source_19_pat_count_0[1:0] }), .Y(_11702_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37465_ ( .A({ _11707_, _11706_, _11705_, _11704_ }), .Y(_11703_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37466_ ( .A(_source_stream_conv2d_16_source_19_pat_count_0[13:10]), .Y(_11704_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37467_ ( .A(_source_stream_conv2d_16_source_19_pat_count_0[9:6]), .Y(_11705_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37468_ ( .A(_source_stream_conv2d_16_source_19_pat_count_0[21:18]), .Y(_11706_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37469_ ( .A(_source_stream_conv2d_16_source_19_pat_count_0[17:14]), .Y(_11707_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37470_ ( .A(_source_stream_conv2d_16_source_19_pat_count_0[5:2]), .Y(_11708_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _37471_ ( .A(_source_stream_conv2d_16_source_19_pat_count_0[32:30]), .Y(_11709_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37472_ ( .A(_source_stream_conv2d_16_source_19_pat_count_0[29:26]), .Y(_11710_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37473_ ( .A(_source_stream_conv2d_16_source_19_pat_count_0[25:22]), .Y(_11711_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37474_ ( .A({ _11712_, _06697_ }), .Y(_06698_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37475_ ( .A({ _11722_, _11720_, _11713_ }), .Y(_11712_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37476_ ( .A({ _11719_, _11714_, _source_stream_conv2d_16_source_19_pat_count_1[1:0] }), .Y(_11713_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37477_ ( .A({ _11718_, _11717_, _11716_, _11715_ }), .Y(_11714_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37478_ ( .A(_source_stream_conv2d_16_source_19_pat_count_1[13:10]), .Y(_11715_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37479_ ( .A(_source_stream_conv2d_16_source_19_pat_count_1[9:6]), .Y(_11716_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37480_ ( .A(_source_stream_conv2d_16_source_19_pat_count_1[21:18]), .Y(_11717_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37481_ ( .A(_source_stream_conv2d_16_source_19_pat_count_1[17:14]), .Y(_11718_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37482_ ( .A(_source_stream_conv2d_16_source_19_pat_count_1[5:2]), .Y(_11719_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37483_ ( .A({ _11721_, _source_stream_conv2d_16_source_19_pat_count_1[32:30] }), .Y(_11720_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37484_ ( .A({ _source_stream_conv2d_16_source_19_pat_count_1[28:27], _source_stream_conv2d_16_source_19_pat_count_1[25], _source_stream_conv2d_16_source_19_pat_count_1[22] }), .Y(_11721_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37485_ ( .A({ _source_stream_conv2d_16_source_19_pat_count_1[29], _source_stream_conv2d_16_source_19_pat_count_1[26], _source_stream_conv2d_16_source_19_pat_count_1[24:23] }), .Y(_11722_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37486_ ( .A({ _11723_, _11712_, _06697_ }), .Y(_06699_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37487_ ( .A({ _11733_, _11728_, _11726_, _11724_ }), .Y(_11723_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37488_ ( .A({ _11725_, _source_stream_conv2d_16_source_19_pat_count_2[32:30] }), .Y(_11724_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37489_ ( .A({ _source_stream_conv2d_16_source_19_pat_count_2[28:27], _source_stream_conv2d_16_source_19_pat_count_2[25], _source_stream_conv2d_16_source_19_pat_count_2[22] }), .Y(_11725_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37490_ ( .A({ _11727_, _source_stream_conv2d_16_source_19_pat_count_2[1:0] }), .Y(_11726_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37491_ ( .A(_source_stream_conv2d_16_source_19_pat_count_2[5:2]), .Y(_11727_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37492_ ( .A({ _11732_, _11731_, _11730_, _11729_ }), .Y(_11728_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37493_ ( .A(_source_stream_conv2d_16_source_19_pat_count_2[13:10]), .Y(_11729_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37494_ ( .A(_source_stream_conv2d_16_source_19_pat_count_2[9:6]), .Y(_11730_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37495_ ( .A(_source_stream_conv2d_16_source_19_pat_count_2[21:18]), .Y(_11731_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37496_ ( .A(_source_stream_conv2d_16_source_19_pat_count_2[17:14]), .Y(_11732_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37497_ ( .A({ _source_stream_conv2d_16_source_19_pat_count_2[29], _source_stream_conv2d_16_source_19_pat_count_2[26], _source_stream_conv2d_16_source_19_pat_count_2[24:23] }), .Y(_11733_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37498_ ( .A({ _06839_, _05983_ }), .Y(_06700_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37499_ ( .A({ _11734_, _11723_, _11712_, _11701_ }), .Y(_06839_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37500_ ( .A({ _11744_, _11739_, _11737_, _11735_ }), .Y(_11734_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37501_ ( .A({ _11736_, _source_stream_conv2d_16_source_19_pat_count_3[32:30] }), .Y(_11735_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37502_ ( .A({ _source_stream_conv2d_16_source_19_pat_count_3[28:27], _source_stream_conv2d_16_source_19_pat_count_3[25], _source_stream_conv2d_16_source_19_pat_count_3[22] }), .Y(_11736_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37503_ ( .A({ _11738_, _source_stream_conv2d_16_source_19_pat_count_3[1:0] }), .Y(_11737_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37504_ ( .A(_source_stream_conv2d_16_source_19_pat_count_3[5:2]), .Y(_11738_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37505_ ( .A({ _11743_, _11742_, _11741_, _11740_ }), .Y(_11739_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37506_ ( .A(_source_stream_conv2d_16_source_19_pat_count_3[13:10]), .Y(_11740_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37507_ ( .A(_source_stream_conv2d_16_source_19_pat_count_3[9:6]), .Y(_11741_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37508_ ( .A(_source_stream_conv2d_16_source_19_pat_count_3[21:18]), .Y(_11742_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37509_ ( .A(_source_stream_conv2d_16_source_19_pat_count_3[17:14]), .Y(_11743_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37510_ ( .A({ _source_stream_conv2d_16_source_19_pat_count_3[29], _source_stream_conv2d_16_source_19_pat_count_3[26], _source_stream_conv2d_16_source_19_pat_count_3[24:23] }), .Y(_11744_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37511_ ( .A({ _11745_, _05982_ }), .Y(_06702_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37512_ ( .A({ _11755_, _11754_, _11753_, _11746_ }), .Y(_11745_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37513_ ( .A({ _11752_, _11747_, _source_stream_conv2d_16_source_20_pat_count_0[1:0] }), .Y(_11746_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37514_ ( .A({ _11751_, _11750_, _11749_, _11748_ }), .Y(_11747_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37515_ ( .A(_source_stream_conv2d_16_source_20_pat_count_0[13:10]), .Y(_11748_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37516_ ( .A(_source_stream_conv2d_16_source_20_pat_count_0[9:6]), .Y(_11749_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37517_ ( .A(_source_stream_conv2d_16_source_20_pat_count_0[21:18]), .Y(_11750_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37518_ ( .A(_source_stream_conv2d_16_source_20_pat_count_0[17:14]), .Y(_11751_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37519_ ( .A(_source_stream_conv2d_16_source_20_pat_count_0[5:2]), .Y(_11752_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _37520_ ( .A(_source_stream_conv2d_16_source_20_pat_count_0[32:30]), .Y(_11753_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37521_ ( .A(_source_stream_conv2d_16_source_20_pat_count_0[29:26]), .Y(_11754_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37522_ ( .A(_source_stream_conv2d_16_source_20_pat_count_0[25:22]), .Y(_11755_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37523_ ( .A({ _11756_, _06702_ }), .Y(_06703_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37524_ ( .A({ _11766_, _11764_, _11757_ }), .Y(_11756_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37525_ ( .A({ _11763_, _11758_, _source_stream_conv2d_16_source_20_pat_count_1[1:0] }), .Y(_11757_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37526_ ( .A({ _11762_, _11761_, _11760_, _11759_ }), .Y(_11758_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37527_ ( .A(_source_stream_conv2d_16_source_20_pat_count_1[13:10]), .Y(_11759_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37528_ ( .A(_source_stream_conv2d_16_source_20_pat_count_1[9:6]), .Y(_11760_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37529_ ( .A(_source_stream_conv2d_16_source_20_pat_count_1[21:18]), .Y(_11761_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37530_ ( .A(_source_stream_conv2d_16_source_20_pat_count_1[17:14]), .Y(_11762_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37531_ ( .A(_source_stream_conv2d_16_source_20_pat_count_1[5:2]), .Y(_11763_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37532_ ( .A({ _11765_, _source_stream_conv2d_16_source_20_pat_count_1[32:30] }), .Y(_11764_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37533_ ( .A({ _source_stream_conv2d_16_source_20_pat_count_1[28:27], _source_stream_conv2d_16_source_20_pat_count_1[25], _source_stream_conv2d_16_source_20_pat_count_1[22] }), .Y(_11765_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37534_ ( .A({ _source_stream_conv2d_16_source_20_pat_count_1[29], _source_stream_conv2d_16_source_20_pat_count_1[26], _source_stream_conv2d_16_source_20_pat_count_1[24:23] }), .Y(_11766_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37535_ ( .A({ _11767_, _11756_, _06702_ }), .Y(_06704_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37536_ ( .A({ _11777_, _11772_, _11770_, _11768_ }), .Y(_11767_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37537_ ( .A({ _11769_, _source_stream_conv2d_16_source_20_pat_count_2[32:30] }), .Y(_11768_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37538_ ( .A({ _source_stream_conv2d_16_source_20_pat_count_2[28:27], _source_stream_conv2d_16_source_20_pat_count_2[25], _source_stream_conv2d_16_source_20_pat_count_2[22] }), .Y(_11769_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37539_ ( .A({ _11771_, _source_stream_conv2d_16_source_20_pat_count_2[1:0] }), .Y(_11770_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37540_ ( .A(_source_stream_conv2d_16_source_20_pat_count_2[5:2]), .Y(_11771_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37541_ ( .A({ _11776_, _11775_, _11774_, _11773_ }), .Y(_11772_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37542_ ( .A(_source_stream_conv2d_16_source_20_pat_count_2[13:10]), .Y(_11773_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37543_ ( .A(_source_stream_conv2d_16_source_20_pat_count_2[9:6]), .Y(_11774_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37544_ ( .A(_source_stream_conv2d_16_source_20_pat_count_2[21:18]), .Y(_11775_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37545_ ( .A(_source_stream_conv2d_16_source_20_pat_count_2[17:14]), .Y(_11776_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37546_ ( .A({ _source_stream_conv2d_16_source_20_pat_count_2[29], _source_stream_conv2d_16_source_20_pat_count_2[26], _source_stream_conv2d_16_source_20_pat_count_2[24:23] }), .Y(_11777_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37547_ ( .A({ _06840_, _05982_ }), .Y(_06705_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37548_ ( .A({ _11778_, _11756_, _11745_ }), .Y(_06840_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37549_ ( .A({ _11788_, _11786_, _11779_, _11767_ }), .Y(_11778_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37550_ ( .A({ _11785_, _11780_, _source_stream_conv2d_16_source_20_pat_count_3[1:0] }), .Y(_11779_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37551_ ( .A({ _11784_, _11783_, _11782_, _11781_ }), .Y(_11780_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37552_ ( .A(_source_stream_conv2d_16_source_20_pat_count_3[13:10]), .Y(_11781_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37553_ ( .A(_source_stream_conv2d_16_source_20_pat_count_3[9:6]), .Y(_11782_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37554_ ( .A(_source_stream_conv2d_16_source_20_pat_count_3[21:18]), .Y(_11783_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37555_ ( .A(_source_stream_conv2d_16_source_20_pat_count_3[17:14]), .Y(_11784_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37556_ ( .A(_source_stream_conv2d_16_source_20_pat_count_3[5:2]), .Y(_11785_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37557_ ( .A({ _11787_, _source_stream_conv2d_16_source_20_pat_count_3[32:30] }), .Y(_11786_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37558_ ( .A({ _source_stream_conv2d_16_source_20_pat_count_3[28:27], _source_stream_conv2d_16_source_20_pat_count_3[25], _source_stream_conv2d_16_source_20_pat_count_3[22] }), .Y(_11787_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37559_ ( .A({ _source_stream_conv2d_16_source_20_pat_count_3[29], _source_stream_conv2d_16_source_20_pat_count_3[26], _source_stream_conv2d_16_source_20_pat_count_3[24:23] }), .Y(_11788_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37560_ ( .A({ _11789_, _05981_ }), .Y(_06707_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37561_ ( .A({ _11799_, _11794_, _11792_, _11790_ }), .Y(_11789_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37562_ ( .A({ _11791_, _source_stream_conv2d_16_source_21_pat_count_0[32:30] }), .Y(_11790_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37563_ ( .A({ _source_stream_conv2d_16_source_21_pat_count_0[28:27], _source_stream_conv2d_16_source_21_pat_count_0[25], _source_stream_conv2d_16_source_21_pat_count_0[22] }), .Y(_11791_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37564_ ( .A({ _11793_, _source_stream_conv2d_16_source_21_pat_count_0[1:0] }), .Y(_11792_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37565_ ( .A(_source_stream_conv2d_16_source_21_pat_count_0[5:2]), .Y(_11793_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37566_ ( .A({ _11798_, _11797_, _11796_, _11795_ }), .Y(_11794_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37567_ ( .A(_source_stream_conv2d_16_source_21_pat_count_0[13:10]), .Y(_11795_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37568_ ( .A(_source_stream_conv2d_16_source_21_pat_count_0[9:6]), .Y(_11796_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37569_ ( .A(_source_stream_conv2d_16_source_21_pat_count_0[21:18]), .Y(_11797_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37570_ ( .A(_source_stream_conv2d_16_source_21_pat_count_0[17:14]), .Y(_11798_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37571_ ( .A({ _source_stream_conv2d_16_source_21_pat_count_0[29], _source_stream_conv2d_16_source_21_pat_count_0[26], _source_stream_conv2d_16_source_21_pat_count_0[24:23] }), .Y(_11799_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37572_ ( .A({ _11800_, _06707_ }), .Y(_06708_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37573_ ( .A({ _11810_, _11808_, _11801_ }), .Y(_11800_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37574_ ( .A({ _11807_, _11802_, _source_stream_conv2d_16_source_21_pat_count_1[1:0] }), .Y(_11801_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37575_ ( .A({ _11806_, _11805_, _11804_, _11803_ }), .Y(_11802_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37576_ ( .A(_source_stream_conv2d_16_source_21_pat_count_1[13:10]), .Y(_11803_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37577_ ( .A(_source_stream_conv2d_16_source_21_pat_count_1[9:6]), .Y(_11804_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37578_ ( .A(_source_stream_conv2d_16_source_21_pat_count_1[21:18]), .Y(_11805_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37579_ ( .A(_source_stream_conv2d_16_source_21_pat_count_1[17:14]), .Y(_11806_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37580_ ( .A(_source_stream_conv2d_16_source_21_pat_count_1[5:2]), .Y(_11807_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37581_ ( .A({ _11809_, _source_stream_conv2d_16_source_21_pat_count_1[32:30] }), .Y(_11808_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37582_ ( .A({ _source_stream_conv2d_16_source_21_pat_count_1[28:27], _source_stream_conv2d_16_source_21_pat_count_1[25], _source_stream_conv2d_16_source_21_pat_count_1[22] }), .Y(_11809_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37583_ ( .A({ _source_stream_conv2d_16_source_21_pat_count_1[29], _source_stream_conv2d_16_source_21_pat_count_1[26], _source_stream_conv2d_16_source_21_pat_count_1[24:23] }), .Y(_11810_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37584_ ( .A({ _11811_, _11800_, _06707_ }), .Y(_06709_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37585_ ( .A({ _11821_, _11816_, _11814_, _11812_ }), .Y(_11811_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37586_ ( .A({ _11813_, _source_stream_conv2d_16_source_21_pat_count_2[32:30] }), .Y(_11812_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37587_ ( .A({ _source_stream_conv2d_16_source_21_pat_count_2[28:27], _source_stream_conv2d_16_source_21_pat_count_2[25], _source_stream_conv2d_16_source_21_pat_count_2[22] }), .Y(_11813_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37588_ ( .A({ _11815_, _source_stream_conv2d_16_source_21_pat_count_2[1:0] }), .Y(_11814_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37589_ ( .A(_source_stream_conv2d_16_source_21_pat_count_2[5:2]), .Y(_11815_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37590_ ( .A({ _11820_, _11819_, _11818_, _11817_ }), .Y(_11816_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37591_ ( .A(_source_stream_conv2d_16_source_21_pat_count_2[13:10]), .Y(_11817_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37592_ ( .A(_source_stream_conv2d_16_source_21_pat_count_2[9:6]), .Y(_11818_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37593_ ( .A(_source_stream_conv2d_16_source_21_pat_count_2[21:18]), .Y(_11819_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37594_ ( .A(_source_stream_conv2d_16_source_21_pat_count_2[17:14]), .Y(_11820_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37595_ ( .A({ _source_stream_conv2d_16_source_21_pat_count_2[29], _source_stream_conv2d_16_source_21_pat_count_2[26], _source_stream_conv2d_16_source_21_pat_count_2[24:23] }), .Y(_11821_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37596_ ( .A({ _06841_, _05981_ }), .Y(_06710_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37597_ ( .A({ _11822_, _11811_, _11789_, _11800_ }), .Y(_06841_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37598_ ( .A({ _11832_, _11827_, _11825_, _11823_ }), .Y(_11822_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37599_ ( .A({ _11824_, _source_stream_conv2d_16_source_21_pat_count_3[32:30] }), .Y(_11823_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37600_ ( .A({ _source_stream_conv2d_16_source_21_pat_count_3[28:27], _source_stream_conv2d_16_source_21_pat_count_3[25], _source_stream_conv2d_16_source_21_pat_count_3[22] }), .Y(_11824_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37601_ ( .A({ _11826_, _source_stream_conv2d_16_source_21_pat_count_3[1:0] }), .Y(_11825_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37602_ ( .A(_source_stream_conv2d_16_source_21_pat_count_3[5:2]), .Y(_11826_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37603_ ( .A({ _11831_, _11830_, _11829_, _11828_ }), .Y(_11827_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37604_ ( .A(_source_stream_conv2d_16_source_21_pat_count_3[13:10]), .Y(_11828_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37605_ ( .A(_source_stream_conv2d_16_source_21_pat_count_3[9:6]), .Y(_11829_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37606_ ( .A(_source_stream_conv2d_16_source_21_pat_count_3[21:18]), .Y(_11830_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37607_ ( .A(_source_stream_conv2d_16_source_21_pat_count_3[17:14]), .Y(_11831_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37608_ ( .A({ _source_stream_conv2d_16_source_21_pat_count_3[29], _source_stream_conv2d_16_source_21_pat_count_3[26], _source_stream_conv2d_16_source_21_pat_count_3[24:23] }), .Y(_11832_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37609_ ( .A({ _11833_, _05979_ }), .Y(_06712_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37610_ ( .A({ _11843_, _11838_, _11836_, _11834_ }), .Y(_11833_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37611_ ( .A({ _11835_, _source_stream_conv2d_16_source_22_pat_count_0[32:30] }), .Y(_11834_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37612_ ( .A({ _source_stream_conv2d_16_source_22_pat_count_0[28:27], _source_stream_conv2d_16_source_22_pat_count_0[25], _source_stream_conv2d_16_source_22_pat_count_0[22] }), .Y(_11835_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37613_ ( .A({ _11837_, _source_stream_conv2d_16_source_22_pat_count_0[1:0] }), .Y(_11836_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37614_ ( .A(_source_stream_conv2d_16_source_22_pat_count_0[5:2]), .Y(_11837_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37615_ ( .A({ _11842_, _11841_, _11840_, _11839_ }), .Y(_11838_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37616_ ( .A(_source_stream_conv2d_16_source_22_pat_count_0[13:10]), .Y(_11839_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37617_ ( .A(_source_stream_conv2d_16_source_22_pat_count_0[9:6]), .Y(_11840_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37618_ ( .A(_source_stream_conv2d_16_source_22_pat_count_0[21:18]), .Y(_11841_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37619_ ( .A(_source_stream_conv2d_16_source_22_pat_count_0[17:14]), .Y(_11842_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37620_ ( .A({ _source_stream_conv2d_16_source_22_pat_count_0[29], _source_stream_conv2d_16_source_22_pat_count_0[26], _source_stream_conv2d_16_source_22_pat_count_0[24:23] }), .Y(_11843_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37621_ ( .A({ _11844_, _06712_ }), .Y(_06713_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37622_ ( .A({ _11854_, _11852_, _11845_ }), .Y(_11844_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37623_ ( .A({ _11851_, _11846_, _source_stream_conv2d_16_source_22_pat_count_1[1:0] }), .Y(_11845_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37624_ ( .A({ _11850_, _11849_, _11848_, _11847_ }), .Y(_11846_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37625_ ( .A(_source_stream_conv2d_16_source_22_pat_count_1[13:10]), .Y(_11847_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37626_ ( .A(_source_stream_conv2d_16_source_22_pat_count_1[9:6]), .Y(_11848_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37627_ ( .A(_source_stream_conv2d_16_source_22_pat_count_1[21:18]), .Y(_11849_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37628_ ( .A(_source_stream_conv2d_16_source_22_pat_count_1[17:14]), .Y(_11850_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37629_ ( .A(_source_stream_conv2d_16_source_22_pat_count_1[5:2]), .Y(_11851_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37630_ ( .A({ _11853_, _source_stream_conv2d_16_source_22_pat_count_1[32:30] }), .Y(_11852_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37631_ ( .A({ _source_stream_conv2d_16_source_22_pat_count_1[28:27], _source_stream_conv2d_16_source_22_pat_count_1[25], _source_stream_conv2d_16_source_22_pat_count_1[22] }), .Y(_11853_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37632_ ( .A({ _source_stream_conv2d_16_source_22_pat_count_1[29], _source_stream_conv2d_16_source_22_pat_count_1[26], _source_stream_conv2d_16_source_22_pat_count_1[24:23] }), .Y(_11854_) );
  \$lut  #( .LUT(8'h40), .WIDTH(3) ) _37633_ ( .A({ _11833_, _11855_, _05979_ }), .Y(_06714_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37634_ ( .A({ _11856_, _11844_ }), .Y(_11855_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37635_ ( .A({ _11866_, _11861_, _11859_, _11857_ }), .Y(_11856_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37636_ ( .A({ _11858_, _source_stream_conv2d_16_source_22_pat_count_2[32:30] }), .Y(_11857_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37637_ ( .A({ _source_stream_conv2d_16_source_22_pat_count_2[28:27], _source_stream_conv2d_16_source_22_pat_count_2[25], _source_stream_conv2d_16_source_22_pat_count_2[22] }), .Y(_11858_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37638_ ( .A({ _11860_, _source_stream_conv2d_16_source_22_pat_count_2[1:0] }), .Y(_11859_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37639_ ( .A(_source_stream_conv2d_16_source_22_pat_count_2[5:2]), .Y(_11860_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37640_ ( .A({ _11865_, _11864_, _11863_, _11862_ }), .Y(_11861_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37641_ ( .A(_source_stream_conv2d_16_source_22_pat_count_2[13:10]), .Y(_11862_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37642_ ( .A(_source_stream_conv2d_16_source_22_pat_count_2[9:6]), .Y(_11863_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37643_ ( .A(_source_stream_conv2d_16_source_22_pat_count_2[21:18]), .Y(_11864_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37644_ ( .A(_source_stream_conv2d_16_source_22_pat_count_2[17:14]), .Y(_11865_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37645_ ( .A({ _source_stream_conv2d_16_source_22_pat_count_2[29], _source_stream_conv2d_16_source_22_pat_count_2[26], _source_stream_conv2d_16_source_22_pat_count_2[24:23] }), .Y(_11866_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37646_ ( .A({ _11867_, _06714_ }), .Y(_06715_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37647_ ( .A({ _11877_, _11875_, _11868_ }), .Y(_11867_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37648_ ( .A({ _11874_, _11869_, _source_stream_conv2d_16_source_22_pat_count_3[1:0] }), .Y(_11868_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37649_ ( .A({ _11873_, _11872_, _11871_, _11870_ }), .Y(_11869_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37650_ ( .A(_source_stream_conv2d_16_source_22_pat_count_3[13:10]), .Y(_11870_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37651_ ( .A(_source_stream_conv2d_16_source_22_pat_count_3[9:6]), .Y(_11871_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37652_ ( .A(_source_stream_conv2d_16_source_22_pat_count_3[21:18]), .Y(_11872_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37653_ ( .A(_source_stream_conv2d_16_source_22_pat_count_3[17:14]), .Y(_11873_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37654_ ( .A(_source_stream_conv2d_16_source_22_pat_count_3[5:2]), .Y(_11874_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37655_ ( .A({ _11876_, _source_stream_conv2d_16_source_22_pat_count_3[32:30] }), .Y(_11875_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37656_ ( .A({ _source_stream_conv2d_16_source_22_pat_count_3[28:27], _source_stream_conv2d_16_source_22_pat_count_3[25], _source_stream_conv2d_16_source_22_pat_count_3[22] }), .Y(_11876_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37657_ ( .A({ _source_stream_conv2d_16_source_22_pat_count_3[29], _source_stream_conv2d_16_source_22_pat_count_3[26], _source_stream_conv2d_16_source_22_pat_count_3[24:23] }), .Y(_11877_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37658_ ( .A({ _11878_, _05977_ }), .Y(_06717_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37659_ ( .A({ _11888_, _11883_, _11881_, _11879_ }), .Y(_11878_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37660_ ( .A({ _11880_, _source_stream_conv2d_16_source_23_pat_count_0[32:30] }), .Y(_11879_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37661_ ( .A({ _source_stream_conv2d_16_source_23_pat_count_0[28:27], _source_stream_conv2d_16_source_23_pat_count_0[25], _source_stream_conv2d_16_source_23_pat_count_0[22] }), .Y(_11880_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37662_ ( .A({ _11882_, _source_stream_conv2d_16_source_23_pat_count_0[1:0] }), .Y(_11881_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37663_ ( .A(_source_stream_conv2d_16_source_23_pat_count_0[5:2]), .Y(_11882_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37664_ ( .A({ _11887_, _11886_, _11885_, _11884_ }), .Y(_11883_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37665_ ( .A(_source_stream_conv2d_16_source_23_pat_count_0[13:10]), .Y(_11884_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37666_ ( .A(_source_stream_conv2d_16_source_23_pat_count_0[9:6]), .Y(_11885_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37667_ ( .A(_source_stream_conv2d_16_source_23_pat_count_0[21:18]), .Y(_11886_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37668_ ( .A(_source_stream_conv2d_16_source_23_pat_count_0[17:14]), .Y(_11887_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37669_ ( .A({ _source_stream_conv2d_16_source_23_pat_count_0[29], _source_stream_conv2d_16_source_23_pat_count_0[26], _source_stream_conv2d_16_source_23_pat_count_0[24:23] }), .Y(_11888_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37670_ ( .A({ _11889_, _06717_ }), .Y(_06718_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37671_ ( .A({ _11899_, _11897_, _11890_ }), .Y(_11889_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37672_ ( .A({ _11896_, _11891_, _source_stream_conv2d_16_source_23_pat_count_1[1:0] }), .Y(_11890_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37673_ ( .A({ _11895_, _11894_, _11893_, _11892_ }), .Y(_11891_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37674_ ( .A(_source_stream_conv2d_16_source_23_pat_count_1[13:10]), .Y(_11892_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37675_ ( .A(_source_stream_conv2d_16_source_23_pat_count_1[9:6]), .Y(_11893_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37676_ ( .A(_source_stream_conv2d_16_source_23_pat_count_1[21:18]), .Y(_11894_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37677_ ( .A(_source_stream_conv2d_16_source_23_pat_count_1[17:14]), .Y(_11895_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37678_ ( .A(_source_stream_conv2d_16_source_23_pat_count_1[5:2]), .Y(_11896_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37679_ ( .A({ _11898_, _source_stream_conv2d_16_source_23_pat_count_1[32:30] }), .Y(_11897_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37680_ ( .A({ _source_stream_conv2d_16_source_23_pat_count_1[28:27], _source_stream_conv2d_16_source_23_pat_count_1[25], _source_stream_conv2d_16_source_23_pat_count_1[22] }), .Y(_11898_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37681_ ( .A({ _source_stream_conv2d_16_source_23_pat_count_1[29], _source_stream_conv2d_16_source_23_pat_count_1[26], _source_stream_conv2d_16_source_23_pat_count_1[24:23] }), .Y(_11899_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37682_ ( .A({ _11900_, _11889_, _06717_ }), .Y(_06719_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37683_ ( .A({ _11910_, _11905_, _11903_, _11901_ }), .Y(_11900_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37684_ ( .A({ _11902_, _source_stream_conv2d_16_source_23_pat_count_2[32:30] }), .Y(_11901_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37685_ ( .A({ _source_stream_conv2d_16_source_23_pat_count_2[28:27], _source_stream_conv2d_16_source_23_pat_count_2[25], _source_stream_conv2d_16_source_23_pat_count_2[22] }), .Y(_11902_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37686_ ( .A({ _11904_, _source_stream_conv2d_16_source_23_pat_count_2[1:0] }), .Y(_11903_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37687_ ( .A(_source_stream_conv2d_16_source_23_pat_count_2[5:2]), .Y(_11904_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37688_ ( .A({ _11909_, _11908_, _11907_, _11906_ }), .Y(_11905_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37689_ ( .A(_source_stream_conv2d_16_source_23_pat_count_2[13:10]), .Y(_11906_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37690_ ( .A(_source_stream_conv2d_16_source_23_pat_count_2[9:6]), .Y(_11907_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37691_ ( .A(_source_stream_conv2d_16_source_23_pat_count_2[21:18]), .Y(_11908_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37692_ ( .A(_source_stream_conv2d_16_source_23_pat_count_2[17:14]), .Y(_11909_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37693_ ( .A({ _source_stream_conv2d_16_source_23_pat_count_2[29], _source_stream_conv2d_16_source_23_pat_count_2[26], _source_stream_conv2d_16_source_23_pat_count_2[24:23] }), .Y(_11910_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37694_ ( .A({ _06843_, _05977_ }), .Y(_06720_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37695_ ( .A({ _11911_, _11900_, _11878_, _11889_ }), .Y(_06843_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37696_ ( .A({ _11921_, _11916_, _11914_, _11912_ }), .Y(_11911_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37697_ ( .A({ _11913_, _source_stream_conv2d_16_source_23_pat_count_3[32:30] }), .Y(_11912_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37698_ ( .A({ _source_stream_conv2d_16_source_23_pat_count_3[28:27], _source_stream_conv2d_16_source_23_pat_count_3[25], _source_stream_conv2d_16_source_23_pat_count_3[22] }), .Y(_11913_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37699_ ( .A({ _11915_, _source_stream_conv2d_16_source_23_pat_count_3[1:0] }), .Y(_11914_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37700_ ( .A(_source_stream_conv2d_16_source_23_pat_count_3[5:2]), .Y(_11915_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37701_ ( .A({ _11920_, _11919_, _11918_, _11917_ }), .Y(_11916_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37702_ ( .A(_source_stream_conv2d_16_source_23_pat_count_3[13:10]), .Y(_11917_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37703_ ( .A(_source_stream_conv2d_16_source_23_pat_count_3[9:6]), .Y(_11918_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37704_ ( .A(_source_stream_conv2d_16_source_23_pat_count_3[21:18]), .Y(_11919_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37705_ ( .A(_source_stream_conv2d_16_source_23_pat_count_3[17:14]), .Y(_11920_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37706_ ( .A({ _source_stream_conv2d_16_source_23_pat_count_3[29], _source_stream_conv2d_16_source_23_pat_count_3[26], _source_stream_conv2d_16_source_23_pat_count_3[24:23] }), .Y(_11921_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37707_ ( .A({ _11922_, _05972_ }), .Y(_06722_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37708_ ( .A({ _11932_, _11931_, _11930_, _11923_ }), .Y(_11922_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37709_ ( .A({ _11929_, _11924_, _source_stream_conv2d_16_source_24_pat_count_0[1:0] }), .Y(_11923_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37710_ ( .A({ _11928_, _11927_, _11926_, _11925_ }), .Y(_11924_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37711_ ( .A(_source_stream_conv2d_16_source_24_pat_count_0[13:10]), .Y(_11925_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37712_ ( .A(_source_stream_conv2d_16_source_24_pat_count_0[9:6]), .Y(_11926_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37713_ ( .A(_source_stream_conv2d_16_source_24_pat_count_0[21:18]), .Y(_11927_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37714_ ( .A(_source_stream_conv2d_16_source_24_pat_count_0[17:14]), .Y(_11928_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37715_ ( .A(_source_stream_conv2d_16_source_24_pat_count_0[5:2]), .Y(_11929_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _37716_ ( .A(_source_stream_conv2d_16_source_24_pat_count_0[32:30]), .Y(_11930_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37717_ ( .A(_source_stream_conv2d_16_source_24_pat_count_0[29:26]), .Y(_11931_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37718_ ( .A(_source_stream_conv2d_16_source_24_pat_count_0[25:22]), .Y(_11932_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37719_ ( .A({ _11933_, _06722_ }), .Y(_06723_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37720_ ( .A({ _11943_, _11941_, _11934_ }), .Y(_11933_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37721_ ( .A({ _11940_, _11935_, _source_stream_conv2d_16_source_24_pat_count_1[1:0] }), .Y(_11934_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37722_ ( .A({ _11939_, _11938_, _11937_, _11936_ }), .Y(_11935_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37723_ ( .A(_source_stream_conv2d_16_source_24_pat_count_1[13:10]), .Y(_11936_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37724_ ( .A(_source_stream_conv2d_16_source_24_pat_count_1[9:6]), .Y(_11937_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37725_ ( .A(_source_stream_conv2d_16_source_24_pat_count_1[21:18]), .Y(_11938_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37726_ ( .A(_source_stream_conv2d_16_source_24_pat_count_1[17:14]), .Y(_11939_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37727_ ( .A(_source_stream_conv2d_16_source_24_pat_count_1[5:2]), .Y(_11940_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37728_ ( .A({ _11942_, _source_stream_conv2d_16_source_24_pat_count_1[32:30] }), .Y(_11941_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37729_ ( .A({ _source_stream_conv2d_16_source_24_pat_count_1[28:27], _source_stream_conv2d_16_source_24_pat_count_1[25], _source_stream_conv2d_16_source_24_pat_count_1[22] }), .Y(_11942_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37730_ ( .A({ _source_stream_conv2d_16_source_24_pat_count_1[29], _source_stream_conv2d_16_source_24_pat_count_1[26], _source_stream_conv2d_16_source_24_pat_count_1[24:23] }), .Y(_11943_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37731_ ( .A({ _11944_, _11933_, _06722_ }), .Y(_06724_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37732_ ( .A({ _11954_, _11949_, _11947_, _11945_ }), .Y(_11944_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37733_ ( .A({ _11946_, _source_stream_conv2d_16_source_24_pat_count_2[32:30] }), .Y(_11945_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37734_ ( .A({ _source_stream_conv2d_16_source_24_pat_count_2[28:27], _source_stream_conv2d_16_source_24_pat_count_2[25], _source_stream_conv2d_16_source_24_pat_count_2[22] }), .Y(_11946_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37735_ ( .A({ _11948_, _source_stream_conv2d_16_source_24_pat_count_2[1:0] }), .Y(_11947_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37736_ ( .A(_source_stream_conv2d_16_source_24_pat_count_2[5:2]), .Y(_11948_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37737_ ( .A({ _11953_, _11952_, _11951_, _11950_ }), .Y(_11949_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37738_ ( .A(_source_stream_conv2d_16_source_24_pat_count_2[13:10]), .Y(_11950_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37739_ ( .A(_source_stream_conv2d_16_source_24_pat_count_2[9:6]), .Y(_11951_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37740_ ( .A(_source_stream_conv2d_16_source_24_pat_count_2[21:18]), .Y(_11952_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37741_ ( .A(_source_stream_conv2d_16_source_24_pat_count_2[17:14]), .Y(_11953_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37742_ ( .A({ _source_stream_conv2d_16_source_24_pat_count_2[29], _source_stream_conv2d_16_source_24_pat_count_2[26], _source_stream_conv2d_16_source_24_pat_count_2[24:23] }), .Y(_11954_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37743_ ( .A({ _06844_, _05972_ }), .Y(_06725_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37744_ ( .A({ _11955_, _11944_, _11933_, _11922_ }), .Y(_06844_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37745_ ( .A({ _11965_, _11960_, _11958_, _11956_ }), .Y(_11955_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37746_ ( .A({ _11957_, _source_stream_conv2d_16_source_24_pat_count_3[32:30] }), .Y(_11956_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37747_ ( .A({ _source_stream_conv2d_16_source_24_pat_count_3[28:27], _source_stream_conv2d_16_source_24_pat_count_3[25], _source_stream_conv2d_16_source_24_pat_count_3[22] }), .Y(_11957_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37748_ ( .A({ _11959_, _source_stream_conv2d_16_source_24_pat_count_3[1:0] }), .Y(_11958_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37749_ ( .A(_source_stream_conv2d_16_source_24_pat_count_3[5:2]), .Y(_11959_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37750_ ( .A({ _11964_, _11963_, _11962_, _11961_ }), .Y(_11960_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37751_ ( .A(_source_stream_conv2d_16_source_24_pat_count_3[13:10]), .Y(_11961_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37752_ ( .A(_source_stream_conv2d_16_source_24_pat_count_3[9:6]), .Y(_11962_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37753_ ( .A(_source_stream_conv2d_16_source_24_pat_count_3[21:18]), .Y(_11963_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37754_ ( .A(_source_stream_conv2d_16_source_24_pat_count_3[17:14]), .Y(_11964_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37755_ ( .A({ _source_stream_conv2d_16_source_24_pat_count_3[29], _source_stream_conv2d_16_source_24_pat_count_3[26], _source_stream_conv2d_16_source_24_pat_count_3[24:23] }), .Y(_11965_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37756_ ( .A({ _11966_, _05974_ }), .Y(_06727_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37757_ ( .A({ _11976_, _11971_, _11969_, _11967_ }), .Y(_11966_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37758_ ( .A({ _11968_, _source_stream_conv2d_16_source_25_pat_count_0[32:30] }), .Y(_11967_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37759_ ( .A({ _source_stream_conv2d_16_source_25_pat_count_0[28:27], _source_stream_conv2d_16_source_25_pat_count_0[25], _source_stream_conv2d_16_source_25_pat_count_0[22] }), .Y(_11968_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37760_ ( .A({ _11970_, _source_stream_conv2d_16_source_25_pat_count_0[1:0] }), .Y(_11969_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37761_ ( .A(_source_stream_conv2d_16_source_25_pat_count_0[5:2]), .Y(_11970_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37762_ ( .A({ _11975_, _11974_, _11973_, _11972_ }), .Y(_11971_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37763_ ( .A(_source_stream_conv2d_16_source_25_pat_count_0[13:10]), .Y(_11972_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37764_ ( .A(_source_stream_conv2d_16_source_25_pat_count_0[9:6]), .Y(_11973_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37765_ ( .A(_source_stream_conv2d_16_source_25_pat_count_0[21:18]), .Y(_11974_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37766_ ( .A(_source_stream_conv2d_16_source_25_pat_count_0[17:14]), .Y(_11975_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37767_ ( .A({ _source_stream_conv2d_16_source_25_pat_count_0[29], _source_stream_conv2d_16_source_25_pat_count_0[26], _source_stream_conv2d_16_source_25_pat_count_0[24:23] }), .Y(_11976_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37768_ ( .A({ _11977_, _06727_ }), .Y(_06728_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37769_ ( .A({ _11987_, _11985_, _11978_ }), .Y(_11977_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37770_ ( .A({ _11984_, _11979_, _source_stream_conv2d_16_source_25_pat_count_1[1:0] }), .Y(_11978_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37771_ ( .A({ _11983_, _11982_, _11981_, _11980_ }), .Y(_11979_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37772_ ( .A(_source_stream_conv2d_16_source_25_pat_count_1[13:10]), .Y(_11980_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37773_ ( .A(_source_stream_conv2d_16_source_25_pat_count_1[9:6]), .Y(_11981_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37774_ ( .A(_source_stream_conv2d_16_source_25_pat_count_1[21:18]), .Y(_11982_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37775_ ( .A(_source_stream_conv2d_16_source_25_pat_count_1[17:14]), .Y(_11983_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37776_ ( .A(_source_stream_conv2d_16_source_25_pat_count_1[5:2]), .Y(_11984_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37777_ ( .A({ _11986_, _source_stream_conv2d_16_source_25_pat_count_1[32:30] }), .Y(_11985_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37778_ ( .A({ _source_stream_conv2d_16_source_25_pat_count_1[28:27], _source_stream_conv2d_16_source_25_pat_count_1[25], _source_stream_conv2d_16_source_25_pat_count_1[22] }), .Y(_11986_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37779_ ( .A({ _source_stream_conv2d_16_source_25_pat_count_1[29], _source_stream_conv2d_16_source_25_pat_count_1[26], _source_stream_conv2d_16_source_25_pat_count_1[24:23] }), .Y(_11987_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37780_ ( .A({ _11988_, _11977_, _06727_ }), .Y(_06729_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37781_ ( .A({ _11998_, _11993_, _11991_, _11989_ }), .Y(_11988_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37782_ ( .A({ _11990_, _source_stream_conv2d_16_source_25_pat_count_2[32:30] }), .Y(_11989_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37783_ ( .A({ _source_stream_conv2d_16_source_25_pat_count_2[28:27], _source_stream_conv2d_16_source_25_pat_count_2[25], _source_stream_conv2d_16_source_25_pat_count_2[22] }), .Y(_11990_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37784_ ( .A({ _11992_, _source_stream_conv2d_16_source_25_pat_count_2[1:0] }), .Y(_11991_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37785_ ( .A(_source_stream_conv2d_16_source_25_pat_count_2[5:2]), .Y(_11992_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37786_ ( .A({ _11997_, _11996_, _11995_, _11994_ }), .Y(_11993_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37787_ ( .A(_source_stream_conv2d_16_source_25_pat_count_2[13:10]), .Y(_11994_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37788_ ( .A(_source_stream_conv2d_16_source_25_pat_count_2[9:6]), .Y(_11995_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37789_ ( .A(_source_stream_conv2d_16_source_25_pat_count_2[21:18]), .Y(_11996_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37790_ ( .A(_source_stream_conv2d_16_source_25_pat_count_2[17:14]), .Y(_11997_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37791_ ( .A({ _source_stream_conv2d_16_source_25_pat_count_2[29], _source_stream_conv2d_16_source_25_pat_count_2[26], _source_stream_conv2d_16_source_25_pat_count_2[24:23] }), .Y(_11998_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37792_ ( .A({ _06845_, _05974_ }), .Y(_06730_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37793_ ( .A({ _11999_, _11988_, _11966_, _11977_ }), .Y(_06845_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37794_ ( .A({ _12009_, _12004_, _12002_, _12000_ }), .Y(_11999_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37795_ ( .A({ _12001_, _source_stream_conv2d_16_source_25_pat_count_3[32:30] }), .Y(_12000_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37796_ ( .A({ _source_stream_conv2d_16_source_25_pat_count_3[28:27], _source_stream_conv2d_16_source_25_pat_count_3[25], _source_stream_conv2d_16_source_25_pat_count_3[22] }), .Y(_12001_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37797_ ( .A({ _12003_, _source_stream_conv2d_16_source_25_pat_count_3[1:0] }), .Y(_12002_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37798_ ( .A(_source_stream_conv2d_16_source_25_pat_count_3[5:2]), .Y(_12003_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37799_ ( .A({ _12008_, _12007_, _12006_, _12005_ }), .Y(_12004_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37800_ ( .A(_source_stream_conv2d_16_source_25_pat_count_3[13:10]), .Y(_12005_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37801_ ( .A(_source_stream_conv2d_16_source_25_pat_count_3[9:6]), .Y(_12006_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37802_ ( .A(_source_stream_conv2d_16_source_25_pat_count_3[21:18]), .Y(_12007_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37803_ ( .A(_source_stream_conv2d_16_source_25_pat_count_3[17:14]), .Y(_12008_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37804_ ( .A({ _source_stream_conv2d_16_source_25_pat_count_3[29], _source_stream_conv2d_16_source_25_pat_count_3[26], _source_stream_conv2d_16_source_25_pat_count_3[24:23] }), .Y(_12009_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37805_ ( .A({ _12010_, _05971_ }), .Y(_06732_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37806_ ( .A({ _12020_, _12015_, _12013_, _12011_ }), .Y(_12010_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37807_ ( .A({ _12012_, _source_stream_conv2d_16_source_26_pat_count_0[32:30] }), .Y(_12011_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37808_ ( .A({ _source_stream_conv2d_16_source_26_pat_count_0[28:27], _source_stream_conv2d_16_source_26_pat_count_0[25], _source_stream_conv2d_16_source_26_pat_count_0[22] }), .Y(_12012_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37809_ ( .A({ _12014_, _source_stream_conv2d_16_source_26_pat_count_0[1:0] }), .Y(_12013_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37810_ ( .A(_source_stream_conv2d_16_source_26_pat_count_0[5:2]), .Y(_12014_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37811_ ( .A({ _12019_, _12018_, _12017_, _12016_ }), .Y(_12015_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37812_ ( .A(_source_stream_conv2d_16_source_26_pat_count_0[13:10]), .Y(_12016_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37813_ ( .A(_source_stream_conv2d_16_source_26_pat_count_0[9:6]), .Y(_12017_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37814_ ( .A(_source_stream_conv2d_16_source_26_pat_count_0[21:18]), .Y(_12018_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37815_ ( .A(_source_stream_conv2d_16_source_26_pat_count_0[17:14]), .Y(_12019_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37816_ ( .A({ _source_stream_conv2d_16_source_26_pat_count_0[29], _source_stream_conv2d_16_source_26_pat_count_0[26], _source_stream_conv2d_16_source_26_pat_count_0[24:23] }), .Y(_12020_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37817_ ( .A({ _12021_, _06732_ }), .Y(_06733_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37818_ ( .A({ _12031_, _12029_, _12022_ }), .Y(_12021_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37819_ ( .A({ _12028_, _12023_, _source_stream_conv2d_16_source_26_pat_count_1[1:0] }), .Y(_12022_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37820_ ( .A({ _12027_, _12026_, _12025_, _12024_ }), .Y(_12023_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37821_ ( .A(_source_stream_conv2d_16_source_26_pat_count_1[13:10]), .Y(_12024_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37822_ ( .A(_source_stream_conv2d_16_source_26_pat_count_1[9:6]), .Y(_12025_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37823_ ( .A(_source_stream_conv2d_16_source_26_pat_count_1[21:18]), .Y(_12026_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37824_ ( .A(_source_stream_conv2d_16_source_26_pat_count_1[17:14]), .Y(_12027_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37825_ ( .A(_source_stream_conv2d_16_source_26_pat_count_1[5:2]), .Y(_12028_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37826_ ( .A({ _12030_, _source_stream_conv2d_16_source_26_pat_count_1[32:30] }), .Y(_12029_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37827_ ( .A({ _source_stream_conv2d_16_source_26_pat_count_1[28:27], _source_stream_conv2d_16_source_26_pat_count_1[25], _source_stream_conv2d_16_source_26_pat_count_1[22] }), .Y(_12030_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37828_ ( .A({ _source_stream_conv2d_16_source_26_pat_count_1[29], _source_stream_conv2d_16_source_26_pat_count_1[26], _source_stream_conv2d_16_source_26_pat_count_1[24:23] }), .Y(_12031_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37829_ ( .A({ _12032_, _12021_, _06732_ }), .Y(_06734_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37830_ ( .A({ _12042_, _12037_, _12035_, _12033_ }), .Y(_12032_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37831_ ( .A({ _12034_, _source_stream_conv2d_16_source_26_pat_count_2[32:30] }), .Y(_12033_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37832_ ( .A({ _source_stream_conv2d_16_source_26_pat_count_2[28:27], _source_stream_conv2d_16_source_26_pat_count_2[25], _source_stream_conv2d_16_source_26_pat_count_2[22] }), .Y(_12034_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37833_ ( .A({ _12036_, _source_stream_conv2d_16_source_26_pat_count_2[1:0] }), .Y(_12035_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37834_ ( .A(_source_stream_conv2d_16_source_26_pat_count_2[5:2]), .Y(_12036_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37835_ ( .A({ _12041_, _12040_, _12039_, _12038_ }), .Y(_12037_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37836_ ( .A(_source_stream_conv2d_16_source_26_pat_count_2[13:10]), .Y(_12038_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37837_ ( .A(_source_stream_conv2d_16_source_26_pat_count_2[9:6]), .Y(_12039_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37838_ ( .A(_source_stream_conv2d_16_source_26_pat_count_2[21:18]), .Y(_12040_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37839_ ( .A(_source_stream_conv2d_16_source_26_pat_count_2[17:14]), .Y(_12041_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37840_ ( .A({ _source_stream_conv2d_16_source_26_pat_count_2[29], _source_stream_conv2d_16_source_26_pat_count_2[26], _source_stream_conv2d_16_source_26_pat_count_2[24:23] }), .Y(_12042_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37841_ ( .A({ _06846_, _05971_ }), .Y(_06735_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37842_ ( .A({ _12032_, _12043_, _12021_ }), .Y(_06846_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37843_ ( .A({ _12053_, _12051_, _12044_, _12010_ }), .Y(_12043_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37844_ ( .A({ _12050_, _12045_, _source_stream_conv2d_16_source_26_pat_count_3[1:0] }), .Y(_12044_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37845_ ( .A({ _12049_, _12048_, _12047_, _12046_ }), .Y(_12045_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37846_ ( .A(_source_stream_conv2d_16_source_26_pat_count_3[13:10]), .Y(_12046_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37847_ ( .A(_source_stream_conv2d_16_source_26_pat_count_3[9:6]), .Y(_12047_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37848_ ( .A(_source_stream_conv2d_16_source_26_pat_count_3[21:18]), .Y(_12048_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37849_ ( .A(_source_stream_conv2d_16_source_26_pat_count_3[17:14]), .Y(_12049_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37850_ ( .A(_source_stream_conv2d_16_source_26_pat_count_3[5:2]), .Y(_12050_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37851_ ( .A({ _12052_, _source_stream_conv2d_16_source_26_pat_count_3[32:30] }), .Y(_12051_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37852_ ( .A({ _source_stream_conv2d_16_source_26_pat_count_3[28:27], _source_stream_conv2d_16_source_26_pat_count_3[25], _source_stream_conv2d_16_source_26_pat_count_3[22] }), .Y(_12052_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37853_ ( .A({ _source_stream_conv2d_16_source_26_pat_count_3[29], _source_stream_conv2d_16_source_26_pat_count_3[26], _source_stream_conv2d_16_source_26_pat_count_3[24:23] }), .Y(_12053_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37854_ ( .A({ _12054_, _05968_ }), .Y(_06737_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37855_ ( .A({ _12064_, _12059_, _12057_, _12055_ }), .Y(_12054_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37856_ ( .A({ _12056_, _source_stream_conv2d_16_source_27_pat_count_0[32:30] }), .Y(_12055_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37857_ ( .A({ _source_stream_conv2d_16_source_27_pat_count_0[28:27], _source_stream_conv2d_16_source_27_pat_count_0[25], _source_stream_conv2d_16_source_27_pat_count_0[22] }), .Y(_12056_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37858_ ( .A({ _12058_, _source_stream_conv2d_16_source_27_pat_count_0[1:0] }), .Y(_12057_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37859_ ( .A(_source_stream_conv2d_16_source_27_pat_count_0[5:2]), .Y(_12058_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37860_ ( .A({ _12063_, _12062_, _12061_, _12060_ }), .Y(_12059_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37861_ ( .A(_source_stream_conv2d_16_source_27_pat_count_0[13:10]), .Y(_12060_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37862_ ( .A(_source_stream_conv2d_16_source_27_pat_count_0[9:6]), .Y(_12061_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37863_ ( .A(_source_stream_conv2d_16_source_27_pat_count_0[21:18]), .Y(_12062_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37864_ ( .A(_source_stream_conv2d_16_source_27_pat_count_0[17:14]), .Y(_12063_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37865_ ( .A({ _source_stream_conv2d_16_source_27_pat_count_0[29], _source_stream_conv2d_16_source_27_pat_count_0[26], _source_stream_conv2d_16_source_27_pat_count_0[24:23] }), .Y(_12064_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37866_ ( .A({ _12065_, _06737_ }), .Y(_06738_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37867_ ( .A({ _12075_, _12073_, _12066_ }), .Y(_12065_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37868_ ( .A({ _12072_, _12067_, _source_stream_conv2d_16_source_27_pat_count_1[1:0] }), .Y(_12066_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37869_ ( .A({ _12071_, _12070_, _12069_, _12068_ }), .Y(_12067_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37870_ ( .A(_source_stream_conv2d_16_source_27_pat_count_1[13:10]), .Y(_12068_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37871_ ( .A(_source_stream_conv2d_16_source_27_pat_count_1[9:6]), .Y(_12069_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37872_ ( .A(_source_stream_conv2d_16_source_27_pat_count_1[21:18]), .Y(_12070_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37873_ ( .A(_source_stream_conv2d_16_source_27_pat_count_1[17:14]), .Y(_12071_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37874_ ( .A(_source_stream_conv2d_16_source_27_pat_count_1[5:2]), .Y(_12072_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37875_ ( .A({ _12074_, _source_stream_conv2d_16_source_27_pat_count_1[32:30] }), .Y(_12073_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37876_ ( .A({ _source_stream_conv2d_16_source_27_pat_count_1[28:27], _source_stream_conv2d_16_source_27_pat_count_1[25], _source_stream_conv2d_16_source_27_pat_count_1[22] }), .Y(_12074_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37877_ ( .A({ _source_stream_conv2d_16_source_27_pat_count_1[29], _source_stream_conv2d_16_source_27_pat_count_1[26], _source_stream_conv2d_16_source_27_pat_count_1[24:23] }), .Y(_12075_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37878_ ( .A({ _12076_, _12065_, _06737_ }), .Y(_06739_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37879_ ( .A({ _12086_, _12081_, _12079_, _12077_ }), .Y(_12076_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37880_ ( .A({ _12078_, _source_stream_conv2d_16_source_27_pat_count_2[32:30] }), .Y(_12077_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37881_ ( .A({ _source_stream_conv2d_16_source_27_pat_count_2[28:27], _source_stream_conv2d_16_source_27_pat_count_2[25], _source_stream_conv2d_16_source_27_pat_count_2[22] }), .Y(_12078_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37882_ ( .A({ _12080_, _source_stream_conv2d_16_source_27_pat_count_2[1:0] }), .Y(_12079_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37883_ ( .A(_source_stream_conv2d_16_source_27_pat_count_2[5:2]), .Y(_12080_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37884_ ( .A({ _12085_, _12084_, _12083_, _12082_ }), .Y(_12081_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37885_ ( .A(_source_stream_conv2d_16_source_27_pat_count_2[13:10]), .Y(_12082_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37886_ ( .A(_source_stream_conv2d_16_source_27_pat_count_2[9:6]), .Y(_12083_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37887_ ( .A(_source_stream_conv2d_16_source_27_pat_count_2[21:18]), .Y(_12084_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37888_ ( .A(_source_stream_conv2d_16_source_27_pat_count_2[17:14]), .Y(_12085_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37889_ ( .A({ _source_stream_conv2d_16_source_27_pat_count_2[29], _source_stream_conv2d_16_source_27_pat_count_2[26], _source_stream_conv2d_16_source_27_pat_count_2[24:23] }), .Y(_12086_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37890_ ( .A({ _06847_, _05968_ }), .Y(_06740_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37891_ ( .A({ _12087_, _12076_, _12054_, _12065_ }), .Y(_06847_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37892_ ( .A({ _12097_, _12092_, _12090_, _12088_ }), .Y(_12087_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37893_ ( .A({ _12089_, _source_stream_conv2d_16_source_27_pat_count_3[32:30] }), .Y(_12088_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37894_ ( .A({ _source_stream_conv2d_16_source_27_pat_count_3[28:27], _source_stream_conv2d_16_source_27_pat_count_3[25], _source_stream_conv2d_16_source_27_pat_count_3[22] }), .Y(_12089_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37895_ ( .A({ _12091_, _source_stream_conv2d_16_source_27_pat_count_3[1:0] }), .Y(_12090_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37896_ ( .A(_source_stream_conv2d_16_source_27_pat_count_3[5:2]), .Y(_12091_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37897_ ( .A({ _12096_, _12095_, _12094_, _12093_ }), .Y(_12092_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37898_ ( .A(_source_stream_conv2d_16_source_27_pat_count_3[13:10]), .Y(_12093_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37899_ ( .A(_source_stream_conv2d_16_source_27_pat_count_3[9:6]), .Y(_12094_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37900_ ( .A(_source_stream_conv2d_16_source_27_pat_count_3[21:18]), .Y(_12095_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37901_ ( .A(_source_stream_conv2d_16_source_27_pat_count_3[17:14]), .Y(_12096_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37902_ ( .A({ _source_stream_conv2d_16_source_27_pat_count_3[29], _source_stream_conv2d_16_source_27_pat_count_3[26], _source_stream_conv2d_16_source_27_pat_count_3[24:23] }), .Y(_12097_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37903_ ( .A({ _12098_, _05966_ }), .Y(_06742_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37904_ ( .A({ _12108_, _12107_, _12106_, _12099_ }), .Y(_12098_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37905_ ( .A({ _12105_, _12100_, _source_stream_conv2d_16_source_28_pat_count_0[1:0] }), .Y(_12099_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37906_ ( .A({ _12104_, _12103_, _12102_, _12101_ }), .Y(_12100_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37907_ ( .A(_source_stream_conv2d_16_source_28_pat_count_0[13:10]), .Y(_12101_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37908_ ( .A(_source_stream_conv2d_16_source_28_pat_count_0[9:6]), .Y(_12102_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37909_ ( .A(_source_stream_conv2d_16_source_28_pat_count_0[21:18]), .Y(_12103_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37910_ ( .A(_source_stream_conv2d_16_source_28_pat_count_0[17:14]), .Y(_12104_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37911_ ( .A(_source_stream_conv2d_16_source_28_pat_count_0[5:2]), .Y(_12105_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _37912_ ( .A(_source_stream_conv2d_16_source_28_pat_count_0[32:30]), .Y(_12106_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37913_ ( .A(_source_stream_conv2d_16_source_28_pat_count_0[29:26]), .Y(_12107_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37914_ ( .A(_source_stream_conv2d_16_source_28_pat_count_0[25:22]), .Y(_12108_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37915_ ( .A({ _12109_, _06742_ }), .Y(_06743_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37916_ ( .A({ _12119_, _12117_, _12110_ }), .Y(_12109_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37917_ ( .A({ _12116_, _12111_, _source_stream_conv2d_16_source_28_pat_count_1[1:0] }), .Y(_12110_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37918_ ( .A({ _12115_, _12114_, _12113_, _12112_ }), .Y(_12111_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37919_ ( .A(_source_stream_conv2d_16_source_28_pat_count_1[13:10]), .Y(_12112_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37920_ ( .A(_source_stream_conv2d_16_source_28_pat_count_1[9:6]), .Y(_12113_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37921_ ( .A(_source_stream_conv2d_16_source_28_pat_count_1[21:18]), .Y(_12114_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37922_ ( .A(_source_stream_conv2d_16_source_28_pat_count_1[17:14]), .Y(_12115_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37923_ ( .A(_source_stream_conv2d_16_source_28_pat_count_1[5:2]), .Y(_12116_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37924_ ( .A({ _12118_, _source_stream_conv2d_16_source_28_pat_count_1[32:30] }), .Y(_12117_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37925_ ( .A({ _source_stream_conv2d_16_source_28_pat_count_1[28:27], _source_stream_conv2d_16_source_28_pat_count_1[25], _source_stream_conv2d_16_source_28_pat_count_1[22] }), .Y(_12118_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37926_ ( .A({ _source_stream_conv2d_16_source_28_pat_count_1[29], _source_stream_conv2d_16_source_28_pat_count_1[26], _source_stream_conv2d_16_source_28_pat_count_1[24:23] }), .Y(_12119_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37927_ ( .A({ _12120_, _06742_ }), .Y(_06744_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37928_ ( .A({ _12127_, _12121_, _12109_ }), .Y(_12120_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37929_ ( .A({ _12126_, _12124_, _12122_ }), .Y(_12121_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37930_ ( .A({ _12123_, _source_stream_conv2d_16_source_28_pat_count_2[17], _source_stream_conv2d_16_source_28_pat_count_2[14], _source_stream_conv2d_16_source_28_pat_count_2[4] }), .Y(_12122_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37931_ ( .A({ _source_stream_conv2d_16_source_28_pat_count_2[21], _source_stream_conv2d_16_source_28_pat_count_2[18], _source_stream_conv2d_16_source_28_pat_count_2[16:15] }), .Y(_12123_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37932_ ( .A({ _12125_, _source_stream_conv2d_16_source_28_pat_count_2[27], _source_stream_conv2d_16_source_28_pat_count_2[20], _source_stream_conv2d_16_source_28_pat_count_2[1] }), .Y(_12124_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37933_ ( .A({ _source_stream_conv2d_16_source_28_pat_count_2[28], _source_stream_conv2d_16_source_28_pat_count_2[22], _source_stream_conv2d_16_source_28_pat_count_2[19], _source_stream_conv2d_16_source_28_pat_count_2[3] }), .Y(_12125_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37934_ ( .A({ _source_stream_conv2d_16_source_28_pat_count_2[12:11], _source_stream_conv2d_16_source_28_pat_count_2[9], _source_stream_conv2d_16_source_28_pat_count_2[6] }), .Y(_12126_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37935_ ( .A({ _12131_, _12128_, _source_stream_conv2d_16_source_28_pat_count_2[2], _source_stream_conv2d_16_source_28_pat_count_2[0] }), .Y(_12127_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37936_ ( .A({ _12130_, _12129_, _source_stream_conv2d_16_source_28_pat_count_2[10], _source_stream_conv2d_16_source_28_pat_count_2[5] }), .Y(_12128_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _37937_ ( .A(_source_stream_conv2d_16_source_28_pat_count_2[25:23]), .Y(_12129_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _37938_ ( .A({ _source_stream_conv2d_16_source_28_pat_count_2[13], _source_stream_conv2d_16_source_28_pat_count_2[8:7] }), .Y(_12130_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37939_ ( .A({ _12132_, _source_stream_conv2d_16_source_28_pat_count_2[29], _source_stream_conv2d_16_source_28_pat_count_2[26] }), .Y(_12131_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _37940_ ( .A(_source_stream_conv2d_16_source_28_pat_count_2[32:30]), .Y(_12132_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37941_ ( .A({ _12133_, _06744_ }), .Y(_06745_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37942_ ( .A({ _12143_, _12141_, _12134_ }), .Y(_12133_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37943_ ( .A({ _12140_, _12135_, _source_stream_conv2d_16_source_28_pat_count_3[1:0] }), .Y(_12134_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37944_ ( .A({ _12139_, _12138_, _12137_, _12136_ }), .Y(_12135_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37945_ ( .A(_source_stream_conv2d_16_source_28_pat_count_3[13:10]), .Y(_12136_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37946_ ( .A(_source_stream_conv2d_16_source_28_pat_count_3[9:6]), .Y(_12137_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37947_ ( .A(_source_stream_conv2d_16_source_28_pat_count_3[21:18]), .Y(_12138_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37948_ ( .A(_source_stream_conv2d_16_source_28_pat_count_3[17:14]), .Y(_12139_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37949_ ( .A(_source_stream_conv2d_16_source_28_pat_count_3[5:2]), .Y(_12140_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37950_ ( .A({ _12142_, _source_stream_conv2d_16_source_28_pat_count_3[32:30] }), .Y(_12141_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37951_ ( .A({ _source_stream_conv2d_16_source_28_pat_count_3[28:27], _source_stream_conv2d_16_source_28_pat_count_3[25], _source_stream_conv2d_16_source_28_pat_count_3[22] }), .Y(_12142_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37952_ ( .A({ _source_stream_conv2d_16_source_28_pat_count_3[29], _source_stream_conv2d_16_source_28_pat_count_3[26], _source_stream_conv2d_16_source_28_pat_count_3[24:23] }), .Y(_12143_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _37953_ ( .A({ _12144_, _05965_ }), .Y(_06747_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37954_ ( .A({ _12154_, _12153_, _12152_, _12145_ }), .Y(_12144_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37955_ ( .A({ _12151_, _12146_, _source_stream_conv2d_16_source_29_pat_count_0[1:0] }), .Y(_12145_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37956_ ( .A({ _12150_, _12149_, _12148_, _12147_ }), .Y(_12146_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37957_ ( .A(_source_stream_conv2d_16_source_29_pat_count_0[13:10]), .Y(_12147_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37958_ ( .A(_source_stream_conv2d_16_source_29_pat_count_0[9:6]), .Y(_12148_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37959_ ( .A(_source_stream_conv2d_16_source_29_pat_count_0[21:18]), .Y(_12149_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37960_ ( .A(_source_stream_conv2d_16_source_29_pat_count_0[17:14]), .Y(_12150_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37961_ ( .A(_source_stream_conv2d_16_source_29_pat_count_0[5:2]), .Y(_12151_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _37962_ ( .A(_source_stream_conv2d_16_source_29_pat_count_0[32:30]), .Y(_12152_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37963_ ( .A(_source_stream_conv2d_16_source_29_pat_count_0[29:26]), .Y(_12153_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37964_ ( .A(_source_stream_conv2d_16_source_29_pat_count_0[25:22]), .Y(_12154_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37965_ ( .A({ _12155_, _06747_ }), .Y(_06748_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37966_ ( .A({ _12165_, _12163_, _12156_ }), .Y(_12155_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37967_ ( .A({ _12162_, _12157_, _source_stream_conv2d_16_source_29_pat_count_1[1:0] }), .Y(_12156_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37968_ ( .A({ _12161_, _12160_, _12159_, _12158_ }), .Y(_12157_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37969_ ( .A(_source_stream_conv2d_16_source_29_pat_count_1[13:10]), .Y(_12158_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37970_ ( .A(_source_stream_conv2d_16_source_29_pat_count_1[9:6]), .Y(_12159_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37971_ ( .A(_source_stream_conv2d_16_source_29_pat_count_1[21:18]), .Y(_12160_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37972_ ( .A(_source_stream_conv2d_16_source_29_pat_count_1[17:14]), .Y(_12161_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37973_ ( .A(_source_stream_conv2d_16_source_29_pat_count_1[5:2]), .Y(_12162_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37974_ ( .A({ _12164_, _source_stream_conv2d_16_source_29_pat_count_1[32:30] }), .Y(_12163_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37975_ ( .A({ _source_stream_conv2d_16_source_29_pat_count_1[28:27], _source_stream_conv2d_16_source_29_pat_count_1[25], _source_stream_conv2d_16_source_29_pat_count_1[22] }), .Y(_12164_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37976_ ( .A({ _source_stream_conv2d_16_source_29_pat_count_1[29], _source_stream_conv2d_16_source_29_pat_count_1[26], _source_stream_conv2d_16_source_29_pat_count_1[24:23] }), .Y(_12165_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37977_ ( .A({ _12166_, _06747_ }), .Y(_06749_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37978_ ( .A({ _12173_, _12167_, _12155_ }), .Y(_12166_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37979_ ( .A({ _12172_, _12170_, _12168_ }), .Y(_12167_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37980_ ( .A({ _12169_, _source_stream_conv2d_16_source_29_pat_count_2[17], _source_stream_conv2d_16_source_29_pat_count_2[14], _source_stream_conv2d_16_source_29_pat_count_2[4] }), .Y(_12168_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37981_ ( .A({ _source_stream_conv2d_16_source_29_pat_count_2[21], _source_stream_conv2d_16_source_29_pat_count_2[18], _source_stream_conv2d_16_source_29_pat_count_2[16:15] }), .Y(_12169_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _37982_ ( .A({ _12171_, _source_stream_conv2d_16_source_29_pat_count_2[27], _source_stream_conv2d_16_source_29_pat_count_2[20], _source_stream_conv2d_16_source_29_pat_count_2[1] }), .Y(_12170_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37983_ ( .A({ _source_stream_conv2d_16_source_29_pat_count_2[28], _source_stream_conv2d_16_source_29_pat_count_2[22], _source_stream_conv2d_16_source_29_pat_count_2[19], _source_stream_conv2d_16_source_29_pat_count_2[3] }), .Y(_12171_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37984_ ( .A({ _source_stream_conv2d_16_source_29_pat_count_2[12:11], _source_stream_conv2d_16_source_29_pat_count_2[9], _source_stream_conv2d_16_source_29_pat_count_2[6] }), .Y(_12172_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37985_ ( .A({ _12177_, _12174_, _source_stream_conv2d_16_source_29_pat_count_2[2], _source_stream_conv2d_16_source_29_pat_count_2[0] }), .Y(_12173_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37986_ ( .A({ _12176_, _12175_, _source_stream_conv2d_16_source_29_pat_count_2[10], _source_stream_conv2d_16_source_29_pat_count_2[5] }), .Y(_12174_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _37987_ ( .A(_source_stream_conv2d_16_source_29_pat_count_2[25:23]), .Y(_12175_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _37988_ ( .A({ _source_stream_conv2d_16_source_29_pat_count_2[13], _source_stream_conv2d_16_source_29_pat_count_2[8:7] }), .Y(_12176_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _37989_ ( .A({ _12178_, _source_stream_conv2d_16_source_29_pat_count_2[29], _source_stream_conv2d_16_source_29_pat_count_2[26] }), .Y(_12177_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _37990_ ( .A(_source_stream_conv2d_16_source_29_pat_count_2[32:30]), .Y(_12178_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _37991_ ( .A({ _12179_, _06749_ }), .Y(_06750_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _37992_ ( .A({ _12189_, _12187_, _12180_ }), .Y(_12179_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _37993_ ( .A({ _12186_, _12181_, _source_stream_conv2d_16_source_29_pat_count_3[1:0] }), .Y(_12180_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _37994_ ( .A({ _12185_, _12184_, _12183_, _12182_ }), .Y(_12181_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37995_ ( .A(_source_stream_conv2d_16_source_29_pat_count_3[13:10]), .Y(_12182_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37996_ ( .A(_source_stream_conv2d_16_source_29_pat_count_3[9:6]), .Y(_12183_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37997_ ( .A(_source_stream_conv2d_16_source_29_pat_count_3[21:18]), .Y(_12184_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37998_ ( .A(_source_stream_conv2d_16_source_29_pat_count_3[17:14]), .Y(_12185_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _37999_ ( .A(_source_stream_conv2d_16_source_29_pat_count_3[5:2]), .Y(_12186_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38000_ ( .A({ _12188_, _source_stream_conv2d_16_source_29_pat_count_3[32:30] }), .Y(_12187_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38001_ ( .A({ _source_stream_conv2d_16_source_29_pat_count_3[28:27], _source_stream_conv2d_16_source_29_pat_count_3[25], _source_stream_conv2d_16_source_29_pat_count_3[22] }), .Y(_12188_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38002_ ( .A({ _source_stream_conv2d_16_source_29_pat_count_3[29], _source_stream_conv2d_16_source_29_pat_count_3[26], _source_stream_conv2d_16_source_29_pat_count_3[24:23] }), .Y(_12189_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38003_ ( .A({ _12190_, _05960_ }), .Y(_06752_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38004_ ( .A({ _12200_, _12199_, _12198_, _12191_ }), .Y(_12190_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38005_ ( .A({ _12197_, _12192_, _source_stream_conv2d_16_source_30_pat_count_0[1:0] }), .Y(_12191_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38006_ ( .A({ _12196_, _12195_, _12194_, _12193_ }), .Y(_12192_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38007_ ( .A(_source_stream_conv2d_16_source_30_pat_count_0[13:10]), .Y(_12193_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38008_ ( .A(_source_stream_conv2d_16_source_30_pat_count_0[9:6]), .Y(_12194_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38009_ ( .A(_source_stream_conv2d_16_source_30_pat_count_0[21:18]), .Y(_12195_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38010_ ( .A(_source_stream_conv2d_16_source_30_pat_count_0[17:14]), .Y(_12196_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38011_ ( .A(_source_stream_conv2d_16_source_30_pat_count_0[5:2]), .Y(_12197_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38012_ ( .A(_source_stream_conv2d_16_source_30_pat_count_0[32:30]), .Y(_12198_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38013_ ( .A(_source_stream_conv2d_16_source_30_pat_count_0[29:26]), .Y(_12199_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38014_ ( .A(_source_stream_conv2d_16_source_30_pat_count_0[25:22]), .Y(_12200_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38015_ ( .A({ _12201_, _06752_ }), .Y(_06753_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38016_ ( .A({ _12211_, _12209_, _12202_ }), .Y(_12201_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38017_ ( .A({ _12208_, _12203_, _source_stream_conv2d_16_source_30_pat_count_1[1:0] }), .Y(_12202_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38018_ ( .A({ _12207_, _12206_, _12205_, _12204_ }), .Y(_12203_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38019_ ( .A(_source_stream_conv2d_16_source_30_pat_count_1[13:10]), .Y(_12204_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38020_ ( .A(_source_stream_conv2d_16_source_30_pat_count_1[9:6]), .Y(_12205_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38021_ ( .A(_source_stream_conv2d_16_source_30_pat_count_1[21:18]), .Y(_12206_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38022_ ( .A(_source_stream_conv2d_16_source_30_pat_count_1[17:14]), .Y(_12207_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38023_ ( .A(_source_stream_conv2d_16_source_30_pat_count_1[5:2]), .Y(_12208_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38024_ ( .A({ _12210_, _source_stream_conv2d_16_source_30_pat_count_1[32:30] }), .Y(_12209_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38025_ ( .A({ _source_stream_conv2d_16_source_30_pat_count_1[28:27], _source_stream_conv2d_16_source_30_pat_count_1[25], _source_stream_conv2d_16_source_30_pat_count_1[22] }), .Y(_12210_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38026_ ( .A({ _source_stream_conv2d_16_source_30_pat_count_1[29], _source_stream_conv2d_16_source_30_pat_count_1[26], _source_stream_conv2d_16_source_30_pat_count_1[24:23] }), .Y(_12211_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38027_ ( .A({ _12212_, _06752_ }), .Y(_06754_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38028_ ( .A({ _12222_, _12219_, _12213_, _12201_ }), .Y(_12212_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38029_ ( .A({ _12218_, _12216_, _12214_ }), .Y(_12213_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38030_ ( .A({ _12215_, _source_stream_conv2d_16_source_30_pat_count_2[17], _source_stream_conv2d_16_source_30_pat_count_2[14], _source_stream_conv2d_16_source_30_pat_count_2[4] }), .Y(_12214_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38031_ ( .A({ _source_stream_conv2d_16_source_30_pat_count_2[21], _source_stream_conv2d_16_source_30_pat_count_2[18], _source_stream_conv2d_16_source_30_pat_count_2[16:15] }), .Y(_12215_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38032_ ( .A({ _12217_, _source_stream_conv2d_16_source_30_pat_count_2[10], _source_stream_conv2d_16_source_30_pat_count_2[5] }), .Y(_12216_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38033_ ( .A({ _source_stream_conv2d_16_source_30_pat_count_2[13], _source_stream_conv2d_16_source_30_pat_count_2[8:7] }), .Y(_12217_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38034_ ( .A({ _source_stream_conv2d_16_source_30_pat_count_2[12:11], _source_stream_conv2d_16_source_30_pat_count_2[9], _source_stream_conv2d_16_source_30_pat_count_2[6] }), .Y(_12218_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38035_ ( .A({ _12220_, _source_stream_conv2d_16_source_30_pat_count_2[2], _source_stream_conv2d_16_source_30_pat_count_2[0] }), .Y(_12219_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38036_ ( .A({ _12221_, _source_stream_conv2d_16_source_30_pat_count_2[29], _source_stream_conv2d_16_source_30_pat_count_2[26] }), .Y(_12220_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38037_ ( .A(_source_stream_conv2d_16_source_30_pat_count_2[32:30]), .Y(_12221_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38038_ ( .A({ _12223_, _source_stream_conv2d_16_source_30_pat_count_2[25:23] }), .Y(_12222_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38039_ ( .A({ _12224_, _source_stream_conv2d_16_source_30_pat_count_2[27], _source_stream_conv2d_16_source_30_pat_count_2[20], _source_stream_conv2d_16_source_30_pat_count_2[1] }), .Y(_12223_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38040_ ( .A({ _source_stream_conv2d_16_source_30_pat_count_2[28], _source_stream_conv2d_16_source_30_pat_count_2[22], _source_stream_conv2d_16_source_30_pat_count_2[19], _source_stream_conv2d_16_source_30_pat_count_2[3] }), .Y(_12224_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38041_ ( .A({ _12225_, _06754_ }), .Y(_06755_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38042_ ( .A({ _12235_, _12233_, _12226_ }), .Y(_12225_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38043_ ( .A({ _12232_, _12227_, _source_stream_conv2d_16_source_30_pat_count_3[1:0] }), .Y(_12226_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38044_ ( .A({ _12231_, _12230_, _12229_, _12228_ }), .Y(_12227_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38045_ ( .A(_source_stream_conv2d_16_source_30_pat_count_3[13:10]), .Y(_12228_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38046_ ( .A(_source_stream_conv2d_16_source_30_pat_count_3[9:6]), .Y(_12229_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38047_ ( .A(_source_stream_conv2d_16_source_30_pat_count_3[21:18]), .Y(_12230_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38048_ ( .A(_source_stream_conv2d_16_source_30_pat_count_3[17:14]), .Y(_12231_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38049_ ( .A(_source_stream_conv2d_16_source_30_pat_count_3[5:2]), .Y(_12232_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38050_ ( .A({ _12234_, _source_stream_conv2d_16_source_30_pat_count_3[32:30] }), .Y(_12233_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38051_ ( .A({ _source_stream_conv2d_16_source_30_pat_count_3[28:27], _source_stream_conv2d_16_source_30_pat_count_3[25], _source_stream_conv2d_16_source_30_pat_count_3[22] }), .Y(_12234_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38052_ ( .A({ _source_stream_conv2d_16_source_30_pat_count_3[29], _source_stream_conv2d_16_source_30_pat_count_3[26], _source_stream_conv2d_16_source_30_pat_count_3[24:23] }), .Y(_12235_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38053_ ( .A({ _12236_, _05962_ }), .Y(_06757_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38054_ ( .A({ _12246_, _12245_, _12244_, _12237_ }), .Y(_12236_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38055_ ( .A({ _12243_, _12238_, _source_stream_conv2d_16_source_31_pat_count_0[1:0] }), .Y(_12237_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38056_ ( .A({ _12242_, _12241_, _12240_, _12239_ }), .Y(_12238_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38057_ ( .A(_source_stream_conv2d_16_source_31_pat_count_0[13:10]), .Y(_12239_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38058_ ( .A(_source_stream_conv2d_16_source_31_pat_count_0[9:6]), .Y(_12240_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38059_ ( .A(_source_stream_conv2d_16_source_31_pat_count_0[21:18]), .Y(_12241_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38060_ ( .A(_source_stream_conv2d_16_source_31_pat_count_0[17:14]), .Y(_12242_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38061_ ( .A(_source_stream_conv2d_16_source_31_pat_count_0[5:2]), .Y(_12243_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38062_ ( .A(_source_stream_conv2d_16_source_31_pat_count_0[32:30]), .Y(_12244_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38063_ ( .A(_source_stream_conv2d_16_source_31_pat_count_0[29:26]), .Y(_12245_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38064_ ( .A(_source_stream_conv2d_16_source_31_pat_count_0[25:22]), .Y(_12246_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38065_ ( .A({ _12247_, _06757_ }), .Y(_06758_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38066_ ( .A({ _12257_, _12255_, _12248_ }), .Y(_12247_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38067_ ( .A({ _12254_, _12249_, _source_stream_conv2d_16_source_31_pat_count_1[1:0] }), .Y(_12248_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38068_ ( .A({ _12253_, _12252_, _12251_, _12250_ }), .Y(_12249_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38069_ ( .A(_source_stream_conv2d_16_source_31_pat_count_1[13:10]), .Y(_12250_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38070_ ( .A(_source_stream_conv2d_16_source_31_pat_count_1[9:6]), .Y(_12251_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38071_ ( .A(_source_stream_conv2d_16_source_31_pat_count_1[21:18]), .Y(_12252_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38072_ ( .A(_source_stream_conv2d_16_source_31_pat_count_1[17:14]), .Y(_12253_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38073_ ( .A(_source_stream_conv2d_16_source_31_pat_count_1[5:2]), .Y(_12254_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38074_ ( .A({ _12256_, _source_stream_conv2d_16_source_31_pat_count_1[32:30] }), .Y(_12255_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38075_ ( .A({ _source_stream_conv2d_16_source_31_pat_count_1[28:27], _source_stream_conv2d_16_source_31_pat_count_1[25], _source_stream_conv2d_16_source_31_pat_count_1[22] }), .Y(_12256_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38076_ ( .A({ _source_stream_conv2d_16_source_31_pat_count_1[29], _source_stream_conv2d_16_source_31_pat_count_1[26], _source_stream_conv2d_16_source_31_pat_count_1[24:23] }), .Y(_12257_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38077_ ( .A({ _12258_, _06757_ }), .Y(_06759_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38078_ ( .A({ _12268_, _12265_, _12259_, _12247_ }), .Y(_12258_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38079_ ( .A({ _12264_, _12262_, _12260_ }), .Y(_12259_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38080_ ( .A({ _12261_, _source_stream_conv2d_16_source_31_pat_count_2[17], _source_stream_conv2d_16_source_31_pat_count_2[14], _source_stream_conv2d_16_source_31_pat_count_2[4] }), .Y(_12260_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38081_ ( .A({ _source_stream_conv2d_16_source_31_pat_count_2[21], _source_stream_conv2d_16_source_31_pat_count_2[18], _source_stream_conv2d_16_source_31_pat_count_2[16:15] }), .Y(_12261_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38082_ ( .A({ _12263_, _source_stream_conv2d_16_source_31_pat_count_2[10], _source_stream_conv2d_16_source_31_pat_count_2[5] }), .Y(_12262_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38083_ ( .A({ _source_stream_conv2d_16_source_31_pat_count_2[13], _source_stream_conv2d_16_source_31_pat_count_2[8:7] }), .Y(_12263_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38084_ ( .A({ _source_stream_conv2d_16_source_31_pat_count_2[12:11], _source_stream_conv2d_16_source_31_pat_count_2[9], _source_stream_conv2d_16_source_31_pat_count_2[6] }), .Y(_12264_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38085_ ( .A({ _12266_, _source_stream_conv2d_16_source_31_pat_count_2[2], _source_stream_conv2d_16_source_31_pat_count_2[0] }), .Y(_12265_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38086_ ( .A({ _12267_, _source_stream_conv2d_16_source_31_pat_count_2[29], _source_stream_conv2d_16_source_31_pat_count_2[26] }), .Y(_12266_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38087_ ( .A(_source_stream_conv2d_16_source_31_pat_count_2[32:30]), .Y(_12267_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38088_ ( .A({ _12269_, _source_stream_conv2d_16_source_31_pat_count_2[25:23] }), .Y(_12268_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38089_ ( .A({ _12270_, _source_stream_conv2d_16_source_31_pat_count_2[27], _source_stream_conv2d_16_source_31_pat_count_2[20], _source_stream_conv2d_16_source_31_pat_count_2[1] }), .Y(_12269_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38090_ ( .A({ _source_stream_conv2d_16_source_31_pat_count_2[28], _source_stream_conv2d_16_source_31_pat_count_2[22], _source_stream_conv2d_16_source_31_pat_count_2[19], _source_stream_conv2d_16_source_31_pat_count_2[3] }), .Y(_12270_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38091_ ( .A({ _12271_, _06759_ }), .Y(_06760_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38092_ ( .A({ _12281_, _12279_, _12272_ }), .Y(_12271_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38093_ ( .A({ _12278_, _12273_, _source_stream_conv2d_16_source_31_pat_count_3[1:0] }), .Y(_12272_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38094_ ( .A({ _12277_, _12276_, _12275_, _12274_ }), .Y(_12273_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38095_ ( .A(_source_stream_conv2d_16_source_31_pat_count_3[13:10]), .Y(_12274_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38096_ ( .A(_source_stream_conv2d_16_source_31_pat_count_3[9:6]), .Y(_12275_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38097_ ( .A(_source_stream_conv2d_16_source_31_pat_count_3[21:18]), .Y(_12276_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38098_ ( .A(_source_stream_conv2d_16_source_31_pat_count_3[17:14]), .Y(_12277_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38099_ ( .A(_source_stream_conv2d_16_source_31_pat_count_3[5:2]), .Y(_12278_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38100_ ( .A({ _12280_, _source_stream_conv2d_16_source_31_pat_count_3[32:30] }), .Y(_12279_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38101_ ( .A({ _source_stream_conv2d_16_source_31_pat_count_3[28:27], _source_stream_conv2d_16_source_31_pat_count_3[25], _source_stream_conv2d_16_source_31_pat_count_3[22] }), .Y(_12280_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38102_ ( .A({ _source_stream_conv2d_16_source_31_pat_count_3[29], _source_stream_conv2d_16_source_31_pat_count_3[26], _source_stream_conv2d_16_source_31_pat_count_3[24:23] }), .Y(_12281_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38103_ ( .A({ _12282_, _05959_ }), .Y(_06762_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38104_ ( .A({ _12292_, _12291_, _12290_, _12283_ }), .Y(_12282_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38105_ ( .A({ _12289_, _12284_, _source_stream_conv2d_16_source_32_pat_count_0[1:0] }), .Y(_12283_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38106_ ( .A({ _12288_, _12287_, _12286_, _12285_ }), .Y(_12284_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38107_ ( .A(_source_stream_conv2d_16_source_32_pat_count_0[13:10]), .Y(_12285_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38108_ ( .A(_source_stream_conv2d_16_source_32_pat_count_0[9:6]), .Y(_12286_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38109_ ( .A(_source_stream_conv2d_16_source_32_pat_count_0[21:18]), .Y(_12287_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38110_ ( .A(_source_stream_conv2d_16_source_32_pat_count_0[17:14]), .Y(_12288_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38111_ ( .A(_source_stream_conv2d_16_source_32_pat_count_0[5:2]), .Y(_12289_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38112_ ( .A(_source_stream_conv2d_16_source_32_pat_count_0[32:30]), .Y(_12290_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38113_ ( .A(_source_stream_conv2d_16_source_32_pat_count_0[29:26]), .Y(_12291_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38114_ ( .A(_source_stream_conv2d_16_source_32_pat_count_0[25:22]), .Y(_12292_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38115_ ( .A({ _12293_, _05959_ }), .Y(_06763_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38116_ ( .A({ _12303_, _12301_, _12294_, _12282_ }), .Y(_12293_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38117_ ( .A({ _12300_, _12295_, _source_stream_conv2d_16_source_32_pat_count_1[1:0] }), .Y(_12294_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38118_ ( .A({ _12299_, _12298_, _12297_, _12296_ }), .Y(_12295_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38119_ ( .A(_source_stream_conv2d_16_source_32_pat_count_1[13:10]), .Y(_12296_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38120_ ( .A(_source_stream_conv2d_16_source_32_pat_count_1[9:6]), .Y(_12297_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38121_ ( .A(_source_stream_conv2d_16_source_32_pat_count_1[21:18]), .Y(_12298_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38122_ ( .A(_source_stream_conv2d_16_source_32_pat_count_1[17:14]), .Y(_12299_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38123_ ( .A(_source_stream_conv2d_16_source_32_pat_count_1[5:2]), .Y(_12300_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38124_ ( .A({ _12302_, _source_stream_conv2d_16_source_32_pat_count_1[32:30] }), .Y(_12301_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38125_ ( .A({ _source_stream_conv2d_16_source_32_pat_count_1[28:27], _source_stream_conv2d_16_source_32_pat_count_1[25], _source_stream_conv2d_16_source_32_pat_count_1[22] }), .Y(_12302_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38126_ ( .A({ _source_stream_conv2d_16_source_32_pat_count_1[29], _source_stream_conv2d_16_source_32_pat_count_1[26], _source_stream_conv2d_16_source_32_pat_count_1[24:23] }), .Y(_12303_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38127_ ( .A({ _12304_, _06763_ }), .Y(_06764_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38128_ ( .A({ _12314_, _12309_, _12307_, _12305_ }), .Y(_12304_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38129_ ( .A({ _12306_, _source_stream_conv2d_16_source_32_pat_count_2[32:30] }), .Y(_12305_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38130_ ( .A({ _source_stream_conv2d_16_source_32_pat_count_2[28:27], _source_stream_conv2d_16_source_32_pat_count_2[25], _source_stream_conv2d_16_source_32_pat_count_2[22] }), .Y(_12306_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38131_ ( .A({ _12308_, _source_stream_conv2d_16_source_32_pat_count_2[1:0] }), .Y(_12307_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38132_ ( .A(_source_stream_conv2d_16_source_32_pat_count_2[5:2]), .Y(_12308_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38133_ ( .A({ _12313_, _12312_, _12311_, _12310_ }), .Y(_12309_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38134_ ( .A(_source_stream_conv2d_16_source_32_pat_count_2[13:10]), .Y(_12310_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38135_ ( .A(_source_stream_conv2d_16_source_32_pat_count_2[9:6]), .Y(_12311_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38136_ ( .A(_source_stream_conv2d_16_source_32_pat_count_2[21:18]), .Y(_12312_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38137_ ( .A(_source_stream_conv2d_16_source_32_pat_count_2[17:14]), .Y(_12313_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38138_ ( .A({ _source_stream_conv2d_16_source_32_pat_count_2[29], _source_stream_conv2d_16_source_32_pat_count_2[26], _source_stream_conv2d_16_source_32_pat_count_2[24:23] }), .Y(_12314_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38139_ ( .A({ _12315_, _06763_ }), .Y(_06765_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38140_ ( .A({ _12326_, _12325_, _12304_, _12316_ }), .Y(_12315_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38141_ ( .A({ _12324_, _12322_, _12317_ }), .Y(_12316_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38142_ ( .A({ _12321_, _12320_, _12318_ }), .Y(_12317_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38143_ ( .A({ _12319_, _source_stream_conv2d_16_source_32_pat_count_3[1:0] }), .Y(_12318_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38144_ ( .A(_source_stream_conv2d_16_source_32_pat_count_3[5:2]), .Y(_12319_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38145_ ( .A({ _source_stream_conv2d_16_source_32_pat_count_3[13], _source_stream_conv2d_16_source_32_pat_count_3[10], _source_stream_conv2d_16_source_32_pat_count_3[8:7] }), .Y(_12320_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38146_ ( .A({ _source_stream_conv2d_16_source_32_pat_count_3[20:19], _source_stream_conv2d_16_source_32_pat_count_3[17], _source_stream_conv2d_16_source_32_pat_count_3[14] }), .Y(_12321_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38147_ ( .A({ _12323_, _source_stream_conv2d_16_source_32_pat_count_3[32:30] }), .Y(_12322_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38148_ ( .A({ _source_stream_conv2d_16_source_32_pat_count_3[28:27], _source_stream_conv2d_16_source_32_pat_count_3[25], _source_stream_conv2d_16_source_32_pat_count_3[22] }), .Y(_12323_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38149_ ( .A({ _source_stream_conv2d_16_source_32_pat_count_3[29], _source_stream_conv2d_16_source_32_pat_count_3[26], _source_stream_conv2d_16_source_32_pat_count_3[24:23] }), .Y(_12324_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38150_ ( .A({ _source_stream_conv2d_16_source_32_pat_count_3[12:11], _source_stream_conv2d_16_source_32_pat_count_3[9], _source_stream_conv2d_16_source_32_pat_count_3[6] }), .Y(_12325_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38151_ ( .A({ _source_stream_conv2d_16_source_32_pat_count_3[21], _source_stream_conv2d_16_source_32_pat_count_3[18], _source_stream_conv2d_16_source_32_pat_count_3[16:15] }), .Y(_12326_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38152_ ( .A({ _12327_, _05956_ }), .Y(_06767_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38153_ ( .A({ _12337_, _12336_, _12335_, _12328_ }), .Y(_12327_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38154_ ( .A({ _12334_, _12329_, _source_stream_conv2d_16_source_33_pat_count_0[1:0] }), .Y(_12328_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38155_ ( .A({ _12333_, _12332_, _12331_, _12330_ }), .Y(_12329_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38156_ ( .A(_source_stream_conv2d_16_source_33_pat_count_0[13:10]), .Y(_12330_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38157_ ( .A(_source_stream_conv2d_16_source_33_pat_count_0[9:6]), .Y(_12331_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38158_ ( .A(_source_stream_conv2d_16_source_33_pat_count_0[21:18]), .Y(_12332_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38159_ ( .A(_source_stream_conv2d_16_source_33_pat_count_0[17:14]), .Y(_12333_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38160_ ( .A(_source_stream_conv2d_16_source_33_pat_count_0[5:2]), .Y(_12334_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38161_ ( .A(_source_stream_conv2d_16_source_33_pat_count_0[32:30]), .Y(_12335_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38162_ ( .A(_source_stream_conv2d_16_source_33_pat_count_0[29:26]), .Y(_12336_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38163_ ( .A(_source_stream_conv2d_16_source_33_pat_count_0[25:22]), .Y(_12337_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38164_ ( .A({ _12338_, _06767_ }), .Y(_06768_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38165_ ( .A({ _12348_, _12346_, _12339_ }), .Y(_12338_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38166_ ( .A({ _12345_, _12340_, _source_stream_conv2d_16_source_33_pat_count_1[1:0] }), .Y(_12339_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38167_ ( .A({ _12344_, _12343_, _12342_, _12341_ }), .Y(_12340_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38168_ ( .A(_source_stream_conv2d_16_source_33_pat_count_1[13:10]), .Y(_12341_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38169_ ( .A(_source_stream_conv2d_16_source_33_pat_count_1[9:6]), .Y(_12342_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38170_ ( .A(_source_stream_conv2d_16_source_33_pat_count_1[21:18]), .Y(_12343_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38171_ ( .A(_source_stream_conv2d_16_source_33_pat_count_1[17:14]), .Y(_12344_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38172_ ( .A(_source_stream_conv2d_16_source_33_pat_count_1[5:2]), .Y(_12345_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38173_ ( .A({ _12347_, _source_stream_conv2d_16_source_33_pat_count_1[32:30] }), .Y(_12346_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38174_ ( .A({ _source_stream_conv2d_16_source_33_pat_count_1[28:27], _source_stream_conv2d_16_source_33_pat_count_1[25], _source_stream_conv2d_16_source_33_pat_count_1[22] }), .Y(_12347_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38175_ ( .A({ _source_stream_conv2d_16_source_33_pat_count_1[29], _source_stream_conv2d_16_source_33_pat_count_1[26], _source_stream_conv2d_16_source_33_pat_count_1[24:23] }), .Y(_12348_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38176_ ( .A({ _12349_, _06767_ }), .Y(_06769_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38177_ ( .A({ _12350_, _12338_ }), .Y(_12349_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38178_ ( .A({ _12360_, _12359_, _12358_, _12351_ }), .Y(_12350_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38179_ ( .A({ _12357_, _12352_, _source_stream_conv2d_16_source_33_pat_count_2[1:0] }), .Y(_12351_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38180_ ( .A({ _12356_, _12355_, _12354_, _12353_ }), .Y(_12352_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38181_ ( .A(_source_stream_conv2d_16_source_33_pat_count_2[13:10]), .Y(_12353_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38182_ ( .A(_source_stream_conv2d_16_source_33_pat_count_2[9:6]), .Y(_12354_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38183_ ( .A(_source_stream_conv2d_16_source_33_pat_count_2[21:18]), .Y(_12355_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38184_ ( .A(_source_stream_conv2d_16_source_33_pat_count_2[17:14]), .Y(_12356_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38185_ ( .A(_source_stream_conv2d_16_source_33_pat_count_2[5:2]), .Y(_12357_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38186_ ( .A(_source_stream_conv2d_16_source_33_pat_count_2[32:30]), .Y(_12358_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38187_ ( .A(_source_stream_conv2d_16_source_33_pat_count_2[29:26]), .Y(_12359_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38188_ ( .A(_source_stream_conv2d_16_source_33_pat_count_2[25:22]), .Y(_12360_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38189_ ( .A({ _12361_, _06769_ }), .Y(_06770_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38190_ ( .A({ _12371_, _12369_, _12362_ }), .Y(_12361_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38191_ ( .A({ _12368_, _12363_, _source_stream_conv2d_16_source_33_pat_count_3[1:0] }), .Y(_12362_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38192_ ( .A({ _12367_, _12366_, _12365_, _12364_ }), .Y(_12363_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38193_ ( .A(_source_stream_conv2d_16_source_33_pat_count_3[13:10]), .Y(_12364_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38194_ ( .A(_source_stream_conv2d_16_source_33_pat_count_3[9:6]), .Y(_12365_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38195_ ( .A(_source_stream_conv2d_16_source_33_pat_count_3[21:18]), .Y(_12366_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38196_ ( .A(_source_stream_conv2d_16_source_33_pat_count_3[17:14]), .Y(_12367_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38197_ ( .A(_source_stream_conv2d_16_source_33_pat_count_3[5:2]), .Y(_12368_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38198_ ( .A({ _12370_, _source_stream_conv2d_16_source_33_pat_count_3[32:30] }), .Y(_12369_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38199_ ( .A({ _source_stream_conv2d_16_source_33_pat_count_3[28:27], _source_stream_conv2d_16_source_33_pat_count_3[25], _source_stream_conv2d_16_source_33_pat_count_3[22] }), .Y(_12370_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38200_ ( .A({ _source_stream_conv2d_16_source_33_pat_count_3[29], _source_stream_conv2d_16_source_33_pat_count_3[26], _source_stream_conv2d_16_source_33_pat_count_3[24:23] }), .Y(_12371_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38201_ ( .A({ _12372_, _05954_ }), .Y(_06772_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38202_ ( .A({ _12382_, _12381_, _12380_, _12373_ }), .Y(_12372_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38203_ ( .A({ _12379_, _12374_, _source_stream_conv2d_16_source_34_pat_count_0[1:0] }), .Y(_12373_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38204_ ( .A({ _12378_, _12377_, _12376_, _12375_ }), .Y(_12374_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38205_ ( .A(_source_stream_conv2d_16_source_34_pat_count_0[13:10]), .Y(_12375_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38206_ ( .A(_source_stream_conv2d_16_source_34_pat_count_0[9:6]), .Y(_12376_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38207_ ( .A(_source_stream_conv2d_16_source_34_pat_count_0[21:18]), .Y(_12377_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38208_ ( .A(_source_stream_conv2d_16_source_34_pat_count_0[17:14]), .Y(_12378_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38209_ ( .A(_source_stream_conv2d_16_source_34_pat_count_0[5:2]), .Y(_12379_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38210_ ( .A(_source_stream_conv2d_16_source_34_pat_count_0[32:30]), .Y(_12380_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38211_ ( .A(_source_stream_conv2d_16_source_34_pat_count_0[29:26]), .Y(_12381_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38212_ ( .A(_source_stream_conv2d_16_source_34_pat_count_0[25:22]), .Y(_12382_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38213_ ( .A({ _12383_, _05954_ }), .Y(_06773_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38214_ ( .A({ _12393_, _12391_, _12384_, _12372_ }), .Y(_12383_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38215_ ( .A({ _12390_, _12385_, _source_stream_conv2d_16_source_34_pat_count_1[1:0] }), .Y(_12384_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38216_ ( .A({ _12389_, _12388_, _12387_, _12386_ }), .Y(_12385_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38217_ ( .A(_source_stream_conv2d_16_source_34_pat_count_1[13:10]), .Y(_12386_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38218_ ( .A(_source_stream_conv2d_16_source_34_pat_count_1[9:6]), .Y(_12387_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38219_ ( .A(_source_stream_conv2d_16_source_34_pat_count_1[21:18]), .Y(_12388_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38220_ ( .A(_source_stream_conv2d_16_source_34_pat_count_1[17:14]), .Y(_12389_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38221_ ( .A(_source_stream_conv2d_16_source_34_pat_count_1[5:2]), .Y(_12390_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38222_ ( .A({ _12392_, _source_stream_conv2d_16_source_34_pat_count_1[32:30] }), .Y(_12391_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38223_ ( .A({ _source_stream_conv2d_16_source_34_pat_count_1[28:27], _source_stream_conv2d_16_source_34_pat_count_1[25], _source_stream_conv2d_16_source_34_pat_count_1[22] }), .Y(_12392_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38224_ ( .A({ _source_stream_conv2d_16_source_34_pat_count_1[29], _source_stream_conv2d_16_source_34_pat_count_1[26], _source_stream_conv2d_16_source_34_pat_count_1[24:23] }), .Y(_12393_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38225_ ( .A({ _12394_, _06773_ }), .Y(_06774_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38226_ ( .A({ _12404_, _12399_, _12397_, _12395_ }), .Y(_12394_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38227_ ( .A({ _12396_, _source_stream_conv2d_16_source_34_pat_count_2[32:30] }), .Y(_12395_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38228_ ( .A({ _source_stream_conv2d_16_source_34_pat_count_2[28:27], _source_stream_conv2d_16_source_34_pat_count_2[25], _source_stream_conv2d_16_source_34_pat_count_2[22] }), .Y(_12396_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38229_ ( .A({ _12398_, _source_stream_conv2d_16_source_34_pat_count_2[1:0] }), .Y(_12397_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38230_ ( .A(_source_stream_conv2d_16_source_34_pat_count_2[5:2]), .Y(_12398_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38231_ ( .A({ _12403_, _12402_, _12401_, _12400_ }), .Y(_12399_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38232_ ( .A(_source_stream_conv2d_16_source_34_pat_count_2[13:10]), .Y(_12400_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38233_ ( .A(_source_stream_conv2d_16_source_34_pat_count_2[9:6]), .Y(_12401_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38234_ ( .A(_source_stream_conv2d_16_source_34_pat_count_2[21:18]), .Y(_12402_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38235_ ( .A(_source_stream_conv2d_16_source_34_pat_count_2[17:14]), .Y(_12403_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38236_ ( .A({ _source_stream_conv2d_16_source_34_pat_count_2[29], _source_stream_conv2d_16_source_34_pat_count_2[26], _source_stream_conv2d_16_source_34_pat_count_2[24:23] }), .Y(_12404_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38237_ ( .A({ _12405_, _06773_ }), .Y(_06775_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38238_ ( .A({ _12416_, _12415_, _12394_, _12406_ }), .Y(_12405_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38239_ ( .A({ _12414_, _12412_, _12407_ }), .Y(_12406_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38240_ ( .A({ _12411_, _12410_, _12408_ }), .Y(_12407_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38241_ ( .A({ _12409_, _source_stream_conv2d_16_source_34_pat_count_3[1:0] }), .Y(_12408_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38242_ ( .A(_source_stream_conv2d_16_source_34_pat_count_3[5:2]), .Y(_12409_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38243_ ( .A({ _source_stream_conv2d_16_source_34_pat_count_3[13], _source_stream_conv2d_16_source_34_pat_count_3[10], _source_stream_conv2d_16_source_34_pat_count_3[8:7] }), .Y(_12410_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38244_ ( .A({ _source_stream_conv2d_16_source_34_pat_count_3[20:19], _source_stream_conv2d_16_source_34_pat_count_3[17], _source_stream_conv2d_16_source_34_pat_count_3[14] }), .Y(_12411_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38245_ ( .A({ _12413_, _source_stream_conv2d_16_source_34_pat_count_3[32:30] }), .Y(_12412_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38246_ ( .A({ _source_stream_conv2d_16_source_34_pat_count_3[28:27], _source_stream_conv2d_16_source_34_pat_count_3[25], _source_stream_conv2d_16_source_34_pat_count_3[22] }), .Y(_12413_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38247_ ( .A({ _source_stream_conv2d_16_source_34_pat_count_3[29], _source_stream_conv2d_16_source_34_pat_count_3[26], _source_stream_conv2d_16_source_34_pat_count_3[24:23] }), .Y(_12414_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38248_ ( .A({ _source_stream_conv2d_16_source_34_pat_count_3[12:11], _source_stream_conv2d_16_source_34_pat_count_3[9], _source_stream_conv2d_16_source_34_pat_count_3[6] }), .Y(_12415_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38249_ ( .A({ _source_stream_conv2d_16_source_34_pat_count_3[21], _source_stream_conv2d_16_source_34_pat_count_3[18], _source_stream_conv2d_16_source_34_pat_count_3[16:15] }), .Y(_12416_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38250_ ( .A({ _12417_, _05952_ }), .Y(_06777_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38251_ ( .A({ _12427_, _12426_, _12425_, _12418_ }), .Y(_12417_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38252_ ( .A({ _12424_, _12419_, _source_stream_conv2d_16_source_35_pat_count_0[1:0] }), .Y(_12418_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38253_ ( .A({ _12423_, _12422_, _12421_, _12420_ }), .Y(_12419_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38254_ ( .A(_source_stream_conv2d_16_source_35_pat_count_0[13:10]), .Y(_12420_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38255_ ( .A(_source_stream_conv2d_16_source_35_pat_count_0[9:6]), .Y(_12421_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38256_ ( .A(_source_stream_conv2d_16_source_35_pat_count_0[21:18]), .Y(_12422_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38257_ ( .A(_source_stream_conv2d_16_source_35_pat_count_0[17:14]), .Y(_12423_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38258_ ( .A(_source_stream_conv2d_16_source_35_pat_count_0[5:2]), .Y(_12424_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38259_ ( .A(_source_stream_conv2d_16_source_35_pat_count_0[32:30]), .Y(_12425_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38260_ ( .A(_source_stream_conv2d_16_source_35_pat_count_0[29:26]), .Y(_12426_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38261_ ( .A(_source_stream_conv2d_16_source_35_pat_count_0[25:22]), .Y(_12427_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38262_ ( .A({ _12428_, _06777_ }), .Y(_06778_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38263_ ( .A({ _12438_, _12436_, _12429_ }), .Y(_12428_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38264_ ( .A({ _12435_, _12430_, _source_stream_conv2d_16_source_35_pat_count_1[1:0] }), .Y(_12429_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38265_ ( .A({ _12434_, _12433_, _12432_, _12431_ }), .Y(_12430_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38266_ ( .A(_source_stream_conv2d_16_source_35_pat_count_1[13:10]), .Y(_12431_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38267_ ( .A(_source_stream_conv2d_16_source_35_pat_count_1[9:6]), .Y(_12432_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38268_ ( .A(_source_stream_conv2d_16_source_35_pat_count_1[21:18]), .Y(_12433_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38269_ ( .A(_source_stream_conv2d_16_source_35_pat_count_1[17:14]), .Y(_12434_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38270_ ( .A(_source_stream_conv2d_16_source_35_pat_count_1[5:2]), .Y(_12435_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38271_ ( .A({ _12437_, _source_stream_conv2d_16_source_35_pat_count_1[32:30] }), .Y(_12436_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38272_ ( .A({ _source_stream_conv2d_16_source_35_pat_count_1[28:27], _source_stream_conv2d_16_source_35_pat_count_1[25], _source_stream_conv2d_16_source_35_pat_count_1[22] }), .Y(_12437_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38273_ ( .A({ _source_stream_conv2d_16_source_35_pat_count_1[29], _source_stream_conv2d_16_source_35_pat_count_1[26], _source_stream_conv2d_16_source_35_pat_count_1[24:23] }), .Y(_12438_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38274_ ( .A({ _12439_, _06777_ }), .Y(_06779_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38275_ ( .A({ _12440_, _12428_ }), .Y(_12439_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38276_ ( .A({ _12450_, _12449_, _12448_, _12441_ }), .Y(_12440_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38277_ ( .A({ _12447_, _12442_, _source_stream_conv2d_16_source_35_pat_count_2[1:0] }), .Y(_12441_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38278_ ( .A({ _12446_, _12445_, _12444_, _12443_ }), .Y(_12442_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38279_ ( .A(_source_stream_conv2d_16_source_35_pat_count_2[13:10]), .Y(_12443_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38280_ ( .A(_source_stream_conv2d_16_source_35_pat_count_2[9:6]), .Y(_12444_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38281_ ( .A(_source_stream_conv2d_16_source_35_pat_count_2[21:18]), .Y(_12445_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38282_ ( .A(_source_stream_conv2d_16_source_35_pat_count_2[17:14]), .Y(_12446_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38283_ ( .A(_source_stream_conv2d_16_source_35_pat_count_2[5:2]), .Y(_12447_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38284_ ( .A(_source_stream_conv2d_16_source_35_pat_count_2[32:30]), .Y(_12448_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38285_ ( .A(_source_stream_conv2d_16_source_35_pat_count_2[29:26]), .Y(_12449_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38286_ ( .A(_source_stream_conv2d_16_source_35_pat_count_2[25:22]), .Y(_12450_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38287_ ( .A({ _12451_, _06779_ }), .Y(_06780_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38288_ ( .A({ _12461_, _12459_, _12452_ }), .Y(_12451_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38289_ ( .A({ _12458_, _12453_, _source_stream_conv2d_16_source_35_pat_count_3[1:0] }), .Y(_12452_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38290_ ( .A({ _12457_, _12456_, _12455_, _12454_ }), .Y(_12453_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38291_ ( .A(_source_stream_conv2d_16_source_35_pat_count_3[13:10]), .Y(_12454_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38292_ ( .A(_source_stream_conv2d_16_source_35_pat_count_3[9:6]), .Y(_12455_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38293_ ( .A(_source_stream_conv2d_16_source_35_pat_count_3[21:18]), .Y(_12456_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38294_ ( .A(_source_stream_conv2d_16_source_35_pat_count_3[17:14]), .Y(_12457_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38295_ ( .A(_source_stream_conv2d_16_source_35_pat_count_3[5:2]), .Y(_12458_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38296_ ( .A({ _12460_, _source_stream_conv2d_16_source_35_pat_count_3[32:30] }), .Y(_12459_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38297_ ( .A({ _source_stream_conv2d_16_source_35_pat_count_3[28:27], _source_stream_conv2d_16_source_35_pat_count_3[25], _source_stream_conv2d_16_source_35_pat_count_3[22] }), .Y(_12460_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38298_ ( .A({ _source_stream_conv2d_16_source_35_pat_count_3[29], _source_stream_conv2d_16_source_35_pat_count_3[26], _source_stream_conv2d_16_source_35_pat_count_3[24:23] }), .Y(_12461_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38299_ ( .A({ _12462_, _05949_ }), .Y(_06782_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38300_ ( .A({ _12472_, _12471_, _12470_, _12463_ }), .Y(_12462_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38301_ ( .A({ _12469_, _12464_, _source_stream_conv2d_16_source_36_pat_count_0[1:0] }), .Y(_12463_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38302_ ( .A({ _12468_, _12467_, _12466_, _12465_ }), .Y(_12464_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38303_ ( .A(_source_stream_conv2d_16_source_36_pat_count_0[13:10]), .Y(_12465_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38304_ ( .A(_source_stream_conv2d_16_source_36_pat_count_0[9:6]), .Y(_12466_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38305_ ( .A(_source_stream_conv2d_16_source_36_pat_count_0[21:18]), .Y(_12467_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38306_ ( .A(_source_stream_conv2d_16_source_36_pat_count_0[17:14]), .Y(_12468_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38307_ ( .A(_source_stream_conv2d_16_source_36_pat_count_0[5:2]), .Y(_12469_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38308_ ( .A(_source_stream_conv2d_16_source_36_pat_count_0[32:30]), .Y(_12470_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38309_ ( .A(_source_stream_conv2d_16_source_36_pat_count_0[29:26]), .Y(_12471_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38310_ ( .A(_source_stream_conv2d_16_source_36_pat_count_0[25:22]), .Y(_12472_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38311_ ( .A({ _12473_, _06782_ }), .Y(_06783_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38312_ ( .A({ _12483_, _12481_, _12474_ }), .Y(_12473_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38313_ ( .A({ _12480_, _12475_, _source_stream_conv2d_16_source_36_pat_count_1[1:0] }), .Y(_12474_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38314_ ( .A({ _12479_, _12478_, _12477_, _12476_ }), .Y(_12475_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38315_ ( .A(_source_stream_conv2d_16_source_36_pat_count_1[13:10]), .Y(_12476_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38316_ ( .A(_source_stream_conv2d_16_source_36_pat_count_1[9:6]), .Y(_12477_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38317_ ( .A(_source_stream_conv2d_16_source_36_pat_count_1[21:18]), .Y(_12478_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38318_ ( .A(_source_stream_conv2d_16_source_36_pat_count_1[17:14]), .Y(_12479_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38319_ ( .A(_source_stream_conv2d_16_source_36_pat_count_1[5:2]), .Y(_12480_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38320_ ( .A({ _12482_, _source_stream_conv2d_16_source_36_pat_count_1[32:30] }), .Y(_12481_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38321_ ( .A({ _source_stream_conv2d_16_source_36_pat_count_1[28:27], _source_stream_conv2d_16_source_36_pat_count_1[25], _source_stream_conv2d_16_source_36_pat_count_1[22] }), .Y(_12482_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38322_ ( .A({ _source_stream_conv2d_16_source_36_pat_count_1[29], _source_stream_conv2d_16_source_36_pat_count_1[26], _source_stream_conv2d_16_source_36_pat_count_1[24:23] }), .Y(_12483_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38323_ ( .A({ _12484_, _06782_ }), .Y(_06784_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38324_ ( .A({ _12494_, _12491_, _12485_, _12473_ }), .Y(_12484_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38325_ ( .A({ _12490_, _12488_, _12486_ }), .Y(_12485_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38326_ ( .A({ _12487_, _source_stream_conv2d_16_source_36_pat_count_2[17], _source_stream_conv2d_16_source_36_pat_count_2[14], _source_stream_conv2d_16_source_36_pat_count_2[4] }), .Y(_12486_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38327_ ( .A({ _source_stream_conv2d_16_source_36_pat_count_2[21], _source_stream_conv2d_16_source_36_pat_count_2[18], _source_stream_conv2d_16_source_36_pat_count_2[16:15] }), .Y(_12487_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38328_ ( .A({ _12489_, _source_stream_conv2d_16_source_36_pat_count_2[10], _source_stream_conv2d_16_source_36_pat_count_2[5] }), .Y(_12488_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38329_ ( .A({ _source_stream_conv2d_16_source_36_pat_count_2[13], _source_stream_conv2d_16_source_36_pat_count_2[8:7] }), .Y(_12489_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38330_ ( .A({ _source_stream_conv2d_16_source_36_pat_count_2[12:11], _source_stream_conv2d_16_source_36_pat_count_2[9], _source_stream_conv2d_16_source_36_pat_count_2[6] }), .Y(_12490_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38331_ ( .A({ _12492_, _source_stream_conv2d_16_source_36_pat_count_2[2], _source_stream_conv2d_16_source_36_pat_count_2[0] }), .Y(_12491_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38332_ ( .A({ _12493_, _source_stream_conv2d_16_source_36_pat_count_2[29], _source_stream_conv2d_16_source_36_pat_count_2[26] }), .Y(_12492_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38333_ ( .A(_source_stream_conv2d_16_source_36_pat_count_2[32:30]), .Y(_12493_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38334_ ( .A({ _12495_, _source_stream_conv2d_16_source_36_pat_count_2[25:23] }), .Y(_12494_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38335_ ( .A({ _12496_, _source_stream_conv2d_16_source_36_pat_count_2[27], _source_stream_conv2d_16_source_36_pat_count_2[20], _source_stream_conv2d_16_source_36_pat_count_2[1] }), .Y(_12495_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38336_ ( .A({ _source_stream_conv2d_16_source_36_pat_count_2[28], _source_stream_conv2d_16_source_36_pat_count_2[22], _source_stream_conv2d_16_source_36_pat_count_2[19], _source_stream_conv2d_16_source_36_pat_count_2[3] }), .Y(_12496_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38337_ ( .A({ _12497_, _06784_ }), .Y(_06785_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38338_ ( .A({ _12507_, _12505_, _12498_ }), .Y(_12497_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38339_ ( .A({ _12504_, _12499_, _source_stream_conv2d_16_source_36_pat_count_3[1:0] }), .Y(_12498_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38340_ ( .A({ _12503_, _12502_, _12501_, _12500_ }), .Y(_12499_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38341_ ( .A(_source_stream_conv2d_16_source_36_pat_count_3[13:10]), .Y(_12500_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38342_ ( .A(_source_stream_conv2d_16_source_36_pat_count_3[9:6]), .Y(_12501_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38343_ ( .A(_source_stream_conv2d_16_source_36_pat_count_3[21:18]), .Y(_12502_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38344_ ( .A(_source_stream_conv2d_16_source_36_pat_count_3[17:14]), .Y(_12503_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38345_ ( .A(_source_stream_conv2d_16_source_36_pat_count_3[5:2]), .Y(_12504_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38346_ ( .A({ _12506_, _source_stream_conv2d_16_source_36_pat_count_3[32:30] }), .Y(_12505_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38347_ ( .A({ _source_stream_conv2d_16_source_36_pat_count_3[28:27], _source_stream_conv2d_16_source_36_pat_count_3[25], _source_stream_conv2d_16_source_36_pat_count_3[22] }), .Y(_12506_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38348_ ( .A({ _source_stream_conv2d_16_source_36_pat_count_3[29], _source_stream_conv2d_16_source_36_pat_count_3[26], _source_stream_conv2d_16_source_36_pat_count_3[24:23] }), .Y(_12507_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38349_ ( .A({ __delay_data_1614, _07016_ }), .Y(_06787_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38350_ ( .A({ _stream_conv2d_16_start_flag, _05687_ }), .Y(_tmp_713) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38351_ ( .A({ _12508_, _05932_ }), .Y(_06789_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38352_ ( .A({ _12518_, _12517_, _12516_, _12509_ }), .Y(_12508_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38353_ ( .A({ _12515_, _12510_, _source_stream_max_pool_serial_18_source_1_pat_count_0[1:0] }), .Y(_12509_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38354_ ( .A({ _12514_, _12513_, _12512_, _12511_ }), .Y(_12510_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38355_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_0[13:10]), .Y(_12511_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38356_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_0[9:6]), .Y(_12512_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38357_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_0[21:18]), .Y(_12513_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38358_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_0[17:14]), .Y(_12514_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38359_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_0[5:2]), .Y(_12515_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38360_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_0[32:30]), .Y(_12516_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38361_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_0[29:26]), .Y(_12517_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38362_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_0[25:22]), .Y(_12518_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38363_ ( .A({ _12519_, _06789_ }), .Y(_06790_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38364_ ( .A({ _12529_, _12527_, _12520_ }), .Y(_12519_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38365_ ( .A({ _12526_, _12521_, _source_stream_max_pool_serial_18_source_1_pat_count_1[1:0] }), .Y(_12520_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38366_ ( .A({ _12525_, _12524_, _12523_, _12522_ }), .Y(_12521_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38367_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_1[13:10]), .Y(_12522_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38368_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_1[9:6]), .Y(_12523_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38369_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_1[21:18]), .Y(_12524_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38370_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_1[17:14]), .Y(_12525_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38371_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_1[5:2]), .Y(_12526_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38372_ ( .A({ _12528_, _source_stream_max_pool_serial_18_source_1_pat_count_1[32:30] }), .Y(_12527_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38373_ ( .A({ _source_stream_max_pool_serial_18_source_1_pat_count_1[28:27], _source_stream_max_pool_serial_18_source_1_pat_count_1[25], _source_stream_max_pool_serial_18_source_1_pat_count_1[22] }), .Y(_12528_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38374_ ( .A({ _source_stream_max_pool_serial_18_source_1_pat_count_1[29], _source_stream_max_pool_serial_18_source_1_pat_count_1[26], _source_stream_max_pool_serial_18_source_1_pat_count_1[24:23] }), .Y(_12529_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38375_ ( .A({ _12530_, _12519_, _06789_ }), .Y(_06791_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38376_ ( .A({ _12540_, _12535_, _12533_, _12531_ }), .Y(_12530_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38377_ ( .A({ _12532_, _source_stream_max_pool_serial_18_source_1_pat_count_2[32:30] }), .Y(_12531_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38378_ ( .A({ _source_stream_max_pool_serial_18_source_1_pat_count_2[28:27], _source_stream_max_pool_serial_18_source_1_pat_count_2[25], _source_stream_max_pool_serial_18_source_1_pat_count_2[22] }), .Y(_12532_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38379_ ( .A({ _12534_, _source_stream_max_pool_serial_18_source_1_pat_count_2[1:0] }), .Y(_12533_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38380_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_2[5:2]), .Y(_12534_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38381_ ( .A({ _12539_, _12538_, _12537_, _12536_ }), .Y(_12535_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38382_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_2[13:10]), .Y(_12536_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38383_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_2[9:6]), .Y(_12537_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38384_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_2[21:18]), .Y(_12538_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38385_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_2[17:14]), .Y(_12539_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38386_ ( .A({ _source_stream_max_pool_serial_18_source_1_pat_count_2[29], _source_stream_max_pool_serial_18_source_1_pat_count_2[26], _source_stream_max_pool_serial_18_source_1_pat_count_2[24:23] }), .Y(_12540_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38387_ ( .A({ _06864_, _05932_ }), .Y(_06792_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38388_ ( .A({ _12541_, _12530_, _12519_, _12508_ }), .Y(_06864_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38389_ ( .A({ _12551_, _12546_, _12544_, _12542_ }), .Y(_12541_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38390_ ( .A({ _12543_, _source_stream_max_pool_serial_18_source_1_pat_count_3[32:30] }), .Y(_12542_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38391_ ( .A({ _source_stream_max_pool_serial_18_source_1_pat_count_3[28:27], _source_stream_max_pool_serial_18_source_1_pat_count_3[25], _source_stream_max_pool_serial_18_source_1_pat_count_3[22] }), .Y(_12543_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38392_ ( .A({ _12545_, _source_stream_max_pool_serial_18_source_1_pat_count_3[1:0] }), .Y(_12544_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38393_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_3[5:2]), .Y(_12545_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38394_ ( .A({ _12550_, _12549_, _12548_, _12547_ }), .Y(_12546_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38395_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_3[13:10]), .Y(_12547_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38396_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_3[9:6]), .Y(_12548_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38397_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_3[21:18]), .Y(_12549_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38398_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_3[17:14]), .Y(_12550_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38399_ ( .A({ _source_stream_max_pool_serial_18_source_1_pat_count_3[29], _source_stream_max_pool_serial_18_source_1_pat_count_3[26], _source_stream_max_pool_serial_18_source_1_pat_count_3[24:23] }), .Y(_12551_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38400_ ( .A({ __substreamoutput_data_794, _stream_max_pool_serial_18_sink_3_sink_fsm_1[0], _24040_ }), .Y(_06794_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38401_ ( .A({ _stream_max_pool_serial_18_start_flag, _05686_ }), .Y(_tmp_1040) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38402_ ( .A({ _12552_, _05912_ }), .Y(_06796_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38403_ ( .A({ _12562_, _12561_, _12560_, _12553_ }), .Y(_12552_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38404_ ( .A({ _12559_, _12554_, _source_stream_matmul_29_source_6_pat_count_0[1:0] }), .Y(_12553_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38405_ ( .A({ _12558_, _12557_, _12556_, _12555_ }), .Y(_12554_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38406_ ( .A(_source_stream_matmul_29_source_6_pat_count_0[13:10]), .Y(_12555_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38407_ ( .A(_source_stream_matmul_29_source_6_pat_count_0[9:6]), .Y(_12556_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38408_ ( .A(_source_stream_matmul_29_source_6_pat_count_0[21:18]), .Y(_12557_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38409_ ( .A(_source_stream_matmul_29_source_6_pat_count_0[17:14]), .Y(_12558_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38410_ ( .A(_source_stream_matmul_29_source_6_pat_count_0[5:2]), .Y(_12559_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38411_ ( .A(_source_stream_matmul_29_source_6_pat_count_0[32:30]), .Y(_12560_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38412_ ( .A(_source_stream_matmul_29_source_6_pat_count_0[29:26]), .Y(_12561_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38413_ ( .A(_source_stream_matmul_29_source_6_pat_count_0[25:22]), .Y(_12562_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38414_ ( .A({ _12563_, _06796_ }), .Y(_06797_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38415_ ( .A({ _12573_, _12571_, _12564_ }), .Y(_12563_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38416_ ( .A({ _12570_, _12565_, _source_stream_matmul_29_source_6_pat_count_1[1:0] }), .Y(_12564_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38417_ ( .A({ _12569_, _12568_, _12567_, _12566_ }), .Y(_12565_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38418_ ( .A(_source_stream_matmul_29_source_6_pat_count_1[13:10]), .Y(_12566_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38419_ ( .A(_source_stream_matmul_29_source_6_pat_count_1[9:6]), .Y(_12567_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38420_ ( .A(_source_stream_matmul_29_source_6_pat_count_1[21:18]), .Y(_12568_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38421_ ( .A(_source_stream_matmul_29_source_6_pat_count_1[17:14]), .Y(_12569_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38422_ ( .A(_source_stream_matmul_29_source_6_pat_count_1[5:2]), .Y(_12570_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38423_ ( .A({ _12572_, _source_stream_matmul_29_source_6_pat_count_1[32:30] }), .Y(_12571_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38424_ ( .A({ _source_stream_matmul_29_source_6_pat_count_1[28:27], _source_stream_matmul_29_source_6_pat_count_1[25], _source_stream_matmul_29_source_6_pat_count_1[22] }), .Y(_12572_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38425_ ( .A({ _source_stream_matmul_29_source_6_pat_count_1[29], _source_stream_matmul_29_source_6_pat_count_1[26], _source_stream_matmul_29_source_6_pat_count_1[24:23] }), .Y(_12573_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38426_ ( .A({ _12574_, _06796_ }), .Y(_06798_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38427_ ( .A({ _12584_, _12581_, _12575_, _12563_ }), .Y(_12574_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38428_ ( .A({ _12580_, _12578_, _12576_ }), .Y(_12575_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38429_ ( .A({ _12577_, _source_stream_matmul_29_source_6_pat_count_2[17], _source_stream_matmul_29_source_6_pat_count_2[14], _source_stream_matmul_29_source_6_pat_count_2[4] }), .Y(_12576_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38430_ ( .A({ _source_stream_matmul_29_source_6_pat_count_2[21], _source_stream_matmul_29_source_6_pat_count_2[18], _source_stream_matmul_29_source_6_pat_count_2[16:15] }), .Y(_12577_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38431_ ( .A({ _12579_, _source_stream_matmul_29_source_6_pat_count_2[10], _source_stream_matmul_29_source_6_pat_count_2[5] }), .Y(_12578_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38432_ ( .A({ _source_stream_matmul_29_source_6_pat_count_2[13], _source_stream_matmul_29_source_6_pat_count_2[8:7] }), .Y(_12579_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38433_ ( .A({ _source_stream_matmul_29_source_6_pat_count_2[12:11], _source_stream_matmul_29_source_6_pat_count_2[9], _source_stream_matmul_29_source_6_pat_count_2[6] }), .Y(_12580_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38434_ ( .A({ _12582_, _source_stream_matmul_29_source_6_pat_count_2[2], _source_stream_matmul_29_source_6_pat_count_2[0] }), .Y(_12581_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38435_ ( .A({ _12583_, _source_stream_matmul_29_source_6_pat_count_2[29], _source_stream_matmul_29_source_6_pat_count_2[26] }), .Y(_12582_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38436_ ( .A(_source_stream_matmul_29_source_6_pat_count_2[32:30]), .Y(_12583_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38437_ ( .A({ _12585_, _source_stream_matmul_29_source_6_pat_count_2[25:23] }), .Y(_12584_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38438_ ( .A({ _12586_, _source_stream_matmul_29_source_6_pat_count_2[27], _source_stream_matmul_29_source_6_pat_count_2[20], _source_stream_matmul_29_source_6_pat_count_2[1] }), .Y(_12585_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38439_ ( .A({ _source_stream_matmul_29_source_6_pat_count_2[28], _source_stream_matmul_29_source_6_pat_count_2[22], _source_stream_matmul_29_source_6_pat_count_2[19], _source_stream_matmul_29_source_6_pat_count_2[3] }), .Y(_12586_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38440_ ( .A({ _12587_, _06798_ }), .Y(_06799_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38441_ ( .A({ _12597_, _12595_, _12588_ }), .Y(_12587_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38442_ ( .A({ _12594_, _12589_, _source_stream_matmul_29_source_6_pat_count_3[1:0] }), .Y(_12588_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38443_ ( .A({ _12593_, _12592_, _12591_, _12590_ }), .Y(_12589_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38444_ ( .A(_source_stream_matmul_29_source_6_pat_count_3[13:10]), .Y(_12590_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38445_ ( .A(_source_stream_matmul_29_source_6_pat_count_3[9:6]), .Y(_12591_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38446_ ( .A(_source_stream_matmul_29_source_6_pat_count_3[21:18]), .Y(_12592_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38447_ ( .A(_source_stream_matmul_29_source_6_pat_count_3[17:14]), .Y(_12593_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38448_ ( .A(_source_stream_matmul_29_source_6_pat_count_3[5:2]), .Y(_12594_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38449_ ( .A({ _12596_, _source_stream_matmul_29_source_6_pat_count_3[32:30] }), .Y(_12595_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38450_ ( .A({ _source_stream_matmul_29_source_6_pat_count_3[28:27], _source_stream_matmul_29_source_6_pat_count_3[25], _source_stream_matmul_29_source_6_pat_count_3[22] }), .Y(_12596_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38451_ ( .A({ _source_stream_matmul_29_source_6_pat_count_3[29], _source_stream_matmul_29_source_6_pat_count_3[26], _source_stream_matmul_29_source_6_pat_count_3[24:23] }), .Y(_12597_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38452_ ( .A({ _12598_, _05911_ }), .Y(_06801_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38453_ ( .A({ _12608_, _12607_, _12606_, _12599_ }), .Y(_12598_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38454_ ( .A({ _12605_, _12600_, _source_stream_matmul_29_source_8_pat_count_0[1:0] }), .Y(_12599_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38455_ ( .A({ _12604_, _12603_, _12602_, _12601_ }), .Y(_12600_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38456_ ( .A(_source_stream_matmul_29_source_8_pat_count_0[13:10]), .Y(_12601_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38457_ ( .A(_source_stream_matmul_29_source_8_pat_count_0[9:6]), .Y(_12602_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38458_ ( .A(_source_stream_matmul_29_source_8_pat_count_0[21:18]), .Y(_12603_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38459_ ( .A(_source_stream_matmul_29_source_8_pat_count_0[17:14]), .Y(_12604_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38460_ ( .A(_source_stream_matmul_29_source_8_pat_count_0[5:2]), .Y(_12605_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38461_ ( .A(_source_stream_matmul_29_source_8_pat_count_0[32:30]), .Y(_12606_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38462_ ( .A(_source_stream_matmul_29_source_8_pat_count_0[29:26]), .Y(_12607_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38463_ ( .A(_source_stream_matmul_29_source_8_pat_count_0[25:22]), .Y(_12608_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38464_ ( .A({ _12609_, _06801_ }), .Y(_06802_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38465_ ( .A({ _12619_, _12617_, _12610_ }), .Y(_12609_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38466_ ( .A({ _12616_, _12611_, _source_stream_matmul_29_source_8_pat_count_1[1:0] }), .Y(_12610_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38467_ ( .A({ _12615_, _12614_, _12613_, _12612_ }), .Y(_12611_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38468_ ( .A(_source_stream_matmul_29_source_8_pat_count_1[13:10]), .Y(_12612_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38469_ ( .A(_source_stream_matmul_29_source_8_pat_count_1[9:6]), .Y(_12613_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38470_ ( .A(_source_stream_matmul_29_source_8_pat_count_1[21:18]), .Y(_12614_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38471_ ( .A(_source_stream_matmul_29_source_8_pat_count_1[17:14]), .Y(_12615_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38472_ ( .A(_source_stream_matmul_29_source_8_pat_count_1[5:2]), .Y(_12616_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38473_ ( .A({ _12618_, _source_stream_matmul_29_source_8_pat_count_1[32:30] }), .Y(_12617_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38474_ ( .A({ _source_stream_matmul_29_source_8_pat_count_1[28:27], _source_stream_matmul_29_source_8_pat_count_1[25], _source_stream_matmul_29_source_8_pat_count_1[22] }), .Y(_12618_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38475_ ( .A({ _source_stream_matmul_29_source_8_pat_count_1[29], _source_stream_matmul_29_source_8_pat_count_1[26], _source_stream_matmul_29_source_8_pat_count_1[24:23] }), .Y(_12619_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38476_ ( .A({ _12620_, _06801_ }), .Y(_06803_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38477_ ( .A({ _12630_, _12627_, _12621_, _12609_ }), .Y(_12620_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38478_ ( .A({ _12626_, _12624_, _12622_ }), .Y(_12621_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38479_ ( .A({ _12623_, _source_stream_matmul_29_source_8_pat_count_2[17], _source_stream_matmul_29_source_8_pat_count_2[14], _source_stream_matmul_29_source_8_pat_count_2[4] }), .Y(_12622_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38480_ ( .A({ _source_stream_matmul_29_source_8_pat_count_2[21], _source_stream_matmul_29_source_8_pat_count_2[18], _source_stream_matmul_29_source_8_pat_count_2[16:15] }), .Y(_12623_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38481_ ( .A({ _12625_, _source_stream_matmul_29_source_8_pat_count_2[10], _source_stream_matmul_29_source_8_pat_count_2[5] }), .Y(_12624_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38482_ ( .A({ _source_stream_matmul_29_source_8_pat_count_2[13], _source_stream_matmul_29_source_8_pat_count_2[8:7] }), .Y(_12625_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38483_ ( .A({ _source_stream_matmul_29_source_8_pat_count_2[12:11], _source_stream_matmul_29_source_8_pat_count_2[9], _source_stream_matmul_29_source_8_pat_count_2[6] }), .Y(_12626_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38484_ ( .A({ _12628_, _source_stream_matmul_29_source_8_pat_count_2[2], _source_stream_matmul_29_source_8_pat_count_2[0] }), .Y(_12627_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38485_ ( .A({ _12629_, _source_stream_matmul_29_source_8_pat_count_2[29], _source_stream_matmul_29_source_8_pat_count_2[26] }), .Y(_12628_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38486_ ( .A(_source_stream_matmul_29_source_8_pat_count_2[32:30]), .Y(_12629_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38487_ ( .A({ _12631_, _source_stream_matmul_29_source_8_pat_count_2[25:23] }), .Y(_12630_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38488_ ( .A({ _12632_, _source_stream_matmul_29_source_8_pat_count_2[27], _source_stream_matmul_29_source_8_pat_count_2[20], _source_stream_matmul_29_source_8_pat_count_2[1] }), .Y(_12631_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38489_ ( .A({ _source_stream_matmul_29_source_8_pat_count_2[28], _source_stream_matmul_29_source_8_pat_count_2[22], _source_stream_matmul_29_source_8_pat_count_2[19], _source_stream_matmul_29_source_8_pat_count_2[3] }), .Y(_12632_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38490_ ( .A({ _12633_, _06803_ }), .Y(_06804_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38491_ ( .A({ _12643_, _12641_, _12634_ }), .Y(_12633_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38492_ ( .A({ _12640_, _12635_, _source_stream_matmul_29_source_8_pat_count_3[1:0] }), .Y(_12634_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38493_ ( .A({ _12639_, _12638_, _12637_, _12636_ }), .Y(_12635_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38494_ ( .A(_source_stream_matmul_29_source_8_pat_count_3[13:10]), .Y(_12636_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38495_ ( .A(_source_stream_matmul_29_source_8_pat_count_3[9:6]), .Y(_12637_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38496_ ( .A(_source_stream_matmul_29_source_8_pat_count_3[21:18]), .Y(_12638_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38497_ ( .A(_source_stream_matmul_29_source_8_pat_count_3[17:14]), .Y(_12639_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38498_ ( .A(_source_stream_matmul_29_source_8_pat_count_3[5:2]), .Y(_12640_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38499_ ( .A({ _12642_, _source_stream_matmul_29_source_8_pat_count_3[32:30] }), .Y(_12641_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38500_ ( .A({ _source_stream_matmul_29_source_8_pat_count_3[28:27], _source_stream_matmul_29_source_8_pat_count_3[25], _source_stream_matmul_29_source_8_pat_count_3[22] }), .Y(_12642_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38501_ ( .A({ _source_stream_matmul_29_source_8_pat_count_3[29], _source_stream_matmul_29_source_8_pat_count_3[26], _source_stream_matmul_29_source_8_pat_count_3[24:23] }), .Y(_12643_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38502_ ( .A({ _12644_, _05913_ }), .Y(_06806_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38503_ ( .A({ _12654_, _12653_, _12652_, _12645_ }), .Y(_12644_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38504_ ( .A({ _12651_, _12646_, _source_stream_matmul_29_source_19_pat_count_0[1:0] }), .Y(_12645_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38505_ ( .A({ _12650_, _12649_, _12648_, _12647_ }), .Y(_12646_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38506_ ( .A(_source_stream_matmul_29_source_19_pat_count_0[13:10]), .Y(_12647_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38507_ ( .A(_source_stream_matmul_29_source_19_pat_count_0[9:6]), .Y(_12648_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38508_ ( .A(_source_stream_matmul_29_source_19_pat_count_0[21:18]), .Y(_12649_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38509_ ( .A(_source_stream_matmul_29_source_19_pat_count_0[17:14]), .Y(_12650_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38510_ ( .A(_source_stream_matmul_29_source_19_pat_count_0[5:2]), .Y(_12651_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38511_ ( .A(_source_stream_matmul_29_source_19_pat_count_0[32:30]), .Y(_12652_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38512_ ( .A(_source_stream_matmul_29_source_19_pat_count_0[29:26]), .Y(_12653_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38513_ ( .A(_source_stream_matmul_29_source_19_pat_count_0[25:22]), .Y(_12654_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38514_ ( .A({ _12655_, _06806_ }), .Y(_06807_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38515_ ( .A({ _12665_, _12663_, _12656_ }), .Y(_12655_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38516_ ( .A({ _12662_, _12657_, _source_stream_matmul_29_source_19_pat_count_1[1:0] }), .Y(_12656_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38517_ ( .A({ _12661_, _12660_, _12659_, _12658_ }), .Y(_12657_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38518_ ( .A(_source_stream_matmul_29_source_19_pat_count_1[13:10]), .Y(_12658_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38519_ ( .A(_source_stream_matmul_29_source_19_pat_count_1[9:6]), .Y(_12659_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38520_ ( .A(_source_stream_matmul_29_source_19_pat_count_1[21:18]), .Y(_12660_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38521_ ( .A(_source_stream_matmul_29_source_19_pat_count_1[17:14]), .Y(_12661_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38522_ ( .A(_source_stream_matmul_29_source_19_pat_count_1[5:2]), .Y(_12662_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38523_ ( .A({ _12664_, _source_stream_matmul_29_source_19_pat_count_1[32:30] }), .Y(_12663_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38524_ ( .A({ _source_stream_matmul_29_source_19_pat_count_1[28:27], _source_stream_matmul_29_source_19_pat_count_1[25], _source_stream_matmul_29_source_19_pat_count_1[22] }), .Y(_12664_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38525_ ( .A({ _source_stream_matmul_29_source_19_pat_count_1[29], _source_stream_matmul_29_source_19_pat_count_1[26], _source_stream_matmul_29_source_19_pat_count_1[24:23] }), .Y(_12665_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38526_ ( .A({ _12666_, _06806_ }), .Y(_06808_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38527_ ( .A({ _12676_, _12673_, _12667_, _12655_ }), .Y(_12666_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38528_ ( .A({ _12672_, _12670_, _12668_ }), .Y(_12667_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38529_ ( .A({ _12669_, _source_stream_matmul_29_source_19_pat_count_2[17], _source_stream_matmul_29_source_19_pat_count_2[14], _source_stream_matmul_29_source_19_pat_count_2[4] }), .Y(_12668_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38530_ ( .A({ _source_stream_matmul_29_source_19_pat_count_2[21], _source_stream_matmul_29_source_19_pat_count_2[18], _source_stream_matmul_29_source_19_pat_count_2[16:15] }), .Y(_12669_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38531_ ( .A({ _12671_, _source_stream_matmul_29_source_19_pat_count_2[10], _source_stream_matmul_29_source_19_pat_count_2[5] }), .Y(_12670_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38532_ ( .A({ _source_stream_matmul_29_source_19_pat_count_2[13], _source_stream_matmul_29_source_19_pat_count_2[8:7] }), .Y(_12671_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38533_ ( .A({ _source_stream_matmul_29_source_19_pat_count_2[12:11], _source_stream_matmul_29_source_19_pat_count_2[9], _source_stream_matmul_29_source_19_pat_count_2[6] }), .Y(_12672_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38534_ ( .A({ _12674_, _source_stream_matmul_29_source_19_pat_count_2[2], _source_stream_matmul_29_source_19_pat_count_2[0] }), .Y(_12673_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38535_ ( .A({ _12675_, _source_stream_matmul_29_source_19_pat_count_2[29], _source_stream_matmul_29_source_19_pat_count_2[26] }), .Y(_12674_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38536_ ( .A(_source_stream_matmul_29_source_19_pat_count_2[32:30]), .Y(_12675_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38537_ ( .A({ _12677_, _source_stream_matmul_29_source_19_pat_count_2[25:23] }), .Y(_12676_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38538_ ( .A({ _12678_, _source_stream_matmul_29_source_19_pat_count_2[27], _source_stream_matmul_29_source_19_pat_count_2[20], _source_stream_matmul_29_source_19_pat_count_2[1] }), .Y(_12677_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38539_ ( .A({ _source_stream_matmul_29_source_19_pat_count_2[28], _source_stream_matmul_29_source_19_pat_count_2[22], _source_stream_matmul_29_source_19_pat_count_2[19], _source_stream_matmul_29_source_19_pat_count_2[3] }), .Y(_12678_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38540_ ( .A({ _12679_, _06808_ }), .Y(_06809_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38541_ ( .A({ _12689_, _12687_, _12680_ }), .Y(_12679_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38542_ ( .A({ _12686_, _12681_, _source_stream_matmul_29_source_19_pat_count_3[1:0] }), .Y(_12680_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38543_ ( .A({ _12685_, _12684_, _12683_, _12682_ }), .Y(_12681_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38544_ ( .A(_source_stream_matmul_29_source_19_pat_count_3[13:10]), .Y(_12682_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38545_ ( .A(_source_stream_matmul_29_source_19_pat_count_3[9:6]), .Y(_12683_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38546_ ( .A(_source_stream_matmul_29_source_19_pat_count_3[21:18]), .Y(_12684_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38547_ ( .A(_source_stream_matmul_29_source_19_pat_count_3[17:14]), .Y(_12685_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38548_ ( .A(_source_stream_matmul_29_source_19_pat_count_3[5:2]), .Y(_12686_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38549_ ( .A({ _12688_, _source_stream_matmul_29_source_19_pat_count_3[32:30] }), .Y(_12687_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38550_ ( .A({ _source_stream_matmul_29_source_19_pat_count_3[28:27], _source_stream_matmul_29_source_19_pat_count_3[25], _source_stream_matmul_29_source_19_pat_count_3[22] }), .Y(_12688_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38551_ ( .A({ _source_stream_matmul_29_source_19_pat_count_3[29], _source_stream_matmul_29_source_19_pat_count_3[26], _source_stream_matmul_29_source_19_pat_count_3[24:23] }), .Y(_12689_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38552_ ( .A({ _12690_, _05909_ }), .Y(_06811_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38553_ ( .A({ _12700_, _12695_, _12693_, _12691_ }), .Y(_12690_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38554_ ( .A({ _12692_, _source_stream_matmul_29_source_20_pat_count_0[32:30] }), .Y(_12691_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38555_ ( .A({ _source_stream_matmul_29_source_20_pat_count_0[28:27], _source_stream_matmul_29_source_20_pat_count_0[25], _source_stream_matmul_29_source_20_pat_count_0[22] }), .Y(_12692_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38556_ ( .A({ _12694_, _source_stream_matmul_29_source_20_pat_count_0[1:0] }), .Y(_12693_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38557_ ( .A(_source_stream_matmul_29_source_20_pat_count_0[5:2]), .Y(_12694_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38558_ ( .A({ _12699_, _12698_, _12697_, _12696_ }), .Y(_12695_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38559_ ( .A(_source_stream_matmul_29_source_20_pat_count_0[13:10]), .Y(_12696_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38560_ ( .A(_source_stream_matmul_29_source_20_pat_count_0[9:6]), .Y(_12697_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38561_ ( .A(_source_stream_matmul_29_source_20_pat_count_0[21:18]), .Y(_12698_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38562_ ( .A(_source_stream_matmul_29_source_20_pat_count_0[17:14]), .Y(_12699_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38563_ ( .A({ _source_stream_matmul_29_source_20_pat_count_0[29], _source_stream_matmul_29_source_20_pat_count_0[26], _source_stream_matmul_29_source_20_pat_count_0[24:23] }), .Y(_12700_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38564_ ( .A({ _12701_, _06811_ }), .Y(_06812_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38565_ ( .A({ _12711_, _12709_, _12702_ }), .Y(_12701_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38566_ ( .A({ _12708_, _12703_, _source_stream_matmul_29_source_20_pat_count_1[1:0] }), .Y(_12702_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38567_ ( .A({ _12707_, _12706_, _12705_, _12704_ }), .Y(_12703_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38568_ ( .A(_source_stream_matmul_29_source_20_pat_count_1[13:10]), .Y(_12704_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38569_ ( .A(_source_stream_matmul_29_source_20_pat_count_1[9:6]), .Y(_12705_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38570_ ( .A(_source_stream_matmul_29_source_20_pat_count_1[21:18]), .Y(_12706_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38571_ ( .A(_source_stream_matmul_29_source_20_pat_count_1[17:14]), .Y(_12707_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38572_ ( .A(_source_stream_matmul_29_source_20_pat_count_1[5:2]), .Y(_12708_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38573_ ( .A({ _12710_, _source_stream_matmul_29_source_20_pat_count_1[32:30] }), .Y(_12709_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38574_ ( .A({ _source_stream_matmul_29_source_20_pat_count_1[28:27], _source_stream_matmul_29_source_20_pat_count_1[25], _source_stream_matmul_29_source_20_pat_count_1[22] }), .Y(_12710_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38575_ ( .A({ _source_stream_matmul_29_source_20_pat_count_1[29], _source_stream_matmul_29_source_20_pat_count_1[26], _source_stream_matmul_29_source_20_pat_count_1[24:23] }), .Y(_12711_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38576_ ( .A({ _12712_, _12701_, _06811_ }), .Y(_06813_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38577_ ( .A({ _12722_, _12717_, _12715_, _12713_ }), .Y(_12712_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38578_ ( .A({ _12714_, _source_stream_matmul_29_source_20_pat_count_2[32:30] }), .Y(_12713_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38579_ ( .A({ _source_stream_matmul_29_source_20_pat_count_2[28:27], _source_stream_matmul_29_source_20_pat_count_2[25], _source_stream_matmul_29_source_20_pat_count_2[22] }), .Y(_12714_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38580_ ( .A({ _12716_, _source_stream_matmul_29_source_20_pat_count_2[1:0] }), .Y(_12715_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38581_ ( .A(_source_stream_matmul_29_source_20_pat_count_2[5:2]), .Y(_12716_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38582_ ( .A({ _12721_, _12720_, _12719_, _12718_ }), .Y(_12717_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38583_ ( .A(_source_stream_matmul_29_source_20_pat_count_2[13:10]), .Y(_12718_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38584_ ( .A(_source_stream_matmul_29_source_20_pat_count_2[9:6]), .Y(_12719_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38585_ ( .A(_source_stream_matmul_29_source_20_pat_count_2[21:18]), .Y(_12720_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38586_ ( .A(_source_stream_matmul_29_source_20_pat_count_2[17:14]), .Y(_12721_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38587_ ( .A({ _source_stream_matmul_29_source_20_pat_count_2[29], _source_stream_matmul_29_source_20_pat_count_2[26], _source_stream_matmul_29_source_20_pat_count_2[24:23] }), .Y(_12722_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38588_ ( .A({ _06872_, _05909_ }), .Y(_06814_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38589_ ( .A({ _12723_, _12712_, _12690_, _12701_ }), .Y(_06872_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38590_ ( .A({ _12733_, _12728_, _12726_, _12724_ }), .Y(_12723_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38591_ ( .A({ _12725_, _source_stream_matmul_29_source_20_pat_count_3[32:30] }), .Y(_12724_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38592_ ( .A({ _source_stream_matmul_29_source_20_pat_count_3[28:27], _source_stream_matmul_29_source_20_pat_count_3[25], _source_stream_matmul_29_source_20_pat_count_3[22] }), .Y(_12725_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38593_ ( .A({ _12727_, _source_stream_matmul_29_source_20_pat_count_3[1:0] }), .Y(_12726_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38594_ ( .A(_source_stream_matmul_29_source_20_pat_count_3[5:2]), .Y(_12727_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38595_ ( .A({ _12732_, _12731_, _12730_, _12729_ }), .Y(_12728_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38596_ ( .A(_source_stream_matmul_29_source_20_pat_count_3[13:10]), .Y(_12729_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38597_ ( .A(_source_stream_matmul_29_source_20_pat_count_3[9:6]), .Y(_12730_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38598_ ( .A(_source_stream_matmul_29_source_20_pat_count_3[21:18]), .Y(_12731_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38599_ ( .A(_source_stream_matmul_29_source_20_pat_count_3[17:14]), .Y(_12732_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38600_ ( .A({ _source_stream_matmul_29_source_20_pat_count_3[29], _source_stream_matmul_29_source_20_pat_count_3[26], _source_stream_matmul_29_source_20_pat_count_3[24:23] }), .Y(_12733_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38601_ ( .A({ __delay_data_1616, _stream_matmul_29_sink_21_sink_fsm_4[0], _24030_ }), .Y(_06816_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38602_ ( .A({ _stream_matmul_29_start_flag, _05685_ }), .Y(_tmp_1227) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _38603_ ( .A({ conv2d_16_mux_dma_flag_0, conv2d_16_mux_dma_pad_mask_0 }), .Y(_06879_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _38604_ ( .A({ conv2d_16_mux_dma_flag_1, conv2d_16_mux_dma_pad_mask_1 }), .Y(_06880_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _38605_ ( .A({ conv2d_16_mux_dma_flag_2, conv2d_16_mux_dma_pad_mask_2 }), .Y(_06881_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _38606_ ( .A({ conv2d_16_update_filter, _12734_, _12741_ }), .Y(_06817_) );
  \$lut  #( .LUT(16'hd000), .WIDTH(4) ) _38607_ ( .A({ _12739_, _12740_, _12735_, _04812_ }), .Y(_12734_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38608_ ( .A({ _12738_, _12736_, _04819_, _04808_ }), .Y(_12735_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38609_ ( .A({ _12737_, _04811_, _04810_, _04809_ }), .Y(_12736_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38610_ ( .A({ _04839_, _04838_, _04837_, _04836_ }), .Y(_12737_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38611_ ( .A({ _04835_, _04834_, _04833_, _04830_ }), .Y(_12738_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38612_ ( .A({ _04832_, _04831_, _04829_, _04828_ }), .Y(_12739_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38613_ ( .A({ _04826_, _04825_, _04823_, _04820_ }), .Y(_12740_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38614_ ( .A({ _12743_, _12742_, _04814_, _04813_ }), .Y(_12741_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38615_ ( .A({ _04818_, _04817_, _04816_, _04815_ }), .Y(_12742_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38616_ ( .A({ _04827_, _04824_, _04822_, _04821_ }), .Y(_12743_) );
  \$lut  #( .LUT(16'hbf00), .WIDTH(4) ) _38617_ ( .A({ conv2d_16_mux_next_dma_flag_0, _12748_, _12752_, _12744_ }), .Y(_06818_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _38618_ ( .A({ _04874_, _12745_, _12747_ }), .Y(_12744_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38619_ ( .A({ _12746_, _04873_, _04903_, _04902_ }), .Y(_12745_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38620_ ( .A({ _04901_, _04898_, _04894_, _04883_ }), .Y(_12746_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38621_ ( .A({ _04900_, _04899_, _04897_, _04872_ }), .Y(_12747_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38622_ ( .A({ _12751_, _12749_, _04880_, _04876_ }), .Y(_12748_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38623_ ( .A({ _12750_, _04893_, _04890_, _04881_ }), .Y(_12749_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38624_ ( .A({ _04895_, _04891_, _04889_, _04888_ }), .Y(_12750_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38625_ ( .A({ _04896_, _04892_, _04878_, _04875_ }), .Y(_12751_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38626_ ( .A({ _12753_, _04887_, _04884_, _04877_ }), .Y(_12752_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38627_ ( .A({ _04886_, _04885_, _04882_, _04879_ }), .Y(_12753_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _38628_ ( .A({ conv2d_16_mux_next_dma_flag_1, _12754_, _04906_, _12761_ }), .Y(_06819_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38629_ ( .A({ _12760_, _12759_, _12755_ }), .Y(_12754_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38630_ ( .A({ _12758_, _12757_, _12756_ }), .Y(_12755_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38631_ ( .A({ _04928_, _04927_, _04925_, _04924_ }), .Y(_12756_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38632_ ( .A({ _04923_, _04922_, _04921_, _04920_ }), .Y(_12757_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38633_ ( .A({ _04919_, _04918_, _04917_, _04916_ }), .Y(_12758_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38634_ ( .A({ _04914_, _04913_, _04912_, _04911_ }), .Y(_12759_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38635_ ( .A({ _04910_, _04909_, _04908_, _04907_ }), .Y(_12760_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38636_ ( .A({ _12764_, _12763_, _12762_ }), .Y(_12761_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38637_ ( .A({ _04905_, _04935_, _04934_ }), .Y(_12762_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38638_ ( .A({ _04933_, _04932_, _04931_, _04930_ }), .Y(_12763_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38639_ ( .A({ _04929_, _04926_, _04915_, _04904_ }), .Y(_12764_) );
  \$lut  #( .LUT(16'hbf00), .WIDTH(4) ) _38640_ ( .A({ conv2d_16_mux_next_dma_flag_2, _12769_, _12773_, _12765_ }), .Y(_06820_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _38641_ ( .A({ _04938_, _12766_, _12768_ }), .Y(_12765_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38642_ ( .A({ _12767_, _04937_, _04967_, _04966_ }), .Y(_12766_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38643_ ( .A({ _04965_, _04962_, _04958_, _04947_ }), .Y(_12767_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38644_ ( .A({ _04964_, _04963_, _04961_, _04936_ }), .Y(_12768_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38645_ ( .A({ _12772_, _12770_, _04944_, _04940_ }), .Y(_12769_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38646_ ( .A({ _12771_, _04951_, _04948_, _04941_ }), .Y(_12770_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38647_ ( .A({ _04950_, _04949_, _04946_, _04943_ }), .Y(_12771_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38648_ ( .A({ _04960_, _04956_, _04942_, _04939_ }), .Y(_12772_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38649_ ( .A({ _12774_, _04957_, _04954_, _04945_ }), .Y(_12773_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38650_ ( .A({ _04959_, _04955_, _04953_, _04952_ }), .Y(_12774_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38651_ ( .A({ _12782_, _12781_, _12776_ }), .Y(_12775_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38652_ ( .A({ _12780_, _12779_, _12778_, _12777_ }), .Y(_12776_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38653_ ( .A(conv2d_16_prev_row_count[23:20]), .Y(_12777_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38654_ ( .A(conv2d_16_prev_row_count[19:16]), .Y(_12778_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38655_ ( .A(conv2d_16_prev_row_count[31:28]), .Y(_12779_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38656_ ( .A(conv2d_16_prev_row_count[27:24]), .Y(_12780_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38657_ ( .A(conv2d_16_prev_row_count[15:12]), .Y(_12781_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38658_ ( .A(conv2d_16_prev_row_count[11:8]), .Y(_12782_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _38659_ ( .A({ conv2d_16_prev_row_count[3], cparam_conv2d_16_max_col_count[3], conv2d_16_prev_row_count[4], cparam_conv2d_16_max_col_count[4] }), .Y(_12783_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _38660_ ( .A({ cparam_conv2d_16_max_col_count[0], cparam_conv2d_16_max_col_count[1], conv2d_16_prev_row_count[0], conv2d_16_prev_row_count[1] }), .Y(_12784_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _38661_ ( .A({ cparam_conv2d_16_max_col_count[2], conv2d_16_prev_row_count[2], cparam_conv2d_16_max_col_count[3], conv2d_16_prev_row_count[3] }), .Y(_12785_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38662_ ( .A(conv2d_16_prev_row_count[7:5]), .Y(_12786_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38663_ ( .A({ _12801_, _12787_, _12775_ }), .Y(_06822_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38664_ ( .A({ _12796_, _12791_, _12788_ }), .Y(_12787_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38665_ ( .A({ _12790_, _12789_, _12786_ }), .Y(_12788_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38666_ ( .A({ conv2d_16_skip_write_out, conv2d_16_prev_och_count[31:29] }), .Y(_12789_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38667_ ( .A(conv2d_16_prev_och_count[28:25]), .Y(_12790_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38668_ ( .A({ _12795_, _12794_, _12793_, _12792_ }), .Y(_12791_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38669_ ( .A(conv2d_16_prev_och_count[16:13]), .Y(_12792_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38670_ ( .A(conv2d_16_prev_och_count[12:9]), .Y(_12793_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38671_ ( .A(conv2d_16_prev_och_count[24:21]), .Y(_12794_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38672_ ( .A(conv2d_16_prev_och_count[20:17]), .Y(_12795_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38673_ ( .A({ _12800_, _12799_, _12798_, _12797_ }), .Y(_12796_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38674_ ( .A({ conv2d_16_prev_och_count[0], conv2d_16_prev_bat_count[31:29] }), .Y(_12797_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38675_ ( .A(conv2d_16_prev_bat_count[28:25]), .Y(_12798_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38676_ ( .A(conv2d_16_prev_och_count[8:5]), .Y(_12799_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38677_ ( .A(conv2d_16_prev_och_count[4:1]), .Y(_12800_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38678_ ( .A({ _12810_, _12809_, _12807_, _12802_ }), .Y(_12801_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38679_ ( .A({ _12806_, _12805_, _12804_, _12803_ }), .Y(_12802_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38680_ ( .A({ conv2d_16_prev_bat_count[16], conv2d_16_prev_bat_count[13], conv2d_16_prev_bat_count[11:10] }), .Y(_12803_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38681_ ( .A({ conv2d_16_prev_bat_count[23:22], conv2d_16_prev_bat_count[20], conv2d_16_prev_bat_count[17] }), .Y(_12804_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38682_ ( .A({ conv2d_16_prev_bat_count[0], conv2d_16_prev_row_count[2:0] }), .Y(_12805_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38683_ ( .A({ conv2d_16_prev_bat_count[8], conv2d_16_prev_bat_count[5], conv2d_16_prev_bat_count[3:2] }), .Y(_12806_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38684_ ( .A({ _12808_, conv2d_16_prev_row_count[4:3] }), .Y(_12807_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38685_ ( .A({ conv2d_16_prev_bat_count[7:6], conv2d_16_prev_bat_count[4], conv2d_16_prev_bat_count[1] }), .Y(_12808_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38686_ ( .A({ conv2d_16_prev_bat_count[15:14], conv2d_16_prev_bat_count[12], conv2d_16_prev_bat_count[9] }), .Y(_12809_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38687_ ( .A({ conv2d_16_prev_bat_count[24], conv2d_16_prev_bat_count[21], conv2d_16_prev_bat_count[19:18] }), .Y(_12810_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38688_ ( .A({ _06175_, _12811_ }), .Y(_06823_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38689_ ( .A({ _12817_, _12816_, _12814_, _12812_ }), .Y(_12811_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38690_ ( .A({ _12813_, _04972_, _04971_ }), .Y(_12812_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38691_ ( .A({ _04976_, _04975_, _04974_, _04973_ }), .Y(_12813_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38692_ ( .A({ _12815_, _04993_, _04992_, _04991_ }), .Y(_12814_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38693_ ( .A({ _04989_, _04988_, _04987_, _04986_ }), .Y(_12815_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38694_ ( .A({ _04985_, _04984_, _04983_, _04982_ }), .Y(_12816_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38695_ ( .A({ _04981_, _04980_, _04978_, _04977_ }), .Y(_12817_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _38696_ ( .A({ _10804_, _maxi_read_op_sel[0], _11346_, _maxi_read_op_sel[1] }), .Y(_06824_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _38697_ ( .A({ _maxi_read_op_sel[1], _10804_, _11346_, _maxi_read_op_sel[0] }), .Y(_06826_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38698_ ( .A({ _maxi_read_op_sel[1:0], _11346_, _10804_ }), .Y(_06827_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _38699_ ( .A({ _10804_, _maxi_read_op_sel[0], _11503_, _maxi_read_op_sel[1] }), .Y(_06829_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38700_ ( .A({ _11503_, _10804_, _maxi_read_op_sel[1:0] }), .Y(_06828_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _38701_ ( .A({ _maxi_read_op_sel[1], _10804_, _11503_, _maxi_read_op_sel[0] }), .Y(_06830_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38702_ ( .A({ _maxi_read_op_sel[1:0], _11503_, _10804_ }), .Y(_06831_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38703_ ( .A({ _11352_, _10804_, _maxi_read_op_sel[1:0] }), .Y(_06832_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _38704_ ( .A({ _10804_, _maxi_read_op_sel[0], _11352_, _maxi_read_op_sel[1] }), .Y(_06833_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38705_ ( .A({ maxi_rlast, _10804_ }), .Y(_06825_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38706_ ( .A({ _06825_, _12818_ }), .Y(_06834_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _38707_ ( .A({ _09516_, _09525_, _09522_, _maxi_read_rest_size[8] }), .Y(_12818_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38708_ ( .A({ _12818_, _06825_ }), .Y(_06835_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38709_ ( .A({ _07465_, conv2d_16_skip_comp }), .Y(_06836_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38710_ ( .A({ _stream_conv2d_16_source_6_source_mode[1], _stream_conv2d_16_start }), .Y(_06686_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38711_ ( .A({ _stream_conv2d_16_source_8_source_mode[1], _stream_conv2d_16_start }), .Y(_06691_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38712_ ( .A({ _stream_conv2d_16_source_19_source_mode[1], _stream_conv2d_16_start }), .Y(_06696_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38713_ ( .A({ _stream_conv2d_16_source_20_source_mode[1], _stream_conv2d_16_start }), .Y(_06701_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38714_ ( .A({ _stream_conv2d_16_source_21_source_mode[1], _stream_conv2d_16_start }), .Y(_06706_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38715_ ( .A({ _stream_conv2d_16_source_22_source_mode[1], _stream_conv2d_16_start }), .Y(_06711_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38716_ ( .A({ _11833_, _11867_, _11855_ }), .Y(_06842_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38717_ ( .A({ _stream_conv2d_16_source_23_source_mode[1], _stream_conv2d_16_start }), .Y(_06716_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38718_ ( .A({ _stream_conv2d_16_source_24_source_mode[1], _stream_conv2d_16_start }), .Y(_06721_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38719_ ( .A({ _stream_conv2d_16_source_25_source_mode[1], _stream_conv2d_16_start }), .Y(_06726_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38720_ ( .A({ _stream_conv2d_16_source_26_source_mode[1], _stream_conv2d_16_start }), .Y(_06731_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38721_ ( .A({ _stream_conv2d_16_source_27_source_mode[1], _stream_conv2d_16_start }), .Y(_06736_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38722_ ( .A({ _stream_conv2d_16_source_28_source_mode[1], _stream_conv2d_16_start }), .Y(_06741_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38723_ ( .A({ _12133_, _12098_, _12120_ }), .Y(_06848_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38724_ ( .A({ _stream_conv2d_16_source_29_source_mode[1], _stream_conv2d_16_start }), .Y(_06746_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38725_ ( .A({ _12179_, _12144_, _12166_ }), .Y(_06849_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38726_ ( .A({ _stream_conv2d_16_source_30_source_mode[1], _stream_conv2d_16_start }), .Y(_06751_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38727_ ( .A({ _12225_, _12190_, _12212_ }), .Y(_06850_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38728_ ( .A({ _stream_conv2d_16_source_31_source_mode[1], _stream_conv2d_16_start }), .Y(_06756_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38729_ ( .A({ _12271_, _12236_, _12258_ }), .Y(_06851_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38730_ ( .A({ _stream_conv2d_16_source_32_source_mode[1], _stream_conv2d_16_start }), .Y(_06761_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38731_ ( .A({ _12315_, _12293_ }), .Y(_06852_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38732_ ( .A({ _stream_conv2d_16_source_33_source_mode[1], _stream_conv2d_16_start }), .Y(_06766_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38733_ ( .A({ _12361_, _12327_, _12349_ }), .Y(_06853_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38734_ ( .A({ _stream_conv2d_16_source_34_source_mode[1], _stream_conv2d_16_start }), .Y(_06771_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38735_ ( .A({ _12405_, _12383_ }), .Y(_06854_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38736_ ( .A({ _stream_conv2d_16_source_35_source_mode[1], _stream_conv2d_16_start }), .Y(_06776_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38737_ ( .A({ _12451_, _12417_, _12439_ }), .Y(_06855_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38738_ ( .A({ _stream_conv2d_16_source_36_source_mode[1], _stream_conv2d_16_start }), .Y(_06781_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38739_ ( .A({ _12497_, _12462_, _12484_ }), .Y(_06856_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38740_ ( .A({ _stream_conv2d_16_sink_37_sink_mode[0], __stream_conv2d_16_start_46 }), .Y(_06786_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38741_ ( .A({ _12828_, _12827_, _12826_, _12819_ }), .Y(_06857_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38742_ ( .A({ _12825_, _12820_, _stream_conv2d_16_sink_37_sink_count[2:1] }), .Y(_12819_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38743_ ( .A({ _12824_, _12823_, _12822_, _12821_ }), .Y(_12820_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38744_ ( .A(_stream_conv2d_16_sink_37_sink_count[14:11]), .Y(_12821_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38745_ ( .A(_stream_conv2d_16_sink_37_sink_count[10:7]), .Y(_12822_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38746_ ( .A(_stream_conv2d_16_sink_37_sink_count[22:19]), .Y(_12823_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38747_ ( .A(_stream_conv2d_16_sink_37_sink_count[18:15]), .Y(_12824_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38748_ ( .A(_stream_conv2d_16_sink_37_sink_count[6:3]), .Y(_12825_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38749_ ( .A({ _stream_conv2d_16_sink_37_sink_count[0], __delay_data_1614, _stream_conv2d_16_sink_37_sink_count[32:31] }), .Y(_12826_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38750_ ( .A(_stream_conv2d_16_sink_37_sink_count[30:27]), .Y(_12827_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38751_ ( .A(_stream_conv2d_16_sink_37_sink_count[26:23]), .Y(_12828_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38752_ ( .A({ _06176_, _12829_ }), .Y(_06858_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38753_ ( .A({ _12835_, _12834_, _12832_, _12830_ }), .Y(_12829_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38754_ ( .A({ _12831_, _05069_, _05068_ }), .Y(_12830_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38755_ ( .A({ _05073_, _05072_, _05071_, _05070_ }), .Y(_12831_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38756_ ( .A({ _12833_, _05090_, _05089_, _05088_ }), .Y(_12832_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38757_ ( .A({ _05086_, _05085_, _05084_, _05083_ }), .Y(_12833_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38758_ ( .A({ _05082_, _05081_, _05080_, _05079_ }), .Y(_12834_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38759_ ( .A({ _05078_, _05077_, _05075_, _05074_ }), .Y(_12835_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38760_ ( .A({ _maxi_write_data_done, _12836_ }), .Y(_06859_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _38761_ ( .A({ _09464_, _09473_, _09470_, _maxi_write_rest_size[8] }), .Y(_12836_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38762_ ( .A({ _maxi_write_data_done, _12836_ }), .Y(_06860_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38763_ ( .A({ _12851_, _12837_ }), .Y(_06862_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38764_ ( .A({ _12850_, _12849_, _12848_, _12838_ }), .Y(_12837_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38765_ ( .A({ _12847_, _12846_, _12844_, _12839_ }), .Y(_12838_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38766_ ( .A({ _12843_, _12842_, _12841_, _12840_ }), .Y(_12839_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38767_ ( .A(max_pool_serial_18_prev_bat_count[16:13]), .Y(_12840_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38768_ ( .A(max_pool_serial_18_prev_bat_count[12:9]), .Y(_12841_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38769_ ( .A(max_pool_serial_18_prev_bat_count[24:21]), .Y(_12842_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38770_ ( .A(max_pool_serial_18_prev_bat_count[20:17]), .Y(_12843_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38771_ ( .A({ _12845_, max_pool_serial_18_prev_row_count[1:0] }), .Y(_12844_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38772_ ( .A({ max_pool_serial_18_prev_bat_count[0], max_pool_serial_18_prev_row_count[4:2] }), .Y(_12845_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38773_ ( .A(max_pool_serial_18_prev_bat_count[8:5]), .Y(_12846_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38774_ ( .A(max_pool_serial_18_prev_bat_count[4:1]), .Y(_12847_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _38775_ ( .A(max_pool_serial_18_prev_row_count[7:5]), .Y(_12848_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _38776_ ( .A({ max_pool_serial_18_skip_write_out, max_pool_serial_18_prev_bat_count[31:29] }), .Y(_12849_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38777_ ( .A(max_pool_serial_18_prev_bat_count[28:25]), .Y(_12850_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38778_ ( .A({ _12858_, _12857_, _12852_ }), .Y(_12851_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38779_ ( .A({ _12856_, _12855_, _12854_, _12853_ }), .Y(_12852_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38780_ ( .A(max_pool_serial_18_prev_row_count[23:20]), .Y(_12853_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38781_ ( .A(max_pool_serial_18_prev_row_count[19:16]), .Y(_12854_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38782_ ( .A(max_pool_serial_18_prev_row_count[31:28]), .Y(_12855_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38783_ ( .A(max_pool_serial_18_prev_row_count[27:24]), .Y(_12856_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38784_ ( .A(max_pool_serial_18_prev_row_count[15:12]), .Y(_12857_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38785_ ( .A(max_pool_serial_18_prev_row_count[11:8]), .Y(_12858_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _38786_ ( .A({ max_pool_serial_18_skip_write_out, _12851_, _12859_ }), .Y(_06861_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _38787_ ( .A({ _12848_, _13140_, cparam_max_pool_serial_18_max_col_count[4], max_pool_serial_18_prev_row_count[4] }), .Y(_12859_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _38788_ ( .A({ max_pool_serial_18_prev_row_count[3], cparam_max_pool_serial_18_max_col_count[3], max_pool_serial_18_prev_row_count[4], cparam_max_pool_serial_18_max_col_count[4] }), .Y(_12860_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _38789_ ( .A({ cparam_max_pool_serial_18_max_col_count[0], cparam_max_pool_serial_18_max_col_count[1], max_pool_serial_18_prev_row_count[0], max_pool_serial_18_prev_row_count[1] }), .Y(_12861_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38790_ ( .A({ _07097_, max_pool_serial_18_skip_comp }), .Y(_06863_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38791_ ( .A({ _stream_max_pool_serial_18_source_1_source_mode[1], _stream_max_pool_serial_18_start }), .Y(_06788_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38792_ ( .A({ _stream_max_pool_serial_18_sink_3_sink_mode[0], __stream_max_pool_serial_18_start_10 }), .Y(_06793_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38793_ ( .A({ _12871_, _12870_, _12869_, _12862_ }), .Y(_06865_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38794_ ( .A({ _12868_, _12863_, _stream_max_pool_serial_18_sink_3_sink_count[2:1] }), .Y(_12862_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38795_ ( .A({ _12867_, _12866_, _12865_, _12864_ }), .Y(_12863_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38796_ ( .A(_stream_max_pool_serial_18_sink_3_sink_count[14:11]), .Y(_12864_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38797_ ( .A(_stream_max_pool_serial_18_sink_3_sink_count[10:7]), .Y(_12865_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38798_ ( .A(_stream_max_pool_serial_18_sink_3_sink_count[22:19]), .Y(_12866_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38799_ ( .A(_stream_max_pool_serial_18_sink_3_sink_count[18:15]), .Y(_12867_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38800_ ( .A(_stream_max_pool_serial_18_sink_3_sink_count[6:3]), .Y(_12868_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38801_ ( .A({ _stream_max_pool_serial_18_sink_3_sink_count[0], __substreamoutput_data_794, _stream_max_pool_serial_18_sink_3_sink_count[32:31] }), .Y(_12869_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38802_ ( .A(_stream_max_pool_serial_18_sink_3_sink_count[30:27]), .Y(_12870_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38803_ ( .A(_stream_max_pool_serial_18_sink_3_sink_count[26:23]), .Y(_12871_) );
  \$lut  #( .LUT(4'hb), .WIDTH(2) ) _38804_ ( .A({ matmul_29_mux_dma_flag_0, matmul_29_mux_dma_pad_mask_0 }), .Y(_06882_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38805_ ( .A({ _12895_, _12887_, _12872_ }), .Y(_06866_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38806_ ( .A({ _12882_, _12877_, _12873_ }), .Y(_12872_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38807_ ( .A({ _12876_, _12875_, _12874_ }), .Y(_12873_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38808_ ( .A({ matmul_29_skip_write_out, matmul_29_prev_och_count[7:6] }), .Y(_12874_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38809_ ( .A(matmul_29_prev_och_count[5:2]), .Y(_12875_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38810_ ( .A({ matmul_29_prev_och_count[1:0], matmul_29_prev_bat_count[31:30] }), .Y(_12876_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38811_ ( .A({ _12881_, _12880_, _12879_, _12878_ }), .Y(_12877_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38812_ ( .A(matmul_29_prev_bat_count[21:18]), .Y(_12878_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38813_ ( .A(matmul_29_prev_bat_count[17:14]), .Y(_12879_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38814_ ( .A(matmul_29_prev_bat_count[29:26]), .Y(_12880_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38815_ ( .A(matmul_29_prev_bat_count[25:22]), .Y(_12881_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38816_ ( .A({ _12886_, _12885_, _12884_, _12883_ }), .Y(_12882_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38817_ ( .A(matmul_29_prev_bat_count[5:2]), .Y(_12883_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38818_ ( .A({ matmul_29_prev_bat_count[1:0], matmul_29_prev_row_count[31:30] }), .Y(_12884_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38819_ ( .A(matmul_29_prev_bat_count[13:10]), .Y(_12885_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38820_ ( .A(matmul_29_prev_bat_count[9:6]), .Y(_12886_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38821_ ( .A({ _12894_, _12893_, _12888_ }), .Y(_12887_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38822_ ( .A({ _12892_, _12891_, _12890_, _12889_ }), .Y(_12888_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38823_ ( .A(matmul_29_prev_och_count[23:20]), .Y(_12889_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38824_ ( .A(matmul_29_prev_och_count[19:16]), .Y(_12890_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38825_ ( .A(matmul_29_prev_och_count[31:28]), .Y(_12891_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38826_ ( .A(matmul_29_prev_och_count[27:24]), .Y(_12892_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38827_ ( .A(matmul_29_prev_och_count[15:12]), .Y(_12893_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38828_ ( .A(matmul_29_prev_och_count[11:8]), .Y(_12894_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38829_ ( .A({ _12904_, _12903_, _12901_, _12896_ }), .Y(_12895_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38830_ ( .A({ _12900_, _12899_, _12898_, _12897_ }), .Y(_12896_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38831_ ( .A({ matmul_29_prev_row_count[21], matmul_29_prev_row_count[18], matmul_29_prev_row_count[16:15] }), .Y(_12897_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38832_ ( .A({ matmul_29_prev_row_count[28:27], matmul_29_prev_row_count[25], matmul_29_prev_row_count[22] }), .Y(_12898_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38833_ ( .A({ matmul_29_prev_row_count[5], matmul_29_prev_row_count[2:0] }), .Y(_12899_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38834_ ( .A({ matmul_29_prev_row_count[13], matmul_29_prev_row_count[10], matmul_29_prev_row_count[8:7] }), .Y(_12900_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _38835_ ( .A({ _12902_, matmul_29_prev_row_count[4:3] }), .Y(_12901_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38836_ ( .A({ matmul_29_prev_row_count[12:11], matmul_29_prev_row_count[9], matmul_29_prev_row_count[6] }), .Y(_12902_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38837_ ( .A({ matmul_29_prev_row_count[20:19], matmul_29_prev_row_count[17], matmul_29_prev_row_count[14] }), .Y(_12903_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38838_ ( .A({ matmul_29_prev_row_count[29], matmul_29_prev_row_count[26], matmul_29_prev_row_count[24:23] }), .Y(_12904_) );
  \$lut  #( .LUT(8'h0d), .WIDTH(3) ) _38839_ ( .A({ matmul_29_skip_write_out, _12905_, _12915_ }), .Y(_06867_) );
  \$lut  #( .LUT(16'h000b), .WIDTH(4) ) _38840_ ( .A({ _12914_, _12906_, _12908_, _12910_ }), .Y(_12905_) );
  \$lut  #( .LUT(16'hf400), .WIDTH(4) ) _38841_ ( .A({ _12907_, _12913_, _12911_, _12912_ }), .Y(_12906_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _38842_ ( .A({ _12910_, _12908_, matmul_29_prev_och_count[4], cparam_matmul_29_max_och_count[4] }), .Y(_12907_) );
  \$lut  #( .LUT(8'h90), .WIDTH(3) ) _38843_ ( .A({ _12909_, cparam_matmul_29_max_och_count[6], matmul_29_prev_och_count[6] }), .Y(_12908_) );
  \$lut  #( .LUT(16'hb00b), .WIDTH(4) ) _38844_ ( .A({ cparam_matmul_29_max_och_count[7], matmul_29_prev_och_count[7], matmul_29_prev_och_count[5], cparam_matmul_29_max_och_count[5] }), .Y(_12909_) );
  \$lut  #( .LUT(16'hb0bb), .WIDTH(4) ) _38845_ ( .A({ cparam_matmul_29_max_och_count[4], matmul_29_prev_och_count[4], cparam_matmul_29_max_och_count[5], matmul_29_prev_och_count[5] }), .Y(_12910_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _38846_ ( .A({ cparam_matmul_29_max_och_count[3], matmul_29_prev_och_count[3], cparam_matmul_29_max_och_count[2], matmul_29_prev_och_count[2] }), .Y(_12911_) );
  \$lut  #( .LUT(16'h2b22), .WIDTH(4) ) _38847_ ( .A({ matmul_29_prev_och_count[0], cparam_matmul_29_max_och_count[0], cparam_matmul_29_max_och_count[1], matmul_29_prev_och_count[1] }), .Y(_12912_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _38848_ ( .A({ cparam_matmul_29_max_och_count[2], cparam_matmul_29_max_och_count[3], matmul_29_prev_och_count[2], matmul_29_prev_och_count[3] }), .Y(_12913_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _38849_ ( .A({ cparam_matmul_29_max_och_count[6], cparam_matmul_29_max_och_count[7], matmul_29_prev_och_count[6], matmul_29_prev_och_count[7] }), .Y(_12914_) );
  \$lut  #( .LUT(16'h7f00), .WIDTH(4) ) _38850_ ( .A({ _12887_, _12911_, _12907_, _12916_ }), .Y(_12915_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _38851_ ( .A({ cparam_matmul_29_max_och_count[1], matmul_29_prev_och_count[1], cparam_matmul_29_max_och_count[0], matmul_29_prev_och_count[0] }), .Y(_12916_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _38852_ ( .A({ _08068_, matmul_29_skip_comp }), .Y(_06868_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38853_ ( .A({ _stream_matmul_29_source_6_source_mode[1], _stream_matmul_29_start }), .Y(_06795_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38854_ ( .A({ _12587_, _12552_, _12574_ }), .Y(_06869_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38855_ ( .A({ _stream_matmul_29_source_8_source_mode[1], _stream_matmul_29_start }), .Y(_06800_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38856_ ( .A({ _12633_, _12598_, _12620_ }), .Y(_06870_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38857_ ( .A({ _stream_matmul_29_source_19_source_mode[1], _stream_matmul_29_start }), .Y(_06805_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _38858_ ( .A({ _12679_, _12644_, _12666_ }), .Y(_06871_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38859_ ( .A({ _stream_matmul_29_source_20_source_mode[1], _stream_matmul_29_start }), .Y(_06810_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38860_ ( .A({ _stream_matmul_29_sink_21_sink_mode[0], __stream_matmul_29_start_42 }), .Y(_06815_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38861_ ( .A({ _12926_, _12925_, _12924_, _12917_ }), .Y(_06873_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38862_ ( .A({ _12923_, _12918_, _stream_matmul_29_sink_21_sink_count[2:1] }), .Y(_12917_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _38863_ ( .A({ _12922_, _12921_, _12920_, _12919_ }), .Y(_12918_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38864_ ( .A(_stream_matmul_29_sink_21_sink_count[14:11]), .Y(_12919_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38865_ ( .A(_stream_matmul_29_sink_21_sink_count[10:7]), .Y(_12920_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38866_ ( .A(_stream_matmul_29_sink_21_sink_count[22:19]), .Y(_12921_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38867_ ( .A(_stream_matmul_29_sink_21_sink_count[18:15]), .Y(_12922_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38868_ ( .A(_stream_matmul_29_sink_21_sink_count[6:3]), .Y(_12923_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _38869_ ( .A({ _stream_matmul_29_sink_21_sink_count[0], __delay_data_1616, _stream_matmul_29_sink_21_sink_count[32:31] }), .Y(_12924_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38870_ ( .A(_stream_matmul_29_sink_21_sink_count[30:27]), .Y(_12925_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38871_ ( .A(_stream_matmul_29_sink_21_sink_count[26:23]), .Y(_12926_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _38872_ ( .A(__variable_wdata_192), .Y(_06173_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _38873_ ( .A(__variable_wdata_175), .Y(_06172_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _38874_ ( .A(__variable_wdata_158), .Y(_06171_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _38875_ ( .A(__variable_wdata_141), .Y(_06170_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _38876_ ( .A(__variable_wdata_124), .Y(_06169_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _38877_ ( .A(__variable_wdata_107), .Y(_06168_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _38878_ ( .A(__variable_wdata_90), .Y(_06167_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _38879_ ( .A(__variable_wdata_73), .Y(_06166_) );
  \$lut  #( .LUT(16'hfffe), .WIDTH(4) ) _38880_ ( .A(__variable_wdata_56), .Y(_06165_) );
  \$lut  #( .LUT(8'hef), .WIDTH(3) ) _38881_ ( .A({ _12927_, __variable_wdata_1[1:0] }), .Y(_06163_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _38882_ ( .A(__variable_wdata_1[5:2]), .Y(_12927_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38883_ ( .A({ conv2d_16_bat_count[0], _06930_ }), .Y(_21159_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38884_ ( .A({ conv2d_16_bat_count[1], _06930_ }), .Y(_21170_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38885_ ( .A({ conv2d_16_bat_count[2], _06930_ }), .Y(_21181_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38886_ ( .A({ conv2d_16_bat_count[3], _06930_ }), .Y(_21184_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38887_ ( .A({ conv2d_16_bat_count[4], _06930_ }), .Y(_21185_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38888_ ( .A({ conv2d_16_bat_count[5], _06930_ }), .Y(_21186_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38889_ ( .A({ conv2d_16_bat_count[6], _06930_ }), .Y(_21187_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38890_ ( .A({ conv2d_16_bat_count[7], _06930_ }), .Y(_21188_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38891_ ( .A({ conv2d_16_bat_count[8], _06930_ }), .Y(_21189_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38892_ ( .A({ conv2d_16_bat_count[9], _06930_ }), .Y(_21190_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38893_ ( .A({ conv2d_16_bat_count[10], _06930_ }), .Y(_21160_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38894_ ( .A({ conv2d_16_bat_count[11], _06930_ }), .Y(_21161_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38895_ ( .A({ conv2d_16_bat_count[12], _06930_ }), .Y(_21162_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38896_ ( .A({ conv2d_16_bat_count[13], _06930_ }), .Y(_21163_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38897_ ( .A({ conv2d_16_bat_count[14], _06930_ }), .Y(_21164_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38898_ ( .A({ conv2d_16_bat_count[15], _06930_ }), .Y(_21165_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38899_ ( .A({ conv2d_16_bat_count[16], _06930_ }), .Y(_21166_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38900_ ( .A({ conv2d_16_bat_count[17], _06930_ }), .Y(_21167_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38901_ ( .A({ conv2d_16_bat_count[18], _06930_ }), .Y(_21168_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38902_ ( .A({ conv2d_16_bat_count[19], _06930_ }), .Y(_21169_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38903_ ( .A({ conv2d_16_bat_count[20], _06930_ }), .Y(_21171_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38904_ ( .A({ conv2d_16_bat_count[21], _06930_ }), .Y(_21172_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38905_ ( .A({ conv2d_16_bat_count[22], _06930_ }), .Y(_21173_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38906_ ( .A({ conv2d_16_bat_count[23], _06930_ }), .Y(_21174_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38907_ ( .A({ conv2d_16_bat_count[24], _06930_ }), .Y(_21175_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38908_ ( .A({ conv2d_16_bat_count[25], _06930_ }), .Y(_21176_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38909_ ( .A({ conv2d_16_bat_count[26], _06930_ }), .Y(_21177_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38910_ ( .A({ conv2d_16_bat_count[27], _06930_ }), .Y(_21178_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38911_ ( .A({ conv2d_16_bat_count[28], _06930_ }), .Y(_21179_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38912_ ( .A({ conv2d_16_bat_count[29], _06930_ }), .Y(_21180_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38913_ ( .A({ conv2d_16_bat_count[30], _06930_ }), .Y(_21182_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38914_ ( .A({ conv2d_16_bat_count[31], _06930_ }), .Y(_21183_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38915_ ( .A({ _04776_, _07066_ }), .Y(_21547_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38916_ ( .A({ _04787_, _07066_ }), .Y(_21558_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38917_ ( .A({ _04798_, _07066_ }), .Y(_21569_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38918_ ( .A({ _04801_, _07066_ }), .Y(_21572_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38919_ ( .A({ _04802_, _07066_ }), .Y(_21573_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38920_ ( .A({ _04803_, _07066_ }), .Y(_21574_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38921_ ( .A({ _04804_, _07066_ }), .Y(_21575_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38922_ ( .A({ _04805_, _07066_ }), .Y(_21576_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38923_ ( .A({ _04806_, _07066_ }), .Y(_21577_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38924_ ( .A({ _04807_, _07066_ }), .Y(_21578_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38925_ ( .A({ _04777_, _07066_ }), .Y(_21548_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38926_ ( .A({ _04778_, _07066_ }), .Y(_21549_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38927_ ( .A({ _04779_, _07066_ }), .Y(_21550_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38928_ ( .A({ _04780_, _07066_ }), .Y(_21551_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38929_ ( .A({ _04781_, _07066_ }), .Y(_21552_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38930_ ( .A({ _04782_, _07066_ }), .Y(_21553_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38931_ ( .A({ _04783_, _07066_ }), .Y(_21554_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38932_ ( .A({ _04784_, _07066_ }), .Y(_21555_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38933_ ( .A({ _04785_, _07066_ }), .Y(_21556_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38934_ ( .A({ _04786_, _07066_ }), .Y(_21557_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38935_ ( .A({ _04788_, _07066_ }), .Y(_21559_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38936_ ( .A({ _04789_, _07066_ }), .Y(_21560_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38937_ ( .A({ _04790_, _07066_ }), .Y(_21561_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38938_ ( .A({ _04791_, _07066_ }), .Y(_21562_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38939_ ( .A({ _04792_, _07066_ }), .Y(_21563_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38940_ ( .A({ _04793_, _07066_ }), .Y(_21564_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38941_ ( .A({ _04794_, _07066_ }), .Y(_21565_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38942_ ( .A({ _04795_, _07066_ }), .Y(_21566_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38943_ ( .A({ _04796_, _07066_ }), .Y(_21567_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38944_ ( .A({ _04797_, _07066_ }), .Y(_21568_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38945_ ( .A({ _04799_, _07066_ }), .Y(_21570_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38946_ ( .A({ _04800_, _07066_ }), .Y(_21571_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38947_ ( .A({ _21581_, _06930_ }), .Y(_21613_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38948_ ( .A({ _21592_, _06930_ }), .Y(_21624_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38949_ ( .A({ _21603_, _06930_ }), .Y(_21635_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38950_ ( .A({ _21606_, _06930_ }), .Y(_21638_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38951_ ( .A({ _21607_, _06930_ }), .Y(_21639_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38952_ ( .A({ _21608_, _06930_ }), .Y(_21640_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38953_ ( .A({ _21609_, _06930_ }), .Y(_21641_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38954_ ( .A({ _21610_, _06930_ }), .Y(_21642_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38955_ ( .A({ _21611_, _06930_ }), .Y(_21643_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38956_ ( .A({ _21612_, _06930_ }), .Y(_21644_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38957_ ( .A({ _21582_, _06930_ }), .Y(_21614_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38958_ ( .A({ _21583_, _06930_ }), .Y(_21615_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38959_ ( .A({ _21584_, _06930_ }), .Y(_21616_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38960_ ( .A({ _21585_, _06930_ }), .Y(_21617_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38961_ ( .A({ _21586_, _06930_ }), .Y(_21618_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38962_ ( .A({ _21587_, _06930_ }), .Y(_21619_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38963_ ( .A({ _21588_, _06930_ }), .Y(_21620_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38964_ ( .A({ _21589_, _06930_ }), .Y(_21621_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38965_ ( .A({ _21590_, _06930_ }), .Y(_21622_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38966_ ( .A({ _21591_, _06930_ }), .Y(_21623_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38967_ ( .A({ _21593_, _06930_ }), .Y(_21625_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38968_ ( .A({ _21594_, _06930_ }), .Y(_21626_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38969_ ( .A({ _21595_, _06930_ }), .Y(_21627_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38970_ ( .A({ _21596_, _06930_ }), .Y(_21628_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38971_ ( .A({ _21597_, _06930_ }), .Y(_21629_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38972_ ( .A({ _21598_, _06930_ }), .Y(_21630_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38973_ ( .A({ _21599_, _06930_ }), .Y(_21631_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38974_ ( .A({ _21600_, _06930_ }), .Y(_21632_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38975_ ( .A({ _21601_, _06930_ }), .Y(_21633_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38976_ ( .A({ _21602_, _06930_ }), .Y(_21634_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38977_ ( .A({ _21604_, _06930_ }), .Y(_21636_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38978_ ( .A({ _21605_, _06930_ }), .Y(_21637_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38979_ ( .A({ conv2d_16_row_count[0], _06930_ }), .Y(_21191_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38980_ ( .A({ conv2d_16_row_count[1], _06930_ }), .Y(_21202_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38981_ ( .A({ conv2d_16_row_count[2], _06930_ }), .Y(_21213_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38982_ ( .A({ conv2d_16_row_count[3], _06930_ }), .Y(_21216_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38983_ ( .A({ conv2d_16_row_count[4], _06930_ }), .Y(_21217_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38984_ ( .A({ conv2d_16_row_count[5], _06930_ }), .Y(_21218_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38985_ ( .A({ conv2d_16_row_count[6], _06930_ }), .Y(_21219_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38986_ ( .A({ conv2d_16_row_count[7], _06930_ }), .Y(_21220_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38987_ ( .A({ conv2d_16_row_count[8], _06930_ }), .Y(_21221_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38988_ ( .A({ conv2d_16_row_count[9], _06930_ }), .Y(_21222_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38989_ ( .A({ conv2d_16_row_count[10], _06930_ }), .Y(_21192_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38990_ ( .A({ conv2d_16_row_count[11], _06930_ }), .Y(_21193_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38991_ ( .A({ conv2d_16_row_count[12], _06930_ }), .Y(_21194_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38992_ ( .A({ conv2d_16_row_count[13], _06930_ }), .Y(_21195_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38993_ ( .A({ conv2d_16_row_count[14], _06930_ }), .Y(_21196_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38994_ ( .A({ conv2d_16_row_count[15], _06930_ }), .Y(_21197_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38995_ ( .A({ conv2d_16_row_count[16], _06930_ }), .Y(_21198_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38996_ ( .A({ conv2d_16_row_count[17], _06930_ }), .Y(_21199_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38997_ ( .A({ conv2d_16_row_count[18], _06930_ }), .Y(_21200_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38998_ ( .A({ conv2d_16_row_count[19], _06930_ }), .Y(_21201_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _38999_ ( .A({ conv2d_16_row_count[20], _06930_ }), .Y(_21203_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39000_ ( .A({ conv2d_16_row_count[21], _06930_ }), .Y(_21204_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39001_ ( .A({ conv2d_16_row_count[22], _06930_ }), .Y(_21205_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39002_ ( .A({ conv2d_16_row_count[23], _06930_ }), .Y(_21206_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39003_ ( .A({ conv2d_16_row_count[24], _06930_ }), .Y(_21207_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39004_ ( .A({ conv2d_16_row_count[25], _06930_ }), .Y(_21208_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39005_ ( .A({ conv2d_16_row_count[26], _06930_ }), .Y(_21209_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39006_ ( .A({ conv2d_16_row_count[27], _06930_ }), .Y(_21210_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39007_ ( .A({ conv2d_16_row_count[28], _06930_ }), .Y(_21211_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39008_ ( .A({ conv2d_16_row_count[29], _06930_ }), .Y(_21212_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39009_ ( .A({ conv2d_16_row_count[30], _06930_ }), .Y(_21214_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39010_ ( .A({ conv2d_16_row_count[31], _06930_ }), .Y(_21215_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39011_ ( .A({ _21645_, _06930_ }), .Y(_21677_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39012_ ( .A({ _21656_, _06930_ }), .Y(_21688_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39013_ ( .A({ _21667_, _06930_ }), .Y(_21699_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39014_ ( .A({ _21670_, _06930_ }), .Y(_21702_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39015_ ( .A({ _21671_, _06930_ }), .Y(_21703_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39016_ ( .A({ _21672_, _06930_ }), .Y(_21704_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39017_ ( .A({ _21673_, _06930_ }), .Y(_21705_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39018_ ( .A({ _21674_, _06930_ }), .Y(_21706_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39019_ ( .A({ _21675_, _06930_ }), .Y(_21707_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39020_ ( .A({ _21676_, _06930_ }), .Y(_21708_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39021_ ( .A({ _21646_, _06930_ }), .Y(_21678_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39022_ ( .A({ _21647_, _06930_ }), .Y(_21679_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39023_ ( .A({ _21648_, _06930_ }), .Y(_21680_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39024_ ( .A({ _21649_, _06930_ }), .Y(_21681_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39025_ ( .A({ _21650_, _06930_ }), .Y(_21682_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39026_ ( .A({ _21651_, _06930_ }), .Y(_21683_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39027_ ( .A({ _21652_, _06930_ }), .Y(_21684_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39028_ ( .A({ _21653_, _06930_ }), .Y(_21685_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39029_ ( .A({ _21654_, _06930_ }), .Y(_21686_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39030_ ( .A({ _21655_, _06930_ }), .Y(_21687_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39031_ ( .A({ _21657_, _06930_ }), .Y(_21689_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39032_ ( .A({ _21658_, _06930_ }), .Y(_21690_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39033_ ( .A({ _21659_, _06930_ }), .Y(_21691_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39034_ ( .A({ _21660_, _06930_ }), .Y(_21692_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39035_ ( .A({ _21661_, _06930_ }), .Y(_21693_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39036_ ( .A({ _21662_, _06930_ }), .Y(_21694_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39037_ ( .A({ _21663_, _06930_ }), .Y(_21695_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39038_ ( .A({ _21664_, _06930_ }), .Y(_21696_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39039_ ( .A({ _21665_, _06930_ }), .Y(_21697_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39040_ ( .A({ _21666_, _06930_ }), .Y(_21698_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39041_ ( .A({ _21668_, _06930_ }), .Y(_21700_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39042_ ( .A({ _21669_, _06930_ }), .Y(_21701_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39043_ ( .A({ _21709_, _06930_ }), .Y(_21741_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39044_ ( .A({ _21720_, _06930_ }), .Y(_21752_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39045_ ( .A({ _21731_, _06930_ }), .Y(_21763_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39046_ ( .A({ _21734_, _06930_ }), .Y(_21766_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39047_ ( .A({ _21735_, _06930_ }), .Y(_21767_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39048_ ( .A({ _21736_, _06930_ }), .Y(_21768_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39049_ ( .A({ _21737_, _06930_ }), .Y(_21769_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39050_ ( .A({ _21738_, _06930_ }), .Y(_21770_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39051_ ( .A({ _21739_, _06930_ }), .Y(_21771_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39052_ ( .A({ _21740_, _06930_ }), .Y(_21772_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39053_ ( .A({ _21710_, _06930_ }), .Y(_21742_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39054_ ( .A({ _21711_, _06930_ }), .Y(_21743_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39055_ ( .A({ _21712_, _06930_ }), .Y(_21744_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39056_ ( .A({ _21713_, _06930_ }), .Y(_21745_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39057_ ( .A({ _21714_, _06930_ }), .Y(_21746_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39058_ ( .A({ _21715_, _06930_ }), .Y(_21747_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39059_ ( .A({ _21716_, _06930_ }), .Y(_21748_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39060_ ( .A({ _21717_, _06930_ }), .Y(_21749_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39061_ ( .A({ _21718_, _06930_ }), .Y(_21750_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39062_ ( .A({ _21719_, _06930_ }), .Y(_21751_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39063_ ( .A({ _21721_, _06930_ }), .Y(_21753_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39064_ ( .A({ _21722_, _06930_ }), .Y(_21754_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39065_ ( .A({ _21723_, _06930_ }), .Y(_21755_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39066_ ( .A({ _21724_, _06930_ }), .Y(_21756_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39067_ ( .A({ _21725_, _06930_ }), .Y(_21757_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39068_ ( .A({ _21726_, _06930_ }), .Y(_21758_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39069_ ( .A({ _21727_, _06930_ }), .Y(_21759_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39070_ ( .A({ _21728_, _06930_ }), .Y(_21760_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39071_ ( .A({ _21729_, _06930_ }), .Y(_21761_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39072_ ( .A({ _21730_, _06930_ }), .Y(_21762_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39073_ ( .A({ _21732_, _06930_ }), .Y(_21764_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39074_ ( .A({ _21733_, _06930_ }), .Y(_21765_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39075_ ( .A({ _21059_, _06930_ }), .Y(_21091_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39076_ ( .A({ _21070_, _06930_ }), .Y(_21102_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39077_ ( .A({ _21081_, _06930_ }), .Y(_21113_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39078_ ( .A({ _21084_, _06930_ }), .Y(_21116_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39079_ ( .A({ _21085_, _06930_ }), .Y(_21117_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39080_ ( .A({ _21086_, _06930_ }), .Y(_21118_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39081_ ( .A({ _21087_, _06930_ }), .Y(_21119_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39082_ ( .A({ _21088_, _06930_ }), .Y(_21120_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39083_ ( .A({ _21089_, _06930_ }), .Y(_21121_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39084_ ( .A({ _21090_, _06930_ }), .Y(_21122_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39085_ ( .A({ _21060_, _06930_ }), .Y(_21092_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39086_ ( .A({ _21061_, _06930_ }), .Y(_21093_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39087_ ( .A({ _21062_, _06930_ }), .Y(_21094_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39088_ ( .A({ _21063_, _06930_ }), .Y(_21095_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39089_ ( .A({ _21064_, _06930_ }), .Y(_21096_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39090_ ( .A({ _21065_, _06930_ }), .Y(_21097_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39091_ ( .A({ _21066_, _06930_ }), .Y(_21098_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39092_ ( .A({ _21067_, _06930_ }), .Y(_21099_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39093_ ( .A({ _21068_, _06930_ }), .Y(_21100_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39094_ ( .A({ _21069_, _06930_ }), .Y(_21101_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39095_ ( .A({ _21071_, _06930_ }), .Y(_21103_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39096_ ( .A({ _21072_, _06930_ }), .Y(_21104_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39097_ ( .A({ _21073_, _06930_ }), .Y(_21105_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39098_ ( .A({ _21074_, _06930_ }), .Y(_21106_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39099_ ( .A({ _21075_, _06930_ }), .Y(_21107_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39100_ ( .A({ _21076_, _06930_ }), .Y(_21108_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39101_ ( .A({ _21077_, _06930_ }), .Y(_21109_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39102_ ( .A({ _21078_, _06930_ }), .Y(_21110_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39103_ ( .A({ _21079_, _06930_ }), .Y(_21111_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39104_ ( .A({ _21080_, _06930_ }), .Y(_21112_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39105_ ( .A({ _21082_, _06930_ }), .Y(_21114_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39106_ ( .A({ _21083_, _06930_ }), .Y(_21115_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39107_ ( .A({ _21123_, _06930_ }), .Y(_21125_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39108_ ( .A({ _21124_, _06930_ }), .Y(_21126_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39109_ ( .A({ _16396_, _07085_ }), .Y(_16428_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39110_ ( .A({ _16407_, _07085_ }), .Y(_16439_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39111_ ( .A({ _16418_, _07085_ }), .Y(_16450_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39112_ ( .A({ _16421_, _07085_ }), .Y(_16453_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39113_ ( .A({ _16422_, _07085_ }), .Y(_16454_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39114_ ( .A({ _16423_, _07085_ }), .Y(_16455_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39115_ ( .A({ _16424_, _07085_ }), .Y(_16456_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39116_ ( .A({ _16425_, _07085_ }), .Y(_16457_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39117_ ( .A({ _16426_, _07085_ }), .Y(_16458_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39118_ ( .A({ _16427_, _07085_ }), .Y(_16459_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39119_ ( .A({ _16397_, _07085_ }), .Y(_16429_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39120_ ( .A({ _16398_, _07085_ }), .Y(_16430_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39121_ ( .A({ _16399_, _07085_ }), .Y(_16431_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39122_ ( .A({ _16400_, _07085_ }), .Y(_16432_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39123_ ( .A({ _16401_, _07085_ }), .Y(_16433_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39124_ ( .A({ _16402_, _07085_ }), .Y(_16434_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39125_ ( .A({ _16403_, _07085_ }), .Y(_16435_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39126_ ( .A({ _16404_, _07085_ }), .Y(_16436_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39127_ ( .A({ _16405_, _07085_ }), .Y(_16437_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39128_ ( .A({ _16406_, _07085_ }), .Y(_16438_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39129_ ( .A({ _16408_, _07085_ }), .Y(_16440_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39130_ ( .A({ _16409_, _07085_ }), .Y(_16441_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39131_ ( .A({ _16410_, _07085_ }), .Y(_16442_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39132_ ( .A({ _16411_, _07085_ }), .Y(_16443_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39133_ ( .A({ _16412_, _07085_ }), .Y(_16444_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39134_ ( .A({ _16413_, _07085_ }), .Y(_16445_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39135_ ( .A({ _16414_, _07085_ }), .Y(_16446_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39136_ ( .A({ _16415_, _07085_ }), .Y(_16447_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39137_ ( .A({ _16416_, _07085_ }), .Y(_16448_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39138_ ( .A({ _16417_, _07085_ }), .Y(_16449_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39139_ ( .A({ _16419_, _07085_ }), .Y(_16451_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39140_ ( .A({ _16420_, _07085_ }), .Y(_16452_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39141_ ( .A({ _16332_, _07085_ }), .Y(_16364_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39142_ ( .A({ _16343_, _07085_ }), .Y(_16375_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39143_ ( .A({ _16354_, _07085_ }), .Y(_16386_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39144_ ( .A({ _16357_, _07085_ }), .Y(_16389_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39145_ ( .A({ _16358_, _07085_ }), .Y(_16390_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39146_ ( .A({ _16359_, _07085_ }), .Y(_16391_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39147_ ( .A({ _16360_, _07085_ }), .Y(_16392_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39148_ ( .A({ _16361_, _07085_ }), .Y(_16393_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39149_ ( .A({ _16362_, _07085_ }), .Y(_16394_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39150_ ( .A({ _16363_, _07085_ }), .Y(_16395_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39151_ ( .A({ _16333_, _07085_ }), .Y(_16365_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39152_ ( .A({ _16334_, _07085_ }), .Y(_16366_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39153_ ( .A({ _16335_, _07085_ }), .Y(_16367_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39154_ ( .A({ _16336_, _07085_ }), .Y(_16368_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39155_ ( .A({ _16337_, _07085_ }), .Y(_16369_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39156_ ( .A({ _16338_, _07085_ }), .Y(_16370_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39157_ ( .A({ _16339_, _07085_ }), .Y(_16371_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39158_ ( .A({ _16340_, _07085_ }), .Y(_16372_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39159_ ( .A({ _16341_, _07085_ }), .Y(_16373_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39160_ ( .A({ _16342_, _07085_ }), .Y(_16374_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39161_ ( .A({ _16344_, _07085_ }), .Y(_16376_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39162_ ( .A({ _16345_, _07085_ }), .Y(_16377_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39163_ ( .A({ _16346_, _07085_ }), .Y(_16378_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39164_ ( .A({ _16347_, _07085_ }), .Y(_16379_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39165_ ( .A({ _16348_, _07085_ }), .Y(_16380_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39166_ ( .A({ _16349_, _07085_ }), .Y(_16381_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39167_ ( .A({ _16350_, _07085_ }), .Y(_16382_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39168_ ( .A({ _16351_, _07085_ }), .Y(_16383_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39169_ ( .A({ _16352_, _07085_ }), .Y(_16384_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39170_ ( .A({ _16353_, _07085_ }), .Y(_16385_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39171_ ( .A({ _16355_, _07085_ }), .Y(_16387_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39172_ ( .A({ _16356_, _07085_ }), .Y(_16388_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39173_ ( .A({ _21773_, _06930_ }), .Y(_21805_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39174_ ( .A({ _21784_, _06930_ }), .Y(_21816_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39175_ ( .A({ _21795_, _06930_ }), .Y(_21827_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39176_ ( .A({ _21798_, _06930_ }), .Y(_21830_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39177_ ( .A({ _21799_, _06930_ }), .Y(_21831_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39178_ ( .A({ _21800_, _06930_ }), .Y(_21832_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39179_ ( .A({ _21801_, _06930_ }), .Y(_21833_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39180_ ( .A({ _21802_, _06930_ }), .Y(_21834_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39181_ ( .A({ _21803_, _06930_ }), .Y(_21835_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39182_ ( .A({ _21804_, _06930_ }), .Y(_21836_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39183_ ( .A({ _21774_, _06930_ }), .Y(_21806_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39184_ ( .A({ _21775_, _06930_ }), .Y(_21807_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39185_ ( .A({ _21776_, _06930_ }), .Y(_21808_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39186_ ( .A({ _21777_, _06930_ }), .Y(_21809_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39187_ ( .A({ _21778_, _06930_ }), .Y(_21810_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39188_ ( .A({ _21779_, _06930_ }), .Y(_21811_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39189_ ( .A({ _21780_, _06930_ }), .Y(_21812_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39190_ ( .A({ _21781_, _06930_ }), .Y(_21813_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39191_ ( .A({ _21782_, _06930_ }), .Y(_21814_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39192_ ( .A({ _21783_, _06930_ }), .Y(_21815_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39193_ ( .A({ _21785_, _06930_ }), .Y(_21817_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39194_ ( .A({ _21786_, _06930_ }), .Y(_21818_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39195_ ( .A({ _21787_, _06930_ }), .Y(_21819_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39196_ ( .A({ _21788_, _06930_ }), .Y(_21820_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39197_ ( .A({ _21789_, _06930_ }), .Y(_21821_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39198_ ( .A({ _21790_, _06930_ }), .Y(_21822_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39199_ ( .A({ _21791_, _06930_ }), .Y(_21823_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39200_ ( .A({ _21792_, _06930_ }), .Y(_21824_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39201_ ( .A({ _21793_, _06930_ }), .Y(_21825_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39202_ ( .A({ _21794_, _06930_ }), .Y(_21826_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39203_ ( .A({ _21796_, _06930_ }), .Y(_21828_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39204_ ( .A({ _21797_, _06930_ }), .Y(_21829_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39205_ ( .A({ _16268_, _07085_ }), .Y(_16300_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39206_ ( .A({ _16279_, _07085_ }), .Y(_16311_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39207_ ( .A({ _16290_, _07085_ }), .Y(_16322_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39208_ ( .A({ _16293_, _07085_ }), .Y(_16325_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39209_ ( .A({ _16294_, _07085_ }), .Y(_16326_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39210_ ( .A({ _16295_, _07085_ }), .Y(_16327_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39211_ ( .A({ _16296_, _07085_ }), .Y(_16328_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39212_ ( .A({ _16297_, _07085_ }), .Y(_16329_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39213_ ( .A({ _16298_, _07085_ }), .Y(_16330_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39214_ ( .A({ _16299_, _07085_ }), .Y(_16331_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39215_ ( .A({ _16269_, _07085_ }), .Y(_16301_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39216_ ( .A({ _16270_, _07085_ }), .Y(_16302_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39217_ ( .A({ _16271_, _07085_ }), .Y(_16303_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39218_ ( .A({ _16272_, _07085_ }), .Y(_16304_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39219_ ( .A({ _16273_, _07085_ }), .Y(_16305_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39220_ ( .A({ _16274_, _07085_ }), .Y(_16306_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39221_ ( .A({ _16275_, _07085_ }), .Y(_16307_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39222_ ( .A({ _16276_, _07085_ }), .Y(_16308_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39223_ ( .A({ _16277_, _07085_ }), .Y(_16309_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39224_ ( .A({ _16278_, _07085_ }), .Y(_16310_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39225_ ( .A({ _16280_, _07085_ }), .Y(_16312_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39226_ ( .A({ _16281_, _07085_ }), .Y(_16313_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39227_ ( .A({ _16282_, _07085_ }), .Y(_16314_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39228_ ( .A({ _16283_, _07085_ }), .Y(_16315_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39229_ ( .A({ _16284_, _07085_ }), .Y(_16316_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39230_ ( .A({ _16285_, _07085_ }), .Y(_16317_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39231_ ( .A({ _16286_, _07085_ }), .Y(_16318_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39232_ ( .A({ _16287_, _07085_ }), .Y(_16319_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39233_ ( .A({ _16288_, _07085_ }), .Y(_16320_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39234_ ( .A({ _16289_, _07085_ }), .Y(_16321_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39235_ ( .A({ _16291_, _07085_ }), .Y(_16323_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39236_ ( .A({ _16292_, _07085_ }), .Y(_16324_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39237_ ( .A({ _16140_, _07085_ }), .Y(_16172_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39238_ ( .A({ _16151_, _07085_ }), .Y(_16183_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39239_ ( .A({ _16162_, _07085_ }), .Y(_16194_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39240_ ( .A({ _16165_, _07085_ }), .Y(_16197_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39241_ ( .A({ _16166_, _07085_ }), .Y(_16198_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39242_ ( .A({ _16167_, _07085_ }), .Y(_16199_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39243_ ( .A({ _16168_, _07085_ }), .Y(_16200_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39244_ ( .A({ _16169_, _07085_ }), .Y(_16201_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39245_ ( .A({ _16170_, _07085_ }), .Y(_16202_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39246_ ( .A({ _16171_, _07085_ }), .Y(_16203_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39247_ ( .A({ _16141_, _07085_ }), .Y(_16173_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39248_ ( .A({ _16142_, _07085_ }), .Y(_16174_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39249_ ( .A({ _16143_, _07085_ }), .Y(_16175_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39250_ ( .A({ _16144_, _07085_ }), .Y(_16176_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39251_ ( .A({ _16145_, _07085_ }), .Y(_16177_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39252_ ( .A({ _16146_, _07085_ }), .Y(_16178_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39253_ ( .A({ _16147_, _07085_ }), .Y(_16179_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39254_ ( .A({ _16148_, _07085_ }), .Y(_16180_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39255_ ( .A({ _16149_, _07085_ }), .Y(_16181_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39256_ ( .A({ _16150_, _07085_ }), .Y(_16182_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39257_ ( .A({ _16152_, _07085_ }), .Y(_16184_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39258_ ( .A({ _16153_, _07085_ }), .Y(_16185_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39259_ ( .A({ _16154_, _07085_ }), .Y(_16186_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39260_ ( .A({ _16155_, _07085_ }), .Y(_16187_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39261_ ( .A({ _16156_, _07085_ }), .Y(_16188_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39262_ ( .A({ _16157_, _07085_ }), .Y(_16189_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39263_ ( .A({ _16158_, _07085_ }), .Y(_16190_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39264_ ( .A({ _16159_, _07085_ }), .Y(_16191_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39265_ ( .A({ _16160_, _07085_ }), .Y(_16192_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39266_ ( .A({ _16161_, _07085_ }), .Y(_16193_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39267_ ( .A({ _16163_, _07085_ }), .Y(_16195_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39268_ ( .A({ _16164_, _07085_ }), .Y(_16196_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39269_ ( .A({ _16204_, _07085_ }), .Y(_16236_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39270_ ( .A({ _16215_, _07085_ }), .Y(_16247_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39271_ ( .A({ _16226_, _07085_ }), .Y(_16258_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39272_ ( .A({ _16229_, _07085_ }), .Y(_16261_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39273_ ( .A({ _16230_, _07085_ }), .Y(_16262_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39274_ ( .A({ _16231_, _07085_ }), .Y(_16263_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39275_ ( .A({ _16232_, _07085_ }), .Y(_16264_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39276_ ( .A({ _16233_, _07085_ }), .Y(_16265_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39277_ ( .A({ _16234_, _07085_ }), .Y(_16266_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39278_ ( .A({ _16235_, _07085_ }), .Y(_16267_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39279_ ( .A({ _16205_, _07085_ }), .Y(_16237_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39280_ ( .A({ _16206_, _07085_ }), .Y(_16238_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39281_ ( .A({ _16207_, _07085_ }), .Y(_16239_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39282_ ( .A({ _16208_, _07085_ }), .Y(_16240_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39283_ ( .A({ _16209_, _07085_ }), .Y(_16241_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39284_ ( .A({ _16210_, _07085_ }), .Y(_16242_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39285_ ( .A({ _16211_, _07085_ }), .Y(_16243_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39286_ ( .A({ _16212_, _07085_ }), .Y(_16244_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39287_ ( .A({ _16213_, _07085_ }), .Y(_16245_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39288_ ( .A({ _16214_, _07085_ }), .Y(_16246_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39289_ ( .A({ _16216_, _07085_ }), .Y(_16248_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39290_ ( .A({ _16217_, _07085_ }), .Y(_16249_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39291_ ( .A({ _16218_, _07085_ }), .Y(_16250_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39292_ ( .A({ _16219_, _07085_ }), .Y(_16251_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39293_ ( .A({ _16220_, _07085_ }), .Y(_16252_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39294_ ( .A({ _16221_, _07085_ }), .Y(_16253_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39295_ ( .A({ _16222_, _07085_ }), .Y(_16254_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39296_ ( .A({ _16223_, _07085_ }), .Y(_16255_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39297_ ( .A({ _16224_, _07085_ }), .Y(_16256_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39298_ ( .A({ _16225_, _07085_ }), .Y(_16257_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39299_ ( .A({ _16227_, _07085_ }), .Y(_16259_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39300_ ( .A({ _16228_, _07085_ }), .Y(_16260_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39301_ ( .A({ _21287_, _06930_ }), .Y(_21319_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39302_ ( .A({ _21298_, _06930_ }), .Y(_21330_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39303_ ( .A({ _21309_, _06930_ }), .Y(_21341_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39304_ ( .A({ _21312_, _06930_ }), .Y(_21344_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39305_ ( .A({ _21313_, _06930_ }), .Y(_21345_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39306_ ( .A({ _21314_, _06930_ }), .Y(_21346_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39307_ ( .A({ _21315_, _06930_ }), .Y(_21347_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39308_ ( .A({ _21316_, _06930_ }), .Y(_21348_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39309_ ( .A({ _21317_, _06930_ }), .Y(_21349_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39310_ ( .A({ _21318_, _06930_ }), .Y(_21350_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39311_ ( .A({ _21288_, _06930_ }), .Y(_21320_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39312_ ( .A({ _21289_, _06930_ }), .Y(_21321_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39313_ ( .A({ _21290_, _06930_ }), .Y(_21322_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39314_ ( .A({ _21291_, _06930_ }), .Y(_21323_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39315_ ( .A({ _21292_, _06930_ }), .Y(_21324_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39316_ ( .A({ _21293_, _06930_ }), .Y(_21325_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39317_ ( .A({ _21294_, _06930_ }), .Y(_21326_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39318_ ( .A({ _21295_, _06930_ }), .Y(_21327_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39319_ ( .A({ _21296_, _06930_ }), .Y(_21328_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39320_ ( .A({ _21297_, _06930_ }), .Y(_21329_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39321_ ( .A({ _21299_, _06930_ }), .Y(_21331_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39322_ ( .A({ _21300_, _06930_ }), .Y(_21332_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39323_ ( .A({ _21301_, _06930_ }), .Y(_21333_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39324_ ( .A({ _21302_, _06930_ }), .Y(_21334_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39325_ ( .A({ _21303_, _06930_ }), .Y(_21335_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39326_ ( .A({ _21304_, _06930_ }), .Y(_21336_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39327_ ( .A({ _21305_, _06930_ }), .Y(_21337_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39328_ ( .A({ _21306_, _06930_ }), .Y(_21338_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39329_ ( .A({ _21307_, _06930_ }), .Y(_21339_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39330_ ( .A({ _21308_, _06930_ }), .Y(_21340_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39331_ ( .A({ _21310_, _06930_ }), .Y(_21342_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39332_ ( .A({ _21311_, _06930_ }), .Y(_21343_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39333_ ( .A({ _16076_, _07085_ }), .Y(_16108_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39334_ ( .A({ _16087_, _07085_ }), .Y(_16119_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39335_ ( .A({ _16098_, _07085_ }), .Y(_16130_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39336_ ( .A({ _16101_, _07085_ }), .Y(_16133_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39337_ ( .A({ _16102_, _07085_ }), .Y(_16134_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39338_ ( .A({ _16103_, _07085_ }), .Y(_16135_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39339_ ( .A({ _16104_, _07085_ }), .Y(_16136_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39340_ ( .A({ _16105_, _07085_ }), .Y(_16137_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39341_ ( .A({ _16106_, _07085_ }), .Y(_16138_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39342_ ( .A({ _16107_, _07085_ }), .Y(_16139_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39343_ ( .A({ _16077_, _07085_ }), .Y(_16109_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39344_ ( .A({ _16078_, _07085_ }), .Y(_16110_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39345_ ( .A({ _16079_, _07085_ }), .Y(_16111_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39346_ ( .A({ _16080_, _07085_ }), .Y(_16112_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39347_ ( .A({ _16081_, _07085_ }), .Y(_16113_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39348_ ( .A({ _16082_, _07085_ }), .Y(_16114_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39349_ ( .A({ _16083_, _07085_ }), .Y(_16115_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39350_ ( .A({ _16084_, _07085_ }), .Y(_16116_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39351_ ( .A({ _16085_, _07085_ }), .Y(_16117_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39352_ ( .A({ _16086_, _07085_ }), .Y(_16118_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39353_ ( .A({ _16088_, _07085_ }), .Y(_16120_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39354_ ( .A({ _16089_, _07085_ }), .Y(_16121_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39355_ ( .A({ _16090_, _07085_ }), .Y(_16122_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39356_ ( .A({ _16091_, _07085_ }), .Y(_16123_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39357_ ( .A({ _16092_, _07085_ }), .Y(_16124_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39358_ ( .A({ _16093_, _07085_ }), .Y(_16125_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39359_ ( .A({ _16094_, _07085_ }), .Y(_16126_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39360_ ( .A({ _16095_, _07085_ }), .Y(_16127_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39361_ ( .A({ _16096_, _07085_ }), .Y(_16128_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39362_ ( .A({ _16097_, _07085_ }), .Y(_16129_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39363_ ( .A({ _16099_, _07085_ }), .Y(_16131_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39364_ ( .A({ _16100_, _07085_ }), .Y(_16132_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39365_ ( .A({ max_pool_serial_18_row_count[0], _07085_ }), .Y(_16044_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39366_ ( .A({ max_pool_serial_18_row_count[1], _07085_ }), .Y(_16055_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39367_ ( .A({ max_pool_serial_18_row_count[2], _07085_ }), .Y(_16066_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39368_ ( .A({ max_pool_serial_18_row_count[3], _07085_ }), .Y(_16069_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39369_ ( .A({ max_pool_serial_18_row_count[4], _07085_ }), .Y(_16070_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39370_ ( .A({ max_pool_serial_18_row_count[5], _07085_ }), .Y(_16071_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39371_ ( .A({ max_pool_serial_18_row_count[6], _07085_ }), .Y(_16072_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39372_ ( .A({ max_pool_serial_18_row_count[7], _07085_ }), .Y(_16073_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39373_ ( .A({ max_pool_serial_18_row_count[8], _07085_ }), .Y(_16074_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39374_ ( .A({ max_pool_serial_18_row_count[9], _07085_ }), .Y(_16075_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39375_ ( .A({ max_pool_serial_18_row_count[10], _07085_ }), .Y(_16045_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39376_ ( .A({ max_pool_serial_18_row_count[11], _07085_ }), .Y(_16046_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39377_ ( .A({ max_pool_serial_18_row_count[12], _07085_ }), .Y(_16047_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39378_ ( .A({ max_pool_serial_18_row_count[13], _07085_ }), .Y(_16048_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39379_ ( .A({ max_pool_serial_18_row_count[14], _07085_ }), .Y(_16049_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39380_ ( .A({ max_pool_serial_18_row_count[15], _07085_ }), .Y(_16050_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39381_ ( .A({ max_pool_serial_18_row_count[16], _07085_ }), .Y(_16051_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39382_ ( .A({ max_pool_serial_18_row_count[17], _07085_ }), .Y(_16052_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39383_ ( .A({ max_pool_serial_18_row_count[18], _07085_ }), .Y(_16053_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39384_ ( .A({ max_pool_serial_18_row_count[19], _07085_ }), .Y(_16054_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39385_ ( .A({ max_pool_serial_18_row_count[20], _07085_ }), .Y(_16056_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39386_ ( .A({ max_pool_serial_18_row_count[21], _07085_ }), .Y(_16057_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39387_ ( .A({ max_pool_serial_18_row_count[22], _07085_ }), .Y(_16058_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39388_ ( .A({ max_pool_serial_18_row_count[23], _07085_ }), .Y(_16059_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39389_ ( .A({ max_pool_serial_18_row_count[24], _07085_ }), .Y(_16060_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39390_ ( .A({ max_pool_serial_18_row_count[25], _07085_ }), .Y(_16061_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39391_ ( .A({ max_pool_serial_18_row_count[26], _07085_ }), .Y(_16062_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39392_ ( .A({ max_pool_serial_18_row_count[27], _07085_ }), .Y(_16063_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39393_ ( .A({ max_pool_serial_18_row_count[28], _07085_ }), .Y(_16064_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39394_ ( .A({ max_pool_serial_18_row_count[29], _07085_ }), .Y(_16065_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39395_ ( .A({ max_pool_serial_18_row_count[30], _07085_ }), .Y(_16067_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39396_ ( .A({ max_pool_serial_18_row_count[31], _07085_ }), .Y(_16068_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39397_ ( .A({ _21837_, _06930_ }), .Y(_21869_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39398_ ( .A({ _21848_, _06930_ }), .Y(_21880_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39399_ ( .A({ _21859_, _06930_ }), .Y(_21891_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39400_ ( .A({ _21862_, _06930_ }), .Y(_21894_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39401_ ( .A({ _21863_, _06930_ }), .Y(_21895_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39402_ ( .A({ _21864_, _06930_ }), .Y(_21896_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39403_ ( .A({ _21865_, _06930_ }), .Y(_21897_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39404_ ( .A({ _21866_, _06930_ }), .Y(_21898_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39405_ ( .A({ _21867_, _06930_ }), .Y(_21899_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39406_ ( .A({ _21868_, _06930_ }), .Y(_21900_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39407_ ( .A({ _21838_, _06930_ }), .Y(_21870_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39408_ ( .A({ _21839_, _06930_ }), .Y(_21871_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39409_ ( .A({ _21840_, _06930_ }), .Y(_21872_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39410_ ( .A({ _21841_, _06930_ }), .Y(_21873_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39411_ ( .A({ _21842_, _06930_ }), .Y(_21874_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39412_ ( .A({ _21843_, _06930_ }), .Y(_21875_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39413_ ( .A({ _21844_, _06930_ }), .Y(_21876_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39414_ ( .A({ _21845_, _06930_ }), .Y(_21877_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39415_ ( .A({ _21846_, _06930_ }), .Y(_21878_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39416_ ( .A({ _21847_, _06930_ }), .Y(_21879_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39417_ ( .A({ _21849_, _06930_ }), .Y(_21881_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39418_ ( .A({ _21850_, _06930_ }), .Y(_21882_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39419_ ( .A({ _21851_, _06930_ }), .Y(_21883_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39420_ ( .A({ _21852_, _06930_ }), .Y(_21884_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39421_ ( .A({ _21853_, _06930_ }), .Y(_21885_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39422_ ( .A({ _21854_, _06930_ }), .Y(_21886_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39423_ ( .A({ _21855_, _06930_ }), .Y(_21887_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39424_ ( .A({ _21856_, _06930_ }), .Y(_21888_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39425_ ( .A({ _21857_, _06930_ }), .Y(_21889_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39426_ ( .A({ _21858_, _06930_ }), .Y(_21890_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39427_ ( .A({ _21860_, _06930_ }), .Y(_21892_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39428_ ( .A({ _21861_, _06930_ }), .Y(_21893_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39429_ ( .A({ _16010_, _07085_ }), .Y(_16011_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39430_ ( .A({ max_pool_serial_18_bat_count[0], _07085_ }), .Y(_16012_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39431_ ( .A({ max_pool_serial_18_bat_count[1], _07085_ }), .Y(_16023_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39432_ ( .A({ max_pool_serial_18_bat_count[2], _07085_ }), .Y(_16034_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39433_ ( .A({ max_pool_serial_18_bat_count[3], _07085_ }), .Y(_16037_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39434_ ( .A({ max_pool_serial_18_bat_count[4], _07085_ }), .Y(_16038_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39435_ ( .A({ max_pool_serial_18_bat_count[5], _07085_ }), .Y(_16039_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39436_ ( .A({ max_pool_serial_18_bat_count[6], _07085_ }), .Y(_16040_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39437_ ( .A({ max_pool_serial_18_bat_count[7], _07085_ }), .Y(_16041_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39438_ ( .A({ max_pool_serial_18_bat_count[8], _07085_ }), .Y(_16042_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39439_ ( .A({ max_pool_serial_18_bat_count[9], _07085_ }), .Y(_16043_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39440_ ( .A({ max_pool_serial_18_bat_count[10], _07085_ }), .Y(_16013_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39441_ ( .A({ max_pool_serial_18_bat_count[11], _07085_ }), .Y(_16014_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39442_ ( .A({ max_pool_serial_18_bat_count[12], _07085_ }), .Y(_16015_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39443_ ( .A({ max_pool_serial_18_bat_count[13], _07085_ }), .Y(_16016_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39444_ ( .A({ max_pool_serial_18_bat_count[14], _07085_ }), .Y(_16017_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39445_ ( .A({ max_pool_serial_18_bat_count[15], _07085_ }), .Y(_16018_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39446_ ( .A({ max_pool_serial_18_bat_count[16], _07085_ }), .Y(_16019_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39447_ ( .A({ max_pool_serial_18_bat_count[17], _07085_ }), .Y(_16020_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39448_ ( .A({ max_pool_serial_18_bat_count[18], _07085_ }), .Y(_16021_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39449_ ( .A({ max_pool_serial_18_bat_count[19], _07085_ }), .Y(_16022_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39450_ ( .A({ max_pool_serial_18_bat_count[20], _07085_ }), .Y(_16024_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39451_ ( .A({ max_pool_serial_18_bat_count[21], _07085_ }), .Y(_16025_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39452_ ( .A({ max_pool_serial_18_bat_count[22], _07085_ }), .Y(_16026_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39453_ ( .A({ max_pool_serial_18_bat_count[23], _07085_ }), .Y(_16027_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39454_ ( .A({ max_pool_serial_18_bat_count[24], _07085_ }), .Y(_16028_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39455_ ( .A({ max_pool_serial_18_bat_count[25], _07085_ }), .Y(_16029_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39456_ ( .A({ max_pool_serial_18_bat_count[26], _07085_ }), .Y(_16030_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39457_ ( .A({ max_pool_serial_18_bat_count[27], _07085_ }), .Y(_16031_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39458_ ( .A({ max_pool_serial_18_bat_count[28], _07085_ }), .Y(_16032_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39459_ ( .A({ max_pool_serial_18_bat_count[29], _07085_ }), .Y(_16033_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39460_ ( .A({ max_pool_serial_18_bat_count[30], _07085_ }), .Y(_16035_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39461_ ( .A({ max_pool_serial_18_bat_count[31], _07085_ }), .Y(_16036_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39462_ ( .A({ _21351_, _06930_ }), .Y(_21353_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39463_ ( .A({ _21352_, _06930_ }), .Y(_21354_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39464_ ( .A({ _15970_, _07085_ }), .Y(_16002_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39465_ ( .A({ _15946_, _07085_ }), .Y(_15978_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39466_ ( .A({ _15957_, _07085_ }), .Y(_15989_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39467_ ( .A({ _15968_, _07085_ }), .Y(_16000_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39468_ ( .A({ _15971_, _07085_ }), .Y(_16003_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39469_ ( .A({ _15972_, _07085_ }), .Y(_16004_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39470_ ( .A({ _15973_, _07085_ }), .Y(_16005_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39471_ ( .A({ _15974_, _07085_ }), .Y(_16006_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39472_ ( .A({ _15975_, _07085_ }), .Y(_16007_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39473_ ( .A({ _15976_, _07085_ }), .Y(_16008_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39474_ ( .A({ _15977_, _07085_ }), .Y(_16009_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39475_ ( .A({ _15947_, _07085_ }), .Y(_15979_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39476_ ( .A({ _15948_, _07085_ }), .Y(_15980_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39477_ ( .A({ _15949_, _07085_ }), .Y(_15981_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39478_ ( .A({ _15950_, _07085_ }), .Y(_15982_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39479_ ( .A({ _15951_, _07085_ }), .Y(_15983_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39480_ ( .A({ _15952_, _07085_ }), .Y(_15984_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39481_ ( .A({ _15953_, _07085_ }), .Y(_15985_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39482_ ( .A({ _15954_, _07085_ }), .Y(_15986_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39483_ ( .A({ _15955_, _07085_ }), .Y(_15987_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39484_ ( .A({ _15956_, _07085_ }), .Y(_15988_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39485_ ( .A({ _15958_, _07085_ }), .Y(_15990_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39486_ ( .A({ _15959_, _07085_ }), .Y(_15991_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39487_ ( .A({ _15960_, _07085_ }), .Y(_15992_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39488_ ( .A({ _15961_, _07085_ }), .Y(_15993_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39489_ ( .A({ _15962_, _07085_ }), .Y(_15994_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39490_ ( .A({ _15963_, _07085_ }), .Y(_15995_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39491_ ( .A({ _15964_, _07085_ }), .Y(_15996_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39492_ ( .A({ _15965_, _07085_ }), .Y(_15997_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39493_ ( .A({ _15966_, _07085_ }), .Y(_15998_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39494_ ( .A({ _15967_, _07085_ }), .Y(_15999_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39495_ ( .A({ _15969_, _07085_ }), .Y(_16001_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39496_ ( .A({ _15944_, _07085_ }), .Y(_15945_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39497_ ( .A({ _15880_, _07085_ }), .Y(_15912_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39498_ ( .A({ _15891_, _07085_ }), .Y(_15923_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39499_ ( .A({ _15902_, _07085_ }), .Y(_15934_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39500_ ( .A({ _15905_, _07085_ }), .Y(_15937_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39501_ ( .A({ _15906_, _07085_ }), .Y(_15938_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39502_ ( .A({ _15907_, _07085_ }), .Y(_15939_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39503_ ( .A({ _15908_, _07085_ }), .Y(_15940_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39504_ ( .A({ _15909_, _07085_ }), .Y(_15941_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39505_ ( .A({ _15910_, _07085_ }), .Y(_15942_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39506_ ( .A({ _15911_, _07085_ }), .Y(_15943_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39507_ ( .A({ _15881_, _07085_ }), .Y(_15913_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39508_ ( .A({ _15882_, _07085_ }), .Y(_15914_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39509_ ( .A({ _15883_, _07085_ }), .Y(_15915_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39510_ ( .A({ _15884_, _07085_ }), .Y(_15916_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39511_ ( .A({ _15885_, _07085_ }), .Y(_15917_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39512_ ( .A({ _15886_, _07085_ }), .Y(_15918_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39513_ ( .A({ _15887_, _07085_ }), .Y(_15919_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39514_ ( .A({ _15888_, _07085_ }), .Y(_15920_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39515_ ( .A({ _15889_, _07085_ }), .Y(_15921_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39516_ ( .A({ _15890_, _07085_ }), .Y(_15922_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39517_ ( .A({ _15892_, _07085_ }), .Y(_15924_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39518_ ( .A({ _15893_, _07085_ }), .Y(_15925_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39519_ ( .A({ _15894_, _07085_ }), .Y(_15926_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39520_ ( .A({ _15895_, _07085_ }), .Y(_15927_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39521_ ( .A({ _15896_, _07085_ }), .Y(_15928_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39522_ ( .A({ _15897_, _07085_ }), .Y(_15929_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39523_ ( .A({ _15898_, _07085_ }), .Y(_15930_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39524_ ( .A({ _15899_, _07085_ }), .Y(_15931_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39525_ ( .A({ _15900_, _07085_ }), .Y(_15932_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39526_ ( .A({ _15901_, _07085_ }), .Y(_15933_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39527_ ( .A({ _15903_, _07085_ }), .Y(_15935_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39528_ ( .A({ _15904_, _07085_ }), .Y(_15936_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39529_ ( .A({ _15814_, _07085_ }), .Y(_15815_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39530_ ( .A({ _15816_, _07085_ }), .Y(_15848_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39531_ ( .A({ _15827_, _07085_ }), .Y(_15859_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39532_ ( .A({ _15838_, _07085_ }), .Y(_15870_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39533_ ( .A({ _15841_, _07085_ }), .Y(_15873_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39534_ ( .A({ _15842_, _07085_ }), .Y(_15874_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39535_ ( .A({ _15843_, _07085_ }), .Y(_15875_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39536_ ( .A({ _15844_, _07085_ }), .Y(_15876_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39537_ ( .A({ _15845_, _07085_ }), .Y(_15877_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39538_ ( .A({ _15846_, _07085_ }), .Y(_15878_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39539_ ( .A({ _15847_, _07085_ }), .Y(_15879_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39540_ ( .A({ _15817_, _07085_ }), .Y(_15849_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39541_ ( .A({ _15818_, _07085_ }), .Y(_15850_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39542_ ( .A({ _15819_, _07085_ }), .Y(_15851_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39543_ ( .A({ _15820_, _07085_ }), .Y(_15852_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39544_ ( .A({ _15821_, _07085_ }), .Y(_15853_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39545_ ( .A({ _15822_, _07085_ }), .Y(_15854_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39546_ ( .A({ _15823_, _07085_ }), .Y(_15855_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39547_ ( .A({ _15824_, _07085_ }), .Y(_15856_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39548_ ( .A({ _15825_, _07085_ }), .Y(_15857_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39549_ ( .A({ _15826_, _07085_ }), .Y(_15858_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39550_ ( .A({ _15828_, _07085_ }), .Y(_15860_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39551_ ( .A({ _15829_, _07085_ }), .Y(_15861_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39552_ ( .A({ _15830_, _07085_ }), .Y(_15862_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39553_ ( .A({ _15831_, _07085_ }), .Y(_15863_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39554_ ( .A({ _15832_, _07085_ }), .Y(_15864_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39555_ ( .A({ _15833_, _07085_ }), .Y(_15865_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39556_ ( .A({ _15834_, _07085_ }), .Y(_15866_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39557_ ( .A({ _15835_, _07085_ }), .Y(_15867_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39558_ ( .A({ _15836_, _07085_ }), .Y(_15868_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39559_ ( .A({ _15837_, _07085_ }), .Y(_15869_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39560_ ( .A({ _15839_, _07085_ }), .Y(_15871_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39561_ ( .A({ _15840_, _07085_ }), .Y(_15872_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39562_ ( .A({ _21901_, _06930_ }), .Y(_21933_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39563_ ( .A({ _21912_, _06930_ }), .Y(_21944_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39564_ ( .A({ _21923_, _06930_ }), .Y(_21955_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39565_ ( .A({ _21926_, _06930_ }), .Y(_21958_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39566_ ( .A({ _21927_, _06930_ }), .Y(_21959_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39567_ ( .A({ _21928_, _06930_ }), .Y(_21960_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39568_ ( .A({ _21929_, _06930_ }), .Y(_21961_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39569_ ( .A({ _21930_, _06930_ }), .Y(_21962_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39570_ ( .A({ _21931_, _06930_ }), .Y(_21963_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39571_ ( .A({ _21932_, _06930_ }), .Y(_21964_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39572_ ( .A({ _21902_, _06930_ }), .Y(_21934_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39573_ ( .A({ _21903_, _06930_ }), .Y(_21935_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39574_ ( .A({ _21904_, _06930_ }), .Y(_21936_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39575_ ( .A({ _21905_, _06930_ }), .Y(_21937_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39576_ ( .A({ _21906_, _06930_ }), .Y(_21938_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39577_ ( .A({ _21907_, _06930_ }), .Y(_21939_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39578_ ( .A({ _21908_, _06930_ }), .Y(_21940_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39579_ ( .A({ _21909_, _06930_ }), .Y(_21941_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39580_ ( .A({ _21910_, _06930_ }), .Y(_21942_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39581_ ( .A({ _21911_, _06930_ }), .Y(_21943_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39582_ ( .A({ _21913_, _06930_ }), .Y(_21945_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39583_ ( .A({ _21914_, _06930_ }), .Y(_21946_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39584_ ( .A({ _21915_, _06930_ }), .Y(_21947_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39585_ ( .A({ _21916_, _06930_ }), .Y(_21948_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39586_ ( .A({ _21917_, _06930_ }), .Y(_21949_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39587_ ( .A({ _21918_, _06930_ }), .Y(_21950_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39588_ ( .A({ _21919_, _06930_ }), .Y(_21951_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39589_ ( .A({ _21920_, _06930_ }), .Y(_21952_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39590_ ( .A({ _21921_, _06930_ }), .Y(_21953_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39591_ ( .A({ _21922_, _06930_ }), .Y(_21954_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39592_ ( .A({ _21924_, _06930_ }), .Y(_21956_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39593_ ( .A({ _21925_, _06930_ }), .Y(_21957_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39594_ ( .A({ _15812_, _07085_ }), .Y(_15813_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39595_ ( .A({ _05130_, _12928_ }), .Y(_15778_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _39596_ ( .A({ _07084_, _07086_, _07070_ }), .Y(_12928_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39597_ ( .A({ _05141_, _12928_ }), .Y(_15789_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39598_ ( .A({ _05152_, _12928_ }), .Y(_15800_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39599_ ( .A({ _05155_, _12928_ }), .Y(_15803_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39600_ ( .A({ _05156_, _12928_ }), .Y(_15804_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39601_ ( .A({ _05157_, _12928_ }), .Y(_15805_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39602_ ( .A({ _05158_, _12928_ }), .Y(_15806_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39603_ ( .A({ _05159_, _12928_ }), .Y(_15807_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39604_ ( .A({ _05160_, _12928_ }), .Y(_15808_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39605_ ( .A({ _05161_, _12928_ }), .Y(_15809_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39606_ ( .A({ _05131_, _12928_ }), .Y(_15779_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39607_ ( .A({ _05132_, _12928_ }), .Y(_15780_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39608_ ( .A({ _05133_, _12928_ }), .Y(_15781_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39609_ ( .A({ _05134_, _12928_ }), .Y(_15782_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39610_ ( .A({ _05135_, _12928_ }), .Y(_15783_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39611_ ( .A({ _05136_, _12928_ }), .Y(_15784_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39612_ ( .A({ _05137_, _12928_ }), .Y(_15785_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39613_ ( .A({ _05138_, _12928_ }), .Y(_15786_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39614_ ( .A({ _05139_, _12928_ }), .Y(_15787_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39615_ ( .A({ _05140_, _12928_ }), .Y(_15788_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39616_ ( .A({ _05142_, _12928_ }), .Y(_15790_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39617_ ( .A({ _05143_, _12928_ }), .Y(_15791_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39618_ ( .A({ _05144_, _12928_ }), .Y(_15792_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39619_ ( .A({ _05145_, _12928_ }), .Y(_15793_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39620_ ( .A({ _05146_, _12928_ }), .Y(_15794_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39621_ ( .A({ _05147_, _12928_ }), .Y(_15795_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39622_ ( .A({ _05148_, _12928_ }), .Y(_15796_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39623_ ( .A({ _05149_, _12928_ }), .Y(_15797_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39624_ ( .A({ _05150_, _12928_ }), .Y(_15798_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39625_ ( .A({ _05151_, _12928_ }), .Y(_15799_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39626_ ( .A({ _05153_, _12928_ }), .Y(_15801_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39627_ ( .A({ _05154_, _12928_ }), .Y(_15802_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39628_ ( .A({ _20995_, _06930_ }), .Y(_21027_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39629_ ( .A({ _21006_, _06930_ }), .Y(_21038_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39630_ ( .A({ _21017_, _06930_ }), .Y(_21049_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39631_ ( .A({ _21020_, _06930_ }), .Y(_21052_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39632_ ( .A({ _21021_, _06930_ }), .Y(_21053_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39633_ ( .A({ _21022_, _06930_ }), .Y(_21054_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39634_ ( .A({ _21023_, _06930_ }), .Y(_21055_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39635_ ( .A({ _21024_, _06930_ }), .Y(_21056_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39636_ ( .A({ _21025_, _06930_ }), .Y(_21057_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39637_ ( .A({ _21026_, _06930_ }), .Y(_21058_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39638_ ( .A({ _20996_, _06930_ }), .Y(_21028_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39639_ ( .A({ _20997_, _06930_ }), .Y(_21029_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39640_ ( .A({ _20998_, _06930_ }), .Y(_21030_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39641_ ( .A({ _20999_, _06930_ }), .Y(_21031_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39642_ ( .A({ _21000_, _06930_ }), .Y(_21032_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39643_ ( .A({ _21001_, _06930_ }), .Y(_21033_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39644_ ( .A({ _21002_, _06930_ }), .Y(_21034_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39645_ ( .A({ _21003_, _06930_ }), .Y(_21035_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39646_ ( .A({ _21004_, _06930_ }), .Y(_21036_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39647_ ( .A({ _21005_, _06930_ }), .Y(_21037_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39648_ ( .A({ _21007_, _06930_ }), .Y(_21039_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39649_ ( .A({ _21008_, _06930_ }), .Y(_21040_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39650_ ( .A({ _21009_, _06930_ }), .Y(_21041_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39651_ ( .A({ _21010_, _06930_ }), .Y(_21042_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39652_ ( .A({ _21011_, _06930_ }), .Y(_21043_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39653_ ( .A({ _21012_, _06930_ }), .Y(_21044_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39654_ ( .A({ _21013_, _06930_ }), .Y(_21045_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39655_ ( .A({ _21014_, _06930_ }), .Y(_21046_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39656_ ( .A({ _21015_, _06930_ }), .Y(_21047_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39657_ ( .A({ _21016_, _06930_ }), .Y(_21048_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39658_ ( .A({ _21018_, _06930_ }), .Y(_21050_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39659_ ( .A({ _21019_, _06930_ }), .Y(_21051_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39660_ ( .A({ _15714_, _07372_ }), .Y(_15746_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39661_ ( .A({ _15725_, _07372_ }), .Y(_15757_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39662_ ( .A({ _15736_, _07372_ }), .Y(_15768_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39663_ ( .A({ _15739_, _07372_ }), .Y(_15771_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39664_ ( .A({ _15740_, _07372_ }), .Y(_15772_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39665_ ( .A({ _15741_, _07372_ }), .Y(_15773_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39666_ ( .A({ _15742_, _07372_ }), .Y(_15774_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39667_ ( .A({ _15743_, _07372_ }), .Y(_15775_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39668_ ( .A({ _15744_, _07372_ }), .Y(_15776_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39669_ ( .A({ _15745_, _07372_ }), .Y(_15777_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39670_ ( .A({ _15715_, _07372_ }), .Y(_15747_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39671_ ( .A({ _15716_, _07372_ }), .Y(_15748_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39672_ ( .A({ _15717_, _07372_ }), .Y(_15749_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39673_ ( .A({ _15718_, _07372_ }), .Y(_15750_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39674_ ( .A({ _15719_, _07372_ }), .Y(_15751_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39675_ ( .A({ _15720_, _07372_ }), .Y(_15752_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39676_ ( .A({ _15721_, _07372_ }), .Y(_15753_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39677_ ( .A({ _15722_, _07372_ }), .Y(_15754_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39678_ ( .A({ _15723_, _07372_ }), .Y(_15755_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39679_ ( .A({ _15724_, _07372_ }), .Y(_15756_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39680_ ( .A({ _15726_, _07372_ }), .Y(_15758_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39681_ ( .A({ _15727_, _07372_ }), .Y(_15759_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39682_ ( .A({ _15728_, _07372_ }), .Y(_15760_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39683_ ( .A({ _15729_, _07372_ }), .Y(_15761_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39684_ ( .A({ _15730_, _07372_ }), .Y(_15762_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39685_ ( .A({ _15731_, _07372_ }), .Y(_15763_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39686_ ( .A({ _15732_, _07372_ }), .Y(_15764_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39687_ ( .A({ _15733_, _07372_ }), .Y(_15765_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39688_ ( .A({ _15734_, _07372_ }), .Y(_15766_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39689_ ( .A({ _15735_, _07372_ }), .Y(_15767_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39690_ ( .A({ _15737_, _07372_ }), .Y(_15769_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39691_ ( .A({ _15738_, _07372_ }), .Y(_15770_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39692_ ( .A({ _15650_, _07372_ }), .Y(_15682_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39693_ ( .A({ _15661_, _07372_ }), .Y(_15693_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39694_ ( .A({ _15672_, _07372_ }), .Y(_15704_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39695_ ( .A({ _15675_, _07372_ }), .Y(_15707_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39696_ ( .A({ _15676_, _07372_ }), .Y(_15708_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39697_ ( .A({ _15677_, _07372_ }), .Y(_15709_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39698_ ( .A({ _15678_, _07372_ }), .Y(_15710_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39699_ ( .A({ _15679_, _07372_ }), .Y(_15711_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39700_ ( .A({ _15680_, _07372_ }), .Y(_15712_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39701_ ( .A({ _15681_, _07372_ }), .Y(_15713_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39702_ ( .A({ _15651_, _07372_ }), .Y(_15683_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39703_ ( .A({ _15652_, _07372_ }), .Y(_15684_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39704_ ( .A({ _15653_, _07372_ }), .Y(_15685_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39705_ ( .A({ _15654_, _07372_ }), .Y(_15686_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39706_ ( .A({ _15655_, _07372_ }), .Y(_15687_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39707_ ( .A({ _15656_, _07372_ }), .Y(_15688_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39708_ ( .A({ _15657_, _07372_ }), .Y(_15689_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39709_ ( .A({ _15658_, _07372_ }), .Y(_15690_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39710_ ( .A({ _15659_, _07372_ }), .Y(_15691_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39711_ ( .A({ _15660_, _07372_ }), .Y(_15692_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39712_ ( .A({ _15662_, _07372_ }), .Y(_15694_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39713_ ( .A({ _15663_, _07372_ }), .Y(_15695_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39714_ ( .A({ _15664_, _07372_ }), .Y(_15696_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39715_ ( .A({ _15665_, _07372_ }), .Y(_15697_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39716_ ( .A({ _15666_, _07372_ }), .Y(_15698_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39717_ ( .A({ _15667_, _07372_ }), .Y(_15699_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39718_ ( .A({ _15668_, _07372_ }), .Y(_15700_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39719_ ( .A({ _15669_, _07372_ }), .Y(_15701_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39720_ ( .A({ _15670_, _07372_ }), .Y(_15702_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39721_ ( .A({ _15671_, _07372_ }), .Y(_15703_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39722_ ( .A({ _15673_, _07372_ }), .Y(_15705_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39723_ ( .A({ _15674_, _07372_ }), .Y(_15706_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39724_ ( .A({ _21965_, _06930_ }), .Y(_21997_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39725_ ( .A({ _21976_, _06930_ }), .Y(_22008_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39726_ ( .A({ _21987_, _06930_ }), .Y(_22019_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39727_ ( .A({ _21990_, _06930_ }), .Y(_22022_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39728_ ( .A({ _21991_, _06930_ }), .Y(_22023_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39729_ ( .A({ _21992_, _06930_ }), .Y(_22024_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39730_ ( .A({ _21993_, _06930_ }), .Y(_22025_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39731_ ( .A({ _21994_, _06930_ }), .Y(_22026_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39732_ ( .A({ _21995_, _06930_ }), .Y(_22027_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39733_ ( .A({ _21996_, _06930_ }), .Y(_22028_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39734_ ( .A({ _21966_, _06930_ }), .Y(_21998_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39735_ ( .A({ _21967_, _06930_ }), .Y(_21999_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39736_ ( .A({ _21968_, _06930_ }), .Y(_22000_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39737_ ( .A({ _21969_, _06930_ }), .Y(_22001_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39738_ ( .A({ _21970_, _06930_ }), .Y(_22002_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39739_ ( .A({ _21971_, _06930_ }), .Y(_22003_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39740_ ( .A({ _21972_, _06930_ }), .Y(_22004_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39741_ ( .A({ _21973_, _06930_ }), .Y(_22005_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39742_ ( .A({ _21974_, _06930_ }), .Y(_22006_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39743_ ( .A({ _21975_, _06930_ }), .Y(_22007_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39744_ ( .A({ _21977_, _06930_ }), .Y(_22009_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39745_ ( .A({ _21978_, _06930_ }), .Y(_22010_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39746_ ( .A({ _21979_, _06930_ }), .Y(_22011_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39747_ ( .A({ _21980_, _06930_ }), .Y(_22012_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39748_ ( .A({ _21981_, _06930_ }), .Y(_22013_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39749_ ( .A({ _21982_, _06930_ }), .Y(_22014_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39750_ ( .A({ _21983_, _06930_ }), .Y(_22015_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39751_ ( .A({ _21984_, _06930_ }), .Y(_22016_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39752_ ( .A({ _21985_, _06930_ }), .Y(_22017_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39753_ ( .A({ _21986_, _06930_ }), .Y(_22018_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39754_ ( .A({ _21988_, _06930_ }), .Y(_22020_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39755_ ( .A({ _21989_, _06930_ }), .Y(_22021_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39756_ ( .A({ _15586_, _07372_ }), .Y(_15618_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39757_ ( .A({ _15597_, _07372_ }), .Y(_15629_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39758_ ( .A({ _15608_, _07372_ }), .Y(_15640_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39759_ ( .A({ _15611_, _07372_ }), .Y(_15643_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39760_ ( .A({ _15612_, _07372_ }), .Y(_15644_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39761_ ( .A({ _15613_, _07372_ }), .Y(_15645_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39762_ ( .A({ _15614_, _07372_ }), .Y(_15646_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39763_ ( .A({ _15615_, _07372_ }), .Y(_15647_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39764_ ( .A({ _15616_, _07372_ }), .Y(_15648_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39765_ ( .A({ _15617_, _07372_ }), .Y(_15649_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39766_ ( .A({ _15587_, _07372_ }), .Y(_15619_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39767_ ( .A({ _15588_, _07372_ }), .Y(_15620_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39768_ ( .A({ _15589_, _07372_ }), .Y(_15621_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39769_ ( .A({ _15590_, _07372_ }), .Y(_15622_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39770_ ( .A({ _15591_, _07372_ }), .Y(_15623_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39771_ ( .A({ _15592_, _07372_ }), .Y(_15624_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39772_ ( .A({ _15593_, _07372_ }), .Y(_15625_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39773_ ( .A({ _15594_, _07372_ }), .Y(_15626_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39774_ ( .A({ _15595_, _07372_ }), .Y(_15627_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39775_ ( .A({ _15596_, _07372_ }), .Y(_15628_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39776_ ( .A({ _15598_, _07372_ }), .Y(_15630_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39777_ ( .A({ _15599_, _07372_ }), .Y(_15631_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39778_ ( .A({ _15600_, _07372_ }), .Y(_15632_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39779_ ( .A({ _15601_, _07372_ }), .Y(_15633_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39780_ ( .A({ _15602_, _07372_ }), .Y(_15634_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39781_ ( .A({ _15603_, _07372_ }), .Y(_15635_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39782_ ( .A({ _15604_, _07372_ }), .Y(_15636_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39783_ ( .A({ _15605_, _07372_ }), .Y(_15637_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39784_ ( .A({ _15606_, _07372_ }), .Y(_15638_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39785_ ( .A({ _15607_, _07372_ }), .Y(_15639_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39786_ ( .A({ _15609_, _07372_ }), .Y(_15641_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39787_ ( .A({ _15610_, _07372_ }), .Y(_15642_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39788_ ( .A({ conv2d_16_och_count[0], _06930_ }), .Y(_21127_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39789_ ( .A({ conv2d_16_och_count[1], _06930_ }), .Y(_21138_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39790_ ( .A({ conv2d_16_och_count[2], _06930_ }), .Y(_21149_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39791_ ( .A({ conv2d_16_och_count[3], _06930_ }), .Y(_21152_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39792_ ( .A({ conv2d_16_och_count[4], _06930_ }), .Y(_21153_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39793_ ( .A({ conv2d_16_och_count[5], _06930_ }), .Y(_21154_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39794_ ( .A({ conv2d_16_och_count[6], _06930_ }), .Y(_21155_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39795_ ( .A({ conv2d_16_och_count[7], _06930_ }), .Y(_21156_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39796_ ( .A({ conv2d_16_och_count[8], _06930_ }), .Y(_21157_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39797_ ( .A({ conv2d_16_och_count[9], _06930_ }), .Y(_21158_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39798_ ( .A({ conv2d_16_och_count[10], _06930_ }), .Y(_21128_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39799_ ( .A({ conv2d_16_och_count[11], _06930_ }), .Y(_21129_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39800_ ( .A({ conv2d_16_och_count[12], _06930_ }), .Y(_21130_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39801_ ( .A({ conv2d_16_och_count[13], _06930_ }), .Y(_21131_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39802_ ( .A({ conv2d_16_och_count[14], _06930_ }), .Y(_21132_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39803_ ( .A({ conv2d_16_och_count[15], _06930_ }), .Y(_21133_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39804_ ( .A({ conv2d_16_och_count[16], _06930_ }), .Y(_21134_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39805_ ( .A({ conv2d_16_och_count[17], _06930_ }), .Y(_21135_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39806_ ( .A({ conv2d_16_och_count[18], _06930_ }), .Y(_21136_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39807_ ( .A({ conv2d_16_och_count[19], _06930_ }), .Y(_21137_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39808_ ( .A({ conv2d_16_och_count[20], _06930_ }), .Y(_21139_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39809_ ( .A({ conv2d_16_och_count[21], _06930_ }), .Y(_21140_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39810_ ( .A({ conv2d_16_och_count[22], _06930_ }), .Y(_21141_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39811_ ( .A({ conv2d_16_och_count[23], _06930_ }), .Y(_21142_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39812_ ( .A({ conv2d_16_och_count[24], _06930_ }), .Y(_21143_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39813_ ( .A({ conv2d_16_och_count[25], _06930_ }), .Y(_21144_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39814_ ( .A({ conv2d_16_och_count[26], _06930_ }), .Y(_21145_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39815_ ( .A({ conv2d_16_och_count[27], _06930_ }), .Y(_21146_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39816_ ( .A({ conv2d_16_och_count[28], _06930_ }), .Y(_21147_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39817_ ( .A({ conv2d_16_och_count[29], _06930_ }), .Y(_21148_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39818_ ( .A({ conv2d_16_och_count[30], _06930_ }), .Y(_21150_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39819_ ( .A({ conv2d_16_och_count[31], _06930_ }), .Y(_21151_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39820_ ( .A({ _21355_, _06930_ }), .Y(_21387_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39821_ ( .A({ _21366_, _06930_ }), .Y(_21398_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39822_ ( .A({ _21377_, _06930_ }), .Y(_21409_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39823_ ( .A({ _21380_, _06930_ }), .Y(_21412_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39824_ ( .A({ _21381_, _06930_ }), .Y(_21413_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39825_ ( .A({ _21382_, _06930_ }), .Y(_21414_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39826_ ( .A({ _21383_, _06930_ }), .Y(_21415_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39827_ ( .A({ _21384_, _06930_ }), .Y(_21416_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39828_ ( .A({ _21385_, _06930_ }), .Y(_21417_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39829_ ( .A({ _21386_, _06930_ }), .Y(_21418_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39830_ ( .A({ _21356_, _06930_ }), .Y(_21388_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39831_ ( .A({ _21357_, _06930_ }), .Y(_21389_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39832_ ( .A({ _21358_, _06930_ }), .Y(_21390_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39833_ ( .A({ _21359_, _06930_ }), .Y(_21391_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39834_ ( .A({ _21360_, _06930_ }), .Y(_21392_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39835_ ( .A({ _21361_, _06930_ }), .Y(_21393_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39836_ ( .A({ _21362_, _06930_ }), .Y(_21394_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39837_ ( .A({ _21363_, _06930_ }), .Y(_21395_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39838_ ( .A({ _21364_, _06930_ }), .Y(_21396_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39839_ ( .A({ _21365_, _06930_ }), .Y(_21397_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39840_ ( .A({ _21367_, _06930_ }), .Y(_21399_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39841_ ( .A({ _21368_, _06930_ }), .Y(_21400_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39842_ ( .A({ _21369_, _06930_ }), .Y(_21401_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39843_ ( .A({ _21370_, _06930_ }), .Y(_21402_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39844_ ( .A({ _21371_, _06930_ }), .Y(_21403_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39845_ ( .A({ _21372_, _06930_ }), .Y(_21404_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39846_ ( .A({ _21373_, _06930_ }), .Y(_21405_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39847_ ( .A({ _21374_, _06930_ }), .Y(_21406_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39848_ ( .A({ _21375_, _06930_ }), .Y(_21407_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39849_ ( .A({ _21376_, _06930_ }), .Y(_21408_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39850_ ( .A({ _21378_, _06930_ }), .Y(_21410_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39851_ ( .A({ _21379_, _06930_ }), .Y(_21411_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39852_ ( .A({ _21419_, _06930_ }), .Y(_21451_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39853_ ( .A({ _21430_, _06930_ }), .Y(_21462_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39854_ ( .A({ _21441_, _06930_ }), .Y(_21473_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39855_ ( .A({ _21444_, _06930_ }), .Y(_21476_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39856_ ( .A({ _21445_, _06930_ }), .Y(_21477_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39857_ ( .A({ _21446_, _06930_ }), .Y(_21478_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39858_ ( .A({ _21447_, _06930_ }), .Y(_21479_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39859_ ( .A({ _21448_, _06930_ }), .Y(_21480_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39860_ ( .A({ _21449_, _06930_ }), .Y(_21481_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39861_ ( .A({ _21450_, _06930_ }), .Y(_21482_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39862_ ( .A({ _21420_, _06930_ }), .Y(_21452_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39863_ ( .A({ _21421_, _06930_ }), .Y(_21453_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39864_ ( .A({ _21422_, _06930_ }), .Y(_21454_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39865_ ( .A({ _21423_, _06930_ }), .Y(_21455_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39866_ ( .A({ _21424_, _06930_ }), .Y(_21456_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39867_ ( .A({ _21425_, _06930_ }), .Y(_21457_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39868_ ( .A({ _21426_, _06930_ }), .Y(_21458_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39869_ ( .A({ _21427_, _06930_ }), .Y(_21459_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39870_ ( .A({ _21428_, _06930_ }), .Y(_21460_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39871_ ( .A({ _21429_, _06930_ }), .Y(_21461_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39872_ ( .A({ _21431_, _06930_ }), .Y(_21463_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39873_ ( .A({ _21432_, _06930_ }), .Y(_21464_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39874_ ( .A({ _21433_, _06930_ }), .Y(_21465_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39875_ ( .A({ _21434_, _06930_ }), .Y(_21466_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39876_ ( .A({ _21435_, _06930_ }), .Y(_21467_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39877_ ( .A({ _21436_, _06930_ }), .Y(_21468_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39878_ ( .A({ _21437_, _06930_ }), .Y(_21469_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39879_ ( .A({ _21438_, _06930_ }), .Y(_21470_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39880_ ( .A({ _21439_, _06930_ }), .Y(_21471_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39881_ ( .A({ _21440_, _06930_ }), .Y(_21472_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39882_ ( .A({ _21442_, _06930_ }), .Y(_21474_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39883_ ( .A({ _21443_, _06930_ }), .Y(_21475_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39884_ ( .A({ _05194_, _13755_ }), .Y(_14658_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39885_ ( .A({ _05205_, _13755_ }), .Y(_14669_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39886_ ( .A({ _05216_, _13755_ }), .Y(_14680_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39887_ ( .A({ _05219_, _13755_ }), .Y(_14683_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39888_ ( .A({ _05220_, _13755_ }), .Y(_14684_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39889_ ( .A({ _05221_, _13755_ }), .Y(_14685_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39890_ ( .A({ _05222_, _13755_ }), .Y(_14686_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39891_ ( .A({ _05223_, _13755_ }), .Y(_14687_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39892_ ( .A({ _05224_, _13755_ }), .Y(_14688_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39893_ ( .A({ _05225_, _13755_ }), .Y(_14689_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39894_ ( .A({ _05195_, _13755_ }), .Y(_14659_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39895_ ( .A({ _05196_, _13755_ }), .Y(_14660_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39896_ ( .A({ _05197_, _13755_ }), .Y(_14661_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39897_ ( .A({ _05198_, _13755_ }), .Y(_14662_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39898_ ( .A({ _05199_, _13755_ }), .Y(_14663_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39899_ ( .A({ _05200_, _13755_ }), .Y(_14664_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39900_ ( .A({ _05201_, _13755_ }), .Y(_14665_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39901_ ( .A({ _05202_, _13755_ }), .Y(_14666_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39902_ ( .A({ _05203_, _13755_ }), .Y(_14667_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39903_ ( .A({ _05204_, _13755_ }), .Y(_14668_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39904_ ( .A({ _05206_, _13755_ }), .Y(_14670_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39905_ ( .A({ _05207_, _13755_ }), .Y(_14671_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39906_ ( .A({ _05208_, _13755_ }), .Y(_14672_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39907_ ( .A({ _05209_, _13755_ }), .Y(_14673_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39908_ ( .A({ _05210_, _13755_ }), .Y(_14674_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39909_ ( .A({ _05211_, _13755_ }), .Y(_14675_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39910_ ( .A({ _05212_, _13755_ }), .Y(_14676_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39911_ ( .A({ _05213_, _13755_ }), .Y(_14677_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39912_ ( .A({ _05214_, _13755_ }), .Y(_14678_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39913_ ( .A({ _05215_, _13755_ }), .Y(_14679_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39914_ ( .A({ _05217_, _13755_ }), .Y(_14681_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39915_ ( .A({ _05218_, _13755_ }), .Y(_14682_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39916_ ( .A({ _14530_, _13755_ }), .Y(_14562_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39917_ ( .A({ _14541_, _13755_ }), .Y(_14573_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39918_ ( .A({ _14552_, _13755_ }), .Y(_14584_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39919_ ( .A({ _14555_, _13755_ }), .Y(_14587_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39920_ ( .A({ _14556_, _13755_ }), .Y(_14588_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39921_ ( .A({ _14557_, _13755_ }), .Y(_14589_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39922_ ( .A({ _14558_, _13755_ }), .Y(_14590_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39923_ ( .A({ _14559_, _13755_ }), .Y(_14591_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39924_ ( .A({ _14560_, _13755_ }), .Y(_14592_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39925_ ( .A({ _14561_, _13755_ }), .Y(_14593_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39926_ ( .A({ _14531_, _13755_ }), .Y(_14563_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39927_ ( .A({ _14532_, _13755_ }), .Y(_14564_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39928_ ( .A({ _14533_, _13755_ }), .Y(_14565_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39929_ ( .A({ _14534_, _13755_ }), .Y(_14566_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39930_ ( .A({ _14535_, _13755_ }), .Y(_14567_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39931_ ( .A({ _14536_, _13755_ }), .Y(_14568_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39932_ ( .A({ _14537_, _13755_ }), .Y(_14569_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39933_ ( .A({ _14538_, _13755_ }), .Y(_14570_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39934_ ( .A({ _14539_, _13755_ }), .Y(_14571_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39935_ ( .A({ _14540_, _13755_ }), .Y(_14572_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39936_ ( .A({ _14542_, _13755_ }), .Y(_14574_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39937_ ( .A({ _14543_, _13755_ }), .Y(_14575_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39938_ ( .A({ _14544_, _13755_ }), .Y(_14576_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39939_ ( .A({ _14545_, _13755_ }), .Y(_14577_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39940_ ( .A({ _14546_, _13755_ }), .Y(_14578_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39941_ ( .A({ _14547_, _13755_ }), .Y(_14579_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39942_ ( .A({ _14548_, _13755_ }), .Y(_14580_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39943_ ( .A({ _14549_, _13755_ }), .Y(_14581_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39944_ ( .A({ _14550_, _13755_ }), .Y(_14582_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39945_ ( .A({ _14551_, _13755_ }), .Y(_14583_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39946_ ( .A({ _14553_, _13755_ }), .Y(_14585_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39947_ ( .A({ _14554_, _13755_ }), .Y(_14586_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39948_ ( .A({ _14466_, _13755_ }), .Y(_14498_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39949_ ( .A({ _14477_, _13755_ }), .Y(_14509_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39950_ ( .A({ _14488_, _13755_ }), .Y(_14520_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39951_ ( .A({ _14491_, _13755_ }), .Y(_14523_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39952_ ( .A({ _14492_, _13755_ }), .Y(_14524_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39953_ ( .A({ _14493_, _13755_ }), .Y(_14525_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39954_ ( .A({ _14494_, _13755_ }), .Y(_14526_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39955_ ( .A({ _14495_, _13755_ }), .Y(_14527_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39956_ ( .A({ _14496_, _13755_ }), .Y(_14528_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39957_ ( .A({ _14497_, _13755_ }), .Y(_14529_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39958_ ( .A({ _14467_, _13755_ }), .Y(_14499_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39959_ ( .A({ _14468_, _13755_ }), .Y(_14500_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39960_ ( .A({ _14469_, _13755_ }), .Y(_14501_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39961_ ( .A({ _14470_, _13755_ }), .Y(_14502_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39962_ ( .A({ _14471_, _13755_ }), .Y(_14503_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39963_ ( .A({ _14472_, _13755_ }), .Y(_14504_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39964_ ( .A({ _14473_, _13755_ }), .Y(_14505_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39965_ ( .A({ _14474_, _13755_ }), .Y(_14506_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39966_ ( .A({ _14475_, _13755_ }), .Y(_14507_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39967_ ( .A({ _14476_, _13755_ }), .Y(_14508_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39968_ ( .A({ _14478_, _13755_ }), .Y(_14510_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39969_ ( .A({ _14479_, _13755_ }), .Y(_14511_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39970_ ( .A({ _14480_, _13755_ }), .Y(_14512_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39971_ ( .A({ _14481_, _13755_ }), .Y(_14513_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39972_ ( .A({ _14482_, _13755_ }), .Y(_14514_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39973_ ( .A({ _14483_, _13755_ }), .Y(_14515_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39974_ ( .A({ _14484_, _13755_ }), .Y(_14516_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39975_ ( .A({ _14485_, _13755_ }), .Y(_14517_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39976_ ( .A({ _14486_, _13755_ }), .Y(_14518_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39977_ ( .A({ _14487_, _13755_ }), .Y(_14519_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39978_ ( .A({ _14489_, _13755_ }), .Y(_14521_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39979_ ( .A({ _14490_, _13755_ }), .Y(_14522_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39980_ ( .A({ _14402_, _13755_ }), .Y(_14434_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39981_ ( .A({ _14413_, _13755_ }), .Y(_14445_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39982_ ( .A({ _14424_, _13755_ }), .Y(_14456_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39983_ ( .A({ _14427_, _13755_ }), .Y(_14459_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39984_ ( .A({ _14428_, _13755_ }), .Y(_14460_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39985_ ( .A({ _14429_, _13755_ }), .Y(_14461_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39986_ ( .A({ _14430_, _13755_ }), .Y(_14462_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39987_ ( .A({ _14431_, _13755_ }), .Y(_14463_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39988_ ( .A({ _14432_, _13755_ }), .Y(_14464_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39989_ ( .A({ _14433_, _13755_ }), .Y(_14465_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39990_ ( .A({ _14403_, _13755_ }), .Y(_14435_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39991_ ( .A({ _14404_, _13755_ }), .Y(_14436_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39992_ ( .A({ _14405_, _13755_ }), .Y(_14437_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39993_ ( .A({ _14406_, _13755_ }), .Y(_14438_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39994_ ( .A({ _14407_, _13755_ }), .Y(_14439_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39995_ ( .A({ _14408_, _13755_ }), .Y(_14440_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39996_ ( .A({ _14409_, _13755_ }), .Y(_14441_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39997_ ( .A({ _14410_, _13755_ }), .Y(_14442_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39998_ ( .A({ _14411_, _13755_ }), .Y(_14443_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _39999_ ( .A({ _14412_, _13755_ }), .Y(_14444_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40000_ ( .A({ _14414_, _13755_ }), .Y(_14446_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40001_ ( .A({ _14415_, _13755_ }), .Y(_14447_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40002_ ( .A({ _14416_, _13755_ }), .Y(_14448_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40003_ ( .A({ _14417_, _13755_ }), .Y(_14449_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40004_ ( .A({ _14418_, _13755_ }), .Y(_14450_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40005_ ( .A({ _14419_, _13755_ }), .Y(_14451_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40006_ ( .A({ _14420_, _13755_ }), .Y(_14452_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40007_ ( .A({ _14421_, _13755_ }), .Y(_14453_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40008_ ( .A({ _14422_, _13755_ }), .Y(_14454_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40009_ ( .A({ _14423_, _13755_ }), .Y(_14455_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40010_ ( .A({ _14425_, _13755_ }), .Y(_14457_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40011_ ( .A({ _14426_, _13755_ }), .Y(_14458_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40012_ ( .A({ _14338_, _08032_ }), .Y(_14370_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40013_ ( .A({ _14349_, _08032_ }), .Y(_14381_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40014_ ( .A({ _14360_, _08032_ }), .Y(_14392_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40015_ ( .A({ _14363_, _08032_ }), .Y(_14395_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40016_ ( .A({ _14364_, _08032_ }), .Y(_14396_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40017_ ( .A({ _14365_, _08032_ }), .Y(_14397_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40018_ ( .A({ _14366_, _08032_ }), .Y(_14398_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40019_ ( .A({ _14367_, _08032_ }), .Y(_14399_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40020_ ( .A({ _14368_, _08032_ }), .Y(_14400_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40021_ ( .A({ _14369_, _08032_ }), .Y(_14401_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40022_ ( .A({ _14339_, _08032_ }), .Y(_14371_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40023_ ( .A({ _14340_, _08032_ }), .Y(_14372_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40024_ ( .A({ _14341_, _08032_ }), .Y(_14373_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40025_ ( .A({ _14342_, _08032_ }), .Y(_14374_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40026_ ( .A({ _14343_, _08032_ }), .Y(_14375_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40027_ ( .A({ _14344_, _08032_ }), .Y(_14376_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40028_ ( .A({ _14345_, _08032_ }), .Y(_14377_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40029_ ( .A({ _14346_, _08032_ }), .Y(_14378_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40030_ ( .A({ _14347_, _08032_ }), .Y(_14379_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40031_ ( .A({ _14348_, _08032_ }), .Y(_14380_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40032_ ( .A({ _14350_, _08032_ }), .Y(_14382_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40033_ ( .A({ _14351_, _08032_ }), .Y(_14383_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40034_ ( .A({ _14352_, _08032_ }), .Y(_14384_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40035_ ( .A({ _14353_, _08032_ }), .Y(_14385_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40036_ ( .A({ _14354_, _08032_ }), .Y(_14386_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40037_ ( .A({ _14355_, _08032_ }), .Y(_14387_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40038_ ( .A({ _14356_, _08032_ }), .Y(_14388_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40039_ ( .A({ _14357_, _08032_ }), .Y(_14389_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40040_ ( .A({ _14358_, _08032_ }), .Y(_14390_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40041_ ( .A({ _14359_, _08032_ }), .Y(_14391_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40042_ ( .A({ _14361_, _08032_ }), .Y(_14393_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40043_ ( .A({ _14362_, _08032_ }), .Y(_14394_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40044_ ( .A({ _05226_, _13755_ }), .Y(_14306_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40045_ ( .A({ _05237_, _13755_ }), .Y(_14317_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40046_ ( .A({ _05248_, _13755_ }), .Y(_14328_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40047_ ( .A({ _05251_, _13755_ }), .Y(_14331_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40048_ ( .A({ _05252_, _13755_ }), .Y(_14332_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40049_ ( .A({ _05253_, _13755_ }), .Y(_14333_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40050_ ( .A({ _05254_, _13755_ }), .Y(_14334_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40051_ ( .A({ _05255_, _13755_ }), .Y(_14335_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40052_ ( .A({ _05256_, _13755_ }), .Y(_14336_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40053_ ( .A({ _05257_, _13755_ }), .Y(_14337_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40054_ ( .A({ _05227_, _13755_ }), .Y(_14307_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40055_ ( .A({ _05228_, _13755_ }), .Y(_14308_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40056_ ( .A({ _05229_, _13755_ }), .Y(_14309_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40057_ ( .A({ _05230_, _13755_ }), .Y(_14310_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40058_ ( .A({ _05231_, _13755_ }), .Y(_14311_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40059_ ( .A({ _05232_, _13755_ }), .Y(_14312_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40060_ ( .A({ _05233_, _13755_ }), .Y(_14313_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40061_ ( .A({ _05234_, _13755_ }), .Y(_14314_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40062_ ( .A({ _05235_, _13755_ }), .Y(_14315_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40063_ ( .A({ _05236_, _13755_ }), .Y(_14316_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40064_ ( .A({ _05238_, _13755_ }), .Y(_14318_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40065_ ( .A({ _05239_, _13755_ }), .Y(_14319_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40066_ ( .A({ _05240_, _13755_ }), .Y(_14320_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40067_ ( .A({ _05241_, _13755_ }), .Y(_14321_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40068_ ( .A({ _05242_, _13755_ }), .Y(_14322_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40069_ ( .A({ _05243_, _13755_ }), .Y(_14323_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40070_ ( .A({ _05244_, _13755_ }), .Y(_14324_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40071_ ( .A({ _05245_, _13755_ }), .Y(_14325_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40072_ ( .A({ _05246_, _13755_ }), .Y(_14326_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40073_ ( .A({ _05247_, _13755_ }), .Y(_14327_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40074_ ( .A({ _05249_, _13755_ }), .Y(_14329_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40075_ ( .A({ _05250_, _13755_ }), .Y(_14330_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40076_ ( .A({ _14242_, _13755_ }), .Y(_14274_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40077_ ( .A({ _14253_, _13755_ }), .Y(_14285_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40078_ ( .A({ _14264_, _13755_ }), .Y(_14296_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40079_ ( .A({ _14267_, _13755_ }), .Y(_14299_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40080_ ( .A({ _14268_, _13755_ }), .Y(_14300_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40081_ ( .A({ _14269_, _13755_ }), .Y(_14301_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40082_ ( .A({ _14270_, _13755_ }), .Y(_14302_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40083_ ( .A({ _14271_, _13755_ }), .Y(_14303_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40084_ ( .A({ _14272_, _13755_ }), .Y(_14304_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40085_ ( .A({ _14273_, _13755_ }), .Y(_14305_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40086_ ( .A({ _14243_, _13755_ }), .Y(_14275_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40087_ ( .A({ _14244_, _13755_ }), .Y(_14276_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40088_ ( .A({ _14245_, _13755_ }), .Y(_14277_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40089_ ( .A({ _14246_, _13755_ }), .Y(_14278_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40090_ ( .A({ _14247_, _13755_ }), .Y(_14279_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40091_ ( .A({ _14248_, _13755_ }), .Y(_14280_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40092_ ( .A({ _14249_, _13755_ }), .Y(_14281_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40093_ ( .A({ _14250_, _13755_ }), .Y(_14282_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40094_ ( .A({ _14251_, _13755_ }), .Y(_14283_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40095_ ( .A({ _14252_, _13755_ }), .Y(_14284_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40096_ ( .A({ _14254_, _13755_ }), .Y(_14286_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40097_ ( .A({ _14255_, _13755_ }), .Y(_14287_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40098_ ( .A({ _14256_, _13755_ }), .Y(_14288_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40099_ ( .A({ _14257_, _13755_ }), .Y(_14289_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40100_ ( .A({ _14258_, _13755_ }), .Y(_14290_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40101_ ( .A({ _14259_, _13755_ }), .Y(_14291_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40102_ ( .A({ _14260_, _13755_ }), .Y(_14292_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40103_ ( .A({ _14261_, _13755_ }), .Y(_14293_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40104_ ( .A({ _14262_, _13755_ }), .Y(_14294_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40105_ ( .A({ _14263_, _13755_ }), .Y(_14295_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40106_ ( .A({ _14265_, _13755_ }), .Y(_14297_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40107_ ( .A({ _14266_, _13755_ }), .Y(_14298_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40108_ ( .A({ matmul_29_row_count[0], _13755_ }), .Y(_14146_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40109_ ( .A({ matmul_29_row_count[1], _13755_ }), .Y(_14157_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40110_ ( .A({ matmul_29_row_count[2], _13755_ }), .Y(_14168_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40111_ ( .A({ matmul_29_row_count[3], _13755_ }), .Y(_14171_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40112_ ( .A({ matmul_29_row_count[4], _13755_ }), .Y(_14172_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40113_ ( .A({ matmul_29_row_count[5], _13755_ }), .Y(_14173_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40114_ ( .A({ matmul_29_row_count[6], _13755_ }), .Y(_14174_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40115_ ( .A({ matmul_29_row_count[7], _13755_ }), .Y(_14175_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40116_ ( .A({ matmul_29_row_count[8], _13755_ }), .Y(_14176_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40117_ ( .A({ matmul_29_row_count[9], _13755_ }), .Y(_14177_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40118_ ( .A({ matmul_29_row_count[10], _13755_ }), .Y(_14147_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40119_ ( .A({ matmul_29_row_count[11], _13755_ }), .Y(_14148_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40120_ ( .A({ matmul_29_row_count[12], _13755_ }), .Y(_14149_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40121_ ( .A({ matmul_29_row_count[13], _13755_ }), .Y(_14150_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40122_ ( .A({ matmul_29_row_count[14], _13755_ }), .Y(_14151_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40123_ ( .A({ matmul_29_row_count[15], _13755_ }), .Y(_14152_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40124_ ( .A({ matmul_29_row_count[16], _13755_ }), .Y(_14153_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40125_ ( .A({ matmul_29_row_count[17], _13755_ }), .Y(_14154_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40126_ ( .A({ matmul_29_row_count[18], _13755_ }), .Y(_14155_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40127_ ( .A({ matmul_29_row_count[19], _13755_ }), .Y(_14156_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40128_ ( .A({ matmul_29_row_count[20], _13755_ }), .Y(_14158_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40129_ ( .A({ matmul_29_row_count[21], _13755_ }), .Y(_14159_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40130_ ( .A({ matmul_29_row_count[22], _13755_ }), .Y(_14160_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40131_ ( .A({ matmul_29_row_count[23], _13755_ }), .Y(_14161_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40132_ ( .A({ matmul_29_row_count[24], _13755_ }), .Y(_14162_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40133_ ( .A({ matmul_29_row_count[25], _13755_ }), .Y(_14163_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40134_ ( .A({ matmul_29_row_count[26], _13755_ }), .Y(_14164_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40135_ ( .A({ matmul_29_row_count[27], _13755_ }), .Y(_14165_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40136_ ( .A({ matmul_29_row_count[28], _13755_ }), .Y(_14166_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40137_ ( .A({ matmul_29_row_count[29], _13755_ }), .Y(_14167_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40138_ ( .A({ matmul_29_row_count[30], _13755_ }), .Y(_14169_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40139_ ( .A({ matmul_29_row_count[31], _13755_ }), .Y(_14170_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40140_ ( .A({ matmul_29_och_count[0], _13755_ }), .Y(_14082_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40141_ ( .A({ matmul_29_och_count[1], _13755_ }), .Y(_14093_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40142_ ( .A({ matmul_29_och_count[2], _13755_ }), .Y(_14104_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40143_ ( .A({ matmul_29_och_count[3], _13755_ }), .Y(_14107_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40144_ ( .A({ matmul_29_och_count[4], _13755_ }), .Y(_14108_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40145_ ( .A({ matmul_29_och_count[5], _13755_ }), .Y(_14109_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40146_ ( .A({ matmul_29_och_count[6], _13755_ }), .Y(_14110_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40147_ ( .A({ matmul_29_och_count[7], _13755_ }), .Y(_14111_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40148_ ( .A({ matmul_29_och_count[8], _13755_ }), .Y(_14112_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40149_ ( .A({ matmul_29_och_count[9], _13755_ }), .Y(_14113_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40150_ ( .A({ matmul_29_och_count[10], _13755_ }), .Y(_14083_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40151_ ( .A({ matmul_29_och_count[11], _13755_ }), .Y(_14084_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40152_ ( .A({ matmul_29_och_count[12], _13755_ }), .Y(_14085_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40153_ ( .A({ matmul_29_och_count[13], _13755_ }), .Y(_14086_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40154_ ( .A({ matmul_29_och_count[14], _13755_ }), .Y(_14087_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40155_ ( .A({ matmul_29_och_count[15], _13755_ }), .Y(_14088_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40156_ ( .A({ matmul_29_och_count[16], _13755_ }), .Y(_14089_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40157_ ( .A({ matmul_29_och_count[17], _13755_ }), .Y(_14090_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40158_ ( .A({ matmul_29_och_count[18], _13755_ }), .Y(_14091_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40159_ ( .A({ matmul_29_och_count[19], _13755_ }), .Y(_14092_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40160_ ( .A({ matmul_29_och_count[20], _13755_ }), .Y(_14094_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40161_ ( .A({ matmul_29_och_count[21], _13755_ }), .Y(_14095_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40162_ ( .A({ matmul_29_och_count[22], _13755_ }), .Y(_14096_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40163_ ( .A({ matmul_29_och_count[23], _13755_ }), .Y(_14097_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40164_ ( .A({ matmul_29_och_count[24], _13755_ }), .Y(_14098_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40165_ ( .A({ matmul_29_och_count[25], _13755_ }), .Y(_14099_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40166_ ( .A({ matmul_29_och_count[26], _13755_ }), .Y(_14100_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40167_ ( .A({ matmul_29_och_count[27], _13755_ }), .Y(_14101_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40168_ ( .A({ matmul_29_och_count[28], _13755_ }), .Y(_14102_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40169_ ( .A({ matmul_29_och_count[29], _13755_ }), .Y(_14103_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40170_ ( .A({ matmul_29_och_count[30], _13755_ }), .Y(_14105_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40171_ ( .A({ matmul_29_och_count[31], _13755_ }), .Y(_14106_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40172_ ( .A({ matmul_29_bat_count[0], _13755_ }), .Y(_14114_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40173_ ( .A({ matmul_29_bat_count[1], _13755_ }), .Y(_14125_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40174_ ( .A({ matmul_29_bat_count[2], _13755_ }), .Y(_14136_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40175_ ( .A({ matmul_29_bat_count[3], _13755_ }), .Y(_14139_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40176_ ( .A({ matmul_29_bat_count[4], _13755_ }), .Y(_14140_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40177_ ( .A({ matmul_29_bat_count[5], _13755_ }), .Y(_14141_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40178_ ( .A({ matmul_29_bat_count[6], _13755_ }), .Y(_14142_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40179_ ( .A({ matmul_29_bat_count[7], _13755_ }), .Y(_14143_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40180_ ( .A({ matmul_29_bat_count[8], _13755_ }), .Y(_14144_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40181_ ( .A({ matmul_29_bat_count[9], _13755_ }), .Y(_14145_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40182_ ( .A({ matmul_29_bat_count[10], _13755_ }), .Y(_14115_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40183_ ( .A({ matmul_29_bat_count[11], _13755_ }), .Y(_14116_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40184_ ( .A({ matmul_29_bat_count[12], _13755_ }), .Y(_14117_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40185_ ( .A({ matmul_29_bat_count[13], _13755_ }), .Y(_14118_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40186_ ( .A({ matmul_29_bat_count[14], _13755_ }), .Y(_14119_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40187_ ( .A({ matmul_29_bat_count[15], _13755_ }), .Y(_14120_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40188_ ( .A({ matmul_29_bat_count[16], _13755_ }), .Y(_14121_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40189_ ( .A({ matmul_29_bat_count[17], _13755_ }), .Y(_14122_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40190_ ( .A({ matmul_29_bat_count[18], _13755_ }), .Y(_14123_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40191_ ( .A({ matmul_29_bat_count[19], _13755_ }), .Y(_14124_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40192_ ( .A({ matmul_29_bat_count[20], _13755_ }), .Y(_14126_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40193_ ( .A({ matmul_29_bat_count[21], _13755_ }), .Y(_14127_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40194_ ( .A({ matmul_29_bat_count[22], _13755_ }), .Y(_14128_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40195_ ( .A({ matmul_29_bat_count[23], _13755_ }), .Y(_14129_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40196_ ( .A({ matmul_29_bat_count[24], _13755_ }), .Y(_14130_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40197_ ( .A({ matmul_29_bat_count[25], _13755_ }), .Y(_14131_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40198_ ( .A({ matmul_29_bat_count[26], _13755_ }), .Y(_14132_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40199_ ( .A({ matmul_29_bat_count[27], _13755_ }), .Y(_14133_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40200_ ( .A({ matmul_29_bat_count[28], _13755_ }), .Y(_14134_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40201_ ( .A({ matmul_29_bat_count[29], _13755_ }), .Y(_14135_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40202_ ( .A({ matmul_29_bat_count[30], _13755_ }), .Y(_14137_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40203_ ( .A({ matmul_29_bat_count[31], _13755_ }), .Y(_14138_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40204_ ( .A({ _14018_, _13755_ }), .Y(_14050_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40205_ ( .A({ _14029_, _13755_ }), .Y(_14061_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40206_ ( .A({ _14040_, _13755_ }), .Y(_14072_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40207_ ( .A({ _14043_, _13755_ }), .Y(_14075_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40208_ ( .A({ _14044_, _13755_ }), .Y(_14076_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40209_ ( .A({ _14045_, _13755_ }), .Y(_14077_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40210_ ( .A({ _14046_, _13755_ }), .Y(_14078_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40211_ ( .A({ _14047_, _13755_ }), .Y(_14079_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40212_ ( .A({ _14048_, _13755_ }), .Y(_14080_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40213_ ( .A({ _14049_, _13755_ }), .Y(_14081_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40214_ ( .A({ _14019_, _13755_ }), .Y(_14051_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40215_ ( .A({ _14020_, _13755_ }), .Y(_14052_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40216_ ( .A({ _14021_, _13755_ }), .Y(_14053_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40217_ ( .A({ _14022_, _13755_ }), .Y(_14054_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40218_ ( .A({ _14023_, _13755_ }), .Y(_14055_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40219_ ( .A({ _14024_, _13755_ }), .Y(_14056_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40220_ ( .A({ _14025_, _13755_ }), .Y(_14057_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40221_ ( .A({ _14026_, _13755_ }), .Y(_14058_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40222_ ( .A({ _14027_, _13755_ }), .Y(_14059_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40223_ ( .A({ _14028_, _13755_ }), .Y(_14060_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40224_ ( .A({ _14030_, _13755_ }), .Y(_14062_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40225_ ( .A({ _14031_, _13755_ }), .Y(_14063_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40226_ ( .A({ _14032_, _13755_ }), .Y(_14064_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40227_ ( .A({ _14033_, _13755_ }), .Y(_14065_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40228_ ( .A({ _14034_, _13755_ }), .Y(_14066_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40229_ ( .A({ _14035_, _13755_ }), .Y(_14067_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40230_ ( .A({ _14036_, _13755_ }), .Y(_14068_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40231_ ( .A({ _14037_, _13755_ }), .Y(_14069_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40232_ ( .A({ _14038_, _13755_ }), .Y(_14070_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40233_ ( .A({ _14039_, _13755_ }), .Y(_14071_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40234_ ( .A({ _14041_, _13755_ }), .Y(_14073_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40235_ ( .A({ _14042_, _13755_ }), .Y(_14074_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40236_ ( .A({ _13952_, _13755_ }), .Y(_13953_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40237_ ( .A({ _13954_, _13755_ }), .Y(_13986_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40238_ ( .A({ _13965_, _13755_ }), .Y(_13997_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40239_ ( .A({ _13976_, _13755_ }), .Y(_14008_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40240_ ( .A({ _13979_, _13755_ }), .Y(_14011_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40241_ ( .A({ _13980_, _13755_ }), .Y(_14012_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40242_ ( .A({ _13981_, _13755_ }), .Y(_14013_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40243_ ( .A({ _13982_, _13755_ }), .Y(_14014_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40244_ ( .A({ _13983_, _13755_ }), .Y(_14015_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40245_ ( .A({ _13984_, _13755_ }), .Y(_14016_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40246_ ( .A({ _13985_, _13755_ }), .Y(_14017_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40247_ ( .A({ _13955_, _13755_ }), .Y(_13987_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40248_ ( .A({ _13956_, _13755_ }), .Y(_13988_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40249_ ( .A({ _13957_, _13755_ }), .Y(_13989_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40250_ ( .A({ _13958_, _13755_ }), .Y(_13990_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40251_ ( .A({ _13959_, _13755_ }), .Y(_13991_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40252_ ( .A({ _13960_, _13755_ }), .Y(_13992_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40253_ ( .A({ _13961_, _13755_ }), .Y(_13993_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40254_ ( .A({ _13962_, _13755_ }), .Y(_13994_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40255_ ( .A({ _13963_, _13755_ }), .Y(_13995_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40256_ ( .A({ _13964_, _13755_ }), .Y(_13996_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40257_ ( .A({ _13966_, _13755_ }), .Y(_13998_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40258_ ( .A({ _13967_, _13755_ }), .Y(_13999_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40259_ ( .A({ _13968_, _13755_ }), .Y(_14000_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40260_ ( .A({ _13969_, _13755_ }), .Y(_14001_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40261_ ( .A({ _13970_, _13755_ }), .Y(_14002_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40262_ ( .A({ _13971_, _13755_ }), .Y(_14003_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40263_ ( .A({ _13972_, _13755_ }), .Y(_14004_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40264_ ( .A({ _13973_, _13755_ }), .Y(_14005_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40265_ ( .A({ _13974_, _13755_ }), .Y(_14006_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40266_ ( .A({ _13975_, _13755_ }), .Y(_14007_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40267_ ( .A({ _13977_, _13755_ }), .Y(_14009_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40268_ ( .A({ _13978_, _13755_ }), .Y(_14010_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40269_ ( .A({ _13888_, _13755_ }), .Y(_13920_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40270_ ( .A({ _13899_, _13755_ }), .Y(_13931_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40271_ ( .A({ _13910_, _13755_ }), .Y(_13942_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40272_ ( .A({ _13913_, _13755_ }), .Y(_13945_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40273_ ( .A({ _13914_, _13755_ }), .Y(_13946_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40274_ ( .A({ _13915_, _13755_ }), .Y(_13947_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40275_ ( .A({ _13916_, _13755_ }), .Y(_13948_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40276_ ( .A({ _13917_, _13755_ }), .Y(_13949_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40277_ ( .A({ _13918_, _13755_ }), .Y(_13950_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40278_ ( .A({ _13919_, _13755_ }), .Y(_13951_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40279_ ( .A({ _13889_, _13755_ }), .Y(_13921_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40280_ ( .A({ _13890_, _13755_ }), .Y(_13922_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40281_ ( .A({ _13891_, _13755_ }), .Y(_13923_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40282_ ( .A({ _13892_, _13755_ }), .Y(_13924_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40283_ ( .A({ _13893_, _13755_ }), .Y(_13925_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40284_ ( .A({ _13894_, _13755_ }), .Y(_13926_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40285_ ( .A({ _13895_, _13755_ }), .Y(_13927_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40286_ ( .A({ _13896_, _13755_ }), .Y(_13928_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40287_ ( .A({ _13897_, _13755_ }), .Y(_13929_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40288_ ( .A({ _13898_, _13755_ }), .Y(_13930_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40289_ ( .A({ _13900_, _13755_ }), .Y(_13932_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40290_ ( .A({ _13901_, _13755_ }), .Y(_13933_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40291_ ( .A({ _13902_, _13755_ }), .Y(_13934_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40292_ ( .A({ _13903_, _13755_ }), .Y(_13935_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40293_ ( .A({ _13904_, _13755_ }), .Y(_13936_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40294_ ( .A({ _13905_, _13755_ }), .Y(_13937_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40295_ ( .A({ _13906_, _13755_ }), .Y(_13938_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40296_ ( .A({ _13907_, _13755_ }), .Y(_13939_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40297_ ( .A({ _13908_, _13755_ }), .Y(_13940_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40298_ ( .A({ _13909_, _13755_ }), .Y(_13941_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40299_ ( .A({ _13911_, _13755_ }), .Y(_13943_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40300_ ( .A({ _13912_, _13755_ }), .Y(_13944_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40301_ ( .A({ _13824_, _13755_ }), .Y(_13856_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40302_ ( .A({ _13835_, _13755_ }), .Y(_13867_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40303_ ( .A({ _13846_, _13755_ }), .Y(_13878_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40304_ ( .A({ _13849_, _13755_ }), .Y(_13881_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40305_ ( .A({ _13850_, _13755_ }), .Y(_13882_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40306_ ( .A({ _13851_, _13755_ }), .Y(_13883_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40307_ ( .A({ _13852_, _13755_ }), .Y(_13884_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40308_ ( .A({ _13853_, _13755_ }), .Y(_13885_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40309_ ( .A({ _13854_, _13755_ }), .Y(_13886_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40310_ ( .A({ _13855_, _13755_ }), .Y(_13887_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40311_ ( .A({ _13825_, _13755_ }), .Y(_13857_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40312_ ( .A({ _13826_, _13755_ }), .Y(_13858_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40313_ ( .A({ _13827_, _13755_ }), .Y(_13859_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40314_ ( .A({ _13828_, _13755_ }), .Y(_13860_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40315_ ( .A({ _13829_, _13755_ }), .Y(_13861_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40316_ ( .A({ _13830_, _13755_ }), .Y(_13862_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40317_ ( .A({ _13831_, _13755_ }), .Y(_13863_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40318_ ( .A({ _13832_, _13755_ }), .Y(_13864_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40319_ ( .A({ _13833_, _13755_ }), .Y(_13865_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40320_ ( .A({ _13834_, _13755_ }), .Y(_13866_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40321_ ( .A({ _13836_, _13755_ }), .Y(_13868_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40322_ ( .A({ _13837_, _13755_ }), .Y(_13869_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40323_ ( .A({ _13838_, _13755_ }), .Y(_13870_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40324_ ( .A({ _13839_, _13755_ }), .Y(_13871_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40325_ ( .A({ _13840_, _13755_ }), .Y(_13872_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40326_ ( .A({ _13841_, _13755_ }), .Y(_13873_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40327_ ( .A({ _13842_, _13755_ }), .Y(_13874_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40328_ ( .A({ _13843_, _13755_ }), .Y(_13875_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40329_ ( .A({ _13844_, _13755_ }), .Y(_13876_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40330_ ( .A({ _13845_, _13755_ }), .Y(_13877_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40331_ ( .A({ _13847_, _13755_ }), .Y(_13879_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40332_ ( .A({ _13848_, _13755_ }), .Y(_13880_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40333_ ( .A({ _13758_, _13755_ }), .Y(_13759_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40334_ ( .A({ _13756_, _13755_ }), .Y(_13757_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40335_ ( .A({ _21483_, _06930_ }), .Y(_21515_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40336_ ( .A({ _21494_, _06930_ }), .Y(_21526_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40337_ ( .A({ _21505_, _06930_ }), .Y(_21537_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40338_ ( .A({ _21508_, _06930_ }), .Y(_21540_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40339_ ( .A({ _21509_, _06930_ }), .Y(_21541_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40340_ ( .A({ _21510_, _06930_ }), .Y(_21542_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40341_ ( .A({ _21511_, _06930_ }), .Y(_21543_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40342_ ( .A({ _21512_, _06930_ }), .Y(_21544_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40343_ ( .A({ _21513_, _06930_ }), .Y(_21545_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40344_ ( .A({ _21514_, _06930_ }), .Y(_21546_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40345_ ( .A({ _21484_, _06930_ }), .Y(_21516_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40346_ ( .A({ _21485_, _06930_ }), .Y(_21517_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40347_ ( .A({ _21486_, _06930_ }), .Y(_21518_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40348_ ( .A({ _21487_, _06930_ }), .Y(_21519_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40349_ ( .A({ _21488_, _06930_ }), .Y(_21520_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40350_ ( .A({ _21489_, _06930_ }), .Y(_21521_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40351_ ( .A({ _21490_, _06930_ }), .Y(_21522_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40352_ ( .A({ _21491_, _06930_ }), .Y(_21523_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40353_ ( .A({ _21492_, _06930_ }), .Y(_21524_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40354_ ( .A({ _21493_, _06930_ }), .Y(_21525_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40355_ ( .A({ _21495_, _06930_ }), .Y(_21527_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40356_ ( .A({ _21496_, _06930_ }), .Y(_21528_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40357_ ( .A({ _21497_, _06930_ }), .Y(_21529_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40358_ ( .A({ _21498_, _06930_ }), .Y(_21530_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40359_ ( .A({ _21499_, _06930_ }), .Y(_21531_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40360_ ( .A({ _21500_, _06930_ }), .Y(_21532_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40361_ ( .A({ _21501_, _06930_ }), .Y(_21533_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40362_ ( .A({ _21502_, _06930_ }), .Y(_21534_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40363_ ( .A({ _21503_, _06930_ }), .Y(_21535_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40364_ ( .A({ _21504_, _06930_ }), .Y(_21536_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40365_ ( .A({ _21506_, _06930_ }), .Y(_21538_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40366_ ( .A({ _21507_, _06930_ }), .Y(_21539_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40367_ ( .A({ _20018_, _09298_ }), .Y(_20020_) );
  \$lut  #( .LUT(8'hd0), .WIDTH(3) ) _40368_ ( .A({ _12933_, _12929_, _05262_ }), .Y(_24028_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _40369_ ( .A({ _12932_, _12930_, _05269_, _05258_ }), .Y(_12929_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _40370_ ( .A({ _12931_, _05261_, _05260_, _05259_ }), .Y(_12930_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40371_ ( .A({ _05289_, _05288_, _05287_, _05286_ }), .Y(_12931_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40372_ ( .A({ _05285_, _05284_, _05283_, _05280_ }), .Y(_12932_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40373_ ( .A({ _12938_, _12937_, _12936_, _12934_ }), .Y(_12933_) );
  \$lut  #( .LUT(8'h10), .WIDTH(3) ) _40374_ ( .A({ _12935_, _05264_, _05263_ }), .Y(_12934_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40375_ ( .A({ _05268_, _05267_, _05266_, _05265_ }), .Y(_12935_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40376_ ( .A({ _05282_, _05281_, _05279_, _05278_ }), .Y(_12936_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40377_ ( .A({ _05277_, _05276_, _05275_, _05274_ }), .Y(_12937_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40378_ ( .A({ _05273_, _05272_, _05271_, _05270_ }), .Y(_12938_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40379_ ( .A({ _20611_, _06930_ }), .Y(_20643_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40380_ ( .A({ _20622_, _06930_ }), .Y(_20654_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40381_ ( .A({ _20633_, _06930_ }), .Y(_20665_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40382_ ( .A({ _20636_, _06930_ }), .Y(_20668_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40383_ ( .A({ _20637_, _06930_ }), .Y(_20669_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40384_ ( .A({ _20638_, _06930_ }), .Y(_20670_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40385_ ( .A({ _20639_, _06930_ }), .Y(_20671_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40386_ ( .A({ _20640_, _06930_ }), .Y(_20672_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40387_ ( .A({ _20641_, _06930_ }), .Y(_20673_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40388_ ( .A({ _20642_, _06930_ }), .Y(_20674_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40389_ ( .A({ _20612_, _06930_ }), .Y(_20644_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40390_ ( .A({ _20613_, _06930_ }), .Y(_20645_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40391_ ( .A({ _20614_, _06930_ }), .Y(_20646_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40392_ ( .A({ _20615_, _06930_ }), .Y(_20647_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40393_ ( .A({ _20616_, _06930_ }), .Y(_20648_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40394_ ( .A({ _20617_, _06930_ }), .Y(_20649_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40395_ ( .A({ _20618_, _06930_ }), .Y(_20650_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40396_ ( .A({ _20619_, _06930_ }), .Y(_20651_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40397_ ( .A({ _20620_, _06930_ }), .Y(_20652_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40398_ ( .A({ _20621_, _06930_ }), .Y(_20653_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40399_ ( .A({ _20623_, _06930_ }), .Y(_20655_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40400_ ( .A({ _20624_, _06930_ }), .Y(_20656_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40401_ ( .A({ _20625_, _06930_ }), .Y(_20657_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40402_ ( .A({ _20626_, _06930_ }), .Y(_20658_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40403_ ( .A({ _20627_, _06930_ }), .Y(_20659_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40404_ ( .A({ _20628_, _06930_ }), .Y(_20660_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40405_ ( .A({ _20629_, _06930_ }), .Y(_20661_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40406_ ( .A({ _20630_, _06930_ }), .Y(_20662_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40407_ ( .A({ _20631_, _06930_ }), .Y(_20663_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40408_ ( .A({ _20632_, _06930_ }), .Y(_20664_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40409_ ( .A({ _20634_, _06930_ }), .Y(_20666_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40410_ ( .A({ _20635_, _06930_ }), .Y(_20667_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40411_ ( .A({ _19698_, _09298_ }), .Y(_19730_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40412_ ( .A({ _19709_, _09298_ }), .Y(_19741_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40413_ ( .A({ _19720_, _09298_ }), .Y(_19752_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40414_ ( .A({ _19723_, _09298_ }), .Y(_19755_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40415_ ( .A({ _19724_, _09298_ }), .Y(_19756_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40416_ ( .A({ _19725_, _09298_ }), .Y(_19757_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40417_ ( .A({ _19726_, _09298_ }), .Y(_19758_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40418_ ( .A({ _19727_, _09298_ }), .Y(_19759_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40419_ ( .A({ _19728_, _09298_ }), .Y(_19760_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40420_ ( .A({ _19729_, _09298_ }), .Y(_19761_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40421_ ( .A({ _19699_, _09298_ }), .Y(_19731_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40422_ ( .A({ _19700_, _09298_ }), .Y(_19732_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40423_ ( .A({ _19701_, _09298_ }), .Y(_19733_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40424_ ( .A({ _19702_, _09298_ }), .Y(_19734_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40425_ ( .A({ _19703_, _09298_ }), .Y(_19735_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40426_ ( .A({ _19704_, _09298_ }), .Y(_19736_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40427_ ( .A({ _19705_, _09298_ }), .Y(_19737_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40428_ ( .A({ _19706_, _09298_ }), .Y(_19738_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40429_ ( .A({ _19707_, _09298_ }), .Y(_19739_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40430_ ( .A({ _19708_, _09298_ }), .Y(_19740_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40431_ ( .A({ _19710_, _09298_ }), .Y(_19742_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40432_ ( .A({ _19711_, _09298_ }), .Y(_19743_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40433_ ( .A({ _19712_, _09298_ }), .Y(_19744_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40434_ ( .A({ _19713_, _09298_ }), .Y(_19745_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40435_ ( .A({ _19714_, _09298_ }), .Y(_19746_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40436_ ( .A({ _19715_, _09298_ }), .Y(_19747_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40437_ ( .A({ _19716_, _09298_ }), .Y(_19748_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40438_ ( .A({ _19717_, _09298_ }), .Y(_19749_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40439_ ( .A({ _19718_, _09298_ }), .Y(_19750_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40440_ ( .A({ _19719_, _09298_ }), .Y(_19751_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40441_ ( .A({ _19721_, _09298_ }), .Y(_19753_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40442_ ( .A({ _19722_, _09298_ }), .Y(_19754_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40443_ ( .A({ _19570_, _09298_ }), .Y(_19602_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40444_ ( .A({ _19581_, _09298_ }), .Y(_19613_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40445_ ( .A({ _19592_, _09298_ }), .Y(_19624_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40446_ ( .A({ _19595_, _09298_ }), .Y(_19627_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40447_ ( .A({ _19596_, _09298_ }), .Y(_19628_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40448_ ( .A({ _19597_, _09298_ }), .Y(_19629_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40449_ ( .A({ _19598_, _09298_ }), .Y(_19630_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40450_ ( .A({ _19599_, _09298_ }), .Y(_19631_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40451_ ( .A({ _19600_, _09298_ }), .Y(_19632_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40452_ ( .A({ _19601_, _09298_ }), .Y(_19633_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40453_ ( .A({ _19571_, _09298_ }), .Y(_19603_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40454_ ( .A({ _19572_, _09298_ }), .Y(_19604_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40455_ ( .A({ _19573_, _09298_ }), .Y(_19605_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40456_ ( .A({ _19574_, _09298_ }), .Y(_19606_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40457_ ( .A({ _19575_, _09298_ }), .Y(_19607_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40458_ ( .A({ _19576_, _09298_ }), .Y(_19608_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40459_ ( .A({ _19577_, _09298_ }), .Y(_19609_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40460_ ( .A({ _19578_, _09298_ }), .Y(_19610_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40461_ ( .A({ _19579_, _09298_ }), .Y(_19611_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40462_ ( .A({ _19580_, _09298_ }), .Y(_19612_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40463_ ( .A({ _19582_, _09298_ }), .Y(_19614_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40464_ ( .A({ _19583_, _09298_ }), .Y(_19615_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40465_ ( .A({ _19584_, _09298_ }), .Y(_19616_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40466_ ( .A({ _19585_, _09298_ }), .Y(_19617_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40467_ ( .A({ _19586_, _09298_ }), .Y(_19618_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40468_ ( .A({ _19587_, _09298_ }), .Y(_19619_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40469_ ( .A({ _19588_, _09298_ }), .Y(_19620_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40470_ ( .A({ _19589_, _09298_ }), .Y(_19621_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40471_ ( .A({ _19590_, _09298_ }), .Y(_19622_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40472_ ( .A({ _19591_, _09298_ }), .Y(_19623_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40473_ ( .A({ _19593_, _09298_ }), .Y(_19625_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40474_ ( .A({ _19594_, _09298_ }), .Y(_19626_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40475_ ( .A({ _20675_, _06930_ }), .Y(_20707_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40476_ ( .A({ _20686_, _06930_ }), .Y(_20718_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40477_ ( .A({ _20697_, _06930_ }), .Y(_20729_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40478_ ( .A({ _20700_, _06930_ }), .Y(_20732_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40479_ ( .A({ _20701_, _06930_ }), .Y(_20733_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40480_ ( .A({ _20702_, _06930_ }), .Y(_20734_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40481_ ( .A({ _20703_, _06930_ }), .Y(_20735_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40482_ ( .A({ _20704_, _06930_ }), .Y(_20736_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40483_ ( .A({ _20705_, _06930_ }), .Y(_20737_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40484_ ( .A({ _20706_, _06930_ }), .Y(_20738_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40485_ ( .A({ _20676_, _06930_ }), .Y(_20708_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40486_ ( .A({ _20677_, _06930_ }), .Y(_20709_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40487_ ( .A({ _20678_, _06930_ }), .Y(_20710_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40488_ ( .A({ _20679_, _06930_ }), .Y(_20711_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40489_ ( .A({ _20680_, _06930_ }), .Y(_20712_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40490_ ( .A({ _20681_, _06930_ }), .Y(_20713_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40491_ ( .A({ _20682_, _06930_ }), .Y(_20714_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40492_ ( .A({ _20683_, _06930_ }), .Y(_20715_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40493_ ( .A({ _20684_, _06930_ }), .Y(_20716_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40494_ ( .A({ _20685_, _06930_ }), .Y(_20717_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40495_ ( .A({ _20687_, _06930_ }), .Y(_20719_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40496_ ( .A({ _20688_, _06930_ }), .Y(_20720_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40497_ ( .A({ _20689_, _06930_ }), .Y(_20721_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40498_ ( .A({ _20690_, _06930_ }), .Y(_20722_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40499_ ( .A({ _20691_, _06930_ }), .Y(_20723_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40500_ ( .A({ _20692_, _06930_ }), .Y(_20724_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40501_ ( .A({ _20693_, _06930_ }), .Y(_20725_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40502_ ( .A({ _20694_, _06930_ }), .Y(_20726_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40503_ ( .A({ _20695_, _06930_ }), .Y(_20727_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40504_ ( .A({ _20696_, _06930_ }), .Y(_20728_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40505_ ( .A({ _20698_, _06930_ }), .Y(_20730_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40506_ ( .A({ _20699_, _06930_ }), .Y(_20731_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _40507_ ( .A({ __substreamoutput_data_886[7], _12939_ }), .Y(_06174_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _40508_ ( .A({ _12940_, __substreamoutput_data_886[6:4] }), .Y(_12939_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40509_ ( .A(__substreamoutput_data_886[3:0]), .Y(_12940_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40510_ ( .A({ _12942_, _12941_ }), .Y(_24029_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40511_ ( .A(__variable_wdata_207[6:3]), .Y(_12941_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _40512_ ( .A({ __variable_wdata_207[7], __variable_wdata_207[2:0] }), .Y(_12942_) );
  \$lut  #( .LUT(8'h71), .WIDTH(3) ) _40513_ ( .A({ __variable_wdata_207[3], _reducemax_data_211[3], _12944_ }), .Y(_12943_) );
  \$lut  #( .LUT(8'hb2), .WIDTH(3) ) _40514_ ( .A({ _reducemax_data_211[2], __variable_wdata_207[2], _12945_ }), .Y(_12944_) );
  \$lut  #( .LUT(16'hd4dd), .WIDTH(4) ) _40515_ ( .A({ __variable_wdata_207[0], _reducemax_data_211[0], _reducemax_data_211[1], __variable_wdata_207[1] }), .Y(_12945_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40516_ ( .A({ _19375_, _09298_ }), .Y(_19407_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40517_ ( .A({ _19386_, _09298_ }), .Y(_19418_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40518_ ( .A({ _19397_, _09298_ }), .Y(_19429_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40519_ ( .A({ _19400_, _09298_ }), .Y(_19432_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40520_ ( .A({ _19401_, _09298_ }), .Y(_19433_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40521_ ( .A({ _19402_, _09298_ }), .Y(_19434_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40522_ ( .A({ _19403_, _09298_ }), .Y(_19435_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40523_ ( .A({ _19404_, _09298_ }), .Y(_19436_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40524_ ( .A({ _19405_, _09298_ }), .Y(_19437_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40525_ ( .A({ _19406_, _09298_ }), .Y(_19438_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40526_ ( .A({ _19376_, _09298_ }), .Y(_19408_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40527_ ( .A({ _19377_, _09298_ }), .Y(_19409_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40528_ ( .A({ _19378_, _09298_ }), .Y(_19410_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40529_ ( .A({ _19379_, _09298_ }), .Y(_19411_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40530_ ( .A({ _19380_, _09298_ }), .Y(_19412_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40531_ ( .A({ _19381_, _09298_ }), .Y(_19413_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40532_ ( .A({ _19382_, _09298_ }), .Y(_19414_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40533_ ( .A({ _19383_, _09298_ }), .Y(_19415_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40534_ ( .A({ _19384_, _09298_ }), .Y(_19416_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40535_ ( .A({ _19385_, _09298_ }), .Y(_19417_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40536_ ( .A({ _19387_, _09298_ }), .Y(_19419_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40537_ ( .A({ _19388_, _09298_ }), .Y(_19420_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40538_ ( .A({ _19389_, _09298_ }), .Y(_19421_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40539_ ( .A({ _19390_, _09298_ }), .Y(_19422_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40540_ ( .A({ _19391_, _09298_ }), .Y(_19423_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40541_ ( .A({ _19392_, _09298_ }), .Y(_19424_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40542_ ( .A({ _19393_, _09298_ }), .Y(_19425_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40543_ ( .A({ _19394_, _09298_ }), .Y(_19426_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40544_ ( .A({ _19395_, _09298_ }), .Y(_19427_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40545_ ( .A({ _19396_, _09298_ }), .Y(_19428_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40546_ ( .A({ _19398_, _09298_ }), .Y(_19430_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40547_ ( .A({ _19399_, _09298_ }), .Y(_19431_) );
  \$lut  #( .LUT(16'hbf00), .WIDTH(4) ) _40548_ ( .A({ _sra_data_42[39], _12946_, _12953_, _12951_ }), .Y(_06883_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40549_ ( .A({ _12950_, _12949_, _12948_, _12947_ }), .Y(_12946_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40550_ ( .A({ _sra_data_42[20:19], _sra_data_42[16], _sra_data_42[10] }), .Y(_12947_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40551_ ( .A({ _sra_data_42[8], _sra_data_42[38:37], _sra_data_42[34] }), .Y(_12948_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40552_ ( .A({ _sra_data_42[36:35], _sra_data_42[33], _sra_data_42[30] }), .Y(_12949_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40553_ ( .A({ _sra_data_42[29], _sra_data_42[26:25], _sra_data_42[22] }), .Y(_12950_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _40554_ ( .A({ _12952_, _sra_data_42[6], _sra_data_42[4], _sra_data_42[2] }), .Y(_12951_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40555_ ( .A({ _sra_data_42[5], _sra_data_42[3], _sra_data_42[1:0] }), .Y(_12952_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40556_ ( .A({ _12957_, _12956_, _12955_, _12954_ }), .Y(_12953_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40557_ ( .A({ _sra_data_42[17], _sra_data_42[15:13] }), .Y(_12954_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40558_ ( .A({ _sra_data_42[12:11], _sra_data_42[9], _sra_data_42[7] }), .Y(_12955_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40559_ ( .A({ _sra_data_42[32:31], _sra_data_42[28:27] }), .Y(_12956_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40560_ ( .A({ _sra_data_42[24:23], _sra_data_42[21], _sra_data_42[18] }), .Y(_12957_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _40561_ ( .A({ _sra_data_42[39], _12958_, _12963_ }), .Y(_06164_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40562_ ( .A({ _12962_, _12961_, _12960_, _12959_ }), .Y(_12958_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40563_ ( .A({ _sra_data_42[17], _sra_data_42[15:13] }), .Y(_12959_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40564_ ( .A({ _sra_data_42[12:11], _sra_data_42[9], _sra_data_42[7] }), .Y(_12960_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40565_ ( .A({ _sra_data_42[32:31], _sra_data_42[28:27] }), .Y(_12961_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40566_ ( .A({ _sra_data_42[24:23], _sra_data_42[21], _sra_data_42[18] }), .Y(_12962_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _40567_ ( .A({ _12967_, _12966_, _12965_, _12964_ }), .Y(_12963_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40568_ ( .A({ _sra_data_42[20:19], _sra_data_42[16], _sra_data_42[10] }), .Y(_12964_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40569_ ( .A({ _sra_data_42[8], _sra_data_42[38:37], _sra_data_42[34] }), .Y(_12965_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40570_ ( .A({ _sra_data_42[36:35], _sra_data_42[33], _sra_data_42[30] }), .Y(_12966_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _40571_ ( .A({ _sra_data_42[29], _sra_data_42[26:25], _sra_data_42[22] }), .Y(_12967_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40572_ ( .A({ _20739_, _06930_ }), .Y(_20771_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40573_ ( .A({ _20750_, _06930_ }), .Y(_20782_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40574_ ( .A({ _20761_, _06930_ }), .Y(_20793_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40575_ ( .A({ _20764_, _06930_ }), .Y(_20796_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40576_ ( .A({ _20765_, _06930_ }), .Y(_20797_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40577_ ( .A({ _20766_, _06930_ }), .Y(_20798_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40578_ ( .A({ _20767_, _06930_ }), .Y(_20799_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40579_ ( .A({ _20768_, _06930_ }), .Y(_20800_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40580_ ( .A({ _20769_, _06930_ }), .Y(_20801_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40581_ ( .A({ _20770_, _06930_ }), .Y(_20802_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40582_ ( .A({ _20740_, _06930_ }), .Y(_20772_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40583_ ( .A({ _20741_, _06930_ }), .Y(_20773_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40584_ ( .A({ _20742_, _06930_ }), .Y(_20774_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40585_ ( .A({ _20743_, _06930_ }), .Y(_20775_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40586_ ( .A({ _20744_, _06930_ }), .Y(_20776_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40587_ ( .A({ _20745_, _06930_ }), .Y(_20777_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40588_ ( .A({ _20746_, _06930_ }), .Y(_20778_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40589_ ( .A({ _20747_, _06930_ }), .Y(_20779_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40590_ ( .A({ _20748_, _06930_ }), .Y(_20780_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40591_ ( .A({ _20749_, _06930_ }), .Y(_20781_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40592_ ( .A({ _20751_, _06930_ }), .Y(_20783_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40593_ ( .A({ _20752_, _06930_ }), .Y(_20784_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40594_ ( .A({ _20753_, _06930_ }), .Y(_20785_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40595_ ( .A({ _20754_, _06930_ }), .Y(_20786_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40596_ ( .A({ _20755_, _06930_ }), .Y(_20787_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40597_ ( .A({ _20756_, _06930_ }), .Y(_20788_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40598_ ( .A({ _20757_, _06930_ }), .Y(_20789_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40599_ ( .A({ _20758_, _06930_ }), .Y(_20790_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40600_ ( .A({ _20759_, _06930_ }), .Y(_20791_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40601_ ( .A({ _20760_, _06930_ }), .Y(_20792_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40602_ ( .A({ _20762_, _06930_ }), .Y(_20794_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40603_ ( .A({ _20763_, _06930_ }), .Y(_20795_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40604_ ( .A({ _20022_, _09298_ }), .Y(_20054_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40605_ ( .A({ _20033_, _09298_ }), .Y(_20065_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40606_ ( .A({ _20044_, _09298_ }), .Y(_20076_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40607_ ( .A({ _20047_, _09298_ }), .Y(_20079_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40608_ ( .A({ _20048_, _09298_ }), .Y(_20080_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40609_ ( .A({ _20049_, _09298_ }), .Y(_20081_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40610_ ( .A({ _20050_, _09298_ }), .Y(_20082_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40611_ ( .A({ _20051_, _09298_ }), .Y(_20083_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40612_ ( .A({ _20052_, _09298_ }), .Y(_20084_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40613_ ( .A({ _20053_, _09298_ }), .Y(_20085_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40614_ ( .A({ _20023_, _09298_ }), .Y(_20055_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40615_ ( .A({ _20024_, _09298_ }), .Y(_20056_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40616_ ( .A({ _20025_, _09298_ }), .Y(_20057_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40617_ ( .A({ _20026_, _09298_ }), .Y(_20058_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40618_ ( .A({ _20027_, _09298_ }), .Y(_20059_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40619_ ( .A({ _20028_, _09298_ }), .Y(_20060_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40620_ ( .A({ _20029_, _09298_ }), .Y(_20061_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40621_ ( .A({ _20030_, _09298_ }), .Y(_20062_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40622_ ( .A({ _20031_, _09298_ }), .Y(_20063_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40623_ ( .A({ _20032_, _09298_ }), .Y(_20064_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40624_ ( .A({ _20034_, _09298_ }), .Y(_20066_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40625_ ( .A({ _20035_, _09298_ }), .Y(_20067_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40626_ ( .A({ _20036_, _09298_ }), .Y(_20068_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40627_ ( .A({ _20037_, _09298_ }), .Y(_20069_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40628_ ( .A({ _20038_, _09298_ }), .Y(_20070_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40629_ ( .A({ _20039_, _09298_ }), .Y(_20071_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40630_ ( .A({ _20040_, _09298_ }), .Y(_20072_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40631_ ( .A({ _20041_, _09298_ }), .Y(_20073_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40632_ ( .A({ _20042_, _09298_ }), .Y(_20074_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40633_ ( .A({ _20043_, _09298_ }), .Y(_20075_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40634_ ( .A({ _20045_, _09298_ }), .Y(_20077_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40635_ ( .A({ _20046_, _09298_ }), .Y(_20078_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40636_ ( .A({ _20803_, _06930_ }), .Y(_20835_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40637_ ( .A({ _20814_, _06930_ }), .Y(_20846_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40638_ ( .A({ _20825_, _06930_ }), .Y(_20857_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40639_ ( .A({ _20828_, _06930_ }), .Y(_20860_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40640_ ( .A({ _20829_, _06930_ }), .Y(_20861_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40641_ ( .A({ _20830_, _06930_ }), .Y(_20862_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40642_ ( .A({ _20831_, _06930_ }), .Y(_20863_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40643_ ( .A({ _20832_, _06930_ }), .Y(_20864_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40644_ ( .A({ _20833_, _06930_ }), .Y(_20865_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40645_ ( .A({ _20834_, _06930_ }), .Y(_20866_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40646_ ( .A({ _20804_, _06930_ }), .Y(_20836_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40647_ ( .A({ _20805_, _06930_ }), .Y(_20837_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40648_ ( .A({ _20806_, _06930_ }), .Y(_20838_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40649_ ( .A({ _20807_, _06930_ }), .Y(_20839_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40650_ ( .A({ _20808_, _06930_ }), .Y(_20840_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40651_ ( .A({ _20809_, _06930_ }), .Y(_20841_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40652_ ( .A({ _20810_, _06930_ }), .Y(_20842_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40653_ ( .A({ _20811_, _06930_ }), .Y(_20843_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40654_ ( .A({ _20812_, _06930_ }), .Y(_20844_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40655_ ( .A({ _20813_, _06930_ }), .Y(_20845_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40656_ ( .A({ _20815_, _06930_ }), .Y(_20847_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40657_ ( .A({ _20816_, _06930_ }), .Y(_20848_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40658_ ( .A({ _20817_, _06930_ }), .Y(_20849_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40659_ ( .A({ _20818_, _06930_ }), .Y(_20850_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40660_ ( .A({ _20819_, _06930_ }), .Y(_20851_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40661_ ( .A({ _20820_, _06930_ }), .Y(_20852_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40662_ ( .A({ _20821_, _06930_ }), .Y(_20853_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40663_ ( .A({ _20822_, _06930_ }), .Y(_20854_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40664_ ( .A({ _20823_, _06930_ }), .Y(_20855_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40665_ ( .A({ _20824_, _06930_ }), .Y(_20856_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40666_ ( .A({ _20826_, _06930_ }), .Y(_20858_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40667_ ( .A({ _20827_, _06930_ }), .Y(_20859_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40668_ ( .A({ _20867_, _06930_ }), .Y(_20899_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40669_ ( .A({ _20878_, _06930_ }), .Y(_20910_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40670_ ( .A({ _20889_, _06930_ }), .Y(_20921_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40671_ ( .A({ _20892_, _06930_ }), .Y(_20924_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40672_ ( .A({ _20893_, _06930_ }), .Y(_20925_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40673_ ( .A({ _20894_, _06930_ }), .Y(_20926_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40674_ ( .A({ _20895_, _06930_ }), .Y(_20927_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40675_ ( .A({ _20896_, _06930_ }), .Y(_20928_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40676_ ( .A({ _20897_, _06930_ }), .Y(_20929_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40677_ ( .A({ _20898_, _06930_ }), .Y(_20930_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40678_ ( .A({ _20868_, _06930_ }), .Y(_20900_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40679_ ( .A({ _20869_, _06930_ }), .Y(_20901_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40680_ ( .A({ _20870_, _06930_ }), .Y(_20902_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40681_ ( .A({ _20871_, _06930_ }), .Y(_20903_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40682_ ( .A({ _20872_, _06930_ }), .Y(_20904_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40683_ ( .A({ _20873_, _06930_ }), .Y(_20905_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40684_ ( .A({ _20874_, _06930_ }), .Y(_20906_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40685_ ( .A({ _20875_, _06930_ }), .Y(_20907_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40686_ ( .A({ _20876_, _06930_ }), .Y(_20908_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40687_ ( .A({ _20877_, _06930_ }), .Y(_20909_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40688_ ( .A({ _20879_, _06930_ }), .Y(_20911_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40689_ ( .A({ _20880_, _06930_ }), .Y(_20912_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40690_ ( .A({ _20881_, _06930_ }), .Y(_20913_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40691_ ( .A({ _20882_, _06930_ }), .Y(_20914_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40692_ ( .A({ _20883_, _06930_ }), .Y(_20915_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40693_ ( .A({ _20884_, _06930_ }), .Y(_20916_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40694_ ( .A({ _20885_, _06930_ }), .Y(_20917_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40695_ ( .A({ _20886_, _06930_ }), .Y(_20918_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40696_ ( .A({ _20887_, _06930_ }), .Y(_20919_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40697_ ( .A({ _20888_, _06930_ }), .Y(_20920_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40698_ ( .A({ _20890_, _06930_ }), .Y(_20922_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40699_ ( .A({ _20891_, _06930_ }), .Y(_20923_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40700_ ( .A({ _20931_, _06930_ }), .Y(_20963_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40701_ ( .A({ _20942_, _06930_ }), .Y(_20974_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40702_ ( .A({ _20953_, _06930_ }), .Y(_20985_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40703_ ( .A({ _20956_, _06930_ }), .Y(_20988_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40704_ ( .A({ _20957_, _06930_ }), .Y(_20989_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40705_ ( .A({ _20958_, _06930_ }), .Y(_20990_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40706_ ( .A({ _20959_, _06930_ }), .Y(_20991_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40707_ ( .A({ _20960_, _06930_ }), .Y(_20992_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40708_ ( .A({ _20961_, _06930_ }), .Y(_20993_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40709_ ( .A({ _20962_, _06930_ }), .Y(_20994_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40710_ ( .A({ _20932_, _06930_ }), .Y(_20964_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40711_ ( .A({ _20933_, _06930_ }), .Y(_20965_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40712_ ( .A({ _20934_, _06930_ }), .Y(_20966_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40713_ ( .A({ _20935_, _06930_ }), .Y(_20967_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40714_ ( .A({ _20936_, _06930_ }), .Y(_20968_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40715_ ( .A({ _20937_, _06930_ }), .Y(_20969_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40716_ ( .A({ _20938_, _06930_ }), .Y(_20970_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40717_ ( .A({ _20939_, _06930_ }), .Y(_20971_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40718_ ( .A({ _20940_, _06930_ }), .Y(_20972_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40719_ ( .A({ _20941_, _06930_ }), .Y(_20973_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40720_ ( .A({ _20943_, _06930_ }), .Y(_20975_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40721_ ( .A({ _20944_, _06930_ }), .Y(_20976_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40722_ ( .A({ _20945_, _06930_ }), .Y(_20977_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40723_ ( .A({ _20946_, _06930_ }), .Y(_20978_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40724_ ( .A({ _20947_, _06930_ }), .Y(_20979_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40725_ ( .A({ _20948_, _06930_ }), .Y(_20980_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40726_ ( .A({ _20949_, _06930_ }), .Y(_20981_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40727_ ( .A({ _20950_, _06930_ }), .Y(_20982_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40728_ ( .A({ _20951_, _06930_ }), .Y(_20983_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40729_ ( .A({ _20952_, _06930_ }), .Y(_20984_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40730_ ( .A({ _20954_, _06930_ }), .Y(_20986_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40731_ ( .A({ _20955_, _06930_ }), .Y(_20987_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _40732_ ( .A(matmul_29_next_out_write_size[1:0]), .Y(_24027_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _40733_ ( .A(cparam_matmul_29_act_bat_step[1:0]), .Y(_24026_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40734_ ( .A({ _20411_, _06930_ }), .Y(_20412_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40735_ ( .A({ _20413_, _06930_ }), .Y(_20414_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _40736_ ( .A(cparam_matmul_29_filter_read_size[2:0]), .Y(_24025_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _40737_ ( .A({ cparam_matmul_29_bias_num[0], cparam_matmul_29_bias_num[1] }), .Y(_24024_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _40738_ ( .A(conv2d_16_next_out_write_size[1:0]), .Y(_24023_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _40739_ ( .A(cparam_conv2d_16_act_offset_values_2[1:0]), .Y(_24022_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _40740_ ( .A(cparam_conv2d_16_filter_read_size[2:0]), .Y(_24021_) );
  \$lut  #( .LUT(4'h1), .WIDTH(2) ) _40741_ ( .A({ cparam_conv2d_16_bias_num[0], cparam_conv2d_16_bias_num[1] }), .Y(_24020_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40742_ ( .A({ _19890_, _09298_ }), .Y(_19922_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40743_ ( .A({ _19901_, _09298_ }), .Y(_19933_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40744_ ( .A({ _19912_, _09298_ }), .Y(_19944_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40745_ ( .A({ _19915_, _09298_ }), .Y(_19947_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40746_ ( .A({ _19916_, _09298_ }), .Y(_19948_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40747_ ( .A({ _19917_, _09298_ }), .Y(_19949_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40748_ ( .A({ _19918_, _09298_ }), .Y(_19950_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40749_ ( .A({ _19919_, _09298_ }), .Y(_19951_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40750_ ( .A({ _19920_, _09298_ }), .Y(_19952_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40751_ ( .A({ _19921_, _09298_ }), .Y(_19953_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40752_ ( .A({ _19891_, _09298_ }), .Y(_19923_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40753_ ( .A({ _19892_, _09298_ }), .Y(_19924_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40754_ ( .A({ _19893_, _09298_ }), .Y(_19925_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40755_ ( .A({ _19894_, _09298_ }), .Y(_19926_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40756_ ( .A({ _19895_, _09298_ }), .Y(_19927_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40757_ ( .A({ _19896_, _09298_ }), .Y(_19928_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40758_ ( .A({ _19897_, _09298_ }), .Y(_19929_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40759_ ( .A({ _19898_, _09298_ }), .Y(_19930_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40760_ ( .A({ _19899_, _09298_ }), .Y(_19931_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40761_ ( .A({ _19900_, _09298_ }), .Y(_19932_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40762_ ( .A({ _19902_, _09298_ }), .Y(_19934_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40763_ ( .A({ _19903_, _09298_ }), .Y(_19935_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40764_ ( .A({ _19904_, _09298_ }), .Y(_19936_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40765_ ( .A({ _19905_, _09298_ }), .Y(_19937_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40766_ ( .A({ _19906_, _09298_ }), .Y(_19938_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40767_ ( .A({ _19907_, _09298_ }), .Y(_19939_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40768_ ( .A({ _19908_, _09298_ }), .Y(_19940_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40769_ ( .A({ _19909_, _09298_ }), .Y(_19941_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40770_ ( .A({ _19910_, _09298_ }), .Y(_19942_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40771_ ( .A({ _19911_, _09298_ }), .Y(_19943_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40772_ ( .A({ _19913_, _09298_ }), .Y(_19945_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40773_ ( .A({ _19914_, _09298_ }), .Y(_19946_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40774_ ( .A({ _19505_, _09298_ }), .Y(_19537_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40775_ ( .A({ _19516_, _09298_ }), .Y(_19548_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40776_ ( .A({ _19527_, _09298_ }), .Y(_19559_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40777_ ( .A({ _19530_, _09298_ }), .Y(_19562_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40778_ ( .A({ _19531_, _09298_ }), .Y(_19563_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40779_ ( .A({ _19532_, _09298_ }), .Y(_19564_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40780_ ( .A({ _19533_, _09298_ }), .Y(_19565_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40781_ ( .A({ _19534_, _09298_ }), .Y(_19566_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40782_ ( .A({ _19535_, _09298_ }), .Y(_19567_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40783_ ( .A({ _19536_, _09298_ }), .Y(_19568_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40784_ ( .A({ _19506_, _09298_ }), .Y(_19538_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40785_ ( .A({ _19507_, _09298_ }), .Y(_19539_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40786_ ( .A({ _19508_, _09298_ }), .Y(_19540_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40787_ ( .A({ _19509_, _09298_ }), .Y(_19541_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40788_ ( .A({ _19510_, _09298_ }), .Y(_19542_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40789_ ( .A({ _19511_, _09298_ }), .Y(_19543_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40790_ ( .A({ _19512_, _09298_ }), .Y(_19544_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40791_ ( .A({ _19513_, _09298_ }), .Y(_19545_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40792_ ( .A({ _19514_, _09298_ }), .Y(_19546_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40793_ ( .A({ _19515_, _09298_ }), .Y(_19547_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40794_ ( .A({ _19517_, _09298_ }), .Y(_19549_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40795_ ( .A({ _19518_, _09298_ }), .Y(_19550_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40796_ ( .A({ _19519_, _09298_ }), .Y(_19551_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40797_ ( .A({ _19520_, _09298_ }), .Y(_19552_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40798_ ( .A({ _19521_, _09298_ }), .Y(_19553_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40799_ ( .A({ _19522_, _09298_ }), .Y(_19554_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40800_ ( .A({ _19523_, _09298_ }), .Y(_19555_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40801_ ( .A({ _19524_, _09298_ }), .Y(_19556_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40802_ ( .A({ _19525_, _09298_ }), .Y(_19557_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40803_ ( .A({ _19526_, _09298_ }), .Y(_19558_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40804_ ( .A({ _19528_, _09298_ }), .Y(_19560_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40805_ ( .A({ _19529_, _09298_ }), .Y(_19561_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40806_ ( .A({ _20415_, _06930_ }), .Y(_20416_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40807_ ( .A({ _19762_, _09298_ }), .Y(_19794_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40808_ ( .A({ _19773_, _09298_ }), .Y(_19805_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40809_ ( .A({ _19784_, _09298_ }), .Y(_19816_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40810_ ( .A({ _19787_, _09298_ }), .Y(_19819_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40811_ ( .A({ _19788_, _09298_ }), .Y(_19820_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40812_ ( .A({ _19789_, _09298_ }), .Y(_19821_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40813_ ( .A({ _19790_, _09298_ }), .Y(_19822_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40814_ ( .A({ _19791_, _09298_ }), .Y(_19823_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40815_ ( .A({ _19792_, _09298_ }), .Y(_19824_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40816_ ( .A({ _19793_, _09298_ }), .Y(_19825_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40817_ ( .A({ _19763_, _09298_ }), .Y(_19795_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40818_ ( .A({ _19764_, _09298_ }), .Y(_19796_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40819_ ( .A({ _19765_, _09298_ }), .Y(_19797_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40820_ ( .A({ _19766_, _09298_ }), .Y(_19798_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40821_ ( .A({ _19767_, _09298_ }), .Y(_19799_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40822_ ( .A({ _19768_, _09298_ }), .Y(_19800_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40823_ ( .A({ _19769_, _09298_ }), .Y(_19801_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40824_ ( .A({ _19770_, _09298_ }), .Y(_19802_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40825_ ( .A({ _19771_, _09298_ }), .Y(_19803_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40826_ ( .A({ _19772_, _09298_ }), .Y(_19804_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40827_ ( .A({ _19774_, _09298_ }), .Y(_19806_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40828_ ( .A({ _19775_, _09298_ }), .Y(_19807_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40829_ ( .A({ _19776_, _09298_ }), .Y(_19808_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40830_ ( .A({ _19777_, _09298_ }), .Y(_19809_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40831_ ( .A({ _19778_, _09298_ }), .Y(_19810_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40832_ ( .A({ _19779_, _09298_ }), .Y(_19811_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40833_ ( .A({ _19780_, _09298_ }), .Y(_19812_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40834_ ( .A({ _19781_, _09298_ }), .Y(_19813_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40835_ ( .A({ _19782_, _09298_ }), .Y(_19814_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40836_ ( .A({ _19783_, _09298_ }), .Y(_19815_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40837_ ( .A({ _19785_, _09298_ }), .Y(_19817_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40838_ ( .A({ _19786_, _09298_ }), .Y(_19818_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40839_ ( .A({ _19954_, _09298_ }), .Y(_19986_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40840_ ( .A({ _19965_, _09298_ }), .Y(_19997_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40841_ ( .A({ _19976_, _09298_ }), .Y(_20008_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40842_ ( .A({ _19979_, _09298_ }), .Y(_20011_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40843_ ( .A({ _19980_, _09298_ }), .Y(_20012_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40844_ ( .A({ _19981_, _09298_ }), .Y(_20013_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40845_ ( .A({ _19982_, _09298_ }), .Y(_20014_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40846_ ( .A({ _19983_, _09298_ }), .Y(_20015_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40847_ ( .A({ _19984_, _09298_ }), .Y(_20016_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40848_ ( .A({ _19985_, _09298_ }), .Y(_20017_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40849_ ( .A({ _19955_, _09298_ }), .Y(_19987_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40850_ ( .A({ _19956_, _09298_ }), .Y(_19988_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40851_ ( .A({ _19957_, _09298_ }), .Y(_19989_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40852_ ( .A({ _19958_, _09298_ }), .Y(_19990_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40853_ ( .A({ _19959_, _09298_ }), .Y(_19991_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40854_ ( .A({ _19960_, _09298_ }), .Y(_19992_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40855_ ( .A({ _19961_, _09298_ }), .Y(_19993_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40856_ ( .A({ _19962_, _09298_ }), .Y(_19994_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40857_ ( .A({ _19963_, _09298_ }), .Y(_19995_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40858_ ( .A({ _19964_, _09298_ }), .Y(_19996_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40859_ ( .A({ _19966_, _09298_ }), .Y(_19998_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40860_ ( .A({ _19967_, _09298_ }), .Y(_19999_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40861_ ( .A({ _19968_, _09298_ }), .Y(_20000_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40862_ ( .A({ _19969_, _09298_ }), .Y(_20001_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40863_ ( .A({ _19970_, _09298_ }), .Y(_20002_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40864_ ( .A({ _19971_, _09298_ }), .Y(_20003_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40865_ ( .A({ _19972_, _09298_ }), .Y(_20004_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40866_ ( .A({ _19973_, _09298_ }), .Y(_20005_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40867_ ( .A({ _19974_, _09298_ }), .Y(_20006_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40868_ ( .A({ _19975_, _09298_ }), .Y(_20007_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40869_ ( .A({ _19977_, _09298_ }), .Y(_20009_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40870_ ( .A({ _19978_, _09298_ }), .Y(_20010_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40871_ ( .A({ _20545_, _06930_ }), .Y(_20577_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40872_ ( .A({ _20556_, _06930_ }), .Y(_20588_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40873_ ( .A({ _20567_, _06930_ }), .Y(_20599_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40874_ ( .A({ _20570_, _06930_ }), .Y(_20602_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40875_ ( .A({ _20571_, _06930_ }), .Y(_20603_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40876_ ( .A({ _20572_, _06930_ }), .Y(_20604_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40877_ ( .A({ _20573_, _06930_ }), .Y(_20605_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40878_ ( .A({ _20574_, _06930_ }), .Y(_20606_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40879_ ( .A({ _20575_, _06930_ }), .Y(_20607_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40880_ ( .A({ _20576_, _06930_ }), .Y(_20608_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40881_ ( .A({ _20546_, _06930_ }), .Y(_20578_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40882_ ( .A({ _20547_, _06930_ }), .Y(_20579_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40883_ ( .A({ _20548_, _06930_ }), .Y(_20580_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40884_ ( .A({ _20549_, _06930_ }), .Y(_20581_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40885_ ( .A({ _20550_, _06930_ }), .Y(_20582_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40886_ ( .A({ _20551_, _06930_ }), .Y(_20583_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40887_ ( .A({ _20552_, _06930_ }), .Y(_20584_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40888_ ( .A({ _20553_, _06930_ }), .Y(_20585_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40889_ ( .A({ _20554_, _06930_ }), .Y(_20586_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40890_ ( .A({ _20555_, _06930_ }), .Y(_20587_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40891_ ( .A({ _20557_, _06930_ }), .Y(_20589_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40892_ ( .A({ _20558_, _06930_ }), .Y(_20590_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40893_ ( .A({ _20559_, _06930_ }), .Y(_20591_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40894_ ( .A({ _20560_, _06930_ }), .Y(_20592_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40895_ ( .A({ _20561_, _06930_ }), .Y(_20593_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40896_ ( .A({ _20562_, _06930_ }), .Y(_20594_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40897_ ( .A({ _20563_, _06930_ }), .Y(_20595_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40898_ ( .A({ _20564_, _06930_ }), .Y(_20596_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40899_ ( .A({ _20565_, _06930_ }), .Y(_20597_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40900_ ( .A({ _20566_, _06930_ }), .Y(_20598_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40901_ ( .A({ _20568_, _06930_ }), .Y(_20600_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40902_ ( .A({ _20569_, _06930_ }), .Y(_20601_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40903_ ( .A({ _20609_, _06930_ }), .Y(_20610_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40904_ ( .A({ _20481_, _06930_ }), .Y(_20513_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40905_ ( .A({ _20492_, _06930_ }), .Y(_20524_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40906_ ( .A({ _20503_, _06930_ }), .Y(_20535_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40907_ ( .A({ _20506_, _06930_ }), .Y(_20538_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40908_ ( .A({ _20507_, _06930_ }), .Y(_20539_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40909_ ( .A({ _20508_, _06930_ }), .Y(_20540_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40910_ ( .A({ _20509_, _06930_ }), .Y(_20541_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40911_ ( .A({ _20510_, _06930_ }), .Y(_20542_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40912_ ( .A({ _20511_, _06930_ }), .Y(_20543_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40913_ ( .A({ _20512_, _06930_ }), .Y(_20544_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40914_ ( .A({ _20482_, _06930_ }), .Y(_20514_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40915_ ( .A({ _20483_, _06930_ }), .Y(_20515_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40916_ ( .A({ _20484_, _06930_ }), .Y(_20516_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40917_ ( .A({ _20485_, _06930_ }), .Y(_20517_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40918_ ( .A({ _20486_, _06930_ }), .Y(_20518_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40919_ ( .A({ _20487_, _06930_ }), .Y(_20519_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40920_ ( .A({ _20488_, _06930_ }), .Y(_20520_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40921_ ( .A({ _20489_, _06930_ }), .Y(_20521_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40922_ ( .A({ _20490_, _06930_ }), .Y(_20522_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40923_ ( .A({ _20491_, _06930_ }), .Y(_20523_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40924_ ( .A({ _20493_, _06930_ }), .Y(_20525_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40925_ ( .A({ _20494_, _06930_ }), .Y(_20526_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40926_ ( .A({ _20495_, _06930_ }), .Y(_20527_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40927_ ( .A({ _20496_, _06930_ }), .Y(_20528_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40928_ ( .A({ _20497_, _06930_ }), .Y(_20529_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40929_ ( .A({ _20498_, _06930_ }), .Y(_20530_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40930_ ( .A({ _20499_, _06930_ }), .Y(_20531_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40931_ ( .A({ _20500_, _06930_ }), .Y(_20532_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40932_ ( .A({ _20501_, _06930_ }), .Y(_20533_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40933_ ( .A({ _20502_, _06930_ }), .Y(_20534_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40934_ ( .A({ _20504_, _06930_ }), .Y(_20536_) );
  \$lut  #( .LUT(4'h8), .WIDTH(2) ) _40935_ ( .A({ _20505_, _06930_ }), .Y(_20537_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _40936_ ( .A({ _23534_, _05685_ }), .Y(_23533_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _40937_ ( .A({ _23632_, _05686_ }), .Y(_23631_) );
  \$lut  #( .LUT(4'h4), .WIDTH(2) ) _40938_ ( .A({ _23730_, _05687_ }), .Y(_23729_) );
  \$lut  #( .LUT(16'hff80), .WIDTH(4) ) _40939_ ( .A({ _RESETN_inv_2, _saxi_register_6[0], _maxi_read_idle, _maxi_write_idle }), .Y(rst_logic) );
  \$lut  #( .LUT(8'hfe), .WIDTH(3) ) _40940_ ( .A({ _rst_logic_2, _rst_logic_1, rst_logic }), .Y(_00000_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _40941_ ( .A(_sra_data_42[39]), .Y(_06149_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _40942_ ( .A(maxi_rready), .Y(_05995_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _40943_ ( .A(RESETN), .Y(RESETN_inv) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _40944_ ( .A(_06182_), .Y(_06875_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _40945_ ( .A(_06186_), .Y(_06876_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _40946_ ( .A(_06331_), .Y(_06877_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _40947_ ( .A(__variable_wdata_797), .Y(_06142_) );
  \$lut  #( .LUT(2'h1), .WIDTH(1) ) _40948_ ( .A(__variable_wdata_798), .Y(_06143_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40949_ ( .A({ _07096_, _16806_, _16742_, _07084_ }), .Y(_12968_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _40950_ ( .A({ _07069_, _07104_, _12968_, _07095_ }), .Y(_12969_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40951_ ( .A({ _07096_, _16780_, _16716_, _07084_ }), .Y(_12970_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _40952_ ( .A({ _07112_, _07111_, _12970_, _07095_ }), .Y(_12971_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _40953_ ( .A({ _07116_, _07113_, _12975_, _12971_ }), .Y(_16492_) );
  \$lut  #( .LUT(16'h88f0), .WIDTH(4) ) _40954_ ( .A({ control_max_pool_serial_18[0], _07092_, _07081_, _16844_ }), .Y(_12972_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _40955_ ( .A({ _16460_, _05942_, _07103_, _16748_ }), .Y(_12973_) );
  \$lut  #( .LUT(16'h07ff), .WIDTH(4) ) _40956_ ( .A({ _07098_, _07086_, _07090_, _16524_ }), .Y(_12974_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _40957_ ( .A({ _12974_, _12973_, control_max_pool_serial_18[1], _12972_ }), .Y(_12975_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40958_ ( .A({ _07095_, _16791_, _16823_, _07092_ }), .Y(_12976_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _40959_ ( .A({ _07133_, _07132_, _12976_, _07096_ }), .Y(_12977_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40960_ ( .A({ _07084_, _16599_, _07091_, _16631_ }), .Y(_12978_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40961_ ( .A({ _07070_, _12978_, _07098_, _16663_ }), .Y(_12979_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40962_ ( .A({ _07095_, _16802_, _16834_, _07092_ }), .Y(_12980_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _40963_ ( .A({ _07144_, _16706_, _12980_, _07096_ }), .Y(_12981_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _40964_ ( .A({ _16485_, _05942_, _07103_, _16773_ }), .Y(_12982_) );
  \$lut  #( .LUT(16'h07ff), .WIDTH(4) ) _40965_ ( .A({ _07092_, _07080_, _07096_, _16837_ }), .Y(_12983_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40966_ ( .A({ _07090_, _16551_, _16679_, _07082_ }), .Y(_12984_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _40967_ ( .A({ _07156_, _07155_, _12984_, _07098_ }), .Y(_12985_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _40968_ ( .A({ _07160_, _07158_, _07157_, _12985_ }), .Y(_16519_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40969_ ( .A({ _07096_, _16809_, _16745_, _07084_ }), .Y(_12986_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _40970_ ( .A({ _07181_, _07180_, _12986_, _07095_ }), .Y(_12987_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _40971_ ( .A({ _07179_, _07178_, _12990_, _12987_ }), .Y(_16521_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40972_ ( .A({ _07084_, _16617_, _07091_, _16649_ }), .Y(_12988_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40973_ ( .A({ _07070_, _12988_, _07098_, _16681_ }), .Y(_12989_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _40974_ ( .A({ _07177_, _12989_, _07082_ }), .Y(_12990_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40975_ ( .A({ _07090_, _16526_, _16654_, _07082_ }), .Y(_12991_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _40976_ ( .A({ _07183_, _07182_, _12991_, _07098_ }), .Y(_12992_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _40977_ ( .A({ _07186_, _07185_, _07184_, _12992_ }), .Y(_16494_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40978_ ( .A({ _07096_, _16811_, _16747_, _07084_ }), .Y(_12993_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _40979_ ( .A({ _07192_, _07191_, _12993_, _07095_ }), .Y(_12994_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _40980_ ( .A({ _07196_, _07198_, _07197_, _07193_ }), .Y(_12995_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _40981_ ( .A({ _07195_, _07194_, _12995_, _12994_ }), .Y(_16523_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40982_ ( .A({ _07090_, _16525_, _16653_, _07082_ }), .Y(_12996_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40983_ ( .A({ _07096_, _16786_, _16722_, _07084_ }), .Y(_12997_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _40984_ ( .A({ _07206_, _07205_, _12997_, _07095_ }), .Y(_12998_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _40985_ ( .A({ _07210_, _07212_, _07211_, _07207_ }), .Y(_12999_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _40986_ ( .A({ _07209_, _07208_, _12999_, _12998_ }), .Y(_16498_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40987_ ( .A({ _07084_, _16591_, _07091_, _16623_ }), .Y(_13000_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40988_ ( .A({ _07070_, _13000_, _07098_, _16655_ }), .Y(_13001_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _40989_ ( .A({ _07213_, _13001_, _07082_ }), .Y(_13002_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _40990_ ( .A({ _07216_, _07215_, _07214_, _13002_ }), .Y(_16495_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40991_ ( .A({ _07084_, _16592_, _07091_, _16624_ }), .Y(_13003_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40992_ ( .A({ _07070_, _13003_, _07098_, _16656_ }), .Y(_13004_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _40993_ ( .A({ _07221_, _13004_, _07082_ }), .Y(_13005_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _40994_ ( .A({ _07224_, _07223_, _07222_, _13005_ }), .Y(_16496_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40995_ ( .A({ _07090_, _16529_, _16657_, _07082_ }), .Y(_13006_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _40996_ ( .A({ _07230_, _07229_, _13006_, _07098_ }), .Y(_13007_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _40997_ ( .A({ _07233_, _07232_, _07231_, _13007_ }), .Y(_16497_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _40998_ ( .A({ _07096_, _16787_, _16723_, _07084_ }), .Y(_13008_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _40999_ ( .A({ _07245_, _07246_, _13008_, _07095_ }), .Y(_13009_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41000_ ( .A({ _07244_, _07243_, _07238_, _13009_ }), .Y(_16499_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41001_ ( .A({ _07096_, _16788_, _16724_, _07084_ }), .Y(_13010_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _41002_ ( .A({ _07262_, _07261_, _13010_, _07095_ }), .Y(_13011_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _41003_ ( .A({ _07264_, _07266_, _07265_, _07263_ }), .Y(_13012_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41004_ ( .A({ _13012_, _07260_, _07259_, _13011_ }), .Y(_16500_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41005_ ( .A({ _07096_, _16789_, _16725_, _07084_ }), .Y(_13013_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _41006_ ( .A({ _07268_, _07267_, _13013_, _07095_ }), .Y(_13014_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41007_ ( .A({ _07271_, _07270_, _07269_, _13014_ }), .Y(_16501_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41008_ ( .A({ _07096_, _16790_, _16726_, _07084_ }), .Y(_13015_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _41009_ ( .A({ _07280_, _07279_, _13015_, _07095_ }), .Y(_13016_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41010_ ( .A({ _07278_, _07277_, _13019_, _13016_ }), .Y(_16502_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41011_ ( .A({ _07084_, _16598_, _07091_, _16630_ }), .Y(_13017_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41012_ ( .A({ _07070_, _13017_, _07098_, _16662_ }), .Y(_13018_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _41013_ ( .A({ _07276_, _13018_, _07082_ }), .Y(_13019_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41014_ ( .A({ _07095_, _16792_, _16824_, _07092_ }), .Y(_13020_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _41015_ ( .A({ _07284_, _07283_, _13020_, _07096_ }), .Y(_13021_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41016_ ( .A({ _13023_, _07282_, _07281_, _13021_ }), .Y(_16504_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41017_ ( .A({ _07088_, _16696_, _07095_, _16728_ }), .Y(_13022_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _41018_ ( .A({ _07285_, _07286_, _13022_, _07084_ }), .Y(_13023_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41019_ ( .A({ _07096_, _16793_, _16729_, _07084_ }), .Y(_13024_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _41020_ ( .A({ _07291_, _07290_, _13024_, _07095_ }), .Y(_13025_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41021_ ( .A({ _07289_, _07288_, _13028_, _13025_ }), .Y(_16505_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41022_ ( .A({ _07084_, _16601_, _07091_, _16633_ }), .Y(_13026_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41023_ ( .A({ _07070_, _13026_, _07098_, _16665_ }), .Y(_13027_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _41024_ ( .A({ _07287_, _13027_, _07082_ }), .Y(_13028_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41025_ ( .A({ _07096_, _16797_, _16733_, _07084_ }), .Y(_13029_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _41026_ ( .A({ _07293_, _07292_, _13029_, _07095_ }), .Y(_13030_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _41027_ ( .A({ _07297_, _07299_, _07298_, _07294_ }), .Y(_13031_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41028_ ( .A({ _07296_, _07295_, _13031_, _13030_ }), .Y(_16509_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41029_ ( .A({ _07090_, _16539_, _16667_, _07082_ }), .Y(_13032_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _41030_ ( .A({ _07301_, _07300_, _13032_, _07098_ }), .Y(_13033_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _41031_ ( .A({ _07306_, _07307_, _07305_, _07302_ }), .Y(_13034_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41032_ ( .A({ _07304_, _07303_, _13034_, _13033_ }), .Y(_16507_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _41033_ ( .A({ _07084_, _16606_, _07091_, _16638_ }), .Y(_13035_) );
  \$lut  #( .LUT(16'h880f), .WIDTH(4) ) _41034_ ( .A({ control_max_pool_serial_18[2], _13035_, _07080_, _16574_ }), .Y(_13036_) );
  \$lut  #( .LUT(16'h00bf), .WIDTH(4) ) _41035_ ( .A({ _07320_, _13036_, _07070_, control_max_pool_serial_18[3] }), .Y(_13037_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41036_ ( .A({ _07096_, _16799_, _16735_, _07084_ }), .Y(_13038_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _41037_ ( .A({ _07344_, _07343_, _13038_, _07095_ }), .Y(_13039_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41038_ ( .A({ _07342_, _07341_, _13042_, _13039_ }), .Y(_16511_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41039_ ( .A({ _07084_, _16607_, _07091_, _16639_ }), .Y(_13040_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41040_ ( .A({ _07070_, _13040_, _07098_, _16671_ }), .Y(_13041_) );
  \$lut  #( .LUT(8'h07), .WIDTH(3) ) _41041_ ( .A({ _07340_, _13041_, _07082_ }), .Y(_13042_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41042_ ( .A({ _07095_, _16801_, _16833_, _07092_ }), .Y(_13043_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _41043_ ( .A({ _07348_, _07347_, _13043_, _07096_ }), .Y(_13044_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41044_ ( .A({ _07349_, _07346_, _07345_, _13044_ }), .Y(_16513_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41045_ ( .A({ _07090_, _16548_, _16676_, _07082_ }), .Y(_13045_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _41046_ ( .A({ _07911_, _07910_, _07904_, _06012_ }), .Y(_13046_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _41047_ ( .A({ _07906_, _13046_, _22376_, _07460_ }), .Y(_13047_) );
  \$lut  #( .LUT(16'h01ff), .WIDTH(4) ) _41048_ ( .A({ _07905_, _07909_, _07468_, _07490_ }), .Y(_13048_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41049_ ( .A({ _07922_, _07912_, _13048_, _13047_ }), .Y(_22088_) );
  \$lut  #( .LUT(16'hfeff), .WIDTH(4) ) _41050_ ( .A({ _07931_, _07920_, _07909_, _07468_ }), .Y(_13049_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _41051_ ( .A({ _07927_, _07917_, _13049_, _07484_ }), .Y(_13050_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _41052_ ( .A({ _07933_, _06016_, _07929_, _07928_ }), .Y(_13051_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _41053_ ( .A({ _13051_, _13050_, _22407_, _07478_ }), .Y(_13052_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _41054_ ( .A({ _07960_, _07957_, _22758_, _06021_ }), .Y(_13053_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _41055_ ( .A({ _07995_, _07992_, _07993_, _07994_ }), .Y(_13054_) );
  \$lut  #( .LUT(16'h30ea), .WIDTH(4) ) _41056_ ( .A({ control_conv2d_16[3], _07930_, control_conv2d_16[2], _07484_ }), .Y(_13055_) );
  \$lut  #( .LUT(16'hef00), .WIDTH(4) ) _41057_ ( .A({ _08007_, _13055_, control_conv2d_16[1:0] }), .Y(_13056_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _41058_ ( .A({ _08006_, _08001_, _07983_, _13056_ }), .Y(_13057_) );
  \$lut  #( .LUT(8'h7f), .WIDTH(3) ) _41059_ ( .A({ _08014_, _08008_, _13057_ }), .Y(_22061_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _41060_ ( .A({ _08118_, _08117_, _14872_, _08070_ }), .Y(_13058_) );
  \$lut  #( .LUT(16'h035f), .WIDTH(4) ) _41061_ ( .A({ _08057_, _08051_, _08038_, _08053_ }), .Y(_13059_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _41062_ ( .A({ _08116_, _05931_, _13059_, _08040_ }), .Y(_13060_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41063_ ( .A({ _08113_, _08108_, _13060_, _13058_ }), .Y(_14744_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _41064_ ( .A({ _08060_, _15163_, _08043_, _08054_ }), .Y(_13061_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _41065_ ( .A({ _08129_, _08075_, _13061_, _08048_ }), .Y(_13062_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _41066_ ( .A({ _08131_, _08130_, _08128_, _13062_ }), .Y(_13063_) );
  \$lut  #( .LUT(16'h8fff), .WIDTH(4) ) _41067_ ( .A({ _08121_, _13063_, _14907_, _08069_ }), .Y(_14747_) );
  \$lut  #( .LUT(16'h1fff), .WIDTH(4) ) _41068_ ( .A({ _06923_, _06920_, _06928_, _07459_ }), .Y(_13064_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _41069_ ( .A({ _08504_, _07917_, _13064_, _07484_ }), .Y(_24076_) );
  \$lut  #( .LUT(16'h01fc), .WIDTH(4) ) _41070_ ( .A({ _09039_, _06902_, _06896_, _06910_ }), .Y(_13065_) );
  \$lut  #( .LUT(16'hc700), .WIDTH(4) ) _41071_ ( .A({ _09079_, _09039_, _13065_, _06901_ }), .Y(_13066_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _41072_ ( .A({ _09078_, _09077_, _09071_, _13066_ }), .Y(_13067_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _41073_ ( .A({ _09039_, _06908_, _06903_, _06901_ }), .Y(_13068_) );
  \$lut  #( .LUT(16'hf400), .WIDTH(4) ) _41074_ ( .A({ _09047_, _09052_, _13068_, _06886_ }), .Y(_13069_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41075_ ( .A({ _09107_, _09100_, _09091_, _13069_ }), .Y(_23192_) );
  \$lut  #( .LUT(16'h01ff), .WIDTH(4) ) _41076_ ( .A({ _06903_, _06914_, _06911_, _06902_ }), .Y(_13070_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _41077_ ( .A({ _13070_, _09039_, _06902_, _07451_ }), .Y(_13071_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _41078_ ( .A({ _09146_, _09074_, _24081_, _24077_ }), .Y(_13072_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _41079_ ( .A({ _09151_, _09147_, _13072_, _13071_ }), .Y(_13073_) );
  \$lut  #( .LUT(16'h0bff), .WIDTH(4) ) _41080_ ( .A({ _09306_, _09307_, cparam_matmul_29_max_och_count[1], matmul_29_och_count[1] }), .Y(_13074_) );
  \$lut  #( .LUT(16'hb222), .WIDTH(4) ) _41081_ ( .A({ _09308_, _13074_, cparam_matmul_29_max_och_count[4], matmul_29_och_count[4] }), .Y(_13075_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _41082_ ( .A({ _09310_, _09311_, _13075_, _09309_ }), .Y(_13076_) );
  \$lut  #( .LUT(16'h8fff), .WIDTH(4) ) _41083_ ( .A({ _09316_, _13076_, _09307_, _09312_ }), .Y(_06146_) );
  \$lut  #( .LUT(16'h0bff), .WIDTH(4) ) _41084_ ( .A({ _09355_, _09358_, _09356_, _09325_ }), .Y(_13077_) );
  \$lut  #( .LUT(8'hb0), .WIDTH(3) ) _41085_ ( .A({ _09365_, _09342_, _09359_ }), .Y(_13078_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _41086_ ( .A({ _13078_, _09341_, _13077_, _09357_ }), .Y(_06162_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _41087_ ( .A({ max_pool_serial_18_col_count[3], cparam_max_pool_serial_18_max_col_count[3], _09386_, _09385_ }), .Y(_13079_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _41088_ ( .A({ _13079_, cparam_max_pool_serial_18_max_col_count[4], _09382_, max_pool_serial_18_col_count[4] }), .Y(_13080_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _41089_ ( .A({ _09391_, _09387_, _13080_, max_pool_serial_18_col_count[5] }), .Y(_06161_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _41090_ ( .A({ max_pool_serial_18_row_count[3], cparam_max_pool_serial_18_max_col_count[3], _09409_, _09408_ }), .Y(_13081_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _41091_ ( .A({ _13081_, cparam_max_pool_serial_18_max_col_count[4], _09405_, max_pool_serial_18_row_count[4] }), .Y(_13082_) );
  \$lut  #( .LUT(8'hbf), .WIDTH(3) ) _41092_ ( .A({ _09396_, _13082_, max_pool_serial_18_row_count[5] }), .Y(_06160_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _41093_ ( .A({ _09451_, _09433_, _09444_, _09410_ }), .Y(_13083_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _41094_ ( .A({ _09452_, _09446_, _13083_, _09457_ }), .Y(_06159_) );
  \$lut  #( .LUT(16'hffb0), .WIDTH(4) ) _41095_ ( .A({ _09570_, _09569_, _09564_, _09551_ }), .Y(_13084_) );
  \$lut  #( .LUT(16'h07ff), .WIDTH(4) ) _41096_ ( .A({ _09572_, _09571_, _13084_, _09568_ }), .Y(_13085_) );
  \$lut  #( .LUT(16'h70ff), .WIDTH(4) ) _41097_ ( .A({ _09592_, _09586_, _13085_, _09580_ }), .Y(_06153_) );
  \$lut  #( .LUT(8'h81), .WIDTH(3) ) _41098_ ( .A({ _09645_, _pulse_count_213[6], _23984_ }), .Y(_13086_) );
  \$lut  #( .LUT(16'h2bb2), .WIDTH(4) ) _41099_ ( .A({ _13086_, _23984_, _pulse_count_213[7], _23985_ }), .Y(_13087_) );
  \$lut  #( .LUT(8'h81), .WIDTH(3) ) _41100_ ( .A({ _09700_, _pulse_count_19[18], _23932_ }), .Y(_13088_) );
  \$lut  #( .LUT(16'hd44d), .WIDTH(4) ) _41101_ ( .A({ _23932_, _13088_, _pulse_count_19[19], _23933_ }), .Y(_13089_) );
  \$lut  #( .LUT(8'h0b), .WIDTH(3) ) _41102_ ( .A({ _09701_, _09696_, _09698_ }), .Y(_13090_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _41103_ ( .A({ _13090_, _13089_, _09695_ }), .Y(_13091_) );
  \$lut  #( .LUT(8'h01), .WIDTH(3) ) _41104_ ( .A({ _09767_, _09765_, _09754_ }), .Y(_13092_) );
  \$lut  #( .LUT(16'h8eaf), .WIDTH(4) ) _41105_ ( .A({ _13092_, _23948_, _09718_, _reduceadd_count_17[32] }), .Y(_06147_) );
  \$lut  #( .LUT(16'hd42b), .WIDTH(4) ) _41106_ ( .A({ cparam_max_pool_serial_18_act_num_col[5], _09858_, _03906_, cparam_max_pool_serial_18_act_num_col[4] }), .Y(_13093_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _41107_ ( .A({ _09869_, _09863_, _03881_, _03911_ }), .Y(_13094_) );
  \$lut  #( .LUT(16'ha3ff), .WIDTH(4) ) _41108_ ( .A({ _13094_, _13093_, cparam_max_pool_serial_18_act_num_col[5], _03907_ }), .Y(max_pool_serial_18_dma_pad_mask_1) );
  \$lut  #( .LUT(16'h370c), .WIDTH(4) ) _41109_ ( .A({ _09881_, _09882_, _09879_, _09880_ }), .Y(_13095_) );
  \$lut  #( .LUT(16'h2bb2), .WIDTH(4) ) _41110_ ( .A({ _13095_, _09879_, cparam_conv2d_16_act_num_row[4], conv2d_16_out_row_count[4] }), .Y(_13096_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _41111_ ( .A({ _09870_, _13096_, cparam_conv2d_16_act_num_row[5], conv2d_16_out_row_count[5] }), .Y(conv2d_16_dma_out_mask_0) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _41112_ ( .A({ conv2d_16_row_count[12], _05293_, _05294_, conv2d_16_row_count[13] }), .Y(_13097_) );
  \$lut  #( .LUT(16'h2fff), .WIDTH(4) ) _41113_ ( .A({ _10244_, _13097_, _13102_, _10241_ }), .Y(_13098_) );
  \$lut  #( .LUT(16'h70ff), .WIDTH(4) ) _41114_ ( .A({ _10245_, _10255_, _10257_, _13098_ }), .Y(_13099_) );
  \$lut  #( .LUT(16'h80ff), .WIDTH(4) ) _41115_ ( .A({ _13105_, _10270_, _10260_, _13099_ }), .Y(conv2d_16_dma_pad_mask_0) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _41116_ ( .A({ conv2d_16_row_count[9], _05321_, conv2d_16_row_count[8], _05320_ }), .Y(_13100_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _41117_ ( .A({ _10238_, _13100_, _05319_, conv2d_16_row_count[7] }), .Y(_13101_) );
  \$lut  #( .LUT(16'h1f00), .WIDTH(4) ) _41118_ ( .A({ _13101_, _10240_, _10239_, _10231_ }), .Y(_13102_) );
  \$lut  #( .LUT(16'h0bff), .WIDTH(4) ) _41119_ ( .A({ _10262_, _10265_, _10263_, _10266_ }), .Y(_13103_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _41120_ ( .A({ _13103_, _10267_, _10260_, _10268_ }), .Y(_13104_) );
  \$lut  #( .LUT(16'hbf00), .WIDTH(4) ) _41121_ ( .A({ _13104_, _10269_, _09531_, conv2d_16_row_count[0] }), .Y(_13105_) );
  \$lut  #( .LUT(16'hffb0), .WIDTH(4) ) _41122_ ( .A({ _10287_, _10285_, _10281_, _13111_ }), .Y(_13106_) );
  \$lut  #( .LUT(16'h07ff), .WIDTH(4) ) _41123_ ( .A({ _10305_, _10286_, _13106_, _10284_ }), .Y(_13107_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _41124_ ( .A({ _13114_, _10309_, _10314_ }), .Y(_13108_) );
  \$lut  #( .LUT(16'h70ff), .WIDTH(4) ) _41125_ ( .A({ _13108_, _10298_, _13107_, _10288_ }), .Y(conv2d_16_dma_pad_mask_1) );
  \$lut  #( .LUT(16'hff2b), .WIDTH(4) ) _41126_ ( .A({ _10271_, _10272_, _05344_, _05312_ }), .Y(_13109_) );
  \$lut  #( .LUT(16'hff70), .WIDTH(4) ) _41127_ ( .A({ _10274_, _10275_, _13109_, _10273_ }), .Y(_13110_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _41128_ ( .A({ _10276_, _10280_, _13110_, _10279_ }), .Y(_13111_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _41129_ ( .A({ _05338_, _05339_, _05306_, _05307_ }), .Y(_13112_) );
  \$lut  #( .LUT(16'h07ff), .WIDTH(4) ) _41130_ ( .A({ _10300_, _10307_, _13112_, _10304_ }), .Y(_13113_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _41131_ ( .A({ _10308_, _13113_, _10301_, _10303_ }), .Y(_13114_) );
  \$lut  #( .LUT(16'hffb0), .WIDTH(4) ) _41132_ ( .A({ _10345_, _10338_, _10333_, _10319_ }), .Y(_13115_) );
  \$lut  #( .LUT(16'h07ff), .WIDTH(4) ) _41133_ ( .A({ _10339_, _10346_, _13115_, _10337_ }), .Y(_13116_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _41134_ ( .A({ _10347_, _10375_, _13116_, _10369_ }), .Y(conv2d_16_dma_pad_mask_2) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _41135_ ( .A({ _05321_, conv2d_16_col_count[9:8], _05320_ }), .Y(_13117_) );
  \$lut  #( .LUT(16'hb000), .WIDTH(4) ) _41136_ ( .A({ _10387_, _13117_, _05319_, conv2d_16_col_count[7] }), .Y(_13118_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _41137_ ( .A({ _10388_, _13118_, _10391_, _10378_ }), .Y(_13119_) );
  \$lut  #( .LUT(16'h8f00), .WIDTH(4) ) _41138_ ( .A({ _10392_, _10413_, _13119_, _10410_ }), .Y(_13120_) );
  \$lut  #( .LUT(16'h7150), .WIDTH(4) ) _41139_ ( .A({ conv2d_16_row_count_buf[8], conv2d_16_row_count_buf[9], _05320_, _05321_ }), .Y(_13121_) );
  \$lut  #( .LUT(8'h70), .WIDTH(3) ) _41140_ ( .A({ _10440_, _13121_, _10439_ }), .Y(_13122_) );
  \$lut  #( .LUT(16'h4f00), .WIDTH(4) ) _41141_ ( .A({ _13122_, _10441_, _10443_, _10430_ }), .Y(_13123_) );
  \$lut  #( .LUT(16'h9009), .WIDTH(4) ) _41142_ ( .A({ _05298_, _05394_, _05393_, _05297_ }), .Y(_13124_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _41143_ ( .A({ _10516_, _10513_, _13124_ }), .Y(_13125_) );
  \$lut  #( .LUT(8'h80), .WIDTH(3) ) _41144_ ( .A({ _10509_, _10505_, _13125_ }), .Y(_13126_) );
  \$lut  #( .LUT(8'h18), .WIDTH(3) ) _41145_ ( .A({ _10739_, cparam_max_pool_serial_18_act_num_col[3], max_pool_serial_18_col_count[3] }), .Y(_13127_) );
  \$lut  #( .LUT(16'hd44d), .WIDTH(4) ) _41146_ ( .A({ _13127_, max_pool_serial_18_col_count[3], cparam_max_pool_serial_18_act_num_col[4], max_pool_serial_18_col_count[4] }), .Y(_13128_) );
  \$lut  #( .LUT(16'hd42b), .WIDTH(4) ) _41147_ ( .A({ cparam_max_pool_serial_18_act_num_col[5], _10743_, max_pool_serial_18_row_count_buf[4], cparam_max_pool_serial_18_act_num_col[4] }), .Y(_13129_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _41148_ ( .A({ _10754_, _10748_, max_pool_serial_18_row_count_buf[10:9] }), .Y(_13130_) );
  \$lut  #( .LUT(16'h5c00), .WIDTH(4) ) _41149_ ( .A({ _13130_, _13129_, cparam_max_pool_serial_18_act_num_col[5], max_pool_serial_18_row_count_buf[5] }), .Y(_13131_) );
  \$lut  #( .LUT(16'hd42b), .WIDTH(4) ) _41150_ ( .A({ cparam_max_pool_serial_18_act_num_col[5], _10755_, _03938_, cparam_max_pool_serial_18_act_num_col[4] }), .Y(_13132_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _41151_ ( .A({ _10766_, _10760_, _03913_, _03943_ }), .Y(_13133_) );
  \$lut  #( .LUT(16'h5c00), .WIDTH(4) ) _41152_ ( .A({ _13133_, _13132_, cparam_max_pool_serial_18_act_num_col[5], _03939_ }), .Y(_13134_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _41153_ ( .A({ _10779_, _10773_, _03945_, _03975_ }), .Y(_13135_) );
  \$lut  #( .LUT(16'h2b00), .WIDTH(4) ) _41154_ ( .A({ _13135_, _10767_, _03971_, cparam_max_pool_serial_18_act_num_col[5] }), .Y(_13136_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _41155_ ( .A({ _12785_, _12784_, conv2d_16_prev_row_count[2], cparam_conv2d_16_max_col_count[2] }), .Y(_13137_) );
  \$lut  #( .LUT(16'hf444), .WIDTH(4) ) _41156_ ( .A({ _12783_, _13137_, cparam_conv2d_16_max_col_count[4], conv2d_16_prev_row_count[4] }), .Y(_13138_) );
  \$lut  #( .LUT(16'h007f), .WIDTH(4) ) _41157_ ( .A({ conv2d_16_skip_write_out, _12786_, _12775_, _13138_ }), .Y(_06821_) );
  \$lut  #( .LUT(8'h2b), .WIDTH(3) ) _41158_ ( .A({ _12861_, cparam_max_pool_serial_18_max_col_count[2], max_pool_serial_18_prev_row_count[2] }), .Y(_13139_) );
  \$lut  #( .LUT(16'hb0ff), .WIDTH(4) ) _41159_ ( .A({ _12860_, _13139_, cparam_max_pool_serial_18_max_col_count[3], max_pool_serial_18_prev_row_count[3] }), .Y(_13140_) );
  \$lut  #( .LUT(16'h2bd4), .WIDTH(4) ) _41160_ ( .A({ __variable_wdata_207[7], _13143_, _reducemax_data_211[6], __variable_wdata_207[6] }), .Y(_13141_) );
  \$lut  #( .LUT(8'ha3), .WIDTH(3) ) _41161_ ( .A({ _13141_, __variable_wdata_207[7], _reducemax_data_211[7] }), .Y(_06884_) );
  \$lut  #( .LUT(8'h18), .WIDTH(3) ) _41162_ ( .A({ _12943_, _reducemax_data_211[4], __variable_wdata_207[4] }), .Y(_13142_) );
  \$lut  #( .LUT(16'hd44d), .WIDTH(4) ) _41163_ ( .A({ __variable_wdata_207[4], _13142_, _reducemax_data_211[5], __variable_wdata_207[5] }), .Y(_13143_) );
  \$lut  #( .LUT(16'h7077), .WIDTH(4) ) _41164_ ( .A({ _16486_, _05942_, _07103_, _16774_ }), .Y(_13144_) );
  \$lut  #( .LUT(16'h07ff), .WIDTH(4) ) _41165_ ( .A({ _07080_, _07088_, _16870_, _07081_ }), .Y(_13145_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _41166_ ( .A({ _07135_, _07138_, _07137_, _07136_ }), .Y(_13146_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41167_ ( .A({ _07090_, _16546_, _16674_, _07082_ }), .Y(_13147_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _41168_ ( .A({ _07140_, _07139_, _13147_, _07098_ }), .Y(_13148_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _41169_ ( .A({ _07145_, _07148_, _07147_, _07146_ }), .Y(_13149_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41170_ ( .A({ _12981_, _13149_, _07141_, _13148_ }), .Y(_16514_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41171_ ( .A({ _07096_, _16805_, _16741_, _07084_ }), .Y(_13150_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _41172_ ( .A({ _12983_, _12982_, _07151_, _07150_ }), .Y(_13151_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41173_ ( .A({ _07088_, _16685_, _07095_, _16717_ }), .Y(_13152_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _41174_ ( .A({ _07084_, _13152_, _12996_, _07098_ }), .Y(_13153_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _41175_ ( .A({ _07203_, _07204_, _07202_, _07201_ }), .Y(_13154_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41176_ ( .A({ _13154_, _07200_, _07199_, _13153_ }), .Y(_16493_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41177_ ( .A({ _07096_, _16804_, _16740_, _07084_ }), .Y(_13155_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _41178_ ( .A({ _07095_, _13155_, _13045_, _07098_ }), .Y(_13156_) );
  \$lut  #( .LUT(16'h0100), .WIDTH(4) ) _41179_ ( .A({ _07369_, _07371_, _07370_, _07368_ }), .Y(_13157_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41180_ ( .A({ _13157_, _07367_, _07366_, _13156_ }), .Y(_16516_) );
  \$lut  #( .LUT(16'h0cce), .WIDTH(4) ) _41181_ ( .A({ control_conv2d_16[1:0], _07930_, _07905_ }), .Y(_13158_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _41182_ ( .A({ _07952_, _07951_, _06015_, _06013_ }), .Y(_13159_) );
  \$lut  #( .LUT(16'h7000), .WIDTH(4) ) _41183_ ( .A({ _07945_, _13159_, _13158_, _07474_ }), .Y(_13160_) );
  \$lut  #( .LUT(16'h0c0a), .WIDTH(4) ) _41184_ ( .A({ control_conv2d_16[3:2], _07484_, _07918_ }), .Y(_13161_) );
  \$lut  #( .LUT(16'he304), .WIDTH(4) ) _41185_ ( .A({ _13161_, control_conv2d_16[1:0], control_conv2d_16[3] }), .Y(_13162_) );
  \$lut  #( .LUT(8'hd3), .WIDTH(3) ) _41186_ ( .A({ _13162_, _13161_, _07905_ }), .Y(_13163_) );
  \$lut  #( .LUT(16'h8000), .WIDTH(4) ) _41187_ ( .A({ _07986_, _07985_, _06017_, _07982_ }), .Y(_13164_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41188_ ( .A({ _13054_, _07996_, _13164_, _13163_ }), .Y(_22072_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41189_ ( .A({ _07090_, _16550_, _16678_, _07082_ }), .Y(_13165_) );
  \$lut  #( .LUT(16'h0007), .WIDTH(4) ) _41190_ ( .A({ _07108_, _07107_, _13165_, _07098_ }), .Y(_13166_) );
  \$lut  #( .LUT(16'h1000), .WIDTH(4) ) _41191_ ( .A({ _13145_, _13144_, _07110_, _07109_ }), .Y(_13167_) );
  \$lut  #( .LUT(16'hbfff), .WIDTH(4) ) _41192_ ( .A({ _12969_, _13167_, _13166_, _07105_ }), .Y(_16518_) );
  \$lut  #( .LUT(16'h07ff), .WIDTH(4) ) _41193_ ( .A({ _07088_, _07091_, _16695_, _07084_ }), .Y(_13168_) );
  \$lut  #( .LUT(16'h7f00), .WIDTH(4) ) _41194_ ( .A({ _13168_, _07095_, _07084_, _16727_ }), .Y(_13169_) );
  \$lut  #( .LUT(16'h0700), .WIDTH(4) ) _41195_ ( .A({ _07134_, _24044_, _07082_, _12979_ }), .Y(_13170_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41196_ ( .A({ _13146_, _12977_, _13170_, _13169_ }), .Y(_16503_) );
  \$lut  #( .LUT(16'hf888), .WIDTH(4) ) _41197_ ( .A({ _07090_, _16549_, _16677_, _07082_ }), .Y(_13171_) );
  \$lut  #( .LUT(16'h0777), .WIDTH(4) ) _41198_ ( .A({ _07098_, _13171_, _13150_, _07095_ }), .Y(_13172_) );
  \$lut  #( .LUT(16'h0001), .WIDTH(4) ) _41199_ ( .A({ _07154_, _07153_, _07152_, _07149_ }), .Y(_13173_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41200_ ( .A({ _13151_, _13173_, _07145_, _13172_ }), .Y(_16517_) );
  \$lut  #( .LUT(16'hf0ee), .WIDTH(4) ) _41201_ ( .A({ _07490_, _22502_, _07909_, _07468_ }), .Y(_13174_) );
  \$lut  #( .LUT(16'h133f), .WIDTH(4) ) _41202_ ( .A({ _07490_, _13174_, _07905_, _07484_ }), .Y(_13175_) );
  \$lut  #( .LUT(16'h4000), .WIDTH(4) ) _41203_ ( .A({ _07936_, _07955_, _07953_, _07956_ }), .Y(_13176_) );
  \$lut  #( .LUT(16'h7fff), .WIDTH(4) ) _41204_ ( .A({ _13160_, _13053_, _13176_, _13175_ }), .Y(_22086_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41205_ ( .A(max_pool_serial_18_act_base_offset_row), .B(max_pool_serial_18_act_base_offset_bat), .Y(max_pool_serial_18_act_base_offset) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41206_ ( .A(max_pool_serial_18_out_base_offset_row), .B(max_pool_serial_18_out_base_offset_bat), .Y(max_pool_serial_18_out_base_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41207_ ( .A(max_pool_serial_18_row_count), .B(1), .Y({ _03904_, _03903_, _03901_, _03900_, _03899_, _03898_, _03897_, _03896_, _03895_, _03894_, _03893_, _03892_, _03890_, _03889_, _03888_, _03887_, _03886_, _03885_, _03884_, _03883_, _03882_, _03881_, _03911_, _03910_, _03909_, _03908_, _03907_, _03906_, _03905_, _03902_, _03891_, _03880_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41208_ ( .A(max_pool_serial_18_col_count), .B(1), .Y({ _03936_, _03935_, _03933_, _03932_, _03931_, _03930_, _03929_, _03928_, _03927_, _03926_, _03925_, _03924_, _03922_, _03921_, _03920_, _03919_, _03918_, _03917_, _03916_, _03915_, _03914_, _03913_, _03943_, _03942_, _03941_, _03940_, _03939_, _03938_, _03937_, _03934_, _03923_, _03912_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41209_ ( .A(max_pool_serial_18_row_count_buf), .B(1), .Y({ _03968_, _03967_, _03965_, _03964_, _03963_, _03962_, _03961_, _03960_, _03959_, _03958_, _03957_, _03956_, _03954_, _03953_, _03952_, _03951_, _03950_, _03949_, _03948_, _03947_, _03946_, _03945_, _03975_, _03974_, _03973_, _03972_, _03971_, _03970_, _03969_, _03966_, _03955_, _03944_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41210_ ( .A(_stream_max_pool_serial_18_source_1_source_offset_buf), .B(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_0), .Y(_24196_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41211_ ( .A(_24196_), .B(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_1), .Y(_24197_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41212_ ( .A(_24197_), .B(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_2), .Y(_24198_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41213_ ( .A(_24198_), .B(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_3), .Y(_stream_max_pool_serial_18_source_1_source_pat_all_offset) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41214_ ( .A(matmul_29_act_base_offset_row), .B(matmul_29_act_base_offset_bat), .Y(matmul_29_act_base_offset) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41215_ ( .A(matmul_29_out_base_offset_val), .B(matmul_29_out_base_offset_col), .Y(_24199_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41216_ ( .A(_24199_), .B(matmul_29_out_base_offset_row), .Y(_24200_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41217_ ( .A(_24200_), .B(matmul_29_out_base_offset_bat), .Y(_24201_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41218_ ( .A(_24201_), .B(matmul_29_out_base_offset_och), .Y(matmul_29_out_base_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41219_ ( .A(matmul_29_arg_objaddr_0), .B(matmul_29_act_base_offset), .Y(_24202_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41220_ ( .A(_stream_matmul_29_source_6_source_offset_buf), .B(_source_stream_matmul_29_source_6_pat_cur_offset_0), .Y(_24203_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41221_ ( .A(_24203_), .B(_source_stream_matmul_29_source_6_pat_cur_offset_1), .Y(_24204_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41222_ ( .A(_24204_), .B(_source_stream_matmul_29_source_6_pat_cur_offset_2), .Y(_24205_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41223_ ( .A(_24205_), .B(_source_stream_matmul_29_source_6_pat_cur_offset_3), .Y(_stream_matmul_29_source_6_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41224_ ( .A(_stream_matmul_29_source_8_source_offset_buf), .B(_source_stream_matmul_29_source_8_pat_cur_offset_0), .Y(_24206_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41225_ ( .A(_24206_), .B(_source_stream_matmul_29_source_8_pat_cur_offset_1), .Y(_24207_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41226_ ( .A(_24207_), .B(_source_stream_matmul_29_source_8_pat_cur_offset_2), .Y(_24208_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41227_ ( .A(_24208_), .B(_source_stream_matmul_29_source_8_pat_cur_offset_3), .Y(_stream_matmul_29_source_8_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41228_ ( .A(_stream_matmul_29_source_19_source_offset_buf), .B(_source_stream_matmul_29_source_19_pat_cur_offset_0), .Y(_24209_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41229_ ( .A(_24209_), .B(_source_stream_matmul_29_source_19_pat_cur_offset_1), .Y(_24210_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41230_ ( .A(_24210_), .B(_source_stream_matmul_29_source_19_pat_cur_offset_2), .Y(_24211_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41231_ ( .A(_24211_), .B(_source_stream_matmul_29_source_19_pat_cur_offset_3), .Y(_stream_matmul_29_source_19_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41232_ ( .A(_stream_matmul_29_source_20_source_offset_buf), .B(_source_stream_matmul_29_source_20_pat_cur_offset_0), .Y(_24212_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41233_ ( .A(_24212_), .B(_source_stream_matmul_29_source_20_pat_cur_offset_1), .Y(_24213_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41234_ ( .A(_24213_), .B(_source_stream_matmul_29_source_20_pat_cur_offset_2), .Y(_24214_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41235_ ( .A(_24214_), .B(_source_stream_matmul_29_source_20_pat_cur_offset_3), .Y(_stream_matmul_29_source_20_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _41236_ ( .A({ 28'h0000000, cparam_conv2d_16_bias_num[6:2] }), .B({ 1'h0, _29100_ }), .Y(_24215_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41237_ ( .A(conv2d_16_arg_objaddr_1), .B(conv2d_16_filter_base_offset), .Y(_24216_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _41238_ ( .A({ 21'h000000, cparam_conv2d_16_filter_read_size[14:3] }), .B({ 1'h0, _29101_ }), .Y(_24217_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _41239_ ( .A({ 26'h0000000, cparam_conv2d_16_act_offset_values_2[8:2] }), .B({ 1'h0, _29102_ }), .Y(_24218_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41240_ ( .A(conv2d_16_out_laddr_offset), .B(conv2d_16_out_page_dma_offset), .Y(_24219_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41241_ ( .A(conv2d_16_objaddr), .B(conv2d_16_out_base_offset), .Y(_24220_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _41242_ ( .A({ 3'h0, conv2d_16_next_out_write_size[31:2] }), .B({ 1'h0, _29103_ }), .Y(_24221_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41243_ ( .A(max_pool_serial_18_arg_objaddr_0), .B(max_pool_serial_18_act_base_offset), .Y(_24222_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(10), .Y_WIDTH(32) ) _41244_ ( .A(max_pool_serial_18_act_page_dma_offset), .B(10'h200), .Y(_24223_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41245_ ( .A(max_pool_serial_18_act_base_offset), .B(512), .Y(_24224_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41246_ ( .A(max_pool_serial_18_arg_objaddr_0), .B(_24224_), .Y(_24225_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41247_ ( .A(max_pool_serial_18_objaddr), .B(max_pool_serial_18_out_base_offset), .Y(_24226_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _41248_ ( .A({ 26'h0000000, cparam_matmul_29_bias_num[8:2] }), .B({ 1'h0, _29104_ }), .Y(_24227_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41249_ ( .A(matmul_29_arg_objaddr_1), .B(matmul_29_filter_base_offset), .Y(_24228_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _41250_ ( .A({ 23'h000000, cparam_matmul_29_filter_read_size[12:3] }), .B({ 1'h0, _29105_ }), .Y(_24229_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _41251_ ( .A({ 24'h000000, cparam_matmul_29_act_bat_step[10:2] }), .B({ 1'h0, _29106_ }), .Y(_24230_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41252_ ( .A(matmul_29_out_laddr_offset), .B(matmul_29_out_page_dma_offset), .Y(_24231_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41253_ ( .A(matmul_29_objaddr), .B(matmul_29_out_base_offset), .Y(_24232_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _41254_ ( .A({ 3'h0, matmul_29_next_out_write_size[31:2] }), .B({ 1'h0, _29107_ }), .Y(_24233_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41255_ ( .A(_tmp_68), .B(1), .Y(_24234_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41256_ ( .A(ram_w4_l8192_id0_0_1_addr), .B(_maxi_read_local_stride), .Y(_24235_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41257_ ( .A(_tmp_99), .B(1), .Y(_24236_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41258_ ( .A(ram_w4_l8192_id0_1_1_addr), .B(_maxi_read_local_stride), .Y(_24237_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41259_ ( .A(_tmp_130), .B(1), .Y(_24238_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41260_ ( .A(ram_w4_l8192_id0_2_1_addr), .B(_maxi_read_local_stride), .Y(_24239_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41261_ ( .A(_tmp_161), .B(1), .Y(_24240_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41262_ ( .A(ram_w4_l8192_id0_3_1_addr), .B(_maxi_read_local_stride), .Y(_24241_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41263_ ( .A(_tmp_192), .B(1), .Y(_24242_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41264_ ( .A(ram_w4_l8192_id0_4_1_addr), .B(_maxi_read_local_stride), .Y(_24243_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41265_ ( .A(_tmp_223), .B(1), .Y(_24244_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41266_ ( .A(ram_w4_l8192_id0_5_1_addr), .B(_maxi_read_local_stride), .Y(_24245_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41267_ ( .A(_tmp_254), .B(1), .Y(_24246_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41268_ ( .A(ram_w4_l8192_id0_6_1_addr), .B(_maxi_read_local_stride), .Y(_24247_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41269_ ( .A(_tmp_285), .B(1), .Y(_24248_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41270_ ( .A(ram_w4_l8192_id0_7_1_addr), .B(_maxi_read_local_stride), .Y(_24249_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41271_ ( .A(ram_w8_l2048_id0_0_1_addr), .B(_maxi_read_local_stride), .Y(_24250_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41272_ ( .A(ram_w8_l2048_id0_0_1_addr), .B(_maxi_write_local_stride), .Y(_24251_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41273_ ( .A(ram_w8_l2048_id0_1_1_addr), .B(_maxi_read_local_stride), .Y(_24252_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41274_ ( .A(ram_w8_l2048_id0_1_1_addr), .B(_maxi_write_local_stride), .Y(_24253_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41275_ ( .A(ram_w8_l2048_id0_2_1_addr), .B(_maxi_read_local_stride), .Y(_24254_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41276_ ( .A(ram_w8_l2048_id0_2_1_addr), .B(_maxi_write_local_stride), .Y(_24255_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41277_ ( .A(ram_w8_l2048_id0_3_1_addr), .B(_maxi_read_local_stride), .Y(_24256_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41278_ ( .A(ram_w8_l2048_id0_3_1_addr), .B(_maxi_write_local_stride), .Y(_24257_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41279_ ( .A(ram_w8_l2048_id1_0_1_addr), .B(_maxi_read_local_stride), .Y(_24258_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41280_ ( .A(ram_w8_l2048_id1_0_1_addr), .B(_maxi_write_local_stride), .Y(_24259_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41281_ ( .A(ram_w8_l2048_id1_1_1_addr), .B(_maxi_read_local_stride), .Y(_24260_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41282_ ( .A(ram_w8_l2048_id1_1_1_addr), .B(_maxi_write_local_stride), .Y(_24261_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41283_ ( .A(ram_w8_l2048_id1_2_1_addr), .B(_maxi_read_local_stride), .Y(_24262_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41284_ ( .A(ram_w8_l2048_id1_2_1_addr), .B(_maxi_write_local_stride), .Y(_24263_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41285_ ( .A(ram_w8_l2048_id1_3_1_addr), .B(_maxi_read_local_stride), .Y(_24264_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41286_ ( .A(ram_w8_l2048_id1_3_1_addr), .B(_maxi_write_local_stride), .Y(_24265_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41287_ ( .A(_tmp_303), .B(1), .Y(_24266_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41288_ ( .A(ram_w8_l2048_id2_0_1_addr), .B(_maxi_read_local_stride), .Y(_24267_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41289_ ( .A(_tmp_316), .B(1), .Y(_24268_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41290_ ( .A(ram_w8_l2048_id2_1_1_addr), .B(_maxi_read_local_stride), .Y(_24269_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41291_ ( .A(_tmp_329), .B(1), .Y(_24270_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41292_ ( .A(ram_w8_l2048_id2_2_1_addr), .B(_maxi_read_local_stride), .Y(_24271_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41293_ ( .A(_tmp_342), .B(1), .Y(_24272_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41294_ ( .A(ram_w8_l2048_id2_3_1_addr), .B(_maxi_read_local_stride), .Y(_24273_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41295_ ( .A(ram_w8_l2048_id3_0_1_addr), .B(_maxi_read_local_stride), .Y(_24274_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41296_ ( .A(ram_w8_l2048_id3_1_1_addr), .B(_maxi_read_local_stride), .Y(_24275_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41297_ ( .A(ram_w8_l2048_id3_2_1_addr), .B(_maxi_read_local_stride), .Y(_24276_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41298_ ( .A(ram_w8_l2048_id3_3_1_addr), .B(_maxi_read_local_stride), .Y(_24277_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41299_ ( .A(_tmp_360), .B(1), .Y(_24278_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41300_ ( .A(_tmp_373), .B(1), .Y(_24279_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41301_ ( .A(_tmp_386), .B(1), .Y(_24280_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41302_ ( .A(_tmp_399), .B(1), .Y(_24281_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41303_ ( .A(_tmp_417), .B(1), .Y(_24282_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41304_ ( .A(_tmp_430), .B(1), .Y(_24283_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41305_ ( .A(_tmp_443), .B(1), .Y(_24284_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41306_ ( .A(_tmp_456), .B(1), .Y(_24285_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41307_ ( .A(ram_w8_l2048_id11_0_1_addr), .B(_maxi_write_local_stride), .Y(_24286_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41308_ ( .A(ram_w8_l2048_id11_1_1_addr), .B(_maxi_write_local_stride), .Y(_24287_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41309_ ( .A(ram_w8_l2048_id11_2_1_addr), .B(_maxi_write_local_stride), .Y(_24288_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41310_ ( .A(ram_w8_l2048_id11_3_1_addr), .B(_maxi_write_local_stride), .Y(_24289_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41311_ ( .A(_reduceadd_data_17), .B(__variable_wdata_0), .Y(_24290_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _41312_ ( .A(_reduceadd_count_17), .B(1), .Y(_24291_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _41313_ ( .A(_pulse_count_19), .B(1), .Y(_24292_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41314_ ( .A(__delay_data_750), .B(_cond_data_13), .Y(_24293_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41315_ ( .A(__variable_wdata_24), .B(__variable_wdata_25), .Y(_24294_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41316_ ( .A(_24294_), .B(__variable_wdata_26), .Y(_24295_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41317_ ( .A(__variable_wdata_27), .B(__variable_wdata_28), .Y(_24296_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41318_ ( .A(_24296_), .B(__variable_wdata_29), .Y(_24297_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41319_ ( .A(__variable_wdata_30), .B(__variable_wdata_31), .Y(_24298_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41320_ ( .A(_24298_), .B(__variable_wdata_32), .Y(_24299_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41321_ ( .A(__plusn_data_34), .B(__plusn_data_35), .Y(_24300_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41322_ ( .A(_24300_), .B(__plusn_data_36), .Y(_24301_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41323_ ( .A(_reducemax_count_211), .B(1), .Y(_24302_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41324_ ( .A(_pulse_count_213), .B(1), .Y(_24303_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(8) ) _41325_ ( .A(_cond_data_249), .B(__delay_data_947), .Y(_24304_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(8) ) _41326_ ( .A(_cond_data_256), .B(__delay_data_1268), .Y(_24305_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(4), .Y_WIDTH(8) ) _41327_ ( .A(_cond_data_263), .B(__delay_data_1339), .Y(_24306_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(32) ) _41328_ ( .A(__substreamoutput_data_881), .B(__delay_data_1338), .Y(_24307_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41329_ ( .A(_source_stream_conv2d_16_source_6_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_6_pat_stride_buf_0), .Y(_24308_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41330_ ( .A(_source_stream_conv2d_16_source_6_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_6_pat_stride_buf_1), .Y(_24309_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41331_ ( .A(_source_stream_conv2d_16_source_6_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_6_pat_stride_buf_2), .Y(_24310_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41332_ ( .A(_source_stream_conv2d_16_source_6_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_6_pat_stride_buf_3), .Y(_24311_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41333_ ( .A(_source_stream_conv2d_16_source_8_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_8_pat_stride_buf_0), .Y(_24312_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41334_ ( .A(_source_stream_conv2d_16_source_8_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_8_pat_stride_buf_1), .Y(_24313_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41335_ ( .A(_source_stream_conv2d_16_source_8_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_8_pat_stride_buf_2), .Y(_24314_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41336_ ( .A(_source_stream_conv2d_16_source_8_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_8_pat_stride_buf_3), .Y(_24315_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41337_ ( .A(conv2d_16_stream_act_local_0), .B(conv2d_16_act_page_comp_offset_buf_0), .Y(_24316_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41338_ ( .A(_source_stream_conv2d_16_source_19_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_19_pat_stride_buf_0), .Y(_24317_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41339_ ( .A(_source_stream_conv2d_16_source_19_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_19_pat_stride_buf_1), .Y(_24318_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41340_ ( .A(_source_stream_conv2d_16_source_19_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_19_pat_stride_buf_2), .Y(_24319_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41341_ ( .A(_source_stream_conv2d_16_source_19_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_19_pat_stride_buf_3), .Y(_24320_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41342_ ( .A(conv2d_16_stream_act_local_1), .B(conv2d_16_act_page_comp_offset_buf_0), .Y(_24321_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41343_ ( .A(_source_stream_conv2d_16_source_20_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_20_pat_stride_buf_0), .Y(_24322_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41344_ ( .A(_source_stream_conv2d_16_source_20_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_20_pat_stride_buf_1), .Y(_24323_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41345_ ( .A(_source_stream_conv2d_16_source_20_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_20_pat_stride_buf_2), .Y(_24324_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41346_ ( .A(_source_stream_conv2d_16_source_20_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_20_pat_stride_buf_3), .Y(_24325_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41347_ ( .A(conv2d_16_stream_act_local_2), .B(conv2d_16_act_page_comp_offset_buf_0), .Y(_24326_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41348_ ( .A(_source_stream_conv2d_16_source_21_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_21_pat_stride_buf_0), .Y(_24327_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41349_ ( .A(_source_stream_conv2d_16_source_21_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_21_pat_stride_buf_1), .Y(_24328_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41350_ ( .A(_source_stream_conv2d_16_source_21_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_21_pat_stride_buf_2), .Y(_24329_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41351_ ( .A(_source_stream_conv2d_16_source_21_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_21_pat_stride_buf_3), .Y(_24330_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41352_ ( .A(conv2d_16_stream_act_local_3), .B(conv2d_16_act_page_comp_offset_buf_1), .Y(_24331_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41353_ ( .A(_source_stream_conv2d_16_source_22_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_22_pat_stride_buf_0), .Y(_24332_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41354_ ( .A(_source_stream_conv2d_16_source_22_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_22_pat_stride_buf_1), .Y(_24333_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41355_ ( .A(_source_stream_conv2d_16_source_22_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_22_pat_stride_buf_2), .Y(_24334_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41356_ ( .A(_source_stream_conv2d_16_source_22_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_22_pat_stride_buf_3), .Y(_24335_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41357_ ( .A(conv2d_16_stream_act_local_4), .B(conv2d_16_act_page_comp_offset_buf_1), .Y(_24336_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41358_ ( .A(_source_stream_conv2d_16_source_23_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_23_pat_stride_buf_0), .Y(_24337_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41359_ ( .A(_source_stream_conv2d_16_source_23_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_23_pat_stride_buf_1), .Y(_24338_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41360_ ( .A(_source_stream_conv2d_16_source_23_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_23_pat_stride_buf_2), .Y(_24339_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41361_ ( .A(_source_stream_conv2d_16_source_23_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_23_pat_stride_buf_3), .Y(_24340_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41362_ ( .A(conv2d_16_stream_act_local_5), .B(conv2d_16_act_page_comp_offset_buf_1), .Y(_24341_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41363_ ( .A(_source_stream_conv2d_16_source_24_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_24_pat_stride_buf_0), .Y(_24342_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41364_ ( .A(_source_stream_conv2d_16_source_24_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_24_pat_stride_buf_1), .Y(_24343_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41365_ ( .A(_source_stream_conv2d_16_source_24_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_24_pat_stride_buf_2), .Y(_24344_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41366_ ( .A(_source_stream_conv2d_16_source_24_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_24_pat_stride_buf_3), .Y(_24345_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41367_ ( .A(conv2d_16_stream_act_local_6), .B(conv2d_16_act_page_comp_offset_buf_2), .Y(_24346_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41368_ ( .A(_source_stream_conv2d_16_source_25_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_25_pat_stride_buf_0), .Y(_24347_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41369_ ( .A(_source_stream_conv2d_16_source_25_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_25_pat_stride_buf_1), .Y(_24348_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41370_ ( .A(_source_stream_conv2d_16_source_25_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_25_pat_stride_buf_2), .Y(_24349_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41371_ ( .A(_source_stream_conv2d_16_source_25_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_25_pat_stride_buf_3), .Y(_24350_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41372_ ( .A(conv2d_16_stream_act_local_7), .B(conv2d_16_act_page_comp_offset_buf_2), .Y(_24351_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41373_ ( .A(_source_stream_conv2d_16_source_26_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_26_pat_stride_buf_0), .Y(_24352_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41374_ ( .A(_source_stream_conv2d_16_source_26_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_26_pat_stride_buf_1), .Y(_24353_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41375_ ( .A(_source_stream_conv2d_16_source_26_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_26_pat_stride_buf_2), .Y(_24354_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41376_ ( .A(_source_stream_conv2d_16_source_26_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_26_pat_stride_buf_3), .Y(_24355_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41377_ ( .A(conv2d_16_stream_act_local_8), .B(conv2d_16_act_page_comp_offset_buf_2), .Y(_24356_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41378_ ( .A(_source_stream_conv2d_16_source_27_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_27_pat_stride_buf_0), .Y(_24357_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41379_ ( .A(_source_stream_conv2d_16_source_27_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_27_pat_stride_buf_1), .Y(_24358_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41380_ ( .A(_source_stream_conv2d_16_source_27_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_27_pat_stride_buf_2), .Y(_24359_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41381_ ( .A(_source_stream_conv2d_16_source_27_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_27_pat_stride_buf_3), .Y(_24360_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41382_ ( .A(_source_stream_conv2d_16_source_28_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_28_pat_stride_buf_0), .Y(_24361_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41383_ ( .A(_source_stream_conv2d_16_source_28_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_28_pat_stride_buf_1), .Y(_24362_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41384_ ( .A(_source_stream_conv2d_16_source_28_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_28_pat_stride_buf_2), .Y(_24363_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41385_ ( .A(_source_stream_conv2d_16_source_28_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_28_pat_stride_buf_3), .Y(_24364_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41386_ ( .A(_source_stream_conv2d_16_source_29_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_29_pat_stride_buf_0), .Y(_24365_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41387_ ( .A(_source_stream_conv2d_16_source_29_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_29_pat_stride_buf_1), .Y(_24366_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41388_ ( .A(_source_stream_conv2d_16_source_29_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_29_pat_stride_buf_2), .Y(_24367_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41389_ ( .A(_source_stream_conv2d_16_source_29_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_29_pat_stride_buf_3), .Y(_24368_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41390_ ( .A(_source_stream_conv2d_16_source_30_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_30_pat_stride_buf_0), .Y(_24369_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41391_ ( .A(_source_stream_conv2d_16_source_30_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_30_pat_stride_buf_1), .Y(_24370_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41392_ ( .A(_source_stream_conv2d_16_source_30_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_30_pat_stride_buf_2), .Y(_24371_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41393_ ( .A(_source_stream_conv2d_16_source_30_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_30_pat_stride_buf_3), .Y(_24372_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41394_ ( .A(_source_stream_conv2d_16_source_31_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_31_pat_stride_buf_0), .Y(_24373_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41395_ ( .A(_source_stream_conv2d_16_source_31_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_31_pat_stride_buf_1), .Y(_24374_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41396_ ( .A(_source_stream_conv2d_16_source_31_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_31_pat_stride_buf_2), .Y(_24375_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41397_ ( .A(_source_stream_conv2d_16_source_31_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_31_pat_stride_buf_3), .Y(_24376_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41398_ ( .A(_source_stream_conv2d_16_source_32_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_32_pat_stride_buf_0), .Y(_24377_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41399_ ( .A(_source_stream_conv2d_16_source_32_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_32_pat_stride_buf_1), .Y(_24378_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41400_ ( .A(_source_stream_conv2d_16_source_32_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_32_pat_stride_buf_2), .Y(_24379_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41401_ ( .A(_source_stream_conv2d_16_source_32_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_32_pat_stride_buf_3), .Y(_24380_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41402_ ( .A(_source_stream_conv2d_16_source_33_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_33_pat_stride_buf_0), .Y(_24381_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41403_ ( .A(_source_stream_conv2d_16_source_33_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_33_pat_stride_buf_1), .Y(_24382_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41404_ ( .A(_source_stream_conv2d_16_source_33_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_33_pat_stride_buf_2), .Y(_24383_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41405_ ( .A(_source_stream_conv2d_16_source_33_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_33_pat_stride_buf_3), .Y(_24384_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41406_ ( .A(_source_stream_conv2d_16_source_34_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_34_pat_stride_buf_0), .Y(_24385_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41407_ ( .A(_source_stream_conv2d_16_source_34_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_34_pat_stride_buf_1), .Y(_24386_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41408_ ( .A(_source_stream_conv2d_16_source_34_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_34_pat_stride_buf_2), .Y(_24387_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41409_ ( .A(_source_stream_conv2d_16_source_34_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_34_pat_stride_buf_3), .Y(_24388_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41410_ ( .A(_source_stream_conv2d_16_source_35_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_35_pat_stride_buf_0), .Y(_24389_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41411_ ( .A(_source_stream_conv2d_16_source_35_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_35_pat_stride_buf_1), .Y(_24390_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41412_ ( .A(_source_stream_conv2d_16_source_35_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_35_pat_stride_buf_2), .Y(_24391_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41413_ ( .A(_source_stream_conv2d_16_source_35_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_35_pat_stride_buf_3), .Y(_24392_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41414_ ( .A(_source_stream_conv2d_16_source_36_pat_cur_offset_0), .B(_source_stream_conv2d_16_source_36_pat_stride_buf_0), .Y(_24393_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41415_ ( .A(_source_stream_conv2d_16_source_36_pat_cur_offset_1), .B(_source_stream_conv2d_16_source_36_pat_stride_buf_1), .Y(_24394_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41416_ ( .A(_source_stream_conv2d_16_source_36_pat_cur_offset_2), .B(_source_stream_conv2d_16_source_36_pat_stride_buf_2), .Y(_24395_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41417_ ( .A(_source_stream_conv2d_16_source_36_pat_cur_offset_3), .B(_source_stream_conv2d_16_source_36_pat_stride_buf_3), .Y(_24396_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41418_ ( .A(conv2d_16_stream_out_local_col), .B(conv2d_16_out_page_comp_offset_buf), .Y(_24397_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41419_ ( .A(_stream_conv2d_16_sink_37_sink_waddr), .B(_stream_conv2d_16_sink_37_sink_stride_buf), .Y(_24398_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(32) ) _41420_ ( .A(_counter_count_782), .B(2'h1), .Y(_24399_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41421_ ( .A(max_pool_serial_18_stream_act_local), .B(max_pool_serial_18_act_page_comp_offset_buf), .Y(_24400_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41422_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_0), .B(_source_stream_max_pool_serial_18_source_1_pat_stride_buf_0), .Y(_24401_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41423_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_1), .B(_source_stream_max_pool_serial_18_source_1_pat_stride_buf_1), .Y(_24402_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41424_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_2), .B(_source_stream_max_pool_serial_18_source_1_pat_stride_buf_2), .Y(_24403_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41425_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_3), .B(_source_stream_max_pool_serial_18_source_1_pat_stride_buf_3), .Y(_24404_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41426_ ( .A(max_pool_serial_18_stream_out_local), .B(max_pool_serial_18_out_page_comp_offset_buf), .Y(_24405_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41427_ ( .A(_stream_max_pool_serial_18_sink_3_sink_waddr), .B(_stream_max_pool_serial_18_sink_3_sink_stride_buf), .Y(_24406_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(8) ) _41428_ ( .A(_cond_data_831), .B(__delay_data_1422), .Y(_24407_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(8) ) _41429_ ( .A(_cond_data_838), .B(__delay_data_1429), .Y(_24408_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(4), .Y_WIDTH(8) ) _41430_ ( .A(_cond_data_845), .B(__delay_data_1482), .Y(_24409_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(32) ) _41431_ ( .A(__substreamoutput_data_881), .B(__delay_data_1481), .Y(_24410_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41432_ ( .A(_source_stream_matmul_29_source_6_pat_cur_offset_0), .B(_source_stream_matmul_29_source_6_pat_stride_buf_0), .Y(_24411_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41433_ ( .A(_source_stream_matmul_29_source_6_pat_cur_offset_1), .B(_source_stream_matmul_29_source_6_pat_stride_buf_1), .Y(_24412_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41434_ ( .A(_source_stream_matmul_29_source_6_pat_cur_offset_2), .B(_source_stream_matmul_29_source_6_pat_stride_buf_2), .Y(_24413_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41435_ ( .A(_source_stream_matmul_29_source_6_pat_cur_offset_3), .B(_source_stream_matmul_29_source_6_pat_stride_buf_3), .Y(_24414_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41436_ ( .A(_source_stream_matmul_29_source_8_pat_cur_offset_0), .B(_source_stream_matmul_29_source_8_pat_stride_buf_0), .Y(_24415_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41437_ ( .A(_source_stream_matmul_29_source_8_pat_cur_offset_1), .B(_source_stream_matmul_29_source_8_pat_stride_buf_1), .Y(_24416_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41438_ ( .A(_source_stream_matmul_29_source_8_pat_cur_offset_2), .B(_source_stream_matmul_29_source_8_pat_stride_buf_2), .Y(_24417_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41439_ ( .A(_source_stream_matmul_29_source_8_pat_cur_offset_3), .B(_source_stream_matmul_29_source_8_pat_stride_buf_3), .Y(_24418_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41440_ ( .A(matmul_29_stream_act_local_0), .B(matmul_29_act_page_comp_offset_buf_0), .Y(_24419_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41441_ ( .A(_source_stream_matmul_29_source_19_pat_cur_offset_0), .B(_source_stream_matmul_29_source_19_pat_stride_buf_0), .Y(_24420_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41442_ ( .A(_source_stream_matmul_29_source_19_pat_cur_offset_1), .B(_source_stream_matmul_29_source_19_pat_stride_buf_1), .Y(_24421_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41443_ ( .A(_source_stream_matmul_29_source_19_pat_cur_offset_2), .B(_source_stream_matmul_29_source_19_pat_stride_buf_2), .Y(_24422_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41444_ ( .A(_source_stream_matmul_29_source_19_pat_cur_offset_3), .B(_source_stream_matmul_29_source_19_pat_stride_buf_3), .Y(_24423_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41445_ ( .A(_source_stream_matmul_29_source_20_pat_cur_offset_0), .B(_source_stream_matmul_29_source_20_pat_stride_buf_0), .Y(_24424_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41446_ ( .A(_source_stream_matmul_29_source_20_pat_cur_offset_1), .B(_source_stream_matmul_29_source_20_pat_stride_buf_1), .Y(_24425_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41447_ ( .A(_source_stream_matmul_29_source_20_pat_cur_offset_2), .B(_source_stream_matmul_29_source_20_pat_stride_buf_2), .Y(_24426_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41448_ ( .A(_source_stream_matmul_29_source_20_pat_cur_offset_3), .B(_source_stream_matmul_29_source_20_pat_stride_buf_3), .Y(_24427_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41449_ ( .A(matmul_29_stream_out_local_col), .B(matmul_29_out_page_comp_offset_buf), .Y(_24428_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41450_ ( .A(_stream_matmul_29_sink_21_sink_waddr), .B(_stream_matmul_29_sink_21_sink_stride_buf), .Y(_24429_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41451_ ( .A(_saxi_register_13), .B(576), .Y({ _04000_, _03999_, _03997_, _03996_, _03995_, _03994_, _03993_, _03992_, _03991_, _03990_, _03989_, _03988_, _03986_, _03985_, _03984_, _03983_, _03982_, _03981_, _03980_, _03979_, _03978_, _03977_, _04007_, _04006_, _04005_, _04004_, _04003_, _04002_, _04001_, _03998_, _03987_, _03976_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41452_ ( .A(_saxi_register_13), .B(640), .Y({ _04032_, _04031_, _04029_, _04028_, _04027_, _04026_, _04025_, _04024_, _04023_, _04022_, _04021_, _04020_, _04018_, _04017_, _04016_, _04015_, _04014_, _04013_, _04012_, _04011_, _04010_, _04009_, _04039_, _04038_, _04037_, _04036_, _04035_, _04034_, _04033_, _04030_, _04019_, _04008_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41453_ ( .A(_saxi_register_10), .B(16384), .Y({ _04064_, _04063_, _04061_, _04060_, _04059_, _04058_, _04057_, _04056_, _04055_, _04054_, _04053_, _04052_, _04050_, _04049_, _04048_, _04047_, _04046_, _04045_, _04044_, _04043_, _04042_, _04041_, _04071_, _04070_, _04069_, _04068_, _04067_, _04066_, _04065_, _04062_, _04051_, _04040_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41454_ ( .A(_saxi_register_13), .B(704), .Y({ _04128_, _04127_, _04125_, _04124_, _04123_, _04122_, _04121_, _04120_, _04119_, _04118_, _04117_, _04116_, _04114_, _04113_, _04112_, _04111_, _04110_, _04109_, _04108_, _04107_, _04106_, _04105_, _04135_, _04134_, _04133_, _04132_, _04131_, _04130_, _04129_, _04126_, _04115_, _04104_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41455_ ( .A(_saxi_register_13), .B(3008), .Y({ _04160_, _04159_, _04157_, _04156_, _04155_, _04154_, _04153_, _04152_, _04151_, _04150_, _04149_, _04148_, _04146_, _04145_, _04144_, _04143_, _04142_, _04141_, _04140_, _04139_, _04138_, _04137_, _04167_, _04166_, _04165_, _04164_, _04163_, _04162_, _04161_, _04158_, _04147_, _04136_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41456_ ( .A(_saxi_register_13), .B(3072), .Y({ _04192_, _04191_, _04189_, _04188_, _04187_, _04186_, _04185_, _04184_, _04183_, _04182_, _04181_, _04180_, _04178_, _04177_, _04176_, _04175_, _04174_, _04173_, _04172_, _04171_, _04170_, _04169_, _04199_, _04198_, _04197_, _04196_, _04195_, _04194_, _04193_, _04190_, _04179_, _04168_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41457_ ( .A(_saxi_register_10), .B(20480), .Y({ _04096_, _04095_, _04093_, _04092_, _04091_, _04090_, _04089_, _04088_, _04087_, _04086_, _04085_, _04084_, _04082_, _04081_, _04080_, _04079_, _04078_, _04077_, _04076_, _04075_, _04074_, _04073_, _04103_, _04102_, _04101_, _04100_, _04099_, _04098_, _04097_, _04094_, _04083_, _04072_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41458_ ( .A(_saxi_register_10), .B(28672), .Y({ _04224_, _04223_, _04221_, _04220_, _04219_, _04218_, _04217_, _04216_, _04215_, _04214_, _04213_, _04212_, _04210_, _04209_, _04208_, _04207_, _04206_, _04205_, _04204_, _04203_, _04202_, _04201_, _04231_, _04230_, _04229_, _04228_, _04227_, _04226_, _04225_, _04222_, _04211_, _04200_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41459_ ( .A(_saxi_register_13), .B(3136), .Y({ _04288_, _04287_, _04285_, _04284_, _04283_, _04282_, _04281_, _04280_, _04279_, _04278_, _04277_, _04276_, _04274_, _04273_, _04272_, _04271_, _04270_, _04269_, _04268_, _04267_, _04266_, _04265_, _04295_, _04294_, _04293_, _04292_, _04291_, _04290_, _04289_, _04286_, _04275_, _04264_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41460_ ( .A(_saxi_register_13), .B(12352), .Y({ _04320_, _04319_, _04317_, _04316_, _04315_, _04314_, _04313_, _04312_, _04311_, _04310_, _04309_, _04308_, _04306_, _04305_, _04304_, _04303_, _04302_, _04301_, _04300_, _04299_, _04298_, _04297_, _04327_, _04326_, _04325_, _04324_, _04323_, _04322_, _04321_, _04318_, _04307_, _04296_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41461_ ( .A(_saxi_register_13), .B(12416), .Y({ _04352_, _04351_, _04349_, _04348_, _04347_, _04346_, _04345_, _04344_, _04343_, _04342_, _04341_, _04340_, _04338_, _04337_, _04336_, _04335_, _04334_, _04333_, _04332_, _04331_, _04330_, _04329_, _04359_, _04358_, _04357_, _04356_, _04355_, _04354_, _04353_, _04350_, _04339_, _04328_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41462_ ( .A(_saxi_register_10), .B(30720), .Y({ _04256_, _04255_, _04253_, _04252_, _04251_, _04250_, _04249_, _04248_, _04247_, _04246_, _04245_, _04244_, _04242_, _04241_, _04240_, _04239_, _04238_, _04237_, _04236_, _04235_, _04234_, _04233_, _04263_, _04262_, _04261_, _04260_, _04259_, _04258_, _04257_, _04254_, _04243_, _04232_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41463_ ( .A(_saxi_register_10), .B(34816), .Y({ _04384_, _04383_, _04381_, _04380_, _04379_, _04378_, _04377_, _04376_, _04375_, _04374_, _04373_, _04372_, _04370_, _04369_, _04368_, _04367_, _04366_, _04365_, _04364_, _04363_, _04362_, _04361_, _04391_, _04390_, _04389_, _04388_, _04387_, _04386_, _04385_, _04382_, _04371_, _04360_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41464_ ( .A(_saxi_register_13), .B(12480), .Y({ _04448_, _04447_, _04445_, _04444_, _04443_, _04442_, _04441_, _04440_, _04439_, _04438_, _04437_, _04436_, _04434_, _04433_, _04432_, _04431_, _04430_, _04429_, _04428_, _04427_, _04426_, _04425_, _04455_, _04454_, _04453_, _04452_, _04451_, _04450_, _04449_, _04446_, _04435_, _04424_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41465_ ( .A(_saxi_register_13), .B(143552), .Y({ _04480_, _04479_, _04477_, _04476_, _04475_, _04474_, _04473_, _04472_, _04471_, _04470_, _04469_, _04468_, _04466_, _04465_, _04464_, _04463_, _04462_, _04461_, _04460_, _04459_, _04458_, _04457_, _04487_, _04486_, _04485_, _04484_, _04483_, _04482_, _04481_, _04478_, _04467_, _04456_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41466_ ( .A(_saxi_register_13), .B(143808), .Y({ _04512_, _04511_, _04509_, _04508_, _04507_, _04506_, _04505_, _04504_, _04503_, _04502_, _04501_, _04500_, _04498_, _04497_, _04496_, _04495_, _04494_, _04493_, _04492_, _04491_, _04490_, _04489_, _04519_, _04518_, _04517_, _04516_, _04515_, _04514_, _04513_, _04510_, _04499_, _04488_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41467_ ( .A(_saxi_register_10), .B(35840), .Y({ _04416_, _04415_, _04413_, _04412_, _04411_, _04410_, _04409_, _04408_, _04407_, _04406_, _04405_, _04404_, _04402_, _04401_, _04400_, _04399_, _04398_, _04397_, _04396_, _04395_, _04394_, _04393_, _04423_, _04422_, _04421_, _04420_, _04419_, _04418_, _04417_, _04414_, _04403_, _04392_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41468_ ( .A(_saxi_register_13), .B(143872), .Y({ _04576_, _04575_, _04573_, _04572_, _04571_, _04570_, _04569_, _04568_, _04567_, _04566_, _04565_, _04564_, _04562_, _04561_, _04560_, _04559_, _04558_, _04557_, _04556_, _04555_, _04554_, _04553_, _04583_, _04582_, _04581_, _04580_, _04579_, _04578_, _04577_, _04574_, _04563_, _04552_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41469_ ( .A(_saxi_register_13), .B(160256), .Y({ _04608_, _04607_, _04605_, _04604_, _04603_, _04602_, _04601_, _04600_, _04599_, _04598_, _04597_, _04596_, _04594_, _04593_, _04592_, _04591_, _04590_, _04589_, _04588_, _04587_, _04586_, _04585_, _04615_, _04614_, _04613_, _04612_, _04611_, _04610_, _04609_, _04606_, _04595_, _04584_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41470_ ( .A(_saxi_register_13), .B(160384), .Y({ _04640_, _04639_, _04637_, _04636_, _04635_, _04634_, _04633_, _04632_, _04631_, _04630_, _04629_, _04628_, _04626_, _04625_, _04624_, _04623_, _04622_, _04621_, _04620_, _04619_, _04618_, _04617_, _04647_, _04646_, _04645_, _04644_, _04643_, _04642_, _04641_, _04638_, _04627_, _04616_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41471_ ( .A(_saxi_register_10), .B(36096), .Y({ _04544_, _04543_, _04541_, _04540_, _04539_, _04538_, _04537_, _04536_, _04535_, _04534_, _04533_, _04532_, _04530_, _04529_, _04528_, _04527_, _04526_, _04525_, _04524_, _04523_, _04522_, _04521_, _04551_, _04550_, _04549_, _04548_, _04547_, _04546_, _04545_, _04542_, _04531_, _04520_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41472_ ( .A(_saxi_register_13), .B(160448), .Y({ _04672_, _04671_, _04669_, _04668_, _04667_, _04666_, _04665_, _04664_, _04663_, _04662_, _04661_, _04660_, _04658_, _04657_, _04656_, _04655_, _04654_, _04653_, _04652_, _04651_, _04650_, _04649_, _04679_, _04678_, _04677_, _04676_, _04675_, _04674_, _04673_, _04670_, _04659_, _04648_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41473_ ( .A(_saxi_register_13), .B(161088), .Y({ _04704_, _04703_, _04701_, _04700_, _04699_, _04698_, _04697_, _04696_, _04695_, _04694_, _04693_, _04692_, _04690_, _04689_, _04688_, _04687_, _04686_, _04685_, _04684_, _04683_, _04682_, _04681_, _04711_, _04710_, _04709_, _04708_, _04707_, _04706_, _04705_, _04702_, _04691_, _04680_ }) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41474_ ( .A(_saxi_register_13), .B(161152), .Y({ _04736_, _04735_, _04733_, _04732_, _04731_, _04730_, _04729_, _04728_, _04727_, _04726_, _04725_, _04724_, _04722_, _04721_, _04720_, _04719_, _04718_, _04717_, _04716_, _04715_, _04714_, _04713_, _04743_, _04742_, _04741_, _04740_, _04739_, _04738_, _04737_, _04734_, _04723_, _04712_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41475_ ( .A(conv2d_16_out_laddr_offset), .B(conv2d_16_next_out_write_size), .Y(_24430_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41476_ ( .A(conv2d_16_out_ram_select), .B(1), .Y(_24431_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(6), .Y_WIDTH(32) ) _41477_ ( .A(conv2d_16_sync_out_count), .B(cparam_conv2d_16_act_num_row), .Y({ _04768_, _04767_, _04765_, _04764_, _04763_, _04762_, _04761_, _04760_, _04759_, _04758_, _04757_, _04756_, _04754_, _04753_, _04752_, _04751_, _04750_, _04749_, _04748_, _04747_, _04746_, _04745_, _04775_, _04774_, _04773_, _04772_, _04771_, _04770_, _04769_, _04766_, _04755_, _04744_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41478_ ( .A(conv2d_16_sync_out_count), .B({ 26'h0000000, cparam_conv2d_16_act_num_row }), .Y({ _04800_, _04799_, _04797_, _04796_, _04795_, _04794_, _04793_, _04792_, _04791_, _04790_, _04789_, _04788_, _04786_, _04785_, _04784_, _04783_, _04782_, _04781_, _04780_, _04779_, _04778_, _04777_, _04807_, _04806_, _04805_, _04804_, _04803_, _04802_, _04801_, _04798_, _04787_, _04776_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(14), .Y_WIDTH(32) ) _41479_ ( .A(conv2d_16_filter_base_offset), .B(cparam_conv2d_16_filter_base_step), .Y(_24432_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(8), .Y_WIDTH(32) ) _41480_ ( .A(conv2d_16_och_count), .B(cparam_conv2d_16_och_count_step), .Y(_24433_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(12), .Y_WIDTH(32) ) _41481_ ( .A(conv2d_16_filter_page_dma_offset), .B(cparam_conv2d_16_filter_read_step), .Y(_24435_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(12), .Y_WIDTH(32) ) _41482_ ( .A(conv2d_16_filter_page_comp_offset), .B(cparam_conv2d_16_filter_read_step), .Y(_24434_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(12), .Y_WIDTH(32) ) _41483_ ( .A(_24434_), .B(cparam_conv2d_16_filter_read_step), .Y({ _04832_, _04831_, _04829_, _04828_, _04827_, _04826_, _04825_, _04824_, _04823_, _04822_, _04821_, _04820_, _04818_, _04817_, _04816_, _04815_, _04814_, _04813_, _04812_, _04811_, _04810_, _04809_, _04839_, _04838_, _04837_, _04836_, _04835_, _04834_, _04833_, _04830_, _04819_, _04808_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(9), .Y_WIDTH(32) ) _41484_ ( .A(conv2d_16_act_base_offset_row), .B(cparam_conv2d_16_act_offset_values_2[8:0]), .Y(_24436_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(32) ) _41485_ ( .A(conv2d_16_row_count), .B(1'h1), .Y(_24437_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(2) ) _41486_ ( .A(conv2d_16_row_select), .B(1'h1), .Y(_24438_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(32) ) _41487_ ( .A(conv2d_16_row_select), .B(1'h1), .Y({ _04864_, _04863_, _04861_, _04860_, _04859_, _04858_, _04857_, _04856_, _04855_, _04854_, _04853_, _04852_, _04850_, _04849_, _04848_, _04847_, _04846_, _04845_, _04844_, _04843_, _04842_, _04841_, _04871_, _04870_, _04869_, _04868_, _04867_, _04866_, _04865_, _04862_, _04851_, _04840_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _41488_ ( .A(conv2d_16_act_page_dma_offset_0), .B(cparam_conv2d_16_act_read_step), .Y(_24440_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _41489_ ( .A(conv2d_16_act_page_comp_offset_0), .B(cparam_conv2d_16_act_read_step), .Y(_24439_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _41490_ ( .A(_24439_), .B(cparam_conv2d_16_act_read_step), .Y({ _04896_, _04895_, _04893_, _04892_, _04891_, _04890_, _04889_, _04888_, _04887_, _04886_, _04885_, _04884_, _04882_, _04881_, _04880_, _04879_, _04878_, _04877_, _04876_, _04875_, _04874_, _04873_, _04903_, _04902_, _04901_, _04900_, _04899_, _04898_, _04897_, _04894_, _04883_, _04872_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _41491_ ( .A(conv2d_16_act_page_dma_offset_1), .B(cparam_conv2d_16_act_read_step), .Y(_24442_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _41492_ ( .A(conv2d_16_act_page_comp_offset_1), .B(cparam_conv2d_16_act_read_step), .Y(_24441_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _41493_ ( .A(_24441_), .B(cparam_conv2d_16_act_read_step), .Y({ _04928_, _04927_, _04925_, _04924_, _04923_, _04922_, _04921_, _04920_, _04919_, _04918_, _04917_, _04916_, _04914_, _04913_, _04912_, _04911_, _04910_, _04909_, _04908_, _04907_, _04906_, _04905_, _04935_, _04934_, _04933_, _04932_, _04931_, _04930_, _04929_, _04926_, _04915_, _04904_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _41494_ ( .A(conv2d_16_act_page_dma_offset_2), .B(cparam_conv2d_16_act_read_step), .Y(_24444_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _41495_ ( .A(conv2d_16_act_page_comp_offset_2), .B(cparam_conv2d_16_act_read_step), .Y(_24443_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _41496_ ( .A(_24443_), .B(cparam_conv2d_16_act_read_step), .Y({ _04960_, _04959_, _04957_, _04956_, _04955_, _04954_, _04953_, _04952_, _04951_, _04950_, _04949_, _04948_, _04946_, _04945_, _04944_, _04943_, _04942_, _04941_, _04940_, _04939_, _04938_, _04937_, _04967_, _04966_, _04965_, _04964_, _04963_, _04962_, _04961_, _04958_, _04947_, _04936_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41497_ ( .A(conv2d_16_out_row_count), .B(1), .Y(_24446_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _41498_ ( .A(conv2d_16_out_base_offset_och), .B(cparam_conv2d_16_bias_num), .Y(_24447_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(10), .Y_WIDTH(32) ) _41499_ ( .A(conv2d_16_out_base_offset_row), .B(10'h200), .Y(_24445_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41500_ ( .A(_maxi_read_global_addr), .B(_maxi_global_base_addr), .Y(_24448_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _41501_ ( .A({ 21'h000000, _maxi_read_cur_global_addr[11:0] }), .B({ _maxi_read_rest_size[30:0], 2'h0 }), .Y({ _04993_, _04992_, _04991_, _04989_, _04988_, _04987_, _04986_, _04985_, _04984_, _04983_, _04982_, _04981_, _04980_, _04978_, _04977_, _04976_, _04975_, _04974_, _04973_, _04972_, _04971_, _04970_, _04969_, _05000_, _04999_, _04998_, _04997_, _04996_, _04995_, _04994_, _04990_, _04979_, _04968_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41502_ ( .A({ 20'h00000, _maxi_read_cur_global_addr[11:0] }), .B(1024), .Y({ _05025_, _05024_, _05022_, _05021_, _05020_, _05019_, _05018_, _05017_, _05016_, _05015_, _05014_, _05013_, _05011_, _05010_, _05009_, _05008_, _05007_, _05006_, _05005_, _05004_, _05003_, _05002_, _05032_, _05031_, _05030_, _05029_, _05028_, _05027_, _05026_, _05023_, _05012_, _05001_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _41503_ ( .A(_maxi_read_cur_global_addr), .B({ _maxi_read_cur_size[30:0], 2'h0 }), .Y(_24449_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41504_ ( .A(conv2d_16_sync_comp_count), .B(1), .Y(_24450_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(6), .Y_WIDTH(32) ) _41505_ ( .A(conv2d_16_stream_act_local_0), .B(cparam_conv2d_16_inc_act_laddr_large), .Y(_24451_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(6), .Y_WIDTH(32) ) _41506_ ( .A(conv2d_16_stream_act_local_1), .B(cparam_conv2d_16_inc_act_laddr_large), .Y(_24452_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(6), .Y_WIDTH(32) ) _41507_ ( .A(conv2d_16_stream_act_local_2), .B(cparam_conv2d_16_inc_act_laddr_large), .Y(_24453_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(6), .Y_WIDTH(32) ) _41508_ ( .A(conv2d_16_stream_act_local_3), .B(cparam_conv2d_16_inc_act_laddr_large), .Y(_24454_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(6), .Y_WIDTH(32) ) _41509_ ( .A(conv2d_16_stream_act_local_4), .B(cparam_conv2d_16_inc_act_laddr_large), .Y(_24455_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(6), .Y_WIDTH(32) ) _41510_ ( .A(conv2d_16_stream_act_local_5), .B(cparam_conv2d_16_inc_act_laddr_large), .Y(_24456_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(6), .Y_WIDTH(32) ) _41511_ ( .A(conv2d_16_stream_act_local_6), .B(cparam_conv2d_16_inc_act_laddr_large), .Y(_24457_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(6), .Y_WIDTH(32) ) _41512_ ( .A(conv2d_16_stream_act_local_7), .B(cparam_conv2d_16_inc_act_laddr_large), .Y(_24458_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(6), .Y_WIDTH(32) ) _41513_ ( .A(conv2d_16_stream_act_local_8), .B(cparam_conv2d_16_inc_act_laddr_large), .Y(_24459_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41514_ ( .A(conv2d_16_stream_out_local_col), .B(conv2d_16_next_stream_num_ops), .Y(_24460_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(32) ) _41515_ ( .A(conv2d_16_col_count), .B(1'h1), .Y(_24461_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(2) ) _41516_ ( .A(conv2d_16_col_select), .B(1'h1), .Y(_24462_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(32) ) _41517_ ( .A(conv2d_16_col_select), .B(1'h1), .Y({ _05057_, _05056_, _05054_, _05053_, _05052_, _05051_, _05050_, _05049_, _05048_, _05047_, _05046_, _05045_, _05043_, _05042_, _05041_, _05040_, _05039_, _05038_, _05037_, _05036_, _05035_, _05034_, _05064_, _05063_, _05062_, _05061_, _05060_, _05059_, _05058_, _05055_, _05044_, _05033_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41518_ ( .A(_maxi_write_global_addr), .B(_maxi_global_base_addr), .Y(_24463_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _41519_ ( .A({ 21'h000000, _maxi_write_cur_global_addr[11:0] }), .B({ _maxi_write_rest_size[30:0], 2'h0 }), .Y({ _05090_, _05089_, _05088_, _05086_, _05085_, _05084_, _05083_, _05082_, _05081_, _05080_, _05079_, _05078_, _05077_, _05075_, _05074_, _05073_, _05072_, _05071_, _05070_, _05069_, _05068_, _05067_, _05066_, _05097_, _05096_, _05095_, _05094_, _05093_, _05092_, _05091_, _05087_, _05076_, _05065_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41520_ ( .A({ 20'h00000, _maxi_write_cur_global_addr[11:0] }), .B(1024), .Y({ _05122_, _05121_, _05119_, _05118_, _05117_, _05116_, _05115_, _05114_, _05113_, _05112_, _05111_, _05110_, _05108_, _05107_, _05106_, _05105_, _05104_, _05103_, _05102_, _05101_, _05100_, _05099_, _05129_, _05128_, _05127_, _05126_, _05125_, _05124_, _05123_, _05120_, _05109_, _05098_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _41521_ ( .A(_maxi_write_cur_global_addr), .B({ _maxi_write_cur_size[30:0], 2'h0 }), .Y(_24464_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(9), .Y_WIDTH(32) ) _41522_ ( .A(max_pool_serial_18_out_count), .B(9'h100), .Y({ _05154_, _05153_, _05151_, _05150_, _05149_, _05148_, _05147_, _05146_, _05145_, _05144_, _05143_, _05142_, _05140_, _05139_, _05138_, _05137_, _05136_, _05135_, _05134_, _05133_, _05132_, _05131_, _05161_, _05160_, _05159_, _05158_, _05157_, _05156_, _05155_, _05152_, _05141_, _05130_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(11), .Y_WIDTH(32) ) _41523_ ( .A(max_pool_serial_18_act_base_offset_row), .B(11'h400), .Y(_24465_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(32) ) _41524_ ( .A(max_pool_serial_18_row_count), .B(2'h2), .Y(_24466_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(9), .Y_WIDTH(32) ) _41525_ ( .A(max_pool_serial_18_out_base_offset_row), .B(9'h100), .Y(_24467_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _41526_ ( .A(max_pool_serial_18_comp_count), .B(cparam_max_pool_serial_18_inc_out_laddr), .Y(_24468_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(8), .Y_WIDTH(32) ) _41527_ ( .A(max_pool_serial_18_stream_act_local), .B(cparam_max_pool_serial_18_inc_act_laddr), .Y(_24469_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(7), .Y_WIDTH(32) ) _41528_ ( .A(max_pool_serial_18_stream_out_local), .B(cparam_max_pool_serial_18_inc_out_laddr), .Y(_24470_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(32) ) _41529_ ( .A(max_pool_serial_18_col_count), .B(2'h2), .Y(_24471_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41530_ ( .A(matmul_29_out_laddr_offset), .B(matmul_29_next_out_write_size), .Y(_24472_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(9), .Y_WIDTH(32) ) _41531_ ( .A(matmul_29_out_base_offset_col), .B(cparam_matmul_29_out_bat_step), .Y(_24473_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41532_ ( .A(matmul_29_out_ram_select), .B(1), .Y(_24474_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(32) ) _41533_ ( .A(matmul_29_sync_out_count), .B(1'h1), .Y({ _05186_, _05185_, _05183_, _05182_, _05181_, _05180_, _05179_, _05178_, _05177_, _05176_, _05175_, _05174_, _05172_, _05171_, _05170_, _05169_, _05168_, _05167_, _05166_, _05165_, _05164_, _05163_, _05193_, _05192_, _05191_, _05190_, _05189_, _05188_, _05187_, _05184_, _05173_, _05162_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41534_ ( .A(matmul_29_sync_out_count), .B(1), .Y({ _14362_, _14361_, _14359_, _14358_, _14357_, _14356_, _14355_, _14354_, _14353_, _14352_, _14351_, _14350_, _14348_, _14347_, _14346_, _14345_, _14344_, _14343_, _14342_, _14341_, _14340_, _14339_, _14369_, _14368_, _14367_, _14366_, _14365_, _14364_, _14363_, _14360_, _14349_, _14338_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(12), .Y_WIDTH(32) ) _41535_ ( .A(matmul_29_filter_base_offset), .B(cparam_matmul_29_filter_base_step), .Y({ _05218_, _05217_, _05215_, _05214_, _05213_, _05212_, _05211_, _05210_, _05209_, _05208_, _05207_, _05206_, _05204_, _05203_, _05202_, _05201_, _05200_, _05199_, _05198_, _05197_, _05196_, _05195_, _05225_, _05224_, _05223_, _05222_, _05221_, _05220_, _05219_, _05216_, _05205_, _05194_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(6), .Y_WIDTH(32) ) _41536_ ( .A(matmul_29_och_count), .B(cparam_matmul_29_och_count_step), .Y({ _05250_, _05249_, _05247_, _05246_, _05245_, _05244_, _05243_, _05242_, _05241_, _05240_, _05239_, _05238_, _05236_, _05235_, _05234_, _05233_, _05232_, _05231_, _05230_, _05229_, _05228_, _05227_, _05257_, _05256_, _05255_, _05254_, _05253_, _05252_, _05251_, _05248_, _05237_, _05226_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(13), .Y_WIDTH(32) ) _41537_ ( .A(matmul_29_filter_page_dma_offset), .B(cparam_matmul_29_filter_read_size), .Y(_24476_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(13), .Y_WIDTH(32) ) _41538_ ( .A(matmul_29_filter_page_comp_offset), .B(cparam_matmul_29_filter_read_size), .Y(_24475_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(13), .Y_WIDTH(32) ) _41539_ ( .A(_24475_), .B(cparam_matmul_29_filter_read_size), .Y({ _05282_, _05281_, _05279_, _05278_, _05277_, _05276_, _05275_, _05274_, _05273_, _05272_, _05271_, _05270_, _05268_, _05267_, _05266_, _05265_, _05264_, _05263_, _05262_, _05261_, _05260_, _05259_, _05289_, _05288_, _05287_, _05286_, _05285_, _05284_, _05283_, _05280_, _05269_, _05258_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(5), .Y_WIDTH(32) ) _41540_ ( .A(matmul_29_out_base_offset_och), .B(cparam_matmul_29_out_och_step), .Y(_24477_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41541_ ( .A(matmul_29_sync_comp_count), .B(1), .Y(_24478_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41542_ ( .A(conv2d_16_act_base_offset_row), .B(conv2d_16_act_base_offset_bat), .Y(conv2d_16_act_base_offset) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41543_ ( .A(conv2d_16_out_base_offset_val), .B(conv2d_16_out_base_offset_col), .Y(_24479_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41544_ ( .A(_24479_), .B(conv2d_16_out_base_offset_row), .Y(_24480_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41545_ ( .A(_24480_), .B(conv2d_16_out_base_offset_bat), .Y(_24481_) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(32), .Y_WIDTH(32) ) _41546_ ( .A(_24481_), .B(conv2d_16_out_base_offset_och), .Y(conv2d_16_out_base_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41547_ ( .A(_tmp_41), .B(_maxi_read_local_stride), .Y({ _24482_[31:10], _tmp_50 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41548_ ( .A(_tmp_42), .B(_maxi_read_local_stride), .Y({ _24483_[31:10], _tmp_51 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41549_ ( .A(_tmp_43), .B(_maxi_read_local_stride), .Y({ _24484_[31:10], _tmp_52 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41550_ ( .A(_tmp_44), .B(_maxi_read_local_stride), .Y({ _24485_[31:10], _tmp_53 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41551_ ( .A(_tmp_45), .B(_maxi_read_local_stride), .Y({ _24486_[31:10], _tmp_54 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41552_ ( .A(_tmp_46), .B(_maxi_read_local_stride), .Y({ _24487_[31:10], _tmp_55 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41553_ ( .A(_tmp_47), .B(_maxi_read_local_stride), .Y({ _24488_[31:10], _tmp_56 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41554_ ( .A(_tmp_48), .B(_maxi_read_local_stride), .Y({ _24489_[31:10], _tmp_57 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41555_ ( .A(_tmp_49), .B(_maxi_read_local_stride), .Y({ _24490_[31:10], _tmp_58 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41556_ ( .A(_tmp_72), .B(_maxi_read_local_stride), .Y({ _24491_[31:10], _tmp_81 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41557_ ( .A(_tmp_73), .B(_maxi_read_local_stride), .Y({ _24492_[31:10], _tmp_82 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41558_ ( .A(_tmp_74), .B(_maxi_read_local_stride), .Y({ _24493_[31:10], _tmp_83 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41559_ ( .A(_tmp_75), .B(_maxi_read_local_stride), .Y({ _24494_[31:10], _tmp_84 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41560_ ( .A(_tmp_76), .B(_maxi_read_local_stride), .Y({ _24495_[31:10], _tmp_85 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41561_ ( .A(_tmp_77), .B(_maxi_read_local_stride), .Y({ _24496_[31:10], _tmp_86 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41562_ ( .A(_tmp_78), .B(_maxi_read_local_stride), .Y({ _24497_[31:10], _tmp_87 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41563_ ( .A(_tmp_79), .B(_maxi_read_local_stride), .Y({ _24498_[31:10], _tmp_88 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41564_ ( .A(_tmp_80), .B(_maxi_read_local_stride), .Y({ _24499_[31:10], _tmp_89 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41565_ ( .A(_tmp_103), .B(_maxi_read_local_stride), .Y({ _24500_[31:10], _tmp_112 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41566_ ( .A(_tmp_104), .B(_maxi_read_local_stride), .Y({ _24501_[31:10], _tmp_113 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41567_ ( .A(_tmp_105), .B(_maxi_read_local_stride), .Y({ _24502_[31:10], _tmp_114 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41568_ ( .A(_tmp_106), .B(_maxi_read_local_stride), .Y({ _24503_[31:10], _tmp_115 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41569_ ( .A(_tmp_107), .B(_maxi_read_local_stride), .Y({ _24504_[31:10], _tmp_116 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41570_ ( .A(_tmp_108), .B(_maxi_read_local_stride), .Y({ _24505_[31:10], _tmp_117 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41571_ ( .A(_tmp_109), .B(_maxi_read_local_stride), .Y({ _24506_[31:10], _tmp_118 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41572_ ( .A(_tmp_110), .B(_maxi_read_local_stride), .Y({ _24507_[31:10], _tmp_119 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41573_ ( .A(_tmp_111), .B(_maxi_read_local_stride), .Y({ _24508_[31:10], _tmp_120 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41574_ ( .A(_tmp_134), .B(_maxi_read_local_stride), .Y({ _24509_[31:10], _tmp_143 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41575_ ( .A(_tmp_135), .B(_maxi_read_local_stride), .Y({ _24510_[31:10], _tmp_144 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41576_ ( .A(_tmp_136), .B(_maxi_read_local_stride), .Y({ _24511_[31:10], _tmp_145 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41577_ ( .A(_tmp_137), .B(_maxi_read_local_stride), .Y({ _24512_[31:10], _tmp_146 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41578_ ( .A(_tmp_138), .B(_maxi_read_local_stride), .Y({ _24513_[31:10], _tmp_147 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41579_ ( .A(_tmp_139), .B(_maxi_read_local_stride), .Y({ _24514_[31:10], _tmp_148 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41580_ ( .A(_tmp_140), .B(_maxi_read_local_stride), .Y({ _24515_[31:10], _tmp_149 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41581_ ( .A(_tmp_141), .B(_maxi_read_local_stride), .Y({ _24516_[31:10], _tmp_150 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41582_ ( .A(_tmp_142), .B(_maxi_read_local_stride), .Y({ _24517_[31:10], _tmp_151 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41583_ ( .A(_tmp_165), .B(_maxi_read_local_stride), .Y({ _24518_[31:10], _tmp_174 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41584_ ( .A(_tmp_166), .B(_maxi_read_local_stride), .Y({ _24519_[31:10], _tmp_175 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41585_ ( .A(_tmp_167), .B(_maxi_read_local_stride), .Y({ _24520_[31:10], _tmp_176 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41586_ ( .A(_tmp_168), .B(_maxi_read_local_stride), .Y({ _24521_[31:10], _tmp_177 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41587_ ( .A(_tmp_169), .B(_maxi_read_local_stride), .Y({ _24522_[31:10], _tmp_178 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41588_ ( .A(_tmp_170), .B(_maxi_read_local_stride), .Y({ _24523_[31:10], _tmp_179 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41589_ ( .A(_tmp_171), .B(_maxi_read_local_stride), .Y({ _24524_[31:10], _tmp_180 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41590_ ( .A(_tmp_172), .B(_maxi_read_local_stride), .Y({ _24525_[31:10], _tmp_181 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41591_ ( .A(_tmp_173), .B(_maxi_read_local_stride), .Y({ _24526_[31:10], _tmp_182 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41592_ ( .A(_tmp_196), .B(_maxi_read_local_stride), .Y({ _24527_[31:10], _tmp_205 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41593_ ( .A(_tmp_197), .B(_maxi_read_local_stride), .Y({ _24528_[31:10], _tmp_206 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41594_ ( .A(_tmp_198), .B(_maxi_read_local_stride), .Y({ _24529_[31:10], _tmp_207 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41595_ ( .A(_tmp_199), .B(_maxi_read_local_stride), .Y({ _24530_[31:10], _tmp_208 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41596_ ( .A(_tmp_200), .B(_maxi_read_local_stride), .Y({ _24531_[31:10], _tmp_209 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41597_ ( .A(_tmp_201), .B(_maxi_read_local_stride), .Y({ _24532_[31:10], _tmp_210 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41598_ ( .A(_tmp_202), .B(_maxi_read_local_stride), .Y({ _24533_[31:10], _tmp_211 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41599_ ( .A(_tmp_203), .B(_maxi_read_local_stride), .Y({ _24534_[31:10], _tmp_212 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41600_ ( .A(_tmp_204), .B(_maxi_read_local_stride), .Y({ _24535_[31:10], _tmp_213 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41601_ ( .A(_tmp_227), .B(_maxi_read_local_stride), .Y({ _24536_[31:10], _tmp_236 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41602_ ( .A(_tmp_228), .B(_maxi_read_local_stride), .Y({ _24537_[31:10], _tmp_237 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41603_ ( .A(_tmp_229), .B(_maxi_read_local_stride), .Y({ _24538_[31:10], _tmp_238 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41604_ ( .A(_tmp_230), .B(_maxi_read_local_stride), .Y({ _24539_[31:10], _tmp_239 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41605_ ( .A(_tmp_231), .B(_maxi_read_local_stride), .Y({ _24540_[31:10], _tmp_240 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41606_ ( .A(_tmp_232), .B(_maxi_read_local_stride), .Y({ _24541_[31:10], _tmp_241 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41607_ ( .A(_tmp_233), .B(_maxi_read_local_stride), .Y({ _24542_[31:10], _tmp_242 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41608_ ( .A(_tmp_234), .B(_maxi_read_local_stride), .Y({ _24543_[31:10], _tmp_243 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41609_ ( .A(_tmp_235), .B(_maxi_read_local_stride), .Y({ _24544_[31:10], _tmp_244 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41610_ ( .A(_tmp_258), .B(_maxi_read_local_stride), .Y({ _24545_[31:10], _tmp_267 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41611_ ( .A(_tmp_259), .B(_maxi_read_local_stride), .Y({ _24546_[31:10], _tmp_268 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41612_ ( .A(_tmp_260), .B(_maxi_read_local_stride), .Y({ _24547_[31:10], _tmp_269 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41613_ ( .A(_tmp_261), .B(_maxi_read_local_stride), .Y({ _24548_[31:10], _tmp_270 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41614_ ( .A(_tmp_262), .B(_maxi_read_local_stride), .Y({ _24549_[31:10], _tmp_271 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41615_ ( .A(_tmp_263), .B(_maxi_read_local_stride), .Y({ _24550_[31:10], _tmp_272 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41616_ ( .A(_tmp_264), .B(_maxi_read_local_stride), .Y({ _24551_[31:10], _tmp_273 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41617_ ( .A(_tmp_265), .B(_maxi_read_local_stride), .Y({ _24552_[31:10], _tmp_274 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41618_ ( .A(_tmp_266), .B(_maxi_read_local_stride), .Y({ _24553_[31:10], _tmp_275 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41619_ ( .A(conv2d_16_act_base_offset), .B(cparam_conv2d_16_act_offset_values_2), .Y(_24556_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41620_ ( .A(conv2d_16_arg_objaddr_0), .B(_24556_), .Y(_24557_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41621_ ( .A(conv2d_16_arg_objaddr_0), .B(conv2d_16_act_base_offset), .Y(_24558_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41622_ ( .A(conv2d_16_act_base_offset), .B(cparam_conv2d_16_act_offset_values_0), .Y(_24554_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41623_ ( .A(conv2d_16_arg_objaddr_0), .B(_24554_), .Y(_24555_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41624_ ( .A(conv2d_16_row_count), .B(1), .Y({ _05346_, _05345_, _05343_, _05342_, _05341_, _05340_, _05339_, _05338_, _05337_, _05336_, _05335_, _05334_, _05332_, _05331_, _05330_, _05329_, _05328_, _05327_, _05326_, _05325_, _05324_, _05323_, _05353_, _05352_, _05351_, _05350_, _05349_, _05348_, _05347_, _05344_, _05333_, _05322_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41625_ ( .A(conv2d_16_row_count), .B(2), .Y({ _05378_, _05377_, _05375_, _05374_, _05373_, _05372_, _05371_, _05370_, _05369_, _05368_, _05367_, _05366_, _05364_, _05363_, _05362_, _05361_, _05360_, _05359_, _05358_, _05357_, _05356_, _05355_, _05385_, _05384_, _05383_, _05382_, _05381_, _05380_, _05379_, _05376_, _05365_, _05354_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41626_ ( .A(_tmp_294), .B(_maxi_read_local_stride), .Y({ _24559_[31:9], _tmp_297 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41627_ ( .A(_tmp_295), .B(_maxi_read_local_stride), .Y({ _24560_[31:9], _tmp_298 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41628_ ( .A(_tmp_296), .B(_maxi_read_local_stride), .Y({ _24561_[31:9], _tmp_299 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41629_ ( .A(_tmp_307), .B(_maxi_read_local_stride), .Y({ _24562_[31:9], _tmp_310 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41630_ ( .A(_tmp_308), .B(_maxi_read_local_stride), .Y({ _24563_[31:9], _tmp_311 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41631_ ( .A(_tmp_309), .B(_maxi_read_local_stride), .Y({ _24564_[31:9], _tmp_312 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41632_ ( .A(_tmp_320), .B(_maxi_read_local_stride), .Y({ _24565_[31:9], _tmp_323 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41633_ ( .A(_tmp_321), .B(_maxi_read_local_stride), .Y({ _24566_[31:9], _tmp_324 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41634_ ( .A(_tmp_322), .B(_maxi_read_local_stride), .Y({ _24567_[31:9], _tmp_325 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41635_ ( .A(_tmp_333), .B(_maxi_read_local_stride), .Y({ _24568_[31:9], _tmp_336 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41636_ ( .A(_tmp_334), .B(_maxi_read_local_stride), .Y({ _24569_[31:9], _tmp_337 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41637_ ( .A(_tmp_335), .B(_maxi_read_local_stride), .Y({ _24570_[31:9], _tmp_338 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41638_ ( .A(_tmp_351), .B(_maxi_read_local_stride), .Y({ _24571_[31:9], _tmp_354 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41639_ ( .A(_tmp_352), .B(_maxi_read_local_stride), .Y({ _24572_[31:9], _tmp_355 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41640_ ( .A(_tmp_353), .B(_maxi_read_local_stride), .Y({ _24573_[31:9], _tmp_356 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41641_ ( .A(_tmp_364), .B(_maxi_read_local_stride), .Y({ _24574_[31:9], _tmp_367 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41642_ ( .A(_tmp_365), .B(_maxi_read_local_stride), .Y({ _24575_[31:9], _tmp_368 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41643_ ( .A(_tmp_366), .B(_maxi_read_local_stride), .Y({ _24576_[31:9], _tmp_369 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41644_ ( .A(_tmp_377), .B(_maxi_read_local_stride), .Y({ _24577_[31:9], _tmp_380 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41645_ ( .A(_tmp_378), .B(_maxi_read_local_stride), .Y({ _24578_[31:9], _tmp_381 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41646_ ( .A(_tmp_379), .B(_maxi_read_local_stride), .Y({ _24579_[31:9], _tmp_382 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41647_ ( .A(_tmp_390), .B(_maxi_read_local_stride), .Y({ _24580_[31:9], _tmp_393 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41648_ ( .A(_tmp_391), .B(_maxi_read_local_stride), .Y({ _24581_[31:9], _tmp_394 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41649_ ( .A(_tmp_392), .B(_maxi_read_local_stride), .Y({ _24582_[31:9], _tmp_395 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41650_ ( .A(_tmp_408), .B(_maxi_read_local_stride), .Y({ _24583_[31:9], _tmp_411 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41651_ ( .A(_tmp_409), .B(_maxi_read_local_stride), .Y({ _24584_[31:9], _tmp_412 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41652_ ( .A(_tmp_410), .B(_maxi_read_local_stride), .Y({ _24585_[31:9], _tmp_413 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41653_ ( .A(_tmp_421), .B(_maxi_read_local_stride), .Y({ _24586_[31:9], _tmp_424 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41654_ ( .A(_tmp_422), .B(_maxi_read_local_stride), .Y({ _24587_[31:9], _tmp_425 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41655_ ( .A(_tmp_423), .B(_maxi_read_local_stride), .Y({ _24588_[31:9], _tmp_426 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41656_ ( .A(_tmp_434), .B(_maxi_read_local_stride), .Y({ _24589_[31:9], _tmp_437 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41657_ ( .A(_tmp_435), .B(_maxi_read_local_stride), .Y({ _24590_[31:9], _tmp_438 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41658_ ( .A(_tmp_436), .B(_maxi_read_local_stride), .Y({ _24591_[31:9], _tmp_439 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41659_ ( .A(_tmp_447), .B(_maxi_read_local_stride), .Y({ _24592_[31:9], _tmp_450 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41660_ ( .A(_tmp_448), .B(_maxi_read_local_stride), .Y({ _24593_[31:9], _tmp_451 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41661_ ( .A(_tmp_449), .B(_maxi_read_local_stride), .Y({ _24594_[31:9], _tmp_452 }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41662_ ( .A(conv2d_16_row_count_buf), .B(1), .Y({ _05474_, _05473_, _05471_, _05470_, _05469_, _05468_, _05467_, _05466_, _05465_, _05464_, _05463_, _05462_, _05460_, _05459_, _05458_, _05457_, _05456_, _05455_, _05454_, _05453_, _05452_, _05451_, _05481_, _05480_, _05479_, _05478_, _05477_, _05476_, _05475_, _05472_, _05461_, _05450_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41663_ ( .A(conv2d_16_col_count), .B(1), .Y({ _05410_, _05409_, _05407_, _05406_, _05405_, _05404_, _05403_, _05402_, _05401_, _05400_, _05399_, _05398_, _05396_, _05395_, _05394_, _05393_, _05392_, _05391_, _05390_, _05389_, _05388_, _05387_, _05417_, _05416_, _05415_, _05414_, _05413_, _05412_, _05411_, _05408_, _05397_, _05386_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41664_ ( .A(conv2d_16_col_count), .B(2), .Y({ _05442_, _05441_, _05439_, _05438_, _05437_, _05436_, _05435_, _05434_, _05433_, _05432_, _05431_, _05430_, _05428_, _05427_, _05426_, _05425_, _05424_, _05423_, _05422_, _05421_, _05420_, _05419_, _05449_, _05448_, _05447_, _05446_, _05445_, _05444_, _05443_, _05440_, _05429_, _05418_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41665_ ( .A(conv2d_16_row_count_buf), .B(2), .Y({ _05506_, _05505_, _05503_, _05502_, _05501_, _05500_, _05499_, _05498_, _05497_, _05496_, _05495_, _05494_, _05492_, _05491_, _05490_, _05489_, _05488_, _05487_, _05486_, _05485_, _05484_, _05483_, _05513_, _05512_, _05511_, _05510_, _05509_, _05508_, _05507_, _05504_, _05493_, _05482_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(6), .B_SIGNED(0), .B_WIDTH(1), .Y_WIDTH(32) ) _41666_ ( .A(cparam_conv2d_16_act_num_row), .B(1'h1), .Y({ _05314_, _05313_, _05311_, _05310_, _05309_, _05308_, _05307_, _05306_, _05305_, _05304_, _05303_, _05302_, _05300_, _05299_, _05298_, _05297_, _05296_, _05295_, _05294_, _05293_, _05292_, _05291_, _05321_, _05320_, _05319_, _05318_, _05317_, _05316_, _05315_, _05312_, _05301_, _05290_ }) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41667_ ( .A(_stream_conv2d_16_source_6_source_offset_buf), .B(_source_stream_conv2d_16_source_6_pat_cur_offset_0), .Y(_24595_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41668_ ( .A(_24595_), .B(_source_stream_conv2d_16_source_6_pat_cur_offset_1), .Y(_24596_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41669_ ( .A(_24596_), .B(_source_stream_conv2d_16_source_6_pat_cur_offset_2), .Y(_24597_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41670_ ( .A(_24597_), .B(_source_stream_conv2d_16_source_6_pat_cur_offset_3), .Y(_stream_conv2d_16_source_6_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41671_ ( .A(_stream_conv2d_16_source_8_source_offset_buf), .B(_source_stream_conv2d_16_source_8_pat_cur_offset_0), .Y(_24598_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41672_ ( .A(_24598_), .B(_source_stream_conv2d_16_source_8_pat_cur_offset_1), .Y(_24599_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41673_ ( .A(_24599_), .B(_source_stream_conv2d_16_source_8_pat_cur_offset_2), .Y(_24600_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41674_ ( .A(_24600_), .B(_source_stream_conv2d_16_source_8_pat_cur_offset_3), .Y(_stream_conv2d_16_source_8_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41675_ ( .A(_stream_conv2d_16_source_19_source_offset_buf), .B(_source_stream_conv2d_16_source_19_pat_cur_offset_0), .Y(_24601_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41676_ ( .A(_24601_), .B(_source_stream_conv2d_16_source_19_pat_cur_offset_1), .Y(_24602_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41677_ ( .A(_24602_), .B(_source_stream_conv2d_16_source_19_pat_cur_offset_2), .Y(_24603_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41678_ ( .A(_24603_), .B(_source_stream_conv2d_16_source_19_pat_cur_offset_3), .Y(_stream_conv2d_16_source_19_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41679_ ( .A(_stream_conv2d_16_source_20_source_offset_buf), .B(_source_stream_conv2d_16_source_20_pat_cur_offset_0), .Y(_24604_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41680_ ( .A(_24604_), .B(_source_stream_conv2d_16_source_20_pat_cur_offset_1), .Y(_24605_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41681_ ( .A(_24605_), .B(_source_stream_conv2d_16_source_20_pat_cur_offset_2), .Y(_24606_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41682_ ( .A(_24606_), .B(_source_stream_conv2d_16_source_20_pat_cur_offset_3), .Y(_stream_conv2d_16_source_20_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41683_ ( .A(_stream_conv2d_16_source_21_source_offset_buf), .B(_source_stream_conv2d_16_source_21_pat_cur_offset_0), .Y(_24607_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41684_ ( .A(_24607_), .B(_source_stream_conv2d_16_source_21_pat_cur_offset_1), .Y(_24608_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41685_ ( .A(_24608_), .B(_source_stream_conv2d_16_source_21_pat_cur_offset_2), .Y(_24609_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41686_ ( .A(_24609_), .B(_source_stream_conv2d_16_source_21_pat_cur_offset_3), .Y(_stream_conv2d_16_source_21_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41687_ ( .A(_stream_conv2d_16_source_22_source_offset_buf), .B(_source_stream_conv2d_16_source_22_pat_cur_offset_0), .Y(_24610_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41688_ ( .A(_24610_), .B(_source_stream_conv2d_16_source_22_pat_cur_offset_1), .Y(_24611_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41689_ ( .A(_24611_), .B(_source_stream_conv2d_16_source_22_pat_cur_offset_2), .Y(_24612_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41690_ ( .A(_24612_), .B(_source_stream_conv2d_16_source_22_pat_cur_offset_3), .Y(_stream_conv2d_16_source_22_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41691_ ( .A(_stream_conv2d_16_source_23_source_offset_buf), .B(_source_stream_conv2d_16_source_23_pat_cur_offset_0), .Y(_24613_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41692_ ( .A(_24613_), .B(_source_stream_conv2d_16_source_23_pat_cur_offset_1), .Y(_24614_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41693_ ( .A(_24614_), .B(_source_stream_conv2d_16_source_23_pat_cur_offset_2), .Y(_24615_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41694_ ( .A(_24615_), .B(_source_stream_conv2d_16_source_23_pat_cur_offset_3), .Y(_stream_conv2d_16_source_23_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41695_ ( .A(_stream_conv2d_16_source_24_source_offset_buf), .B(_source_stream_conv2d_16_source_24_pat_cur_offset_0), .Y(_24616_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41696_ ( .A(_24616_), .B(_source_stream_conv2d_16_source_24_pat_cur_offset_1), .Y(_24617_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41697_ ( .A(_24617_), .B(_source_stream_conv2d_16_source_24_pat_cur_offset_2), .Y(_24618_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41698_ ( .A(_24618_), .B(_source_stream_conv2d_16_source_24_pat_cur_offset_3), .Y(_stream_conv2d_16_source_24_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41699_ ( .A(_stream_conv2d_16_source_25_source_offset_buf), .B(_source_stream_conv2d_16_source_25_pat_cur_offset_0), .Y(_24619_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41700_ ( .A(_24619_), .B(_source_stream_conv2d_16_source_25_pat_cur_offset_1), .Y(_24620_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41701_ ( .A(_24620_), .B(_source_stream_conv2d_16_source_25_pat_cur_offset_2), .Y(_24621_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41702_ ( .A(_24621_), .B(_source_stream_conv2d_16_source_25_pat_cur_offset_3), .Y(_stream_conv2d_16_source_25_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41703_ ( .A(_stream_conv2d_16_source_26_source_offset_buf), .B(_source_stream_conv2d_16_source_26_pat_cur_offset_0), .Y(_24622_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41704_ ( .A(_24622_), .B(_source_stream_conv2d_16_source_26_pat_cur_offset_1), .Y(_24623_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41705_ ( .A(_24623_), .B(_source_stream_conv2d_16_source_26_pat_cur_offset_2), .Y(_24624_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41706_ ( .A(_24624_), .B(_source_stream_conv2d_16_source_26_pat_cur_offset_3), .Y(_stream_conv2d_16_source_26_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41707_ ( .A(_stream_conv2d_16_source_27_source_offset_buf), .B(_source_stream_conv2d_16_source_27_pat_cur_offset_0), .Y(_24625_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41708_ ( .A(_24625_), .B(_source_stream_conv2d_16_source_27_pat_cur_offset_1), .Y(_24626_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41709_ ( .A(_24626_), .B(_source_stream_conv2d_16_source_27_pat_cur_offset_2), .Y(_24627_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41710_ ( .A(_24627_), .B(_source_stream_conv2d_16_source_27_pat_cur_offset_3), .Y(_stream_conv2d_16_source_27_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41711_ ( .A(_stream_conv2d_16_source_28_source_offset_buf), .B(_source_stream_conv2d_16_source_28_pat_cur_offset_0), .Y(_24628_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41712_ ( .A(_24628_), .B(_source_stream_conv2d_16_source_28_pat_cur_offset_1), .Y(_24629_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41713_ ( .A(_24629_), .B(_source_stream_conv2d_16_source_28_pat_cur_offset_2), .Y(_24630_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41714_ ( .A(_24630_), .B(_source_stream_conv2d_16_source_28_pat_cur_offset_3), .Y(_stream_conv2d_16_source_28_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41715_ ( .A(_stream_conv2d_16_source_29_source_offset_buf), .B(_source_stream_conv2d_16_source_29_pat_cur_offset_0), .Y(_24631_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41716_ ( .A(_24631_), .B(_source_stream_conv2d_16_source_29_pat_cur_offset_1), .Y(_24632_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41717_ ( .A(_24632_), .B(_source_stream_conv2d_16_source_29_pat_cur_offset_2), .Y(_24633_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41718_ ( .A(_24633_), .B(_source_stream_conv2d_16_source_29_pat_cur_offset_3), .Y(_stream_conv2d_16_source_29_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41719_ ( .A(_stream_conv2d_16_source_30_source_offset_buf), .B(_source_stream_conv2d_16_source_30_pat_cur_offset_0), .Y(_24634_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41720_ ( .A(_24634_), .B(_source_stream_conv2d_16_source_30_pat_cur_offset_1), .Y(_24635_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41721_ ( .A(_24635_), .B(_source_stream_conv2d_16_source_30_pat_cur_offset_2), .Y(_24636_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41722_ ( .A(_24636_), .B(_source_stream_conv2d_16_source_30_pat_cur_offset_3), .Y(_stream_conv2d_16_source_30_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41723_ ( .A(_stream_conv2d_16_source_31_source_offset_buf), .B(_source_stream_conv2d_16_source_31_pat_cur_offset_0), .Y(_24637_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41724_ ( .A(_24637_), .B(_source_stream_conv2d_16_source_31_pat_cur_offset_1), .Y(_24638_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41725_ ( .A(_24638_), .B(_source_stream_conv2d_16_source_31_pat_cur_offset_2), .Y(_24639_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41726_ ( .A(_24639_), .B(_source_stream_conv2d_16_source_31_pat_cur_offset_3), .Y(_stream_conv2d_16_source_31_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41727_ ( .A(_stream_conv2d_16_source_32_source_offset_buf), .B(_source_stream_conv2d_16_source_32_pat_cur_offset_0), .Y(_24640_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41728_ ( .A(_24640_), .B(_source_stream_conv2d_16_source_32_pat_cur_offset_1), .Y(_24641_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41729_ ( .A(_24641_), .B(_source_stream_conv2d_16_source_32_pat_cur_offset_2), .Y(_24642_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41730_ ( .A(_24642_), .B(_source_stream_conv2d_16_source_32_pat_cur_offset_3), .Y(_stream_conv2d_16_source_32_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41731_ ( .A(_stream_conv2d_16_source_33_source_offset_buf), .B(_source_stream_conv2d_16_source_33_pat_cur_offset_0), .Y(_24643_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41732_ ( .A(_24643_), .B(_source_stream_conv2d_16_source_33_pat_cur_offset_1), .Y(_24644_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41733_ ( .A(_24644_), .B(_source_stream_conv2d_16_source_33_pat_cur_offset_2), .Y(_24645_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41734_ ( .A(_24645_), .B(_source_stream_conv2d_16_source_33_pat_cur_offset_3), .Y(_stream_conv2d_16_source_33_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41735_ ( .A(_stream_conv2d_16_source_34_source_offset_buf), .B(_source_stream_conv2d_16_source_34_pat_cur_offset_0), .Y(_24646_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41736_ ( .A(_24646_), .B(_source_stream_conv2d_16_source_34_pat_cur_offset_1), .Y(_24647_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41737_ ( .A(_24647_), .B(_source_stream_conv2d_16_source_34_pat_cur_offset_2), .Y(_24648_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41738_ ( .A(_24648_), .B(_source_stream_conv2d_16_source_34_pat_cur_offset_3), .Y(_stream_conv2d_16_source_34_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41739_ ( .A(_stream_conv2d_16_source_35_source_offset_buf), .B(_source_stream_conv2d_16_source_35_pat_cur_offset_0), .Y(_24649_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41740_ ( .A(_24649_), .B(_source_stream_conv2d_16_source_35_pat_cur_offset_1), .Y(_24650_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41741_ ( .A(_24650_), .B(_source_stream_conv2d_16_source_35_pat_cur_offset_2), .Y(_24651_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41742_ ( .A(_24651_), .B(_source_stream_conv2d_16_source_35_pat_cur_offset_3), .Y(_stream_conv2d_16_source_35_source_pat_all_offset) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41743_ ( .A(_stream_conv2d_16_source_36_source_offset_buf), .B(_source_stream_conv2d_16_source_36_pat_cur_offset_0), .Y(_24652_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41744_ ( .A(_24652_), .B(_source_stream_conv2d_16_source_36_pat_cur_offset_1), .Y(_24653_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41745_ ( .A(_24653_), .B(_source_stream_conv2d_16_source_36_pat_cur_offset_2), .Y(_24654_) );
  \$add  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _41746_ ( .A(_24654_), .B(_source_stream_conv2d_16_source_36_pat_cur_offset_3), .Y(_stream_conv2d_16_source_36_source_pat_all_offset) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(12), .B_SIGNED(1), .B_WIDTH(12), .Y_WIDTH(12) ) _54132_ ( .A(\__muladd_madd_103.madd._mul ), .B(\__muladd_madd_103.madd._c ), .Y(\__muladd_madd_103.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(12), .B_SIGNED(1), .B_WIDTH(12), .Y_WIDTH(12) ) _54139_ ( .A(\__muladd_madd_120.madd._mul ), .B(\__muladd_madd_120.madd._c ), .Y(\__muladd_madd_120.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(12), .B_SIGNED(1), .B_WIDTH(12), .Y_WIDTH(12) ) _54146_ ( .A(\__muladd_madd_137.madd._mul ), .B(\__muladd_madd_137.madd._c ), .Y(\__muladd_madd_137.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(12), .B_SIGNED(1), .B_WIDTH(12), .Y_WIDTH(12) ) _54153_ ( .A(\__muladd_madd_154.madd._mul ), .B(\__muladd_madd_154.madd._c ), .Y(\__muladd_madd_154.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(12), .B_SIGNED(1), .B_WIDTH(12), .Y_WIDTH(12) ) _54160_ ( .A(\__muladd_madd_171.madd._mul ), .B(\__muladd_madd_171.madd._c ), .Y(\__muladd_madd_171.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(12), .B_SIGNED(1), .B_WIDTH(12), .Y_WIDTH(12) ) _54167_ ( .A(\__muladd_madd_188.madd._mul ), .B(\__muladd_madd_188.madd._c ), .Y(\__muladd_madd_188.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(12), .B_SIGNED(1), .B_WIDTH(12), .Y_WIDTH(12) ) _54174_ ( .A(\__muladd_madd_205.madd._mul ), .B(\__muladd_madd_205.madd._c ), .Y(\__muladd_madd_205.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(12), .B_SIGNED(1), .B_WIDTH(12), .Y_WIDTH(12) ) _54181_ ( .A(\__muladd_madd_69.madd._mul ), .B(\__muladd_madd_69.madd._c ), .Y(\__muladd_madd_69.madd._madd ) );
  \$add  #( .A_SIGNED(1), .A_WIDTH(12), .B_SIGNED(1), .B_WIDTH(12), .Y_WIDTH(12) ) _54188_ ( .A(\__muladd_madd_86.madd._mul ), .B(\__muladd_madd_86.madd._c ), .Y(\__muladd_madd_86.madd._madd ) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53431_ ( .A(_maxi_read_cur_size), .B(1), .Y(_28532_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53432_ ( .A(_tmp_20), .B(1), .Y(_28533_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53433_ ( .A(_maxi_write_cur_size), .B(1), .Y(_28534_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53434_ ( .A(_tmp_1019), .B(1), .Y(_28535_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(11), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53435_ ( .A(_tmp_38), .B(1), .Y(_28538_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53436_ ( .A(_tmp_39), .B(1), .Y(_28539_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53437_ ( .A(_tmp_1136), .B(1), .Y(_28540_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(11), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53438_ ( .A(_tmp_69), .B(1), .Y(_28541_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53439_ ( .A(_tmp_70), .B(1), .Y(_28542_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53440_ ( .A(_tmp_1138), .B(1), .Y(_28543_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(11), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53441_ ( .A(_tmp_100), .B(1), .Y(_28544_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53442_ ( .A(_tmp_101), .B(1), .Y(_28545_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53443_ ( .A(_tmp_1140), .B(1), .Y(_28546_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(11), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53444_ ( .A(_tmp_131), .B(1), .Y(_28547_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53445_ ( .A(_tmp_132), .B(1), .Y(_28548_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53446_ ( .A(_tmp_1142), .B(1), .Y(_28549_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(11), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53447_ ( .A(_tmp_162), .B(1), .Y(_28550_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53448_ ( .A(_tmp_163), .B(1), .Y(_28551_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53449_ ( .A(_tmp_1144), .B(1), .Y(_28552_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(11), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53450_ ( .A(_tmp_193), .B(1), .Y(_28553_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53451_ ( .A(_tmp_194), .B(1), .Y(_28554_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53452_ ( .A(_tmp_1146), .B(1), .Y(_28555_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(11), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53453_ ( .A(_tmp_224), .B(1), .Y(_28556_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53454_ ( .A(_tmp_225), .B(1), .Y(_28557_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53455_ ( .A(_tmp_1148), .B(1), .Y(_28558_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(11), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53456_ ( .A(_tmp_255), .B(1), .Y(_28559_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53457_ ( .A(_tmp_256), .B(1), .Y(_28560_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53458_ ( .A(req_block_size_33), .B(1), .Y(_28536_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53459_ ( .A(_tmp_1150), .B(1), .Y(_28561_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53460_ ( .A(_tmp_25), .B(1), .Y(_28562_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53461_ ( .A(_tmp_1083), .B(1), .Y(_28564_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53462_ ( .A(_tmp_27), .B(1), .Y(_28565_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53463_ ( .A(_tmp_1095), .B(1), .Y(_28566_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53464_ ( .A(_tmp_29), .B(1), .Y(_28567_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53465_ ( .A(_tmp_1107), .B(1), .Y(_28568_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53466_ ( .A(_tmp_31), .B(1), .Y(_28569_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53467_ ( .A(_tmp_1119), .B(1), .Y(_28570_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53468_ ( .A(_tmp_12), .B(1), .Y(_28571_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53469_ ( .A(_tmp_1320), .B(1), .Y(_28572_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53470_ ( .A(_tmp_14), .B(1), .Y(_28573_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53471_ ( .A(_tmp_1332), .B(1), .Y(_28574_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53472_ ( .A(_tmp_16), .B(1), .Y(_28575_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53473_ ( .A(_tmp_1344), .B(1), .Y(_28576_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53474_ ( .A(_tmp_18), .B(1), .Y(_28577_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53475_ ( .A(_tmp_1356), .B(1), .Y(_28578_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53476_ ( .A(_tmp_291), .B(1), .Y(_28580_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53477_ ( .A(_tmp_292), .B(1), .Y(_28581_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53478_ ( .A(_tmp_1124), .B(1), .Y(_28582_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53479_ ( .A(_tmp_304), .B(1), .Y(_28583_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53480_ ( .A(_tmp_305), .B(1), .Y(_28584_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53481_ ( .A(_tmp_1126), .B(1), .Y(_28585_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53482_ ( .A(_tmp_317), .B(1), .Y(_28586_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53483_ ( .A(_tmp_318), .B(1), .Y(_28587_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53484_ ( .A(_tmp_1128), .B(1), .Y(_28588_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53485_ ( .A(_tmp_330), .B(1), .Y(_28589_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53486_ ( .A(_tmp_331), .B(1), .Y(_28590_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53487_ ( .A(req_block_size_286), .B(1), .Y(_28579_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53488_ ( .A(_tmp_1130), .B(1), .Y(_28591_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53489_ ( .A(_tmp_1155), .B(1), .Y(_28592_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53490_ ( .A(_tmp_1157), .B(1), .Y(_28593_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53491_ ( .A(_tmp_1159), .B(1), .Y(_28594_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53492_ ( .A(_tmp_1161), .B(1), .Y(_28595_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53493_ ( .A(_tmp_348), .B(1), .Y(_28597_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53494_ ( .A(_tmp_349), .B(1), .Y(_28598_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53495_ ( .A(_tmp_361), .B(1), .Y(_28599_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53496_ ( .A(_tmp_362), .B(1), .Y(_28600_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53497_ ( .A(_tmp_374), .B(1), .Y(_28601_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53498_ ( .A(_tmp_375), .B(1), .Y(_28602_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53499_ ( .A(_tmp_387), .B(1), .Y(_28603_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53500_ ( .A(_tmp_388), .B(1), .Y(_28604_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53501_ ( .A(req_block_size_343), .B(1), .Y(_28596_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53502_ ( .A(_tmp_405), .B(1), .Y(_28606_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53503_ ( .A(_tmp_406), .B(1), .Y(_28607_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53504_ ( .A(_tmp_418), .B(1), .Y(_28608_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53505_ ( .A(_tmp_419), .B(1), .Y(_28609_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53506_ ( .A(_tmp_431), .B(1), .Y(_28610_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53507_ ( .A(_tmp_432), .B(1), .Y(_28611_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53508_ ( .A(_maxi_read_local_addr), .B(_maxi_read_local_stride), .Y(_28537_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(10), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53509_ ( .A(_tmp_444), .B(1), .Y(_28612_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53510_ ( .A(_tmp_445), .B(1), .Y(_28613_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(9), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53511_ ( .A(req_block_size_400), .B(1), .Y(_28605_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53512_ ( .A(_tmp_982), .B(1), .Y(_28614_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53513_ ( .A(_tmp_994), .B(1), .Y(_28615_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53514_ ( .A(_tmp_1006), .B(1), .Y(_28616_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53515_ ( .A(_maxi_write_size), .B(1), .Y(_28563_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(34), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(34) ) _53516_ ( .A(_tmp_1018), .B(1), .Y(_28617_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(6), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(6) ) _53517_ ( .A(__variable_wdata_1), .B(2'h1), .Y(_28618_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53518_ ( .A(__variable_wdata_2), .B(1), .Y({ _23948_, _23947_, _23946_, _23944_, _23943_, _23942_, _23941_, _23940_, _23939_, _23938_, _23937_, _23936_, _23935_, _23933_, _23932_, _23931_, _23930_, _23929_, _23928_, _23927_, _23926_, _23925_, _23924_, _23955_, _23954_, _23953_, _23952_, _23951_, _23950_, _23949_, _23945_, _23934_, _23923_ }) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _53519_ ( .A(__variable_wdata_56), .B(2'h1), .Y(_28619_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _53520_ ( .A(__variable_wdata_73), .B(2'h1), .Y(_28620_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _53521_ ( .A(__variable_wdata_90), .B(2'h1), .Y(_28621_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _53522_ ( .A(__variable_wdata_107), .B(2'h1), .Y(_28622_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _53523_ ( .A(__variable_wdata_124), .B(2'h1), .Y(_28623_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _53524_ ( .A(__variable_wdata_141), .B(2'h1), .Y(_28624_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _53525_ ( .A(__variable_wdata_158), .B(2'h1), .Y(_28625_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _53526_ ( .A(__variable_wdata_175), .B(2'h1), .Y(_28626_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(4), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(4) ) _53527_ ( .A(__variable_wdata_192), .B(2'h1), .Y(_28627_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(8), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53528_ ( .A(__variable_wdata_208), .B(1), .Y({ _23980_, _23979_, _23977_, _23976_, _23975_, _23974_, _23973_, _23972_, _23971_, _23970_, _23969_, _23968_, _23966_, _23965_, _23964_, _23963_, _23962_, _23961_, _23960_, _23959_, _23958_, _23957_, _23987_, _23986_, _23985_, _23984_, _23983_, _23982_, _23981_, _23978_, _23967_, _23956_ }) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53529_ ( .A(_source_stream_conv2d_16_source_6_pat_size_0), .B(1), .Y(_28628_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53530_ ( .A(_source_stream_conv2d_16_source_6_pat_size_1), .B(1), .Y(_28629_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53531_ ( .A(_source_stream_conv2d_16_source_6_pat_size_2), .B(1), .Y(_28630_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53532_ ( .A(_source_stream_conv2d_16_source_6_pat_size_3), .B(1), .Y(_28631_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53533_ ( .A(_source_stream_conv2d_16_source_6_pat_count_0), .B(1), .Y(_28632_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53534_ ( .A(_source_stream_conv2d_16_source_6_pat_size_buf_0), .B(1), .Y(_28633_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53535_ ( .A(_source_stream_conv2d_16_source_6_pat_count_1), .B(1), .Y(_28634_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53536_ ( .A(_source_stream_conv2d_16_source_6_pat_size_buf_1), .B(1), .Y(_28635_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53537_ ( .A(_source_stream_conv2d_16_source_6_pat_count_2), .B(1), .Y(_28636_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53538_ ( .A(_source_stream_conv2d_16_source_6_pat_size_buf_2), .B(1), .Y(_28637_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53539_ ( .A(_source_stream_conv2d_16_source_6_pat_count_3), .B(1), .Y(_28638_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53540_ ( .A(_source_stream_conv2d_16_source_6_pat_size_buf_3), .B(1), .Y(_28639_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53541_ ( .A(_source_stream_conv2d_16_source_8_pat_size_0), .B(1), .Y(_28640_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53542_ ( .A(_source_stream_conv2d_16_source_8_pat_size_1), .B(1), .Y(_28641_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53543_ ( .A(_source_stream_conv2d_16_source_8_pat_size_2), .B(1), .Y(_28642_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53544_ ( .A(_source_stream_conv2d_16_source_8_pat_size_3), .B(1), .Y(_28643_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53545_ ( .A(_source_stream_conv2d_16_source_8_pat_count_0), .B(1), .Y(_28644_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53546_ ( .A(_source_stream_conv2d_16_source_8_pat_size_buf_0), .B(1), .Y(_28645_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53547_ ( .A(_source_stream_conv2d_16_source_8_pat_count_1), .B(1), .Y(_28646_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53548_ ( .A(_source_stream_conv2d_16_source_8_pat_size_buf_1), .B(1), .Y(_28647_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53549_ ( .A(_source_stream_conv2d_16_source_8_pat_count_2), .B(1), .Y(_28648_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53550_ ( .A(_source_stream_conv2d_16_source_8_pat_size_buf_2), .B(1), .Y(_28649_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53551_ ( .A(_source_stream_conv2d_16_source_8_pat_count_3), .B(1), .Y(_28650_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53552_ ( .A(_source_stream_conv2d_16_source_8_pat_size_buf_3), .B(1), .Y(_28651_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53553_ ( .A(_source_stream_conv2d_16_source_19_pat_size_0), .B(1), .Y(_28652_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53554_ ( .A(_source_stream_conv2d_16_source_19_pat_size_1), .B(1), .Y(_28653_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53555_ ( .A(_source_stream_conv2d_16_source_19_pat_size_2), .B(1), .Y(_28654_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53556_ ( .A(_source_stream_conv2d_16_source_19_pat_size_3), .B(1), .Y(_28655_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53557_ ( .A(_source_stream_conv2d_16_source_19_pat_count_0), .B(1), .Y(_28656_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53558_ ( .A(_source_stream_conv2d_16_source_19_pat_size_buf_0), .B(1), .Y(_28657_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53559_ ( .A(_source_stream_conv2d_16_source_19_pat_count_1), .B(1), .Y(_28658_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53560_ ( .A(_source_stream_conv2d_16_source_19_pat_size_buf_1), .B(1), .Y(_28659_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53561_ ( .A(_source_stream_conv2d_16_source_19_pat_count_2), .B(1), .Y(_28660_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53562_ ( .A(_source_stream_conv2d_16_source_19_pat_size_buf_2), .B(1), .Y(_28661_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53563_ ( .A(_source_stream_conv2d_16_source_19_pat_count_3), .B(1), .Y(_28662_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53564_ ( .A(_source_stream_conv2d_16_source_19_pat_size_buf_3), .B(1), .Y(_28663_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53565_ ( .A(_source_stream_conv2d_16_source_20_pat_size_0), .B(1), .Y(_28664_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53566_ ( .A(_source_stream_conv2d_16_source_20_pat_size_1), .B(1), .Y(_28665_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53567_ ( .A(_source_stream_conv2d_16_source_20_pat_size_2), .B(1), .Y(_28666_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53568_ ( .A(_source_stream_conv2d_16_source_20_pat_size_3), .B(1), .Y(_28667_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53569_ ( .A(_source_stream_conv2d_16_source_20_pat_count_0), .B(1), .Y(_28668_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53570_ ( .A(_source_stream_conv2d_16_source_20_pat_size_buf_0), .B(1), .Y(_28669_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53571_ ( .A(_source_stream_conv2d_16_source_20_pat_count_1), .B(1), .Y(_28670_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53572_ ( .A(_source_stream_conv2d_16_source_20_pat_size_buf_1), .B(1), .Y(_28671_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53573_ ( .A(_source_stream_conv2d_16_source_20_pat_count_2), .B(1), .Y(_28672_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53574_ ( .A(_source_stream_conv2d_16_source_20_pat_size_buf_2), .B(1), .Y(_28673_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53575_ ( .A(_source_stream_conv2d_16_source_20_pat_count_3), .B(1), .Y(_28674_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53576_ ( .A(_source_stream_conv2d_16_source_20_pat_size_buf_3), .B(1), .Y(_28675_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53577_ ( .A(_source_stream_conv2d_16_source_21_pat_size_0), .B(1), .Y(_28676_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53578_ ( .A(_source_stream_conv2d_16_source_21_pat_size_1), .B(1), .Y(_28677_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53579_ ( .A(_source_stream_conv2d_16_source_21_pat_size_2), .B(1), .Y(_28678_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53580_ ( .A(_source_stream_conv2d_16_source_21_pat_size_3), .B(1), .Y(_28679_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53581_ ( .A(_source_stream_conv2d_16_source_21_pat_count_0), .B(1), .Y(_28680_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53582_ ( .A(_source_stream_conv2d_16_source_21_pat_size_buf_0), .B(1), .Y(_28681_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53583_ ( .A(_source_stream_conv2d_16_source_21_pat_count_1), .B(1), .Y(_28682_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53584_ ( .A(_source_stream_conv2d_16_source_21_pat_size_buf_1), .B(1), .Y(_28683_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53585_ ( .A(_source_stream_conv2d_16_source_21_pat_count_2), .B(1), .Y(_28684_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53586_ ( .A(_source_stream_conv2d_16_source_21_pat_size_buf_2), .B(1), .Y(_28685_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53587_ ( .A(_source_stream_conv2d_16_source_21_pat_count_3), .B(1), .Y(_28686_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53588_ ( .A(_source_stream_conv2d_16_source_21_pat_size_buf_3), .B(1), .Y(_28687_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53589_ ( .A(_source_stream_conv2d_16_source_22_pat_size_0), .B(1), .Y(_28688_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53590_ ( .A(_source_stream_conv2d_16_source_22_pat_size_1), .B(1), .Y(_28689_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53591_ ( .A(_source_stream_conv2d_16_source_22_pat_size_2), .B(1), .Y(_28690_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53592_ ( .A(_source_stream_conv2d_16_source_22_pat_size_3), .B(1), .Y(_28691_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53593_ ( .A(_source_stream_conv2d_16_source_22_pat_count_0), .B(1), .Y(_28692_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53594_ ( .A(_source_stream_conv2d_16_source_22_pat_size_buf_0), .B(1), .Y(_28693_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53595_ ( .A(_source_stream_conv2d_16_source_22_pat_count_1), .B(1), .Y(_28694_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53596_ ( .A(_source_stream_conv2d_16_source_22_pat_size_buf_1), .B(1), .Y(_28695_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53597_ ( .A(_source_stream_conv2d_16_source_22_pat_count_2), .B(1), .Y(_28696_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53598_ ( .A(_source_stream_conv2d_16_source_22_pat_size_buf_2), .B(1), .Y(_28697_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53599_ ( .A(_source_stream_conv2d_16_source_22_pat_count_3), .B(1), .Y(_28698_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53600_ ( .A(_source_stream_conv2d_16_source_22_pat_size_buf_3), .B(1), .Y(_28699_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53601_ ( .A(_source_stream_conv2d_16_source_23_pat_size_0), .B(1), .Y(_28700_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53602_ ( .A(_source_stream_conv2d_16_source_23_pat_size_1), .B(1), .Y(_28701_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53603_ ( .A(_source_stream_conv2d_16_source_23_pat_size_2), .B(1), .Y(_28702_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53604_ ( .A(_source_stream_conv2d_16_source_23_pat_size_3), .B(1), .Y(_28703_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53605_ ( .A(_source_stream_conv2d_16_source_23_pat_count_0), .B(1), .Y(_28704_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53606_ ( .A(_source_stream_conv2d_16_source_23_pat_size_buf_0), .B(1), .Y(_28705_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53607_ ( .A(_source_stream_conv2d_16_source_23_pat_count_1), .B(1), .Y(_28706_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53608_ ( .A(_source_stream_conv2d_16_source_23_pat_size_buf_1), .B(1), .Y(_28707_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53609_ ( .A(_source_stream_conv2d_16_source_23_pat_count_2), .B(1), .Y(_28708_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53610_ ( .A(_source_stream_conv2d_16_source_23_pat_size_buf_2), .B(1), .Y(_28709_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53611_ ( .A(_source_stream_conv2d_16_source_23_pat_count_3), .B(1), .Y(_28710_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53612_ ( .A(_source_stream_conv2d_16_source_23_pat_size_buf_3), .B(1), .Y(_28711_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53613_ ( .A(_source_stream_conv2d_16_source_24_pat_size_0), .B(1), .Y(_28712_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53614_ ( .A(_source_stream_conv2d_16_source_24_pat_size_1), .B(1), .Y(_28713_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53615_ ( .A(_source_stream_conv2d_16_source_24_pat_size_2), .B(1), .Y(_28714_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53616_ ( .A(_source_stream_conv2d_16_source_24_pat_size_3), .B(1), .Y(_28715_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53617_ ( .A(_source_stream_conv2d_16_source_24_pat_count_0), .B(1), .Y(_28716_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53618_ ( .A(_source_stream_conv2d_16_source_24_pat_size_buf_0), .B(1), .Y(_28717_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53619_ ( .A(_source_stream_conv2d_16_source_24_pat_count_1), .B(1), .Y(_28718_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53620_ ( .A(_source_stream_conv2d_16_source_24_pat_size_buf_1), .B(1), .Y(_28719_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53621_ ( .A(_source_stream_conv2d_16_source_24_pat_count_2), .B(1), .Y(_28720_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53622_ ( .A(_source_stream_conv2d_16_source_24_pat_size_buf_2), .B(1), .Y(_28721_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53623_ ( .A(_source_stream_conv2d_16_source_24_pat_count_3), .B(1), .Y(_28722_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53624_ ( .A(_source_stream_conv2d_16_source_24_pat_size_buf_3), .B(1), .Y(_28723_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53625_ ( .A(_source_stream_conv2d_16_source_25_pat_size_0), .B(1), .Y(_28724_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53626_ ( .A(_source_stream_conv2d_16_source_25_pat_size_1), .B(1), .Y(_28725_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53627_ ( .A(_source_stream_conv2d_16_source_25_pat_size_2), .B(1), .Y(_28726_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53628_ ( .A(_source_stream_conv2d_16_source_25_pat_size_3), .B(1), .Y(_28727_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53629_ ( .A(_source_stream_conv2d_16_source_25_pat_count_0), .B(1), .Y(_28728_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53630_ ( .A(_source_stream_conv2d_16_source_25_pat_size_buf_0), .B(1), .Y(_28729_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53631_ ( .A(_source_stream_conv2d_16_source_25_pat_count_1), .B(1), .Y(_28730_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53632_ ( .A(_source_stream_conv2d_16_source_25_pat_size_buf_1), .B(1), .Y(_28731_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53633_ ( .A(_source_stream_conv2d_16_source_25_pat_count_2), .B(1), .Y(_28732_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53634_ ( .A(_source_stream_conv2d_16_source_25_pat_size_buf_2), .B(1), .Y(_28733_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53635_ ( .A(_source_stream_conv2d_16_source_25_pat_count_3), .B(1), .Y(_28734_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53636_ ( .A(_source_stream_conv2d_16_source_25_pat_size_buf_3), .B(1), .Y(_28735_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53637_ ( .A(_source_stream_conv2d_16_source_26_pat_size_0), .B(1), .Y(_28736_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53638_ ( .A(_source_stream_conv2d_16_source_26_pat_size_1), .B(1), .Y(_28737_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53639_ ( .A(_source_stream_conv2d_16_source_26_pat_size_2), .B(1), .Y(_28738_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53640_ ( .A(_source_stream_conv2d_16_source_26_pat_size_3), .B(1), .Y(_28739_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53641_ ( .A(_source_stream_conv2d_16_source_26_pat_count_0), .B(1), .Y(_28740_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53642_ ( .A(_source_stream_conv2d_16_source_26_pat_size_buf_0), .B(1), .Y(_28741_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53643_ ( .A(_source_stream_conv2d_16_source_26_pat_count_1), .B(1), .Y(_28742_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53644_ ( .A(_source_stream_conv2d_16_source_26_pat_size_buf_1), .B(1), .Y(_28743_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53645_ ( .A(_source_stream_conv2d_16_source_26_pat_count_2), .B(1), .Y(_28744_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53646_ ( .A(_source_stream_conv2d_16_source_26_pat_size_buf_2), .B(1), .Y(_28745_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53647_ ( .A(_source_stream_conv2d_16_source_26_pat_count_3), .B(1), .Y(_28746_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53648_ ( .A(_source_stream_conv2d_16_source_26_pat_size_buf_3), .B(1), .Y(_28747_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53649_ ( .A(_source_stream_conv2d_16_source_27_pat_size_0), .B(1), .Y(_28748_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53650_ ( .A(_source_stream_conv2d_16_source_27_pat_size_1), .B(1), .Y(_28749_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53651_ ( .A(_source_stream_conv2d_16_source_27_pat_size_2), .B(1), .Y(_28750_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53652_ ( .A(_source_stream_conv2d_16_source_27_pat_size_3), .B(1), .Y(_28751_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53653_ ( .A(_source_stream_conv2d_16_source_27_pat_count_0), .B(1), .Y(_28752_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53654_ ( .A(_source_stream_conv2d_16_source_27_pat_size_buf_0), .B(1), .Y(_28753_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53655_ ( .A(_source_stream_conv2d_16_source_27_pat_count_1), .B(1), .Y(_28754_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53656_ ( .A(_source_stream_conv2d_16_source_27_pat_size_buf_1), .B(1), .Y(_28755_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53657_ ( .A(_source_stream_conv2d_16_source_27_pat_count_2), .B(1), .Y(_28756_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53658_ ( .A(_source_stream_conv2d_16_source_27_pat_size_buf_2), .B(1), .Y(_28757_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53659_ ( .A(_source_stream_conv2d_16_source_27_pat_count_3), .B(1), .Y(_28758_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53660_ ( .A(_source_stream_conv2d_16_source_27_pat_size_buf_3), .B(1), .Y(_28759_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53661_ ( .A(_source_stream_conv2d_16_source_28_pat_size_0), .B(1), .Y(_28760_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53662_ ( .A(_source_stream_conv2d_16_source_28_pat_size_1), .B(1), .Y(_28761_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53663_ ( .A(_source_stream_conv2d_16_source_28_pat_size_2), .B(1), .Y(_28762_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53664_ ( .A(_source_stream_conv2d_16_source_28_pat_size_3), .B(1), .Y(_28763_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53665_ ( .A(_source_stream_conv2d_16_source_28_pat_count_0), .B(1), .Y(_28764_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53666_ ( .A(_source_stream_conv2d_16_source_28_pat_size_buf_0), .B(1), .Y(_28765_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53667_ ( .A(_source_stream_conv2d_16_source_28_pat_count_1), .B(1), .Y(_28766_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53668_ ( .A(_source_stream_conv2d_16_source_28_pat_size_buf_1), .B(1), .Y(_28767_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53669_ ( .A(_source_stream_conv2d_16_source_28_pat_count_2), .B(1), .Y(_28768_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53670_ ( .A(_source_stream_conv2d_16_source_28_pat_size_buf_2), .B(1), .Y(_28769_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53671_ ( .A(_source_stream_conv2d_16_source_28_pat_count_3), .B(1), .Y(_28770_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53672_ ( .A(_source_stream_conv2d_16_source_28_pat_size_buf_3), .B(1), .Y(_28771_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53673_ ( .A(_source_stream_conv2d_16_source_29_pat_size_0), .B(1), .Y(_28772_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53674_ ( .A(_source_stream_conv2d_16_source_29_pat_size_1), .B(1), .Y(_28773_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53675_ ( .A(_source_stream_conv2d_16_source_29_pat_size_2), .B(1), .Y(_28774_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53676_ ( .A(_source_stream_conv2d_16_source_29_pat_size_3), .B(1), .Y(_28775_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53677_ ( .A(_source_stream_conv2d_16_source_29_pat_count_0), .B(1), .Y(_28776_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53678_ ( .A(_source_stream_conv2d_16_source_29_pat_size_buf_0), .B(1), .Y(_28777_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53679_ ( .A(_source_stream_conv2d_16_source_29_pat_count_1), .B(1), .Y(_28778_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53680_ ( .A(_source_stream_conv2d_16_source_29_pat_size_buf_1), .B(1), .Y(_28779_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53681_ ( .A(_source_stream_conv2d_16_source_29_pat_count_2), .B(1), .Y(_28780_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53682_ ( .A(_source_stream_conv2d_16_source_29_pat_size_buf_2), .B(1), .Y(_28781_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53683_ ( .A(_source_stream_conv2d_16_source_29_pat_count_3), .B(1), .Y(_28782_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53684_ ( .A(_source_stream_conv2d_16_source_29_pat_size_buf_3), .B(1), .Y(_28783_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53685_ ( .A(_source_stream_conv2d_16_source_30_pat_size_0), .B(1), .Y(_28784_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53686_ ( .A(_source_stream_conv2d_16_source_30_pat_size_1), .B(1), .Y(_28785_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53687_ ( .A(_source_stream_conv2d_16_source_30_pat_size_2), .B(1), .Y(_28786_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53688_ ( .A(_source_stream_conv2d_16_source_30_pat_size_3), .B(1), .Y(_28787_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53689_ ( .A(_source_stream_conv2d_16_source_30_pat_count_0), .B(1), .Y(_28788_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53690_ ( .A(_source_stream_conv2d_16_source_30_pat_size_buf_0), .B(1), .Y(_28789_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53691_ ( .A(_source_stream_conv2d_16_source_30_pat_count_1), .B(1), .Y(_28790_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53692_ ( .A(_source_stream_conv2d_16_source_30_pat_size_buf_1), .B(1), .Y(_28791_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53693_ ( .A(_source_stream_conv2d_16_source_30_pat_count_2), .B(1), .Y(_28792_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53694_ ( .A(_source_stream_conv2d_16_source_30_pat_size_buf_2), .B(1), .Y(_28793_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53695_ ( .A(_source_stream_conv2d_16_source_30_pat_count_3), .B(1), .Y(_28794_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53696_ ( .A(_source_stream_conv2d_16_source_30_pat_size_buf_3), .B(1), .Y(_28795_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53697_ ( .A(_source_stream_conv2d_16_source_31_pat_size_0), .B(1), .Y(_28796_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53698_ ( .A(_source_stream_conv2d_16_source_31_pat_size_1), .B(1), .Y(_28797_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53699_ ( .A(_source_stream_conv2d_16_source_31_pat_size_2), .B(1), .Y(_28798_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53700_ ( .A(_source_stream_conv2d_16_source_31_pat_size_3), .B(1), .Y(_28799_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53701_ ( .A(_source_stream_conv2d_16_source_31_pat_count_0), .B(1), .Y(_28800_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53702_ ( .A(_source_stream_conv2d_16_source_31_pat_size_buf_0), .B(1), .Y(_28801_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53703_ ( .A(_source_stream_conv2d_16_source_31_pat_count_1), .B(1), .Y(_28802_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53704_ ( .A(_source_stream_conv2d_16_source_31_pat_size_buf_1), .B(1), .Y(_28803_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53705_ ( .A(_source_stream_conv2d_16_source_31_pat_count_2), .B(1), .Y(_28804_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53706_ ( .A(_source_stream_conv2d_16_source_31_pat_size_buf_2), .B(1), .Y(_28805_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53707_ ( .A(_source_stream_conv2d_16_source_31_pat_count_3), .B(1), .Y(_28806_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53708_ ( .A(_source_stream_conv2d_16_source_31_pat_size_buf_3), .B(1), .Y(_28807_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53709_ ( .A(_source_stream_conv2d_16_source_32_pat_size_0), .B(1), .Y(_28808_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53710_ ( .A(_source_stream_conv2d_16_source_32_pat_size_1), .B(1), .Y(_28809_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53711_ ( .A(_source_stream_conv2d_16_source_32_pat_size_2), .B(1), .Y(_28810_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53712_ ( .A(_source_stream_conv2d_16_source_32_pat_size_3), .B(1), .Y(_28811_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53713_ ( .A(_source_stream_conv2d_16_source_32_pat_count_0), .B(1), .Y(_28812_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53714_ ( .A(_source_stream_conv2d_16_source_32_pat_size_buf_0), .B(1), .Y(_28813_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53715_ ( .A(_source_stream_conv2d_16_source_32_pat_count_1), .B(1), .Y(_28814_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53716_ ( .A(_source_stream_conv2d_16_source_32_pat_size_buf_1), .B(1), .Y(_28815_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53717_ ( .A(_source_stream_conv2d_16_source_32_pat_count_2), .B(1), .Y(_28816_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53718_ ( .A(_source_stream_conv2d_16_source_32_pat_size_buf_2), .B(1), .Y(_28817_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53719_ ( .A(_source_stream_conv2d_16_source_32_pat_count_3), .B(1), .Y(_28818_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53720_ ( .A(_source_stream_conv2d_16_source_32_pat_size_buf_3), .B(1), .Y(_28819_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53721_ ( .A(_source_stream_conv2d_16_source_33_pat_size_0), .B(1), .Y(_28820_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53722_ ( .A(_source_stream_conv2d_16_source_33_pat_size_1), .B(1), .Y(_28821_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53723_ ( .A(_source_stream_conv2d_16_source_33_pat_size_2), .B(1), .Y(_28822_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53724_ ( .A(_source_stream_conv2d_16_source_33_pat_size_3), .B(1), .Y(_28823_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53725_ ( .A(_source_stream_conv2d_16_source_33_pat_count_0), .B(1), .Y(_28824_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53726_ ( .A(_source_stream_conv2d_16_source_33_pat_size_buf_0), .B(1), .Y(_28825_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53727_ ( .A(_source_stream_conv2d_16_source_33_pat_count_1), .B(1), .Y(_28826_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53728_ ( .A(_source_stream_conv2d_16_source_33_pat_size_buf_1), .B(1), .Y(_28827_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53729_ ( .A(_source_stream_conv2d_16_source_33_pat_count_2), .B(1), .Y(_28828_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53730_ ( .A(_source_stream_conv2d_16_source_33_pat_size_buf_2), .B(1), .Y(_28829_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53731_ ( .A(_source_stream_conv2d_16_source_33_pat_count_3), .B(1), .Y(_28830_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53732_ ( .A(_source_stream_conv2d_16_source_33_pat_size_buf_3), .B(1), .Y(_28831_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53733_ ( .A(_source_stream_conv2d_16_source_34_pat_size_0), .B(1), .Y(_28832_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53734_ ( .A(_source_stream_conv2d_16_source_34_pat_size_1), .B(1), .Y(_28833_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53735_ ( .A(_source_stream_conv2d_16_source_34_pat_size_2), .B(1), .Y(_28834_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53736_ ( .A(_source_stream_conv2d_16_source_34_pat_size_3), .B(1), .Y(_28835_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53737_ ( .A(_source_stream_conv2d_16_source_34_pat_count_0), .B(1), .Y(_28836_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53738_ ( .A(_source_stream_conv2d_16_source_34_pat_size_buf_0), .B(1), .Y(_28837_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53739_ ( .A(_source_stream_conv2d_16_source_34_pat_count_1), .B(1), .Y(_28838_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53740_ ( .A(_source_stream_conv2d_16_source_34_pat_size_buf_1), .B(1), .Y(_28839_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53741_ ( .A(_source_stream_conv2d_16_source_34_pat_count_2), .B(1), .Y(_28840_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53742_ ( .A(_source_stream_conv2d_16_source_34_pat_size_buf_2), .B(1), .Y(_28841_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53743_ ( .A(_source_stream_conv2d_16_source_34_pat_count_3), .B(1), .Y(_28842_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53744_ ( .A(_source_stream_conv2d_16_source_34_pat_size_buf_3), .B(1), .Y(_28843_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53745_ ( .A(_source_stream_conv2d_16_source_35_pat_size_0), .B(1), .Y(_28844_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53746_ ( .A(_source_stream_conv2d_16_source_35_pat_size_1), .B(1), .Y(_28845_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53747_ ( .A(_source_stream_conv2d_16_source_35_pat_size_2), .B(1), .Y(_28846_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53748_ ( .A(_source_stream_conv2d_16_source_35_pat_size_3), .B(1), .Y(_28847_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53749_ ( .A(_source_stream_conv2d_16_source_35_pat_count_0), .B(1), .Y(_28848_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53750_ ( .A(_source_stream_conv2d_16_source_35_pat_size_buf_0), .B(1), .Y(_28849_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53751_ ( .A(_source_stream_conv2d_16_source_35_pat_count_1), .B(1), .Y(_28850_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53752_ ( .A(_source_stream_conv2d_16_source_35_pat_size_buf_1), .B(1), .Y(_28851_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53753_ ( .A(_source_stream_conv2d_16_source_35_pat_count_2), .B(1), .Y(_28852_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53754_ ( .A(_source_stream_conv2d_16_source_35_pat_size_buf_2), .B(1), .Y(_28853_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53755_ ( .A(_source_stream_conv2d_16_source_35_pat_count_3), .B(1), .Y(_28854_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53756_ ( .A(_source_stream_conv2d_16_source_35_pat_size_buf_3), .B(1), .Y(_28855_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53757_ ( .A(_source_stream_conv2d_16_source_36_pat_size_0), .B(1), .Y(_28856_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53758_ ( .A(_source_stream_conv2d_16_source_36_pat_size_1), .B(1), .Y(_28857_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53759_ ( .A(_source_stream_conv2d_16_source_36_pat_size_2), .B(1), .Y(_28858_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53760_ ( .A(_source_stream_conv2d_16_source_36_pat_size_3), .B(1), .Y(_28859_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53761_ ( .A(_source_stream_conv2d_16_source_36_pat_count_0), .B(1), .Y(_28860_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53762_ ( .A(_source_stream_conv2d_16_source_36_pat_size_buf_0), .B(1), .Y(_28861_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53763_ ( .A(_source_stream_conv2d_16_source_36_pat_count_1), .B(1), .Y(_28862_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53764_ ( .A(_source_stream_conv2d_16_source_36_pat_size_buf_1), .B(1), .Y(_28863_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53765_ ( .A(_source_stream_conv2d_16_source_36_pat_count_2), .B(1), .Y(_28864_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53766_ ( .A(_source_stream_conv2d_16_source_36_pat_size_buf_2), .B(1), .Y(_28865_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53767_ ( .A(_source_stream_conv2d_16_source_36_pat_count_3), .B(1), .Y(_28866_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53768_ ( .A(_source_stream_conv2d_16_source_36_pat_size_buf_3), .B(1), .Y(_28867_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53769_ ( .A(_stream_conv2d_16_sink_37_sink_offset), .B(_stream_conv2d_16_sink_37_sink_stride), .Y(_28868_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53770_ ( .A(_stream_conv2d_16_sink_37_sink_count), .B(1), .Y(_28869_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(3), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(32) ) _53771_ ( .A(__variable_wdata_777), .B(2'h1), .Y({ _24012_, _24011_, _24009_, _24008_, _24007_, _24006_, _24005_, _24004_, _24003_, _24002_, _24001_, _24000_, _23998_, _23997_, _23996_, _23995_, _23994_, _23993_, _23992_, _23991_, _23990_, _23989_, _24019_, _24018_, _24017_, _24016_, _24015_, _24014_, _24013_, _24010_, _23999_, _23988_ }) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(3), .Y_WIDTH(32) ) _53772_ ( .A(_24399_), .B(__variable_wdata_777), .Y(_28870_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53773_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_0), .B(1), .Y(_28871_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53774_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_1), .B(1), .Y(_28872_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53775_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_2), .B(1), .Y(_28873_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53776_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_3), .B(1), .Y(_28874_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53777_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_0), .B(1), .Y(_28875_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53778_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_buf_0), .B(1), .Y(_28876_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53779_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_1), .B(1), .Y(_28877_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53780_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_buf_1), .B(1), .Y(_28878_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53781_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_2), .B(1), .Y(_28879_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53782_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_buf_2), .B(1), .Y(_28880_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53783_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_3), .B(1), .Y(_28881_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53784_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_buf_3), .B(1), .Y(_28882_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53785_ ( .A(_stream_max_pool_serial_18_sink_3_sink_offset), .B(_stream_max_pool_serial_18_sink_3_sink_stride), .Y(_28883_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53786_ ( .A(_stream_max_pool_serial_18_sink_3_sink_count), .B(1), .Y(_28884_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53787_ ( .A(_source_stream_matmul_29_source_6_pat_size_0), .B(1), .Y(_28885_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53788_ ( .A(_source_stream_matmul_29_source_6_pat_size_1), .B(1), .Y(_28886_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53789_ ( .A(_source_stream_matmul_29_source_6_pat_size_2), .B(1), .Y(_28887_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53790_ ( .A(_source_stream_matmul_29_source_6_pat_size_3), .B(1), .Y(_28888_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53791_ ( .A(_source_stream_matmul_29_source_6_pat_count_0), .B(1), .Y(_28889_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53792_ ( .A(_source_stream_matmul_29_source_6_pat_size_buf_0), .B(1), .Y(_28890_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53793_ ( .A(_source_stream_matmul_29_source_6_pat_count_1), .B(1), .Y(_28891_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53794_ ( .A(_source_stream_matmul_29_source_6_pat_size_buf_1), .B(1), .Y(_28892_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53795_ ( .A(_source_stream_matmul_29_source_6_pat_count_2), .B(1), .Y(_28893_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53796_ ( .A(_source_stream_matmul_29_source_6_pat_size_buf_2), .B(1), .Y(_28894_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53797_ ( .A(_source_stream_matmul_29_source_6_pat_count_3), .B(1), .Y(_28895_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53798_ ( .A(_source_stream_matmul_29_source_6_pat_size_buf_3), .B(1), .Y(_28896_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53799_ ( .A(_source_stream_matmul_29_source_8_pat_size_0), .B(1), .Y(_28897_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53800_ ( .A(_source_stream_matmul_29_source_8_pat_size_1), .B(1), .Y(_28898_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53801_ ( .A(_source_stream_matmul_29_source_8_pat_size_2), .B(1), .Y(_28899_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53802_ ( .A(_source_stream_matmul_29_source_8_pat_size_3), .B(1), .Y(_28900_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53803_ ( .A(_source_stream_matmul_29_source_8_pat_count_0), .B(1), .Y(_28901_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53804_ ( .A(_source_stream_matmul_29_source_8_pat_size_buf_0), .B(1), .Y(_28902_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53805_ ( .A(_source_stream_matmul_29_source_8_pat_count_1), .B(1), .Y(_28903_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53806_ ( .A(_source_stream_matmul_29_source_8_pat_size_buf_1), .B(1), .Y(_28904_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53807_ ( .A(_source_stream_matmul_29_source_8_pat_count_2), .B(1), .Y(_28905_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53808_ ( .A(_source_stream_matmul_29_source_8_pat_size_buf_2), .B(1), .Y(_28906_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53809_ ( .A(_source_stream_matmul_29_source_8_pat_count_3), .B(1), .Y(_28907_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53810_ ( .A(_source_stream_matmul_29_source_8_pat_size_buf_3), .B(1), .Y(_28908_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53811_ ( .A(_source_stream_matmul_29_source_19_pat_size_0), .B(1), .Y(_28909_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53812_ ( .A(_source_stream_matmul_29_source_19_pat_size_1), .B(1), .Y(_28910_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53813_ ( .A(_source_stream_matmul_29_source_19_pat_size_2), .B(1), .Y(_28911_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53814_ ( .A(_source_stream_matmul_29_source_19_pat_size_3), .B(1), .Y(_28912_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53815_ ( .A(_source_stream_matmul_29_source_19_pat_count_0), .B(1), .Y(_28913_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53816_ ( .A(_source_stream_matmul_29_source_19_pat_size_buf_0), .B(1), .Y(_28914_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53817_ ( .A(_source_stream_matmul_29_source_19_pat_count_1), .B(1), .Y(_28915_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53818_ ( .A(_source_stream_matmul_29_source_19_pat_size_buf_1), .B(1), .Y(_28916_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53819_ ( .A(_source_stream_matmul_29_source_19_pat_count_2), .B(1), .Y(_28917_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53820_ ( .A(_source_stream_matmul_29_source_19_pat_size_buf_2), .B(1), .Y(_28918_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53821_ ( .A(_source_stream_matmul_29_source_19_pat_count_3), .B(1), .Y(_28919_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53822_ ( .A(_source_stream_matmul_29_source_19_pat_size_buf_3), .B(1), .Y(_28920_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53823_ ( .A(_source_stream_matmul_29_source_20_pat_size_0), .B(1), .Y(_28921_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53824_ ( .A(_source_stream_matmul_29_source_20_pat_size_1), .B(1), .Y(_28922_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53825_ ( .A(_source_stream_matmul_29_source_20_pat_size_2), .B(1), .Y(_28923_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53826_ ( .A(_source_stream_matmul_29_source_20_pat_size_3), .B(1), .Y(_28924_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53827_ ( .A(_source_stream_matmul_29_source_20_pat_count_0), .B(1), .Y(_28925_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53828_ ( .A(_source_stream_matmul_29_source_20_pat_size_buf_0), .B(1), .Y(_28926_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53829_ ( .A(_source_stream_matmul_29_source_20_pat_count_1), .B(1), .Y(_28927_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53830_ ( .A(_source_stream_matmul_29_source_20_pat_size_buf_1), .B(1), .Y(_28928_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53831_ ( .A(_source_stream_matmul_29_source_20_pat_count_2), .B(1), .Y(_28929_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53832_ ( .A(_source_stream_matmul_29_source_20_pat_size_buf_2), .B(1), .Y(_28930_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53833_ ( .A(_source_stream_matmul_29_source_20_pat_count_3), .B(1), .Y(_28931_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53834_ ( .A(_source_stream_matmul_29_source_20_pat_size_buf_3), .B(1), .Y(_28932_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53835_ ( .A(_stream_matmul_29_sink_21_sink_offset), .B(_stream_matmul_29_sink_21_sink_stride), .Y(_28933_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53836_ ( .A(_stream_matmul_29_sink_21_sink_count), .B(1), .Y(_28934_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(32) ) _53837_ ( .A(conv2d_16_row_select), .B(2), .Y(_28935_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _53838_ ( .A(4096), .B({ 21'h000000, _maxi_read_cur_global_addr[11:0] }), .Y({ _28519_[30:0], _28936_[1:0] }) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _53839_ ( .A(_maxi_read_rest_size), .B({ 2'h0, _28519_[30:0] }), .Y(_28937_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53840_ ( .A(_maxi_read_rest_size), .B(256), .Y(_28938_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(2), .B_SIGNED(0), .B_WIDTH(2), .Y_WIDTH(2) ) _53841_ ( .A(conv2d_16_col_select), .B(2'h2), .Y(_28939_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(32), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _53842_ ( .A(4096), .B({ 21'h000000, _maxi_write_cur_global_addr[11:0] }), .Y({ _28520_[30:0], _28940_[1:0] }) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(33), .Y_WIDTH(33) ) _53843_ ( .A(_maxi_write_rest_size), .B({ 2'h0, _28520_[30:0] }), .Y(_28941_) );
  \$sub  #( .A_SIGNED(0), .A_WIDTH(33), .B_SIGNED(0), .B_WIDTH(32), .Y_WIDTH(33) ) _53844_ ( .A(_maxi_write_rest_size), .B(256), .Y(_28942_) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(4), .Y_WIDTH(12) ) _54133_ ( .A(\__muladd_madd_103.madd._a ), .B(\__muladd_madd_103.madd._b ), .Y(\__muladd_madd_103.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(4), .Y_WIDTH(12) ) _54140_ ( .A(\__muladd_madd_120.madd._a ), .B(\__muladd_madd_120.madd._b ), .Y(\__muladd_madd_120.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(4), .Y_WIDTH(12) ) _54147_ ( .A(\__muladd_madd_137.madd._a ), .B(\__muladd_madd_137.madd._b ), .Y(\__muladd_madd_137.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(4), .Y_WIDTH(12) ) _54154_ ( .A(\__muladd_madd_154.madd._a ), .B(\__muladd_madd_154.madd._b ), .Y(\__muladd_madd_154.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(4), .Y_WIDTH(12) ) _54161_ ( .A(\__muladd_madd_171.madd._a ), .B(\__muladd_madd_171.madd._b ), .Y(\__muladd_madd_171.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(4), .Y_WIDTH(12) ) _54168_ ( .A(\__muladd_madd_188.madd._a ), .B(\__muladd_madd_188.madd._b ), .Y(\__muladd_madd_188.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(4), .Y_WIDTH(12) ) _54175_ ( .A(\__muladd_madd_205.madd._a ), .B(\__muladd_madd_205.madd._b ), .Y(\__muladd_madd_205.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(4), .Y_WIDTH(12) ) _54182_ ( .A(\__muladd_madd_69.madd._a ), .B(\__muladd_madd_69.madd._b ), .Y(\__muladd_madd_69.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(8), .B_SIGNED(1), .B_WIDTH(4), .Y_WIDTH(12) ) _54189_ ( .A(\__muladd_madd_86.madd._a ), .B(\__muladd_madd_86.madd._b ), .Y(\__muladd_madd_86.madd._mul ) );
  \$mul  #( .A_SIGNED(1), .A_WIDTH(32), .B_SIGNED(1), .B_WIDTH(8), .Y_WIDTH(40) ) _54195_ ( .A(\_times_mul_41.mult._a ), .B(\_times_mul_41.mult._b ), .Y(\_times_mul_41.mult._mul ) );
  \$mux  #( .WIDTH(32) ) _45631_ ( .A(_stream_matmul_29_sink_21_sink_fsm_4), .B(0), .S(_06873_), .Y(_24655_) );
  \$mux  #( .WIDTH(32) ) _45632_ ( .A(_24655_), .B(0), .S(_stream_matmul_29_term_sink), .Y({ _13201_, _13200_, _13198_, _13197_, _13196_, _13195_, _13194_, _13193_, _13192_, _13191_, _13190_, _13189_, _13187_, _13186_, _13185_, _13184_, _13183_, _13182_, _13181_, _13180_, _13179_, _13178_, _13208_, _13207_, _13206_, _13205_, _13204_, _13203_, _13202_, _13199_, _13188_, _13177_ }) );
  \$mux  #( .WIDTH(32) ) _45633_ ( .A(_stream_matmul_29_sink_21_sink_fsm_4), .B(1), .S(_06815_), .Y({ _13265_, _13264_, _13262_, _13261_, _13260_, _13259_, _13258_, _13257_, _13256_, _13255_, _13254_, _13253_, _13251_, _13250_, _13249_, _13248_, _13247_, _13246_, _13245_, _13244_, _13243_, _13242_, _13272_, _13271_, _13270_, _13269_, _13268_, _13267_, _13266_, _13263_, _13252_, _13241_ }) );
  \$mux  #( .WIDTH(32) ) _45634_ ( .A(_24656_), .B(0), .S(RST), .Y(_02715_) );
  \$mux  #( .WIDTH(32) ) _45635_ ( .A(_stream_matmul_29_source_20_source_pat_fsm_3), .B(2), .S(_06872_), .Y({ _13329_, _13328_, _13326_, _13325_, _13324_, _13323_, _13322_, _13321_, _13320_, _13319_, _13318_, _13317_, _13315_, _13314_, _13313_, _13312_, _13311_, _13310_, _13309_, _13308_, _13307_, _13306_, _13336_, _13335_, _13334_, _13333_, _13332_, _13331_, _13330_, _13327_, _13316_, _13305_ }) );
  \$mux  #( .WIDTH(32) ) _45636_ ( .A(_stream_matmul_29_source_20_source_pat_fsm_3), .B(1), .S(_06810_), .Y({ _13361_, _13360_, _13358_, _13357_, _13356_, _13355_, _13354_, _13353_, _13352_, _13351_, _13350_, _13349_, _13347_, _13346_, _13345_, _13344_, _13343_, _13342_, _13341_, _13340_, _13339_, _13338_, _13368_, _13367_, _13366_, _13365_, _13364_, _13363_, _13362_, _13359_, _13348_, _13337_ }) );
  \$mux  #( .WIDTH(32) ) _45637_ ( .A(_24657_), .B(0), .S(RST), .Y(_02744_) );
  \$mux  #( .WIDTH(32) ) _45638_ ( .A(_stream_matmul_29_source_19_source_pat_fsm_2), .B(2), .S(_06871_), .Y({ _13425_, _13424_, _13422_, _13421_, _13420_, _13419_, _13418_, _13417_, _13416_, _13415_, _13414_, _13413_, _13411_, _13410_, _13409_, _13408_, _13407_, _13406_, _13405_, _13404_, _13403_, _13402_, _13432_, _13431_, _13430_, _13429_, _13428_, _13427_, _13426_, _13423_, _13412_, _13401_ }) );
  \$mux  #( .WIDTH(32) ) _45639_ ( .A(_stream_matmul_29_source_19_source_pat_fsm_2), .B(1), .S(_06805_), .Y({ _13457_, _13456_, _13454_, _13453_, _13452_, _13451_, _13450_, _13449_, _13448_, _13447_, _13446_, _13445_, _13443_, _13442_, _13441_, _13440_, _13439_, _13438_, _13437_, _13436_, _13435_, _13434_, _13464_, _13463_, _13462_, _13461_, _13460_, _13459_, _13458_, _13455_, _13444_, _13433_ }) );
  \$mux  #( .WIDTH(32) ) _45640_ ( .A(_24658_), .B(0), .S(RST), .Y(_02735_) );
  \$mux  #( .WIDTH(32) ) _45641_ ( .A(_stream_matmul_29_source_8_source_pat_fsm_1), .B(2), .S(_06870_), .Y({ _13521_, _13520_, _13518_, _13517_, _13516_, _13515_, _13514_, _13513_, _13512_, _13511_, _13510_, _13509_, _13507_, _13506_, _13505_, _13504_, _13503_, _13502_, _13501_, _13500_, _13499_, _13498_, _13528_, _13527_, _13526_, _13525_, _13524_, _13523_, _13522_, _13519_, _13508_, _13497_ }) );
  \$mux  #( .WIDTH(32) ) _45642_ ( .A(_stream_matmul_29_source_8_source_pat_fsm_1), .B(1), .S(_06800_), .Y({ _13553_, _13552_, _13550_, _13549_, _13548_, _13547_, _13546_, _13545_, _13544_, _13543_, _13542_, _13541_, _13539_, _13538_, _13537_, _13536_, _13535_, _13534_, _13533_, _13532_, _13531_, _13530_, _13560_, _13559_, _13558_, _13557_, _13556_, _13555_, _13554_, _13551_, _13540_, _13529_ }) );
  \$mux  #( .WIDTH(32) ) _45643_ ( .A(_24659_), .B(0), .S(RST), .Y(_02762_) );
  \$mux  #( .WIDTH(32) ) _45644_ ( .A(_stream_matmul_29_source_6_source_pat_fsm_0), .B(2), .S(_06869_), .Y({ _13617_, _13616_, _13614_, _13613_, _13612_, _13611_, _13610_, _13609_, _13608_, _13607_, _13606_, _13605_, _13603_, _13602_, _13601_, _13600_, _13599_, _13598_, _13597_, _13596_, _13595_, _13594_, _13624_, _13623_, _13622_, _13621_, _13620_, _13619_, _13618_, _13615_, _13604_, _13593_ }) );
  \$mux  #( .WIDTH(32) ) _45645_ ( .A(_stream_matmul_29_source_6_source_pat_fsm_0), .B(1), .S(_06795_), .Y({ _13649_, _13648_, _13646_, _13645_, _13644_, _13643_, _13642_, _13641_, _13640_, _13639_, _13638_, _13637_, _13635_, _13634_, _13633_, _13632_, _13631_, _13630_, _13629_, _13628_, _13627_, _13626_, _13656_, _13655_, _13654_, _13653_, _13652_, _13651_, _13650_, _13647_, _13636_, _13625_ }) );
  \$mux  #( .WIDTH(32) ) _45646_ ( .A(_24660_), .B(0), .S(RST), .Y(_02753_) );
  \$mux  #( .WIDTH(1) ) _45647_ ( .A(matmul_29_stream_pad_mask_0_0), .B(matmul_29_stream_pad_masks), .S(_05916_), .Y(_24661_) );
  \$mux  #( .WIDTH(1) ) _45648_ ( .A(_24661_), .B(1'h0), .S(RST), .Y(_03330_) );
  \$mux  #( .WIDTH(32) ) _45649_ ( .A(matmul_29_och_count), .B(matmul_29_och_count_buf), .S(_05920_), .Y(_24662_) );
  \$mux  #( .WIDTH(32) ) _45650_ ( .A(_24662_), .B(0), .S(RST), .Y(_03303_) );
  \$mux  #( .WIDTH(1) ) _45651_ ( .A(matmul_29_row_select), .B(matmul_29_row_select_buf), .S(_05920_), .Y(_24663_) );
  \$mux  #( .WIDTH(1) ) _45652_ ( .A(_24663_), .B(1'h0), .S(RST), .Y(_03323_) );
  \$mux  #( .WIDTH(32) ) _45653_ ( .A(matmul_29_row_count), .B(matmul_29_row_count_buf), .S(_05920_), .Y(_24664_) );
  \$mux  #( .WIDTH(32) ) _45654_ ( .A(_24664_), .B(0), .S(RST), .Y(_03321_) );
  \$mux  #( .WIDTH(32) ) _45655_ ( .A(matmul_29_out_page_comp_offset), .B(matmul_29_out_page_comp_offset_buf), .S(_05920_), .Y(_24665_) );
  \$mux  #( .WIDTH(32) ) _45656_ ( .A(_24665_), .B(0), .S(RST), .Y(_03312_) );
  \$mux  #( .WIDTH(32) ) _45657_ ( .A(matmul_29_act_page_comp_offset_0), .B(matmul_29_act_page_comp_offset_buf_0), .S(_05920_), .Y(_24666_) );
  \$mux  #( .WIDTH(32) ) _45658_ ( .A(_24666_), .B(0), .S(RST), .Y(_03283_) );
  \$mux  #( .WIDTH(32) ) _45659_ ( .A(matmul_29_filter_page_comp_offset), .B(matmul_29_filter_page_comp_offset_buf), .S(_05920_), .Y(_24667_) );
  \$mux  #( .WIDTH(32) ) _45660_ ( .A(_24667_), .B(0), .S(RST), .Y(_03297_) );
  \$mux  #( .WIDTH(32) ) _45661_ ( .A(5), .B(matmul_29_comp_fsm), .S(_stream_matmul_29_source_busy), .Y({ _13713_, _13712_, _13710_, _13709_, _13708_, _13707_, _13706_, _13705_, _13704_, _13703_, _13702_, _13701_, _13699_, _13698_, _13697_, _13696_, _13695_, _13694_, _13693_, _13692_, _13691_, _13690_, _13720_, _13719_, _13718_, _13717_, _13716_, _13715_, _13714_, _13711_, _13700_, _13689_ }) );
  \$mux  #( .WIDTH(32) ) _45662_ ( .A(matmul_29_comp_fsm), .B(1), .S(_06868_), .Y({ _13745_, _13744_, _13742_, _13741_, _13740_, _13739_, _13738_, _13737_, _13736_, _13735_, _13734_, _13733_, _13731_, _13730_, _13729_, _13728_, _13727_, _13726_, _13725_, _13724_, _13723_, _13722_, _13752_, _13751_, _13750_, _13749_, _13748_, _13747_, _13746_, _13743_, _13732_, _13721_ }) );
  \$mux  #( .WIDTH(32) ) _45663_ ( .A(_24668_), .B(0), .S(RST), .Y(_03292_) );
  \$mux  #( .WIDTH(32) ) _45664_ ( .A(_24669_), .B(0), .S(RST), .Y(_03329_) );
  \$mux  #( .WIDTH(32) ) _45665_ ( .A(_24670_), .B(0), .S(RST), .Y(_03328_) );
  \$mux  #( .WIDTH(1) ) _45666_ ( .A(_24671_), .B(1'h0), .S(RST), .Y(_03291_) );
  \$mux  #( .WIDTH(32) ) _45667_ ( .A(_24672_), .B(0), .S(RST), .Y(_03290_) );
  \$mux  #( .WIDTH(32) ) _45668_ ( .A(matmul_29_sync_comp_count), .B(_24478_), .S(_stream_matmul_29_end_flag), .Y(_24673_) );
  \$mux  #( .WIDTH(32) ) _45669_ ( .A(0), .B(_24673_), .S(_05930_), .Y(_24674_) );
  \$mux  #( .WIDTH(32) ) _45670_ ( .A(_24674_), .B(0), .S(RST), .Y(_03331_) );
  \$mux  #( .WIDTH(32) ) _45671_ ( .A({ 27'h0000000, cparam_matmul_29_out_write_size }), .B(matmul_29_next_stream_num_ops), .S(_05920_), .Y(_24675_) );
  \$mux  #( .WIDTH(32) ) _45672_ ( .A(_24675_), .B(0), .S(RST), .Y(_03300_) );
  \$mux  #( .WIDTH(1) ) _45673_ ( .A(1'h1), .B(_control_matmul_29_cond_32_4_1), .S(_05925_), .Y(_24676_) );
  \$mux  #( .WIDTH(1) ) _45674_ ( .A(_24676_), .B(1'h0), .S(RST), .Y(_01573_) );
  \$mux  #( .WIDTH(1) ) _45675_ ( .A(axim_flag_1308), .B(1'h0), .S(_control_matmul_29_cond_32_4_1), .Y(_24677_) );
  \$mux  #( .WIDTH(1) ) _45676_ ( .A(_24677_), .B(axim_flag_1308), .S(_05918_), .Y(_24678_) );
  \$mux  #( .WIDTH(1) ) _45677_ ( .A(1'h1), .B(_24678_), .S(_05925_), .Y(_24679_) );
  \$mux  #( .WIDTH(1) ) _45678_ ( .A(_24679_), .B(1'h0), .S(RST), .Y(_03198_) );
  \$mux  #( .WIDTH(1) ) _45679_ ( .A(1'h1), .B(_control_matmul_29_cond_22_3_1), .S(_05926_), .Y(_24680_) );
  \$mux  #( .WIDTH(1) ) _45680_ ( .A(_24680_), .B(1'h0), .S(RST), .Y(_01572_) );
  \$mux  #( .WIDTH(1) ) _45681_ ( .A(axim_flag_1152), .B(1'h0), .S(_control_matmul_29_cond_22_3_1), .Y(_24681_) );
  \$mux  #( .WIDTH(1) ) _45682_ ( .A(_24681_), .B(axim_flag_1152), .S(_05919_), .Y(_24682_) );
  \$mux  #( .WIDTH(1) ) _45683_ ( .A(1'h1), .B(_24682_), .S(_05926_), .Y(_24683_) );
  \$mux  #( .WIDTH(1) ) _45684_ ( .A(_24683_), .B(1'h0), .S(RST), .Y(_03197_) );
  \$mux  #( .WIDTH(1) ) _45685_ ( .A(1'h1), .B(_control_matmul_29_cond_14_2_1), .S(_05927_), .Y(_24684_) );
  \$mux  #( .WIDTH(1) ) _45686_ ( .A(_24684_), .B(1'h0), .S(RST), .Y(_01571_) );
  \$mux  #( .WIDTH(1) ) _45687_ ( .A(axim_flag_1133), .B(1'h0), .S(_control_matmul_29_cond_14_2_1), .Y(_24685_) );
  \$mux  #( .WIDTH(1) ) _45688_ ( .A(_24685_), .B(axim_flag_1133), .S(_05921_), .Y(_24686_) );
  \$mux  #( .WIDTH(1) ) _45689_ ( .A(1'h1), .B(_24686_), .S(_05927_), .Y(_24687_) );
  \$mux  #( .WIDTH(1) ) _45690_ ( .A(_24687_), .B(1'h0), .S(RST), .Y(_03196_) );
  \$mux  #( .WIDTH(1) ) _45691_ ( .A(1'h1), .B(_control_matmul_29_cond_8_1_1), .S(_05928_), .Y(_24688_) );
  \$mux  #( .WIDTH(1) ) _45692_ ( .A(_24688_), .B(1'h0), .S(RST), .Y(_01575_) );
  \$mux  #( .WIDTH(1) ) _45693_ ( .A(axim_flag_1132), .B(1'h0), .S(_control_matmul_29_cond_8_1_1), .Y(_24689_) );
  \$mux  #( .WIDTH(1) ) _45694_ ( .A(_24689_), .B(axim_flag_1132), .S(_05922_), .Y(_24690_) );
  \$mux  #( .WIDTH(1) ) _45695_ ( .A(1'h1), .B(_24690_), .S(_05928_), .Y(_24691_) );
  \$mux  #( .WIDTH(1) ) _45696_ ( .A(_24691_), .B(1'h0), .S(RST), .Y(_03195_) );
  \$mux  #( .WIDTH(1) ) _45697_ ( .A(1'h1), .B(_control_matmul_29_cond_3_0_1), .S(_05931_), .Y(_24692_) );
  \$mux  #( .WIDTH(1) ) _45698_ ( .A(_24692_), .B(1'h0), .S(RST), .Y(_01574_) );
  \$mux  #( .WIDTH(32) ) _45699_ ( .A(control_matmul_29), .B(0), .S(RST), .Y(_01584_) );
  \$mux  #( .WIDTH(1) ) _45700_ ( .A(axim_flag_1121), .B(1'h0), .S(_control_matmul_29_cond_3_0_1), .Y(_24693_) );
  \$mux  #( .WIDTH(1) ) _45701_ ( .A(_24693_), .B(axim_flag_1121), .S(_05923_), .Y(_24694_) );
  \$mux  #( .WIDTH(1) ) _45702_ ( .A(1'h1), .B(_24694_), .S(_05931_), .Y(_24695_) );
  \$mux  #( .WIDTH(1) ) _45703_ ( .A(_24695_), .B(1'h0), .S(RST), .Y(_03194_) );
  \$mux  #( .WIDTH(1) ) _45704_ ( .A(matmul_29_skip_write_out), .B(1'h0), .S(_06866_), .Y(_13753_) );
  \$mux  #( .WIDTH(1) ) _45705_ ( .A(_24696_), .B(1'h1), .S(RST), .Y(_03327_) );
  \$mux  #( .WIDTH(1) ) _45706_ ( .A(matmul_29_skip_comp), .B(1'h1), .S(_06146_), .Y(_13756_) );
  \$mux  #( .WIDTH(1) ) _45707_ ( .A(_24697_), .B(1'h0), .S(RST), .Y(_03324_) );
  \$mux  #( .WIDTH(1) ) _45708_ ( .A(_24698_), .B(1'h0), .S(RST), .Y(_03325_) );
  \$mux  #( .WIDTH(1) ) _45709_ ( .A(matmul_29_skip_read_filter), .B(1'h1), .S(_06146_), .Y(_13758_) );
  \$mux  #( .WIDTH(1) ) _45710_ ( .A(_24699_), .B(1'h0), .S(RST), .Y(_03326_) );
  \$mux  #( .WIDTH(32) ) _45711_ ( .A(0), .B(matmul_29_out_laddr_offset), .S(matmul_29_skip_write_out), .Y({ _13784_, _13783_, _13781_, _13780_, _13779_, _13778_, _13777_, _13776_, _13775_, _13774_, _13773_, _13772_, _13770_, _13769_, _13768_, _13767_, _13766_, _13765_, _13764_, _13763_, _13762_, _13761_, _13791_, _13790_, _13789_, _13788_, _13787_, _13786_, _13785_, _13782_, _13771_, _13760_ }) );
  \$mux  #( .WIDTH(32) ) _45712_ ( .A(_24472_), .B(matmul_29_out_laddr_offset), .S(_05724_), .Y({ _13816_, _13815_, _13813_, _13812_, _13811_, _13810_, _13809_, _13808_, _13807_, _13806_, _13805_, _13804_, _13802_, _13801_, _13800_, _13799_, _13798_, _13797_, _13796_, _13795_, _13794_, _13793_, _13823_, _13822_, _13821_, _13820_, _13819_, _13818_, _13817_, _13814_, _13803_, _13792_ }) );
  \$mux  #( .WIDTH(32) ) _45713_ ( .A(_24700_), .B(0), .S(RST), .Y(_03309_) );
  \$mux  #( .WIDTH(32) ) _45714_ ( .A(0), .B(1024), .S(matmul_29_out_page), .Y({ _13848_, _13847_, _13845_, _13844_, _13843_, _13842_, _13841_, _13840_, _13839_, _13838_, _13837_, _13836_, _13834_, _13833_, _13832_, _13831_, _13830_, _13829_, _13828_, _13827_, _13826_, _13825_, _13855_, _13854_, _13853_, _13852_, _13851_, _13850_, _13849_, _13846_, _13835_, _13824_ }) );
  \$mux  #( .WIDTH(32) ) _45715_ ( .A(_24701_), .B(0), .S(RST), .Y(_03313_) );
  \$mux  #( .WIDTH(32) ) _45716_ ( .A(1024), .B(0), .S(matmul_29_out_page), .Y({ _13912_, _13911_, _13909_, _13908_, _13907_, _13906_, _13905_, _13904_, _13903_, _13902_, _13901_, _13900_, _13898_, _13897_, _13896_, _13895_, _13894_, _13893_, _13892_, _13891_, _13890_, _13889_, _13919_, _13918_, _13917_, _13916_, _13915_, _13914_, _13913_, _13910_, _13899_, _13888_ }) );
  \$mux  #( .WIDTH(32) ) _45717_ ( .A(_24702_), .B(0), .S(RST), .Y(_03311_) );
  \$mux  #( .WIDTH(1) ) _45718_ ( .A(1'h1), .B(1'h0), .S(matmul_29_out_page), .Y(_13952_) );
  \$mux  #( .WIDTH(1) ) _45719_ ( .A(_24703_), .B(1'h0), .S(RST), .Y(_03310_) );
  \$mux  #( .WIDTH(32) ) _45720_ ( .A(0), .B(_24476_), .S(_24028_), .Y({ _13978_, _13977_, _13975_, _13974_, _13973_, _13972_, _13971_, _13970_, _13969_, _13968_, _13967_, _13966_, _13964_, _13963_, _13962_, _13961_, _13960_, _13959_, _13958_, _13957_, _13956_, _13955_, _13985_, _13984_, _13983_, _13982_, _13981_, _13980_, _13979_, _13976_, _13965_, _13954_ }) );
  \$mux  #( .WIDTH(32) ) _45721_ ( .A(_24704_), .B(0), .S(RST), .Y(_03298_) );
  \$mux  #( .WIDTH(32) ) _45722_ ( .A(0), .B(_24475_), .S(_24028_), .Y({ _14042_, _14041_, _14039_, _14038_, _14037_, _14036_, _14035_, _14034_, _14033_, _14032_, _14031_, _14030_, _14028_, _14027_, _14026_, _14025_, _14024_, _14023_, _14022_, _14021_, _14020_, _14019_, _14049_, _14048_, _14047_, _14046_, _14045_, _14044_, _14043_, _14040_, _14029_, _14018_ }) );
  \$mux  #( .WIDTH(32) ) _45723_ ( .A(_24705_), .B(0), .S(RST), .Y(_03296_) );
  \$mux  #( .WIDTH(32) ) _45724_ ( .A(_24706_), .B(0), .S(RST), .Y(_03284_) );
  \$mux  #( .WIDTH(32) ) _45725_ ( .A(_24707_), .B(0), .S(RST), .Y(_03282_) );
  \$mux  #( .WIDTH(1) ) _45726_ ( .A(matmul_29_prev_row_select), .B(1'h0), .S(_05515_), .Y(_24708_) );
  \$mux  #( .WIDTH(1) ) _45727_ ( .A(_24708_), .B(1'h0), .S(RST), .Y(_03319_) );
  \$mux  #( .WIDTH(32) ) _45728_ ( .A(_24709_), .B(0), .S(RST), .Y(_03317_) );
  \$mux  #( .WIDTH(32) ) _45729_ ( .A(_24710_), .B(0), .S(RST), .Y(_03316_) );
  \$mux  #( .WIDTH(32) ) _45730_ ( .A(_24711_), .B(0), .S(RST), .Y(_03318_) );
  \$mux  #( .WIDTH(32) ) _45731_ ( .A(0), .B(matmul_29_out_ram_select), .S(matmul_29_skip_write_out), .Y({ _14202_, _14201_, _14199_, _14198_, _14197_, _14196_, _14195_, _14194_, _14193_, _14192_, _14191_, _14190_, _14188_, _14187_, _14186_, _14185_, _14184_, _14183_, _14182_, _14181_, _14180_, _14179_, _14209_, _14208_, _14207_, _14206_, _14205_, _14204_, _14203_, _14200_, _14189_, _14178_ }) );
  \$mux  #( .WIDTH(32) ) _45732_ ( .A(0), .B(_24474_), .S(_05724_), .Y({ _14234_, _14233_, _14231_, _14230_, _14229_, _14228_, _14227_, _14226_, _14225_, _14224_, _14223_, _14222_, _14220_, _14219_, _14218_, _14217_, _14216_, _14215_, _14214_, _14213_, _14212_, _14211_, _14241_, _14240_, _14239_, _14238_, _14237_, _14236_, _14235_, _14232_, _14221_, _14210_ }) );
  \$mux  #( .WIDTH(32) ) _45733_ ( .A(_24712_), .B(0), .S(RST), .Y(_03314_) );
  \$mux  #( .WIDTH(32) ) _45734_ ( .A(0), .B(matmul_29_out_row_count), .S(matmul_29_skip_write_out), .Y({ _14266_, _14265_, _14263_, _14262_, _14261_, _14260_, _14259_, _14258_, _14257_, _14256_, _14255_, _14254_, _14252_, _14251_, _14250_, _14249_, _14248_, _14247_, _14246_, _14245_, _14244_, _14243_, _14273_, _14272_, _14271_, _14270_, _14269_, _14268_, _14267_, _14264_, _14253_, _14242_ }) );
  \$mux  #( .WIDTH(32) ) _45735_ ( .A(_24713_), .B(0), .S(RST), .Y(_03315_) );
  \$mux  #( .WIDTH(1) ) _45736_ ( .A(matmul_29_row_select), .B(1'h0), .S(_05515_), .Y(_24714_) );
  \$mux  #( .WIDTH(1) ) _45737_ ( .A(_24714_), .B(1'h0), .S(RST), .Y(_03322_) );
  \$mux  #( .WIDTH(32) ) _45738_ ( .A(_24715_), .B(0), .S(RST), .Y(_03302_) );
  \$mux  #( .WIDTH(32) ) _45739_ ( .A(_24716_), .B(0), .S(RST), .Y(_03289_) );
  \$mux  #( .WIDTH(32) ) _45740_ ( .A(_24717_), .B(0), .S(RST), .Y(_03320_) );
  \$mux  #( .WIDTH(32) ) _45741_ ( .A(matmul_29_next_out_write_size), .B({ 27'h0000000, cparam_matmul_29_out_write_size }), .S(_05515_), .Y(_24718_) );
  \$mux  #( .WIDTH(32) ) _45742_ ( .A(_24718_), .B(0), .S(RST), .Y(_03299_) );
  \$mux  #( .WIDTH(32) ) _45743_ ( .A(_24719_), .B(0), .S(RST), .Y(_03332_) );
  \$mux  #( .WIDTH(1) ) _45744_ ( .A(matmul_29_dma_flag_0), .B(1'h1), .S(_05515_), .Y(_24720_) );
  \$mux  #( .WIDTH(1) ) _45745_ ( .A(_24720_), .B(1'h0), .S(RST), .Y(_03294_) );
  \$mux  #( .WIDTH(32) ) _45746_ ( .A(_24477_), .B(matmul_29_out_base_offset_och), .S(matmul_29_skip_write_out), .Y({ _14426_, _14425_, _14423_, _14422_, _14421_, _14420_, _14419_, _14418_, _14417_, _14416_, _14415_, _14414_, _14412_, _14411_, _14410_, _14409_, _14408_, _14407_, _14406_, _14405_, _14404_, _14403_, _14433_, _14432_, _14431_, _14430_, _14429_, _14428_, _14427_, _14424_, _14413_, _14402_ }) );
  \$mux  #( .WIDTH(32) ) _45747_ ( .A(_24721_), .B(0), .S(RST), .Y(_03306_) );
  \$mux  #( .WIDTH(32) ) _45748_ ( .A(0), .B(matmul_29_out_base_offset_bat), .S(matmul_29_skip_write_out), .Y({ _14490_, _14489_, _14487_, _14486_, _14485_, _14484_, _14483_, _14482_, _14481_, _14480_, _14479_, _14478_, _14476_, _14475_, _14474_, _14473_, _14472_, _14471_, _14470_, _14469_, _14468_, _14467_, _14497_, _14496_, _14495_, _14494_, _14493_, _14492_, _14491_, _14488_, _14477_, _14466_ }) );
  \$mux  #( .WIDTH(32) ) _45749_ ( .A(_24722_), .B(0), .S(RST), .Y(_03304_) );
  \$mux  #( .WIDTH(32) ) _45750_ ( .A(0), .B(matmul_29_out_base_offset_row), .S(matmul_29_skip_write_out), .Y({ _14554_, _14553_, _14551_, _14550_, _14549_, _14548_, _14547_, _14546_, _14545_, _14544_, _14543_, _14542_, _14540_, _14539_, _14538_, _14537_, _14536_, _14535_, _14534_, _14533_, _14532_, _14531_, _14561_, _14560_, _14559_, _14558_, _14557_, _14556_, _14555_, _14552_, _14541_, _14530_ }) );
  \$mux  #( .WIDTH(32) ) _45751_ ( .A(_24723_), .B(0), .S(RST), .Y(_03307_) );
  \$mux  #( .WIDTH(32) ) _45752_ ( .A(0), .B(matmul_29_out_base_offset_col), .S(matmul_29_skip_write_out), .Y({ _14618_, _14617_, _14615_, _14614_, _14613_, _14612_, _14611_, _14610_, _14609_, _14608_, _14607_, _14606_, _14604_, _14603_, _14602_, _14601_, _14600_, _14599_, _14598_, _14597_, _14596_, _14595_, _14625_, _14624_, _14623_, _14622_, _14621_, _14620_, _14619_, _14616_, _14605_, _14594_ }) );
  \$mux  #( .WIDTH(32) ) _45753_ ( .A(_24473_), .B(matmul_29_out_base_offset_col), .S(cparam_matmul_29_keep_filter), .Y({ _14650_, _14649_, _14647_, _14646_, _14645_, _14644_, _14643_, _14642_, _14641_, _14640_, _14639_, _14638_, _14636_, _14635_, _14634_, _14633_, _14632_, _14631_, _14630_, _14629_, _14628_, _14627_, _14657_, _14656_, _14655_, _14654_, _14653_, _14652_, _14651_, _14648_, _14637_, _14626_ }) );
  \$mux  #( .WIDTH(32) ) _45754_ ( .A(_24724_), .B(0), .S(RST), .Y(_03305_) );
  \$mux  #( .WIDTH(32) ) _45755_ ( .A(0), .B(matmul_29_out_base_offset_val), .S(_05929_), .Y(_24725_) );
  \$mux  #( .WIDTH(32) ) _45756_ ( .A(_24725_), .B(0), .S(RST), .Y(_03308_) );
  \$mux  #( .WIDTH(32) ) _45757_ ( .A(_24726_), .B(0), .S(RST), .Y(_03295_) );
  \$mux  #( .WIDTH(32) ) _45758_ ( .A(_24727_), .B(0), .S(RST), .Y(_03280_) );
  \$mux  #( .WIDTH(32) ) _45759_ ( .A(_24728_), .B(0), .S(RST), .Y(_03281_) );
  \$mux  #( .WIDTH(32) ) _45760_ ( .A(0), .B(control_matmul_29), .S(_05728_), .Y(_24729_) );
  \$mux  #( .WIDTH(32) ) _45761_ ( .A(0), .B(_24729_), .S(_06025_), .Y(_24730_) );
  \$mux  #( .WIDTH(32) ) _45762_ ( .A(0), .B(_24730_), .S(_06023_), .Y({ _14714_, _14713_, _14711_, _14710_, _14709_, _14708_, _14707_, _14706_, _14705_, _14704_, _14703_, _14702_, _14700_, _14699_, _14698_, _14697_, _14696_, _14695_, _14694_, _14693_, _14692_, _14691_, _14721_, _14720_, _14719_, _14718_, _14717_, _14716_, _14715_, _14712_, _14701_, _14690_ }) );
  \$mux  #( .WIDTH(32) ) _45763_ ( .A(control_matmul_29), .B(39), .S(_maxi_write_idle), .Y({ _14778_, _14777_, _14775_, _14774_, _14773_, _14772_, _14771_, _14770_, _14769_, _14768_, _14767_, _14766_, _14764_, _14763_, _14762_, _14761_, _14760_, _14759_, _14758_, _14757_, _14756_, _14755_, _14785_, _14784_, _14783_, _14782_, _14781_, _14780_, _14779_, _14776_, _14765_, _14754_ }) );
  \$mux  #( .WIDTH(32) ) _45764_ ( .A(13), .B(38), .S(_06867_), .Y({ _14810_, _14809_, _14807_, _14806_, _14805_, _14804_, _14803_, _14802_, _14801_, _14800_, _14799_, _14798_, _14796_, _14795_, _14794_, _14793_, _14792_, _14791_, _14790_, _14789_, _14788_, _14787_, _14817_, _14816_, _14815_, _14814_, _14813_, _14812_, _14811_, _14808_, _14797_, _14786_ }) );
  \$mux  #( .WIDTH(32) ) _45765_ ( .A(control_matmul_29), .B(32), .S(_maxi_write_idle), .Y({ _14842_, _14841_, _14839_, _14838_, _14837_, _14836_, _14835_, _14834_, _14833_, _14832_, _14831_, _14830_, _14828_, _14827_, _14826_, _14825_, _14824_, _14823_, _14822_, _14821_, _14820_, _14819_, _14849_, _14848_, _14847_, _14846_, _14845_, _14844_, _14843_, _14840_, _14829_, _14818_ }) );
  \$mux  #( .WIDTH(32) ) _45766_ ( .A(31), .B(35), .S(matmul_29_dma_out_mask_0), .Y({ _14874_, _14873_, _14871_, _14870_, _14869_, _14868_, _14867_, _14866_, _14865_, _14864_, _14863_, _14862_, _14860_, _14859_, _14858_, _14857_, _14856_, _14855_, _14854_, _14853_, _14852_, _14851_, _14881_, _14880_, _14879_, _14878_, _14877_, _14876_, _14875_, _14872_, _14861_, _14850_ }) );
  \$mux  #( .WIDTH(32) ) _45767_ ( .A(control_matmul_29), .B(30), .S(_06162_), .Y(_24732_) );
  \$mux  #( .WIDTH(32) ) _45768_ ( .A(_24732_), .B(37), .S(matmul_29_skip_write_out), .Y({ _14906_, _14905_, _14903_, _14902_, _14901_, _14900_, _14899_, _14898_, _14897_, _14896_, _14895_, _14894_, _14892_, _14891_, _14890_, _14889_, _14888_, _14887_, _14886_, _14885_, _14884_, _14883_, _14913_, _14912_, _14911_, _14910_, _14909_, _14908_, _14907_, _14904_, _14893_, _14882_ }) );
  \$mux  #( .WIDTH(32) ) _45769_ ( .A(29), .B(control_matmul_29), .S(_05725_), .Y({ _14938_, _14937_, _14935_, _14934_, _14933_, _14932_, _14931_, _14930_, _14929_, _14928_, _14927_, _14926_, _14924_, _14923_, _14922_, _14921_, _14920_, _14919_, _14918_, _14917_, _14916_, _14915_, _14945_, _14944_, _14943_, _14942_, _14941_, _14940_, _14939_, _14936_, _14925_, _14914_ }) );
  \$mux  #( .WIDTH(32) ) _45770_ ( .A(control_matmul_29), .B(26), .S(_maxi_read_idle), .Y({ _14970_, _14969_, _14967_, _14966_, _14965_, _14964_, _14963_, _14962_, _14961_, _14960_, _14959_, _14958_, _14956_, _14955_, _14954_, _14953_, _14952_, _14951_, _14950_, _14949_, _14948_, _14947_, _14977_, _14976_, _14975_, _14974_, _14973_, _14972_, _14971_, _14968_, _14957_, _14946_ }) );
  \$mux  #( .WIDTH(32) ) _45771_ ( .A(control_matmul_29), .B(22), .S(_maxi_read_idle), .Y({ _15002_, _15001_, _14999_, _14998_, _14997_, _14996_, _14995_, _14994_, _14993_, _14992_, _14991_, _14990_, _14988_, _14987_, _14986_, _14985_, _14984_, _14983_, _14982_, _14981_, _14980_, _14979_, _15009_, _15008_, _15007_, _15006_, _15005_, _15004_, _15003_, _15000_, _14989_, _14978_ }) );
  \$mux  #( .WIDTH(32) ) _45772_ ( .A(21), .B(26), .S(_06882_), .Y(_24733_) );
  \$mux  #( .WIDTH(32) ) _45773_ ( .A(_24733_), .B(27), .S(matmul_29_skip_read_act), .Y({ _15034_, _15033_, _15031_, _15030_, _15029_, _15028_, _15027_, _15026_, _15025_, _15024_, _15023_, _15022_, _15020_, _15019_, _15018_, _15017_, _15016_, _15015_, _15014_, _15013_, _15012_, _15011_, _15041_, _15040_, _15039_, _15038_, _15037_, _15036_, _15035_, _15032_, _15021_, _15010_ }) );
  \$mux  #( .WIDTH(32) ) _45774_ ( .A(control_matmul_29), .B(18), .S(_maxi_read_idle), .Y({ _15066_, _15065_, _15063_, _15062_, _15061_, _15060_, _15059_, _15058_, _15057_, _15056_, _15055_, _15054_, _15052_, _15051_, _15050_, _15049_, _15048_, _15047_, _15046_, _15045_, _15044_, _15043_, _15073_, _15072_, _15071_, _15070_, _15069_, _15068_, _15067_, _15064_, _15053_, _15042_ }) );
  \$mux  #( .WIDTH(32) ) _45775_ ( .A(control_matmul_29), .B(14), .S(_maxi_read_idle), .Y(_24734_) );
  \$mux  #( .WIDTH(32) ) _45776_ ( .A(_24734_), .B(19), .S(matmul_29_skip_read_filter), .Y({ _15098_, _15097_, _15095_, _15094_, _15093_, _15092_, _15091_, _15090_, _15089_, _15088_, _15087_, _15086_, _15084_, _15083_, _15082_, _15081_, _15080_, _15079_, _15078_, _15077_, _15076_, _15075_, _15105_, _15104_, _15103_, _15102_, _15101_, _15100_, _15099_, _15096_, _15085_, _15074_ }) );
  \$mux  #( .WIDTH(32) ) _45777_ ( .A(control_matmul_29), .B(12), .S(_maxi_read_idle), .Y({ _15130_, _15129_, _15127_, _15126_, _15125_, _15124_, _15123_, _15122_, _15121_, _15120_, _15119_, _15118_, _15116_, _15115_, _15114_, _15113_, _15112_, _15111_, _15110_, _15109_, _15108_, _15107_, _15137_, _15136_, _15135_, _15134_, _15133_, _15132_, _15131_, _15128_, _15117_, _15106_ }) );
  \$mux  #( .WIDTH(32) ) _45778_ ( .A(control_matmul_29), .B(8), .S(_maxi_read_idle), .Y({ _15162_, _15161_, _15159_, _15158_, _15157_, _15156_, _15155_, _15154_, _15153_, _15152_, _15151_, _15150_, _15148_, _15147_, _15146_, _15145_, _15144_, _15143_, _15142_, _15141_, _15140_, _15139_, _15169_, _15168_, _15167_, _15166_, _15165_, _15164_, _15163_, _15160_, _15149_, _15138_ }) );
  \$mux  #( .WIDTH(32) ) _45779_ ( .A(control_matmul_29), .B(7), .S(_maxi_read_idle), .Y({ _15194_, _15193_, _15191_, _15190_, _15189_, _15188_, _15187_, _15186_, _15185_, _15184_, _15183_, _15182_, _15180_, _15179_, _15178_, _15177_, _15176_, _15175_, _15174_, _15173_, _15172_, _15171_, _15201_, _15200_, _15199_, _15198_, _15197_, _15196_, _15195_, _15192_, _15181_, _15170_ }) );
  \$mux  #( .WIDTH(32) ) _45780_ ( .A(control_matmul_29), .B(3), .S(_maxi_read_idle), .Y({ _15226_, _15225_, _15223_, _15222_, _15221_, _15220_, _15219_, _15218_, _15217_, _15216_, _15215_, _15214_, _15212_, _15211_, _15210_, _15209_, _15208_, _15207_, _15206_, _15205_, _15204_, _15203_, _15233_, _15232_, _15231_, _15230_, _15229_, _15228_, _15227_, _15224_, _15213_, _15202_ }) );
  \$mux  #( .WIDTH(32) ) _45781_ ( .A(1), .B(control_matmul_29), .S(_05729_), .Y(_24735_) );
  \$mux  #( .WIDTH(32) ) _45782_ ( .A(1), .B(_24735_), .S(_06026_), .Y(_24736_) );
  \$mux  #( .WIDTH(32) ) _45783_ ( .A(1), .B(_24736_), .S(_06024_), .Y({ _15258_, _15257_, _15255_, _15254_, _15253_, _15252_, _15251_, _15250_, _15249_, _15248_, _15247_, _15246_, _15244_, _15243_, _15242_, _15241_, _15240_, _15239_, _15238_, _15237_, _15236_, _15235_, _15265_, _15264_, _15263_, _15262_, _15261_, _15260_, _15259_, _15256_, _15245_, _15234_ }) );
  \$mux  #( .WIDTH(32) ) _45784_ ( .A(_24731_), .B(0), .S(RST), .Y(_03208_) );
  \$mux  #( .WIDTH(32) ) _45785_ ( .A(_stream_max_pool_serial_18_sink_3_sink_fsm_1), .B(0), .S(_06865_), .Y(_24737_) );
  \$mux  #( .WIDTH(32) ) _45786_ ( .A(_24737_), .B(0), .S(_stream_max_pool_serial_18_term_sink), .Y({ _15290_, _15289_, _15287_, _15286_, _15285_, _15284_, _15283_, _15282_, _15281_, _15280_, _15279_, _15278_, _15276_, _15275_, _15274_, _15273_, _15272_, _15271_, _15270_, _15269_, _15268_, _15267_, _15297_, _15296_, _15295_, _15294_, _15293_, _15292_, _15291_, _15288_, _15277_, _15266_ }) );
  \$mux  #( .WIDTH(32) ) _45787_ ( .A(_stream_max_pool_serial_18_sink_3_sink_fsm_1), .B(1), .S(_06793_), .Y({ _15354_, _15353_, _15351_, _15350_, _15349_, _15348_, _15347_, _15346_, _15345_, _15344_, _15343_, _15342_, _15340_, _15339_, _15338_, _15337_, _15336_, _15335_, _15334_, _15333_, _15332_, _15331_, _15361_, _15360_, _15359_, _15358_, _15357_, _15356_, _15355_, _15352_, _15341_, _15330_ }) );
  \$mux  #( .WIDTH(32) ) _45788_ ( .A(_24738_), .B(0), .S(RST), .Y(_02776_) );
  \$mux  #( .WIDTH(32) ) _45789_ ( .A(_stream_max_pool_serial_18_source_1_source_pat_fsm_0), .B(2), .S(_06864_), .Y({ _15418_, _15417_, _15415_, _15414_, _15413_, _15412_, _15411_, _15410_, _15409_, _15408_, _15407_, _15406_, _15404_, _15403_, _15402_, _15401_, _15400_, _15399_, _15398_, _15397_, _15396_, _15395_, _15425_, _15424_, _15423_, _15422_, _15421_, _15420_, _15419_, _15416_, _15405_, _15394_ }) );
  \$mux  #( .WIDTH(32) ) _45790_ ( .A(_stream_max_pool_serial_18_source_1_source_pat_fsm_0), .B(1), .S(_06788_), .Y({ _15450_, _15449_, _15447_, _15446_, _15445_, _15444_, _15443_, _15442_, _15441_, _15440_, _15439_, _15438_, _15436_, _15435_, _15434_, _15433_, _15432_, _15431_, _15430_, _15429_, _15428_, _15427_, _15457_, _15456_, _15455_, _15454_, _15453_, _15452_, _15451_, _15448_, _15437_, _15426_ }) );
  \$mux  #( .WIDTH(32) ) _45791_ ( .A(_24739_), .B(0), .S(RST), .Y(_02790_) );
  \$mux  #( .WIDTH(4) ) _45792_ ( .A({ max_pool_serial_18_stream_pad_mask_1_1, max_pool_serial_18_stream_pad_mask_1_0, max_pool_serial_18_stream_pad_mask_0_1, max_pool_serial_18_stream_pad_mask_0_0 }), .B(max_pool_serial_18_stream_pad_masks), .S(_05934_), .Y(_24740_) );
  \$mux  #( .WIDTH(4) ) _45793_ ( .A(_24740_), .B(4'h0), .S(RST), .Y(_03362_) );
  \$mux  #( .WIDTH(32) ) _45794_ ( .A(max_pool_serial_18_row_count), .B(max_pool_serial_18_row_count_buf), .S(_05937_), .Y(_24741_) );
  \$mux  #( .WIDTH(32) ) _45795_ ( .A(_24741_), .B(0), .S(RST), .Y(_03356_) );
  \$mux  #( .WIDTH(32) ) _45796_ ( .A(max_pool_serial_18_out_page_comp_offset), .B(max_pool_serial_18_out_page_comp_offset_buf), .S(_05937_), .Y(_24742_) );
  \$mux  #( .WIDTH(32) ) _45797_ ( .A(_24742_), .B(0), .S(RST), .Y(_03351_) );
  \$mux  #( .WIDTH(32) ) _45798_ ( .A(max_pool_serial_18_act_page_comp_offset), .B(max_pool_serial_18_act_page_comp_offset_buf), .S(_05937_), .Y(_24743_) );
  \$mux  #( .WIDTH(32) ) _45799_ ( .A(_24743_), .B(0), .S(RST), .Y(_03337_) );
  \$mux  #( .WIDTH(32) ) _45800_ ( .A(2), .B(0), .S(_06161_), .Y({ _15482_, _15481_, _15479_, _15478_, _15477_, _15476_, _15475_, _15474_, _15473_, _15472_, _15471_, _15470_, _15468_, _15467_, _15466_, _15465_, _15464_, _15463_, _15462_, _15461_, _15460_, _15459_, _15489_, _15488_, _15487_, _15486_, _15485_, _15484_, _15483_, _15480_, _15469_, _15458_ }) );
  \$mux  #( .WIDTH(32) ) _45801_ ( .A(4), .B(max_pool_serial_18_comp_fsm), .S(_stream_max_pool_serial_18_source_busy), .Y({ _15546_, _15545_, _15543_, _15542_, _15541_, _15540_, _15539_, _15538_, _15537_, _15536_, _15535_, _15534_, _15532_, _15531_, _15530_, _15529_, _15528_, _15527_, _15526_, _15525_, _15524_, _15523_, _15553_, _15552_, _15551_, _15550_, _15549_, _15548_, _15547_, _15544_, _15533_, _15522_ }) );
  \$mux  #( .WIDTH(32) ) _45802_ ( .A(max_pool_serial_18_comp_fsm), .B(1), .S(_06863_), .Y({ _15578_, _15577_, _15575_, _15574_, _15573_, _15572_, _15571_, _15570_, _15569_, _15568_, _15567_, _15566_, _15564_, _15563_, _15562_, _15561_, _15560_, _15559_, _15558_, _15557_, _15556_, _15555_, _15585_, _15584_, _15583_, _15582_, _15581_, _15580_, _15579_, _15576_, _15565_, _15554_ }) );
  \$mux  #( .WIDTH(32) ) _45803_ ( .A(_24744_), .B(0), .S(RST), .Y(_03343_) );
  \$mux  #( .WIDTH(32) ) _45804_ ( .A(0), .B(max_pool_serial_18_comp_count), .S(_05945_), .Y(_24745_) );
  \$mux  #( .WIDTH(32) ) _45805_ ( .A(_24745_), .B(_24468_), .S(_stream_max_pool_serial_18_end_flag), .Y(_24746_) );
  \$mux  #( .WIDTH(32) ) _45806_ ( .A(_24746_), .B(0), .S(RST), .Y(_03342_) );
  \$mux  #( .WIDTH(32) ) _45807_ ( .A(_24470_), .B(0), .S(_06161_), .Y({ _15610_, _15609_, _15607_, _15606_, _15605_, _15604_, _15603_, _15602_, _15601_, _15600_, _15599_, _15598_, _15596_, _15595_, _15594_, _15593_, _15592_, _15591_, _15590_, _15589_, _15588_, _15587_, _15617_, _15616_, _15615_, _15614_, _15613_, _15612_, _15611_, _15608_, _15597_, _15586_ }) );
  \$mux  #( .WIDTH(32) ) _45808_ ( .A(_24747_), .B(0), .S(RST), .Y(_03361_) );
  \$mux  #( .WIDTH(32) ) _45809_ ( .A(_24469_), .B(0), .S(_06161_), .Y({ _15674_, _15673_, _15671_, _15670_, _15669_, _15668_, _15667_, _15666_, _15665_, _15664_, _15663_, _15662_, _15660_, _15659_, _15658_, _15657_, _15656_, _15655_, _15654_, _15653_, _15652_, _15651_, _15681_, _15680_, _15679_, _15678_, _15677_, _15676_, _15675_, _15672_, _15661_, _15650_ }) );
  \$mux  #( .WIDTH(32) ) _45810_ ( .A(_24748_), .B(0), .S(RST), .Y(_03360_) );
  \$mux  #( .WIDTH(32) ) _45811_ ( .A(_24471_), .B(0), .S(_06161_), .Y({ _15738_, _15737_, _15735_, _15734_, _15733_, _15732_, _15731_, _15730_, _15729_, _15728_, _15727_, _15726_, _15724_, _15723_, _15722_, _15721_, _15720_, _15719_, _15718_, _15717_, _15716_, _15715_, _15745_, _15744_, _15743_, _15742_, _15741_, _15740_, _15739_, _15736_, _15725_, _15714_ }) );
  \$mux  #( .WIDTH(32) ) _45812_ ( .A(_24749_), .B(0), .S(RST), .Y(_03341_) );
  \$mux  #( .WIDTH(1) ) _45813_ ( .A(1'h1), .B(_control_max_pool_serial_18_cond_19_2_1), .S(_05941_), .Y(_24750_) );
  \$mux  #( .WIDTH(1) ) _45814_ ( .A(_24750_), .B(1'h0), .S(RST), .Y(_01577_) );
  \$mux  #( .WIDTH(1) ) _45815_ ( .A(axim_flag_1071), .B(1'h0), .S(_control_max_pool_serial_18_cond_19_2_1), .Y(_24751_) );
  \$mux  #( .WIDTH(1) ) _45816_ ( .A(_24751_), .B(axim_flag_1071), .S(_05938_), .Y(_24752_) );
  \$mux  #( .WIDTH(1) ) _45817_ ( .A(1'h1), .B(_24752_), .S(_05941_), .Y(_24753_) );
  \$mux  #( .WIDTH(1) ) _45818_ ( .A(_24753_), .B(1'h0), .S(RST), .Y(_03193_) );
  \$mux  #( .WIDTH(1) ) _45819_ ( .A(1'h1), .B(_control_max_pool_serial_18_cond_11_1_1), .S(_05943_), .Y(_24754_) );
  \$mux  #( .WIDTH(1) ) _45820_ ( .A(_24754_), .B(1'h0), .S(RST), .Y(_01576_) );
  \$mux  #( .WIDTH(1) ) _45821_ ( .A(axim_flag_1023), .B(1'h0), .S(_control_max_pool_serial_18_cond_11_1_1), .Y(_24755_) );
  \$mux  #( .WIDTH(1) ) _45822_ ( .A(_24755_), .B(axim_flag_1023), .S(_05939_), .Y(_24756_) );
  \$mux  #( .WIDTH(1) ) _45823_ ( .A(1'h1), .B(_24756_), .S(_05943_), .Y(_24757_) );
  \$mux  #( .WIDTH(1) ) _45824_ ( .A(_24757_), .B(1'h0), .S(RST), .Y(_03192_) );
  \$mux  #( .WIDTH(1) ) _45825_ ( .A(1'h1), .B(_control_max_pool_serial_18_cond_5_0_1), .S(_05944_), .Y(_24758_) );
  \$mux  #( .WIDTH(1) ) _45826_ ( .A(_24758_), .B(1'h0), .S(RST), .Y(_01578_) );
  \$mux  #( .WIDTH(32) ) _45827_ ( .A(control_max_pool_serial_18), .B(0), .S(RST), .Y(_01585_) );
  \$mux  #( .WIDTH(1) ) _45828_ ( .A(axim_flag_1022), .B(1'h0), .S(_control_max_pool_serial_18_cond_5_0_1), .Y(_24759_) );
  \$mux  #( .WIDTH(1) ) _45829_ ( .A(_24759_), .B(axim_flag_1022), .S(_05940_), .Y(_24760_) );
  \$mux  #( .WIDTH(1) ) _45830_ ( .A(1'h1), .B(_24760_), .S(_05944_), .Y(_24761_) );
  \$mux  #( .WIDTH(1) ) _45831_ ( .A(_24761_), .B(1'h0), .S(RST), .Y(_03191_) );
  \$mux  #( .WIDTH(32) ) _45832_ ( .A(_24762_), .B(0), .S(RST), .Y(_03348_) );
  \$mux  #( .WIDTH(1) ) _45833_ ( .A(max_pool_serial_18_skip_write_out), .B(1'h0), .S(_06862_), .Y(_15810_) );
  \$mux  #( .WIDTH(1) ) _45834_ ( .A(_24763_), .B(1'h0), .S(RST), .Y(_03359_) );
  \$mux  #( .WIDTH(1) ) _45835_ ( .A(max_pool_serial_18_skip_comp), .B(1'h1), .S(_06160_), .Y(_15812_) );
  \$mux  #( .WIDTH(1) ) _45836_ ( .A(_24764_), .B(1'h0), .S(RST), .Y(_03357_) );
  \$mux  #( .WIDTH(1) ) _45837_ ( .A(max_pool_serial_18_skip_read_act), .B(1'h1), .S(_06160_), .Y(_15814_) );
  \$mux  #( .WIDTH(1) ) _45838_ ( .A(_24765_), .B(1'h0), .S(RST), .Y(_03358_) );
  \$mux  #( .WIDTH(32) ) _45839_ ( .A(0), .B(1024), .S(max_pool_serial_18_out_page), .Y({ _15840_, _15839_, _15837_, _15836_, _15835_, _15834_, _15833_, _15832_, _15831_, _15830_, _15829_, _15828_, _15826_, _15825_, _15824_, _15823_, _15822_, _15821_, _15820_, _15819_, _15818_, _15817_, _15847_, _15846_, _15845_, _15844_, _15843_, _15842_, _15841_, _15838_, _15827_, _15816_ }) );
  \$mux  #( .WIDTH(32) ) _45840_ ( .A(_24766_), .B(0), .S(RST), .Y(_03352_) );
  \$mux  #( .WIDTH(32) ) _45841_ ( .A(1024), .B(0), .S(max_pool_serial_18_out_page), .Y({ _15904_, _15903_, _15901_, _15900_, _15899_, _15898_, _15897_, _15896_, _15895_, _15894_, _15893_, _15892_, _15890_, _15889_, _15888_, _15887_, _15886_, _15885_, _15884_, _15883_, _15882_, _15881_, _15911_, _15910_, _15909_, _15908_, _15907_, _15906_, _15905_, _15902_, _15891_, _15880_ }) );
  \$mux  #( .WIDTH(32) ) _45842_ ( .A(_24767_), .B(0), .S(RST), .Y(_03350_) );
  \$mux  #( .WIDTH(1) ) _45843_ ( .A(1'h1), .B(1'h0), .S(max_pool_serial_18_out_page), .Y(_15944_) );
  \$mux  #( .WIDTH(1) ) _45844_ ( .A(_24768_), .B(1'h0), .S(RST), .Y(_03349_) );
  \$mux  #( .WIDTH(32) ) _45845_ ( .A(_24769_), .B(0), .S(RST), .Y(_03338_) );
  \$mux  #( .WIDTH(32) ) _45846_ ( .A(1024), .B(0), .S(max_pool_serial_18_act_page), .Y({ _15970_, _15969_, _15967_, _15966_, _15965_, _15964_, _15963_, _15962_, _15961_, _15960_, _15959_, _15958_, _15956_, _15955_, _15954_, _15953_, _15952_, _15951_, _15950_, _15949_, _15948_, _15947_, _15977_, _15976_, _15975_, _15974_, _15973_, _15972_, _15971_, _15968_, _15957_, _15946_ }) );
  \$mux  #( .WIDTH(32) ) _45847_ ( .A(_24770_), .B(0), .S(RST), .Y(_03336_) );
  \$mux  #( .WIDTH(1) ) _45848_ ( .A(1'h1), .B(1'h0), .S(max_pool_serial_18_act_page), .Y(_16010_) );
  \$mux  #( .WIDTH(1) ) _45849_ ( .A(_24771_), .B(1'h0), .S(RST), .Y(_03335_) );
  \$mux  #( .WIDTH(32) ) _45850_ ( .A(_24772_), .B(0), .S(RST), .Y(_03353_) );
  \$mux  #( .WIDTH(32) ) _45851_ ( .A(_24773_), .B(0), .S(RST), .Y(_03354_) );
  \$mux  #( .WIDTH(32) ) _45852_ ( .A(max_pool_serial_18_bat_count), .B(0), .S(_06160_), .Y({ _16100_, _16099_, _16097_, _16096_, _16095_, _16094_, _16093_, _16092_, _16091_, _16090_, _16089_, _16088_, _16086_, _16085_, _16084_, _16083_, _16082_, _16081_, _16080_, _16079_, _16078_, _16077_, _16107_, _16106_, _16105_, _16104_, _16103_, _16102_, _16101_, _16098_, _16087_, _16076_ }) );
  \$mux  #( .WIDTH(32) ) _45853_ ( .A(_24774_), .B(0), .S(RST), .Y(_03340_) );
  \$mux  #( .WIDTH(32) ) _45854_ ( .A(_24466_), .B(0), .S(_06160_), .Y({ _16164_, _16163_, _16161_, _16160_, _16159_, _16158_, _16157_, _16156_, _16155_, _16154_, _16153_, _16152_, _16150_, _16149_, _16148_, _16147_, _16146_, _16145_, _16144_, _16143_, _16142_, _16141_, _16171_, _16170_, _16169_, _16168_, _16167_, _16166_, _16165_, _16162_, _16151_, _16140_ }) );
  \$mux  #( .WIDTH(32) ) _45855_ ( .A(_24775_), .B(0), .S(RST), .Y(_03355_) );
  \$mux  #( .WIDTH(32) ) _45856_ ( .A(max_pool_serial_18_out_base_offset_bat), .B(0), .S(_06861_), .Y({ _16228_, _16227_, _16225_, _16224_, _16223_, _16222_, _16221_, _16220_, _16219_, _16218_, _16217_, _16216_, _16214_, _16213_, _16212_, _16211_, _16210_, _16209_, _16208_, _16207_, _16206_, _16205_, _16235_, _16234_, _16233_, _16232_, _16231_, _16230_, _16229_, _16226_, _16215_, _16204_ }) );
  \$mux  #( .WIDTH(32) ) _45857_ ( .A(_24776_), .B(0), .S(RST), .Y(_03346_) );
  \$mux  #( .WIDTH(32) ) _45858_ ( .A(_24467_), .B(max_pool_serial_18_out_base_offset_row), .S(max_pool_serial_18_skip_write_out), .Y(_24777_) );
  \$mux  #( .WIDTH(32) ) _45859_ ( .A(_24777_), .B(0), .S(_06861_), .Y({ _16292_, _16291_, _16289_, _16288_, _16287_, _16286_, _16285_, _16284_, _16283_, _16282_, _16281_, _16280_, _16278_, _16277_, _16276_, _16275_, _16274_, _16273_, _16272_, _16271_, _16270_, _16269_, _16299_, _16298_, _16297_, _16296_, _16295_, _16294_, _16293_, _16290_, _16279_, _16268_ }) );
  \$mux  #( .WIDTH(32) ) _45860_ ( .A(_24778_), .B(0), .S(RST), .Y(_03347_) );
  \$mux  #( .WIDTH(32) ) _45861_ ( .A(max_pool_serial_18_act_base_offset_bat), .B(0), .S(_06160_), .Y({ _16356_, _16355_, _16353_, _16352_, _16351_, _16350_, _16349_, _16348_, _16347_, _16346_, _16345_, _16344_, _16342_, _16341_, _16340_, _16339_, _16338_, _16337_, _16336_, _16335_, _16334_, _16333_, _16363_, _16362_, _16361_, _16360_, _16359_, _16358_, _16357_, _16354_, _16343_, _16332_ }) );
  \$mux  #( .WIDTH(32) ) _45862_ ( .A(_24779_), .B(0), .S(RST), .Y(_03333_) );
  \$mux  #( .WIDTH(32) ) _45863_ ( .A(_24465_), .B(0), .S(_06160_), .Y({ _16420_, _16419_, _16417_, _16416_, _16415_, _16414_, _16413_, _16412_, _16411_, _16410_, _16409_, _16408_, _16406_, _16405_, _16404_, _16403_, _16402_, _16401_, _16400_, _16399_, _16398_, _16397_, _16427_, _16426_, _16425_, _16424_, _16423_, _16422_, _16421_, _16418_, _16407_, _16396_ }) );
  \$mux  #( .WIDTH(32) ) _45864_ ( .A(_24780_), .B(0), .S(RST), .Y(_03334_) );
  \$mux  #( .WIDTH(32) ) _45865_ ( .A(0), .B(control_max_pool_serial_18), .S(_05738_), .Y(_24781_) );
  \$mux  #( .WIDTH(32) ) _45866_ ( .A(0), .B(_24781_), .S(_05734_), .Y(_24782_) );
  \$mux  #( .WIDTH(32) ) _45867_ ( .A(0), .B(_24782_), .S(_05730_), .Y({ _16484_, _16483_, _16481_, _16480_, _16479_, _16478_, _16477_, _16476_, _16475_, _16474_, _16473_, _16472_, _16470_, _16469_, _16468_, _16467_, _16466_, _16465_, _16464_, _16463_, _16462_, _16461_, _16491_, _16490_, _16489_, _16488_, _16487_, _16486_, _16485_, _16482_, _16471_, _16460_ }) );
  \$mux  #( .WIDTH(32) ) _45868_ ( .A(control_max_pool_serial_18), .B(25), .S(_maxi_write_idle), .Y({ _16548_, _16547_, _16545_, _16544_, _16543_, _16542_, _16541_, _16540_, _16539_, _16538_, _16537_, _16536_, _16534_, _16533_, _16532_, _16531_, _16530_, _16529_, _16528_, _16527_, _16526_, _16525_, _16555_, _16554_, _16553_, _16552_, _16551_, _16550_, _16549_, _16546_, _16535_, _16524_ }) );
  \$mux  #( .WIDTH(32) ) _45869_ ( .A(3), .B(24), .S(_06861_), .Y({ _16580_, _16579_, _16577_, _16576_, _16575_, _16574_, _16573_, _16572_, _16571_, _16570_, _16569_, _16568_, _16566_, _16565_, _16564_, _16563_, _16562_, _16561_, _16560_, _16559_, _16558_, _16557_, _16587_, _16586_, _16585_, _16584_, _16583_, _16582_, _16581_, _16578_, _16567_, _16556_ }) );
  \$mux  #( .WIDTH(32) ) _45870_ ( .A(control_max_pool_serial_18), .B(19), .S(_maxi_write_idle), .Y({ _16612_, _16611_, _16609_, _16608_, _16607_, _16606_, _16605_, _16604_, _16603_, _16602_, _16601_, _16600_, _16598_, _16597_, _16596_, _16595_, _16594_, _16593_, _16592_, _16591_, _16590_, _16589_, _16619_, _16618_, _16617_, _16616_, _16615_, _16614_, _16613_, _16610_, _16599_, _16588_ }) );
  \$mux  #( .WIDTH(32) ) _45871_ ( .A(control_max_pool_serial_18), .B(18), .S(_06159_), .Y(_24784_) );
  \$mux  #( .WIDTH(32) ) _45872_ ( .A(_24784_), .B(23), .S(max_pool_serial_18_skip_write_out), .Y({ _16644_, _16643_, _16641_, _16640_, _16639_, _16638_, _16637_, _16636_, _16635_, _16634_, _16633_, _16632_, _16630_, _16629_, _16628_, _16627_, _16626_, _16625_, _16624_, _16623_, _16622_, _16621_, _16651_, _16650_, _16649_, _16648_, _16647_, _16646_, _16645_, _16642_, _16631_, _16620_ }) );
  \$mux  #( .WIDTH(32) ) _45873_ ( .A(17), .B(control_max_pool_serial_18), .S(_05726_), .Y({ _16676_, _16675_, _16673_, _16672_, _16671_, _16670_, _16669_, _16668_, _16667_, _16666_, _16665_, _16664_, _16662_, _16661_, _16660_, _16659_, _16658_, _16657_, _16656_, _16655_, _16654_, _16653_, _16683_, _16682_, _16681_, _16680_, _16679_, _16678_, _16677_, _16674_, _16663_, _16652_ }) );
  \$mux  #( .WIDTH(32) ) _45874_ ( .A(control_max_pool_serial_18), .B(15), .S(_maxi_read_idle), .Y({ _16708_, _16707_, _16705_, _16704_, _16703_, _16702_, _16701_, _16700_, _16699_, _16698_, _16697_, _16696_, _16694_, _16693_, _16692_, _16691_, _16690_, _16689_, _16688_, _16687_, _16686_, _16685_, _16715_, _16714_, _16713_, _16712_, _16711_, _16710_, _16709_, _16706_, _16695_, _16684_ }) );
  \$mux  #( .WIDTH(32) ) _45875_ ( .A(control_max_pool_serial_18), .B(11), .S(_maxi_read_idle), .Y({ _16740_, _16739_, _16737_, _16736_, _16735_, _16734_, _16733_, _16732_, _16731_, _16730_, _16729_, _16728_, _16726_, _16725_, _16724_, _16723_, _16722_, _16721_, _16720_, _16719_, _16718_, _16717_, _16747_, _16746_, _16745_, _16744_, _16743_, _16742_, _16741_, _16738_, _16727_, _16716_ }) );
  \$mux  #( .WIDTH(32) ) _45876_ ( .A(10), .B(15), .S(max_pool_serial_18_dma_pad_mask_1), .Y({ _16772_, _16771_, _16769_, _16768_, _16767_, _16766_, _16765_, _16764_, _16763_, _16762_, _16761_, _16760_, _16758_, _16757_, _16756_, _16755_, _16754_, _16753_, _16752_, _16751_, _16750_, _16749_, _16779_, _16778_, _16777_, _16776_, _16775_, _16774_, _16773_, _16770_, _16759_, _16748_ }) );
  \$mux  #( .WIDTH(32) ) _45877_ ( .A(control_max_pool_serial_18), .B(9), .S(_maxi_read_idle), .Y({ _16804_, _16803_, _16801_, _16800_, _16799_, _16798_, _16797_, _16796_, _16795_, _16794_, _16793_, _16792_, _16790_, _16789_, _16788_, _16787_, _16786_, _16785_, _16784_, _16783_, _16782_, _16781_, _16811_, _16810_, _16809_, _16808_, _16807_, _16806_, _16805_, _16802_, _16791_, _16780_ }) );
  \$mux  #( .WIDTH(32) ) _45878_ ( .A(control_max_pool_serial_18), .B(5), .S(_maxi_read_idle), .Y({ _16836_, _16835_, _16833_, _16832_, _16831_, _16830_, _16829_, _16828_, _16827_, _16826_, _16825_, _16824_, _16822_, _16821_, _16820_, _16819_, _16818_, _16817_, _16816_, _16815_, _16814_, _16813_, _16843_, _16842_, _16841_, _16840_, _16839_, _16838_, _16837_, _16834_, _16823_, _16812_ }) );
  \$mux  #( .WIDTH(32) ) _45879_ ( .A(4), .B(9), .S(max_pool_serial_18_dma_pad_mask_0), .Y(_24785_) );
  \$mux  #( .WIDTH(32) ) _45880_ ( .A(_24785_), .B(16), .S(max_pool_serial_18_skip_read_act), .Y({ _16868_, _16867_, _16865_, _16864_, _16863_, _16862_, _16861_, _16860_, _16859_, _16858_, _16857_, _16856_, _16854_, _16853_, _16852_, _16851_, _16850_, _16849_, _16848_, _16847_, _16846_, _16845_, _16875_, _16874_, _16873_, _16872_, _16871_, _16870_, _16869_, _16866_, _16855_, _16844_ }) );
  \$mux  #( .WIDTH(32) ) _45881_ ( .A(1), .B(control_max_pool_serial_18), .S(_05739_), .Y(_24786_) );
  \$mux  #( .WIDTH(32) ) _45882_ ( .A(1), .B(_24786_), .S(_05735_), .Y(_24787_) );
  \$mux  #( .WIDTH(32) ) _45883_ ( .A(1), .B(_24787_), .S(_05731_), .Y({ _16900_, _16899_, _16897_, _16896_, _16895_, _16894_, _16893_, _16892_, _16891_, _16890_, _16889_, _16888_, _16886_, _16885_, _16884_, _16883_, _16882_, _16881_, _16880_, _16879_, _16878_, _16877_, _16907_, _16906_, _16905_, _16904_, _16903_, _16902_, _16901_, _16898_, _16887_, _16876_ }) );
  \$mux  #( .WIDTH(32) ) _45884_ ( .A(_24783_), .B(0), .S(RST), .Y(_03209_) );
  \$mux  #( .WIDTH(1) ) _45885_ ( .A(1'h1), .B(__maxi_write_fsm_cond_4_0_1), .S(_05947_), .Y(_24788_) );
  \$mux  #( .WIDTH(1) ) _45886_ ( .A(_24788_), .B(1'h0), .S(_RESETN_inv_2), .Y(_00691_) );
  \$mux  #( .WIDTH(32) ) _45887_ ( .A(_maxi_write_fsm), .B(0), .S(_RESETN_inv_2), .Y(_01582_) );
  \$mux  #( .WIDTH(1) ) _45888_ ( .A(axim_flag_1021), .B(1'h0), .S(__maxi_write_fsm_cond_4_0_1), .Y(_24789_) );
  \$mux  #( .WIDTH(1) ) _45889_ ( .A(_24789_), .B(axim_flag_1021), .S(_05946_), .Y(_24790_) );
  \$mux  #( .WIDTH(1) ) _45890_ ( .A(1'h1), .B(_24790_), .S(_05947_), .Y(_24791_) );
  \$mux  #( .WIDTH(1) ) _45891_ ( .A(_24791_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03190_) );
  \$mux  #( .WIDTH(33) ) _45892_ ( .A(_28942_), .B(_28941_), .S(_06158_), .Y(_24792_) );
  \$mux  #( .WIDTH(33) ) _45893_ ( .A(_24792_), .B(33'h000000000), .S(_06176_), .Y(_24793_) );
  \$mux  #( .WIDTH(33) ) _45894_ ( .A(_24793_), .B(_28941_), .S(_06858_), .Y({ _16933_, _16932_, _16931_, _16929_, _16928_, _16927_, _16926_, _16925_, _16924_, _16923_, _16922_, _16921_, _16920_, _16918_, _16917_, _16916_, _16915_, _16914_, _16913_, _16912_, _16911_, _16910_, _16909_, _16940_, _16939_, _16938_, _16937_, _16936_, _16935_, _16934_, _16930_, _16919_, _16908_ }) );
  \$mux  #( .WIDTH(33) ) _45895_ ( .A(_maxi_write_rest_size), .B(_maxi_write_size), .S(_maxi_write_start), .Y({ _16999_, _16998_, _16997_, _16995_, _16994_, _16993_, _16992_, _16991_, _16990_, _16989_, _16988_, _16987_, _16986_, _16984_, _16983_, _16982_, _16981_, _16980_, _16979_, _16978_, _16977_, _16976_, _16975_, _17006_, _17005_, _17004_, _17003_, _17002_, _17001_, _17000_, _16996_, _16985_, _16974_ }) );
  \$mux  #( .WIDTH(33) ) _45896_ ( .A(_24794_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01797_) );
  \$mux  #( .WIDTH(33) ) _45897_ ( .A(33'h000000100), .B({ 2'h0, _28520_[30:0] }), .S(_06158_), .Y(_24795_) );
  \$mux  #( .WIDTH(33) ) _45898_ ( .A(_24795_), .B(_maxi_write_rest_size), .S(_06176_), .Y(_24796_) );
  \$mux  #( .WIDTH(33) ) _45899_ ( .A(_24796_), .B({ 2'h0, _28520_[30:0] }), .S(_06858_), .Y(_24797_) );
  \$mux  #( .WIDTH(33) ) _45900_ ( .A(_24797_), .B(_maxi_write_cur_size), .S(_05948_), .Y(_24798_) );
  \$mux  #( .WIDTH(33) ) _45901_ ( .A(_24798_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01790_) );
  \$mux  #( .WIDTH(32) ) _45902_ ( .A(_maxi_write_cur_global_addr), .B(_24464_[31:0]), .S(_maxi_write_data_done), .Y({ _17031_, _17030_, _17028_, _17027_, _17026_, _17025_, _17024_, _17023_, _17022_, _17021_, _17020_, _17019_, _17017_, _17016_, _17015_, _17014_, _17013_, _17012_, _17011_, _17010_, _17009_, _17008_, _17038_, _17037_, _17036_, _17035_, _17034_, _17033_, _17032_, _17029_, _17018_, _17007_ }) );
  \$mux  #( .WIDTH(32) ) _45903_ ( .A(_maxi_write_cur_global_addr), .B({ _24463_[31:2], 2'h0 }), .S(_maxi_write_start), .Y({ _17095_, _17094_, _17092_, _17091_, _17090_, _17089_, _17088_, _17087_, _17086_, _17085_, _17084_, _17083_, _17081_, _17080_, _17079_, _17078_, _17077_, _17076_, _17075_, _17074_, _17073_, _17072_, _17102_, _17101_, _17100_, _17099_, _17098_, _17097_, _17096_, _17093_, _17082_, _17071_ }) );
  \$mux  #( .WIDTH(32) ) _45904_ ( .A(_24799_), .B(0), .S(_RESETN_inv_2), .Y(_01789_) );
  \$mux  #( .WIDTH(32) ) _45905_ ( .A(_maxi_write_fsm), .B(1), .S(_06859_), .Y(_24801_) );
  \$mux  #( .WIDTH(32) ) _45906_ ( .A(_24801_), .B(4), .S(_06860_), .Y({ _17159_, _17158_, _17156_, _17155_, _17154_, _17153_, _17152_, _17151_, _17150_, _17149_, _17148_, _17147_, _17145_, _17144_, _17143_, _17142_, _17141_, _17140_, _17139_, _17138_, _17137_, _17136_, _17166_, _17165_, _17164_, _17163_, _17162_, _17161_, _17160_, _17157_, _17146_, _17135_ }) );
  \$mux  #( .WIDTH(32) ) _45907_ ( .A(_maxi_write_fsm), .B(3), .S(_06876_), .Y({ _17191_, _17190_, _17188_, _17187_, _17186_, _17185_, _17184_, _17183_, _17182_, _17181_, _17180_, _17179_, _17177_, _17176_, _17175_, _17174_, _17173_, _17172_, _17171_, _17170_, _17169_, _17168_, _17198_, _17197_, _17196_, _17195_, _17194_, _17193_, _17192_, _17189_, _17178_, _17167_ }) );
  \$mux  #( .WIDTH(32) ) _45908_ ( .A(_maxi_write_fsm), .B(1), .S(_06662_), .Y(_24802_) );
  \$mux  #( .WIDTH(32) ) _45909_ ( .A(_24802_), .B(1), .S(_06488_), .Y(_24803_) );
  \$mux  #( .WIDTH(32) ) _45910_ ( .A(_24803_), .B(1), .S(_06524_), .Y({ _17223_, _17222_, _17220_, _17219_, _17218_, _17217_, _17216_, _17215_, _17214_, _17213_, _17212_, _17211_, _17209_, _17208_, _17207_, _17206_, _17205_, _17204_, _17203_, _17202_, _17201_, _17200_, _17230_, _17229_, _17228_, _17227_, _17226_, _17225_, _17224_, _17221_, _17210_, _17199_ }) );
  \$mux  #( .WIDTH(32) ) _45911_ ( .A(_24800_), .B(0), .S(_RESETN_inv_2), .Y(_01791_) );
  \$mux  #( .WIDTH(32) ) _45912_ ( .A(_stream_conv2d_16_sink_37_sink_fsm_20), .B(0), .S(_06857_), .Y(_24804_) );
  \$mux  #( .WIDTH(32) ) _45913_ ( .A(_24804_), .B(0), .S(_stream_conv2d_16_term_sink), .Y({ _17255_, _17254_, _17252_, _17251_, _17250_, _17249_, _17248_, _17247_, _17246_, _17245_, _17244_, _17243_, _17241_, _17240_, _17239_, _17238_, _17237_, _17236_, _17235_, _17234_, _17233_, _17232_, _17262_, _17261_, _17260_, _17259_, _17258_, _17257_, _17256_, _17253_, _17242_, _17231_ }) );
  \$mux  #( .WIDTH(32) ) _45914_ ( .A(_stream_conv2d_16_sink_37_sink_fsm_20), .B(1), .S(_06786_), .Y({ _17319_, _17318_, _17316_, _17315_, _17314_, _17313_, _17312_, _17311_, _17310_, _17309_, _17308_, _17307_, _17305_, _17304_, _17303_, _17302_, _17301_, _17300_, _17299_, _17298_, _17297_, _17296_, _17326_, _17325_, _17324_, _17323_, _17322_, _17321_, _17320_, _17317_, _17306_, _17295_ }) );
  \$mux  #( .WIDTH(32) ) _45915_ ( .A(_24805_), .B(0), .S(RST), .Y(_02505_) );
  \$mux  #( .WIDTH(32) ) _45916_ ( .A(_stream_conv2d_16_source_36_source_pat_fsm_19), .B(2), .S(_06856_), .Y({ _17383_, _17382_, _17380_, _17379_, _17378_, _17377_, _17376_, _17375_, _17374_, _17373_, _17372_, _17371_, _17369_, _17368_, _17367_, _17366_, _17365_, _17364_, _17363_, _17362_, _17361_, _17360_, _17390_, _17389_, _17388_, _17387_, _17386_, _17385_, _17384_, _17381_, _17370_, _17359_ }) );
  \$mux  #( .WIDTH(32) ) _45917_ ( .A(_stream_conv2d_16_source_36_source_pat_fsm_19), .B(1), .S(_06781_), .Y({ _17415_, _17414_, _17412_, _17411_, _17410_, _17409_, _17408_, _17407_, _17406_, _17405_, _17404_, _17403_, _17401_, _17400_, _17399_, _17398_, _17397_, _17396_, _17395_, _17394_, _17393_, _17392_, _17422_, _17421_, _17420_, _17419_, _17418_, _17417_, _17416_, _17413_, _17402_, _17391_ }) );
  \$mux  #( .WIDTH(32) ) _45918_ ( .A(_24806_), .B(0), .S(RST), .Y(_02678_) );
  \$mux  #( .WIDTH(3) ) _45919_ ( .A(__tmp_697_1), .B(3'h0), .S(RST), .Y(_01287_) );
  \$mux  #( .WIDTH(3) ) _45920_ ( .A(_stream_conv2d_16_source_36_source_ram_raddr[2:0]), .B(3'h0), .S(RST), .Y(_01286_) );
  \$mux  #( .WIDTH(32) ) _45921_ ( .A(_stream_conv2d_16_source_35_source_pat_fsm_18), .B(2), .S(_06855_), .Y({ _17479_, _17478_, _17476_, _17475_, _17474_, _17473_, _17472_, _17471_, _17470_, _17469_, _17468_, _17467_, _17465_, _17464_, _17463_, _17462_, _17461_, _17460_, _17459_, _17458_, _17457_, _17456_, _17486_, _17485_, _17484_, _17483_, _17482_, _17481_, _17480_, _17477_, _17466_, _17455_ }) );
  \$mux  #( .WIDTH(32) ) _45922_ ( .A(_stream_conv2d_16_source_35_source_pat_fsm_18), .B(1), .S(_06776_), .Y({ _17511_, _17510_, _17508_, _17507_, _17506_, _17505_, _17504_, _17503_, _17502_, _17501_, _17500_, _17499_, _17497_, _17496_, _17495_, _17494_, _17493_, _17492_, _17491_, _17490_, _17489_, _17488_, _17518_, _17517_, _17516_, _17515_, _17514_, _17513_, _17512_, _17509_, _17498_, _17487_ }) );
  \$mux  #( .WIDTH(32) ) _45923_ ( .A(_24807_), .B(0), .S(RST), .Y(_02669_) );
  \$mux  #( .WIDTH(3) ) _45924_ ( .A(__tmp_683_1), .B(3'h0), .S(RST), .Y(_01284_) );
  \$mux  #( .WIDTH(3) ) _45925_ ( .A(_stream_conv2d_16_source_35_source_ram_raddr[2:0]), .B(3'h0), .S(RST), .Y(_01283_) );
  \$mux  #( .WIDTH(32) ) _45926_ ( .A(_stream_conv2d_16_source_34_source_pat_fsm_17), .B(2), .S(_06854_), .Y({ _17575_, _17574_, _17572_, _17571_, _17570_, _17569_, _17568_, _17567_, _17566_, _17565_, _17564_, _17563_, _17561_, _17560_, _17559_, _17558_, _17557_, _17556_, _17555_, _17554_, _17553_, _17552_, _17582_, _17581_, _17580_, _17579_, _17578_, _17577_, _17576_, _17573_, _17562_, _17551_ }) );
  \$mux  #( .WIDTH(32) ) _45927_ ( .A(_stream_conv2d_16_source_34_source_pat_fsm_17), .B(1), .S(_06771_), .Y({ _17607_, _17606_, _17604_, _17603_, _17602_, _17601_, _17600_, _17599_, _17598_, _17597_, _17596_, _17595_, _17593_, _17592_, _17591_, _17590_, _17589_, _17588_, _17587_, _17586_, _17585_, _17584_, _17614_, _17613_, _17612_, _17611_, _17610_, _17609_, _17608_, _17605_, _17594_, _17583_ }) );
  \$mux  #( .WIDTH(32) ) _45928_ ( .A(_24808_), .B(0), .S(RST), .Y(_02660_) );
  \$mux  #( .WIDTH(3) ) _45929_ ( .A(__tmp_669_1), .B(3'h0), .S(RST), .Y(_01281_) );
  \$mux  #( .WIDTH(3) ) _45930_ ( .A(_stream_conv2d_16_source_34_source_ram_raddr[2:0]), .B(3'h0), .S(RST), .Y(_01280_) );
  \$mux  #( .WIDTH(32) ) _45931_ ( .A(_stream_conv2d_16_source_33_source_pat_fsm_16), .B(2), .S(_06853_), .Y({ _17671_, _17670_, _17668_, _17667_, _17666_, _17665_, _17664_, _17663_, _17662_, _17661_, _17660_, _17659_, _17657_, _17656_, _17655_, _17654_, _17653_, _17652_, _17651_, _17650_, _17649_, _17648_, _17678_, _17677_, _17676_, _17675_, _17674_, _17673_, _17672_, _17669_, _17658_, _17647_ }) );
  \$mux  #( .WIDTH(32) ) _45932_ ( .A(_stream_conv2d_16_source_33_source_pat_fsm_16), .B(1), .S(_06766_), .Y({ _17703_, _17702_, _17700_, _17699_, _17698_, _17697_, _17696_, _17695_, _17694_, _17693_, _17692_, _17691_, _17689_, _17688_, _17687_, _17686_, _17685_, _17684_, _17683_, _17682_, _17681_, _17680_, _17710_, _17709_, _17708_, _17707_, _17706_, _17705_, _17704_, _17701_, _17690_, _17679_ }) );
  \$mux  #( .WIDTH(32) ) _45933_ ( .A(_24809_), .B(0), .S(RST), .Y(_02651_) );
  \$mux  #( .WIDTH(3) ) _45934_ ( .A(__tmp_655_1), .B(3'h0), .S(RST), .Y(_01278_) );
  \$mux  #( .WIDTH(3) ) _45935_ ( .A(_stream_conv2d_16_source_33_source_ram_raddr[2:0]), .B(3'h0), .S(RST), .Y(_01277_) );
  \$mux  #( .WIDTH(32) ) _45936_ ( .A(_stream_conv2d_16_source_32_source_pat_fsm_15), .B(2), .S(_06852_), .Y({ _17767_, _17766_, _17764_, _17763_, _17762_, _17761_, _17760_, _17759_, _17758_, _17757_, _17756_, _17755_, _17753_, _17752_, _17751_, _17750_, _17749_, _17748_, _17747_, _17746_, _17745_, _17744_, _17774_, _17773_, _17772_, _17771_, _17770_, _17769_, _17768_, _17765_, _17754_, _17743_ }) );
  \$mux  #( .WIDTH(32) ) _45937_ ( .A(_stream_conv2d_16_source_32_source_pat_fsm_15), .B(1), .S(_06761_), .Y({ _17799_, _17798_, _17796_, _17795_, _17794_, _17793_, _17792_, _17791_, _17790_, _17789_, _17788_, _17787_, _17785_, _17784_, _17783_, _17782_, _17781_, _17780_, _17779_, _17778_, _17777_, _17776_, _17806_, _17805_, _17804_, _17803_, _17802_, _17801_, _17800_, _17797_, _17786_, _17775_ }) );
  \$mux  #( .WIDTH(32) ) _45938_ ( .A(_24810_), .B(0), .S(RST), .Y(_02642_) );
  \$mux  #( .WIDTH(3) ) _45939_ ( .A(__tmp_641_1), .B(3'h0), .S(RST), .Y(_01275_) );
  \$mux  #( .WIDTH(3) ) _45940_ ( .A(_stream_conv2d_16_source_32_source_ram_raddr[2:0]), .B(3'h0), .S(RST), .Y(_01274_) );
  \$mux  #( .WIDTH(32) ) _45941_ ( .A(_stream_conv2d_16_source_31_source_pat_fsm_14), .B(2), .S(_06851_), .Y({ _17863_, _17862_, _17860_, _17859_, _17858_, _17857_, _17856_, _17855_, _17854_, _17853_, _17852_, _17851_, _17849_, _17848_, _17847_, _17846_, _17845_, _17844_, _17843_, _17842_, _17841_, _17840_, _17870_, _17869_, _17868_, _17867_, _17866_, _17865_, _17864_, _17861_, _17850_, _17839_ }) );
  \$mux  #( .WIDTH(32) ) _45942_ ( .A(_stream_conv2d_16_source_31_source_pat_fsm_14), .B(1), .S(_06756_), .Y({ _17895_, _17894_, _17892_, _17891_, _17890_, _17889_, _17888_, _17887_, _17886_, _17885_, _17884_, _17883_, _17881_, _17880_, _17879_, _17878_, _17877_, _17876_, _17875_, _17874_, _17873_, _17872_, _17902_, _17901_, _17900_, _17899_, _17898_, _17897_, _17896_, _17893_, _17882_, _17871_ }) );
  \$mux  #( .WIDTH(32) ) _45943_ ( .A(_24811_), .B(0), .S(RST), .Y(_02633_) );
  \$mux  #( .WIDTH(3) ) _45944_ ( .A(__tmp_627_1), .B(3'h0), .S(RST), .Y(_01272_) );
  \$mux  #( .WIDTH(3) ) _45945_ ( .A(_stream_conv2d_16_source_31_source_ram_raddr[2:0]), .B(3'h0), .S(RST), .Y(_01271_) );
  \$mux  #( .WIDTH(32) ) _45946_ ( .A(_stream_conv2d_16_source_30_source_pat_fsm_13), .B(2), .S(_06850_), .Y({ _17959_, _17958_, _17956_, _17955_, _17954_, _17953_, _17952_, _17951_, _17950_, _17949_, _17948_, _17947_, _17945_, _17944_, _17943_, _17942_, _17941_, _17940_, _17939_, _17938_, _17937_, _17936_, _17966_, _17965_, _17964_, _17963_, _17962_, _17961_, _17960_, _17957_, _17946_, _17935_ }) );
  \$mux  #( .WIDTH(32) ) _45947_ ( .A(_stream_conv2d_16_source_30_source_pat_fsm_13), .B(1), .S(_06751_), .Y({ _17991_, _17990_, _17988_, _17987_, _17986_, _17985_, _17984_, _17983_, _17982_, _17981_, _17980_, _17979_, _17977_, _17976_, _17975_, _17974_, _17973_, _17972_, _17971_, _17970_, _17969_, _17968_, _17998_, _17997_, _17996_, _17995_, _17994_, _17993_, _17992_, _17989_, _17978_, _17967_ }) );
  \$mux  #( .WIDTH(32) ) _45948_ ( .A(_24812_), .B(0), .S(RST), .Y(_02624_) );
  \$mux  #( .WIDTH(3) ) _45949_ ( .A(__tmp_613_1), .B(3'h0), .S(RST), .Y(_01269_) );
  \$mux  #( .WIDTH(3) ) _45950_ ( .A(_stream_conv2d_16_source_30_source_ram_raddr[2:0]), .B(3'h0), .S(RST), .Y(_01268_) );
  \$mux  #( .WIDTH(32) ) _45951_ ( .A(_stream_conv2d_16_source_29_source_pat_fsm_12), .B(2), .S(_06849_), .Y({ _18055_, _18054_, _18052_, _18051_, _18050_, _18049_, _18048_, _18047_, _18046_, _18045_, _18044_, _18043_, _18041_, _18040_, _18039_, _18038_, _18037_, _18036_, _18035_, _18034_, _18033_, _18032_, _18062_, _18061_, _18060_, _18059_, _18058_, _18057_, _18056_, _18053_, _18042_, _18031_ }) );
  \$mux  #( .WIDTH(32) ) _45952_ ( .A(_stream_conv2d_16_source_29_source_pat_fsm_12), .B(1), .S(_06746_), .Y({ _18087_, _18086_, _18084_, _18083_, _18082_, _18081_, _18080_, _18079_, _18078_, _18077_, _18076_, _18075_, _18073_, _18072_, _18071_, _18070_, _18069_, _18068_, _18067_, _18066_, _18065_, _18064_, _18094_, _18093_, _18092_, _18091_, _18090_, _18089_, _18088_, _18085_, _18074_, _18063_ }) );
  \$mux  #( .WIDTH(32) ) _45953_ ( .A(_24813_), .B(0), .S(RST), .Y(_02615_) );
  \$mux  #( .WIDTH(3) ) _45954_ ( .A(__tmp_599_1), .B(3'h0), .S(RST), .Y(_01266_) );
  \$mux  #( .WIDTH(3) ) _45955_ ( .A(_stream_conv2d_16_source_29_source_ram_raddr[2:0]), .B(3'h0), .S(RST), .Y(_01265_) );
  \$mux  #( .WIDTH(32) ) _45956_ ( .A(_stream_conv2d_16_source_28_source_pat_fsm_11), .B(2), .S(_06848_), .Y({ _18151_, _18150_, _18148_, _18147_, _18146_, _18145_, _18144_, _18143_, _18142_, _18141_, _18140_, _18139_, _18137_, _18136_, _18135_, _18134_, _18133_, _18132_, _18131_, _18130_, _18129_, _18128_, _18158_, _18157_, _18156_, _18155_, _18154_, _18153_, _18152_, _18149_, _18138_, _18127_ }) );
  \$mux  #( .WIDTH(32) ) _45957_ ( .A(_stream_conv2d_16_source_28_source_pat_fsm_11), .B(1), .S(_06741_), .Y({ _18183_, _18182_, _18180_, _18179_, _18178_, _18177_, _18176_, _18175_, _18174_, _18173_, _18172_, _18171_, _18169_, _18168_, _18167_, _18166_, _18165_, _18164_, _18163_, _18162_, _18161_, _18160_, _18190_, _18189_, _18188_, _18187_, _18186_, _18185_, _18184_, _18181_, _18170_, _18159_ }) );
  \$mux  #( .WIDTH(32) ) _45958_ ( .A(_24814_), .B(0), .S(RST), .Y(_02606_) );
  \$mux  #( .WIDTH(3) ) _45959_ ( .A(__tmp_1211_1), .B(3'h0), .S(RST), .Y(_01149_) );
  \$mux  #( .WIDTH(3) ) _45960_ ( .A(_stream_matmul_29_source_20_source_ram_raddr[2:0]), .B(3'h0), .S(RST), .Y(_01148_) );
  \$mux  #( .WIDTH(3) ) _45961_ ( .A(__tmp_585_1), .B(3'h0), .S(RST), .Y(_01263_) );
  \$mux  #( .WIDTH(3) ) _45962_ ( .A(_stream_conv2d_16_source_28_source_ram_raddr[2:0]), .B(3'h0), .S(RST), .Y(_01262_) );
  \$mux  #( .WIDTH(32) ) _45963_ ( .A(_stream_conv2d_16_source_27_source_pat_fsm_10), .B(2), .S(_06847_), .Y({ _18247_, _18246_, _18244_, _18243_, _18242_, _18241_, _18240_, _18239_, _18238_, _18237_, _18236_, _18235_, _18233_, _18232_, _18231_, _18230_, _18229_, _18228_, _18227_, _18226_, _18225_, _18224_, _18254_, _18253_, _18252_, _18251_, _18250_, _18249_, _18248_, _18245_, _18234_, _18223_ }) );
  \$mux  #( .WIDTH(32) ) _45964_ ( .A(_stream_conv2d_16_source_27_source_pat_fsm_10), .B(1), .S(_06736_), .Y({ _18279_, _18278_, _18276_, _18275_, _18274_, _18273_, _18272_, _18271_, _18270_, _18269_, _18268_, _18267_, _18265_, _18264_, _18263_, _18262_, _18261_, _18260_, _18259_, _18258_, _18257_, _18256_, _18286_, _18285_, _18284_, _18283_, _18282_, _18281_, _18280_, _18277_, _18266_, _18255_ }) );
  \$mux  #( .WIDTH(32) ) _45965_ ( .A(_24815_), .B(0), .S(RST), .Y(_02597_) );
  \$mux  #( .WIDTH(2) ) _45966_ ( .A(__tmp_575_1), .B(2'h0), .S(RST), .Y(_01260_) );
  \$mux  #( .WIDTH(2) ) _45967_ ( .A(_stream_conv2d_16_source_27_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01259_) );
  \$mux  #( .WIDTH(32) ) _45968_ ( .A(_stream_conv2d_16_source_26_source_pat_fsm_9), .B(2), .S(_06846_), .Y({ _18343_, _18342_, _18340_, _18339_, _18338_, _18337_, _18336_, _18335_, _18334_, _18333_, _18332_, _18331_, _18329_, _18328_, _18327_, _18326_, _18325_, _18324_, _18323_, _18322_, _18321_, _18320_, _18350_, _18349_, _18348_, _18347_, _18346_, _18345_, _18344_, _18341_, _18330_, _18319_ }) );
  \$mux  #( .WIDTH(32) ) _45969_ ( .A(_stream_conv2d_16_source_26_source_pat_fsm_9), .B(1), .S(_06731_), .Y({ _18375_, _18374_, _18372_, _18371_, _18370_, _18369_, _18368_, _18367_, _18366_, _18365_, _18364_, _18363_, _18361_, _18360_, _18359_, _18358_, _18357_, _18356_, _18355_, _18354_, _18353_, _18352_, _18382_, _18381_, _18380_, _18379_, _18378_, _18377_, _18376_, _18373_, _18362_, _18351_ }) );
  \$mux  #( .WIDTH(32) ) _45970_ ( .A(_24816_), .B(0), .S(RST), .Y(_02588_) );
  \$mux  #( .WIDTH(2) ) _45971_ ( .A(__tmp_565_1), .B(2'h0), .S(RST), .Y(_01257_) );
  \$mux  #( .WIDTH(2) ) _45972_ ( .A(_stream_conv2d_16_source_26_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01256_) );
  \$mux  #( .WIDTH(32) ) _45973_ ( .A(_stream_conv2d_16_source_25_source_pat_fsm_8), .B(2), .S(_06845_), .Y({ _18439_, _18438_, _18436_, _18435_, _18434_, _18433_, _18432_, _18431_, _18430_, _18429_, _18428_, _18427_, _18425_, _18424_, _18423_, _18422_, _18421_, _18420_, _18419_, _18418_, _18417_, _18416_, _18446_, _18445_, _18444_, _18443_, _18442_, _18441_, _18440_, _18437_, _18426_, _18415_ }) );
  \$mux  #( .WIDTH(32) ) _45974_ ( .A(_stream_conv2d_16_source_25_source_pat_fsm_8), .B(1), .S(_06726_), .Y({ _18471_, _18470_, _18468_, _18467_, _18466_, _18465_, _18464_, _18463_, _18462_, _18461_, _18460_, _18459_, _18457_, _18456_, _18455_, _18454_, _18453_, _18452_, _18451_, _18450_, _18449_, _18448_, _18478_, _18477_, _18476_, _18475_, _18474_, _18473_, _18472_, _18469_, _18458_, _18447_ }) );
  \$mux  #( .WIDTH(32) ) _45975_ ( .A(_24817_), .B(0), .S(RST), .Y(_02579_) );
  \$mux  #( .WIDTH(2) ) _45976_ ( .A(__tmp_555_1), .B(2'h0), .S(RST), .Y(_01254_) );
  \$mux  #( .WIDTH(2) ) _45977_ ( .A(_stream_conv2d_16_source_25_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01253_) );
  \$mux  #( .WIDTH(32) ) _45978_ ( .A(_stream_conv2d_16_source_24_source_pat_fsm_7), .B(2), .S(_06844_), .Y({ _18535_, _18534_, _18532_, _18531_, _18530_, _18529_, _18528_, _18527_, _18526_, _18525_, _18524_, _18523_, _18521_, _18520_, _18519_, _18518_, _18517_, _18516_, _18515_, _18514_, _18513_, _18512_, _18542_, _18541_, _18540_, _18539_, _18538_, _18537_, _18536_, _18533_, _18522_, _18511_ }) );
  \$mux  #( .WIDTH(32) ) _45979_ ( .A(_stream_conv2d_16_source_24_source_pat_fsm_7), .B(1), .S(_06721_), .Y({ _18567_, _18566_, _18564_, _18563_, _18562_, _18561_, _18560_, _18559_, _18558_, _18557_, _18556_, _18555_, _18553_, _18552_, _18551_, _18550_, _18549_, _18548_, _18547_, _18546_, _18545_, _18544_, _18574_, _18573_, _18572_, _18571_, _18570_, _18569_, _18568_, _18565_, _18554_, _18543_ }) );
  \$mux  #( .WIDTH(32) ) _45980_ ( .A(_24818_), .B(0), .S(RST), .Y(_02570_) );
  \$mux  #( .WIDTH(2) ) _45981_ ( .A(__tmp_545_1), .B(2'h0), .S(RST), .Y(_01251_) );
  \$mux  #( .WIDTH(2) ) _45982_ ( .A(_stream_conv2d_16_source_24_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01250_) );
  \$mux  #( .WIDTH(32) ) _45983_ ( .A(_stream_conv2d_16_source_23_source_pat_fsm_6), .B(2), .S(_06843_), .Y({ _18631_, _18630_, _18628_, _18627_, _18626_, _18625_, _18624_, _18623_, _18622_, _18621_, _18620_, _18619_, _18617_, _18616_, _18615_, _18614_, _18613_, _18612_, _18611_, _18610_, _18609_, _18608_, _18638_, _18637_, _18636_, _18635_, _18634_, _18633_, _18632_, _18629_, _18618_, _18607_ }) );
  \$mux  #( .WIDTH(32) ) _45984_ ( .A(_stream_conv2d_16_source_23_source_pat_fsm_6), .B(1), .S(_06716_), .Y({ _18663_, _18662_, _18660_, _18659_, _18658_, _18657_, _18656_, _18655_, _18654_, _18653_, _18652_, _18651_, _18649_, _18648_, _18647_, _18646_, _18645_, _18644_, _18643_, _18642_, _18641_, _18640_, _18670_, _18669_, _18668_, _18667_, _18666_, _18665_, _18664_, _18661_, _18650_, _18639_ }) );
  \$mux  #( .WIDTH(32) ) _45985_ ( .A(_24819_), .B(0), .S(RST), .Y(_02561_) );
  \$mux  #( .WIDTH(2) ) _45986_ ( .A(__tmp_535_1), .B(2'h0), .S(RST), .Y(_01248_) );
  \$mux  #( .WIDTH(2) ) _45987_ ( .A(_stream_conv2d_16_source_23_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01247_) );
  \$mux  #( .WIDTH(32) ) _45988_ ( .A(_stream_conv2d_16_source_22_source_pat_fsm_5), .B(2), .S(_06842_), .Y({ _18727_, _18726_, _18724_, _18723_, _18722_, _18721_, _18720_, _18719_, _18718_, _18717_, _18716_, _18715_, _18713_, _18712_, _18711_, _18710_, _18709_, _18708_, _18707_, _18706_, _18705_, _18704_, _18734_, _18733_, _18732_, _18731_, _18730_, _18729_, _18728_, _18725_, _18714_, _18703_ }) );
  \$mux  #( .WIDTH(32) ) _45989_ ( .A(_stream_conv2d_16_source_22_source_pat_fsm_5), .B(1), .S(_06711_), .Y({ _18759_, _18758_, _18756_, _18755_, _18754_, _18753_, _18752_, _18751_, _18750_, _18749_, _18748_, _18747_, _18745_, _18744_, _18743_, _18742_, _18741_, _18740_, _18739_, _18738_, _18737_, _18736_, _18766_, _18765_, _18764_, _18763_, _18762_, _18761_, _18760_, _18757_, _18746_, _18735_ }) );
  \$mux  #( .WIDTH(32) ) _45990_ ( .A(_24820_), .B(0), .S(RST), .Y(_02552_) );
  \$mux  #( .WIDTH(2) ) _45991_ ( .A(__tmp_525_1), .B(2'h0), .S(RST), .Y(_01245_) );
  \$mux  #( .WIDTH(2) ) _45992_ ( .A(_stream_conv2d_16_source_22_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01244_) );
  \$mux  #( .WIDTH(32) ) _45993_ ( .A(_stream_conv2d_16_source_21_source_pat_fsm_4), .B(2), .S(_06841_), .Y({ _18823_, _18822_, _18820_, _18819_, _18818_, _18817_, _18816_, _18815_, _18814_, _18813_, _18812_, _18811_, _18809_, _18808_, _18807_, _18806_, _18805_, _18804_, _18803_, _18802_, _18801_, _18800_, _18830_, _18829_, _18828_, _18827_, _18826_, _18825_, _18824_, _18821_, _18810_, _18799_ }) );
  \$mux  #( .WIDTH(32) ) _45994_ ( .A(_stream_conv2d_16_source_21_source_pat_fsm_4), .B(1), .S(_06706_), .Y({ _18855_, _18854_, _18852_, _18851_, _18850_, _18849_, _18848_, _18847_, _18846_, _18845_, _18844_, _18843_, _18841_, _18840_, _18839_, _18838_, _18837_, _18836_, _18835_, _18834_, _18833_, _18832_, _18862_, _18861_, _18860_, _18859_, _18858_, _18857_, _18856_, _18853_, _18842_, _18831_ }) );
  \$mux  #( .WIDTH(32) ) _45995_ ( .A(_24821_), .B(0), .S(RST), .Y(_02543_) );
  \$mux  #( .WIDTH(2) ) _45996_ ( .A(__tmp_515_1), .B(2'h0), .S(RST), .Y(_01242_) );
  \$mux  #( .WIDTH(2) ) _45997_ ( .A(_stream_conv2d_16_source_21_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01241_) );
  \$mux  #( .WIDTH(32) ) _45998_ ( .A(_stream_conv2d_16_source_20_source_pat_fsm_3), .B(2), .S(_06840_), .Y({ _18919_, _18918_, _18916_, _18915_, _18914_, _18913_, _18912_, _18911_, _18910_, _18909_, _18908_, _18907_, _18905_, _18904_, _18903_, _18902_, _18901_, _18900_, _18899_, _18898_, _18897_, _18896_, _18926_, _18925_, _18924_, _18923_, _18922_, _18921_, _18920_, _18917_, _18906_, _18895_ }) );
  \$mux  #( .WIDTH(32) ) _45999_ ( .A(_stream_conv2d_16_source_20_source_pat_fsm_3), .B(1), .S(_06701_), .Y({ _18951_, _18950_, _18948_, _18947_, _18946_, _18945_, _18944_, _18943_, _18942_, _18941_, _18940_, _18939_, _18937_, _18936_, _18935_, _18934_, _18933_, _18932_, _18931_, _18930_, _18929_, _18928_, _18958_, _18957_, _18956_, _18955_, _18954_, _18953_, _18952_, _18949_, _18938_, _18927_ }) );
  \$mux  #( .WIDTH(32) ) _46000_ ( .A(_24822_), .B(0), .S(RST), .Y(_02534_) );
  \$mux  #( .WIDTH(2) ) _46001_ ( .A(__tmp_1201_1), .B(2'h0), .S(RST), .Y(_01146_) );
  \$mux  #( .WIDTH(2) ) _46002_ ( .A(_stream_matmul_29_source_19_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01145_) );
  \$mux  #( .WIDTH(2) ) _46003_ ( .A(__tmp_505_1), .B(2'h0), .S(RST), .Y(_01239_) );
  \$mux  #( .WIDTH(2) ) _46004_ ( .A(_stream_conv2d_16_source_20_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01238_) );
  \$mux  #( .WIDTH(32) ) _46005_ ( .A(_stream_conv2d_16_source_19_source_pat_fsm_2), .B(2), .S(_06839_), .Y({ _19015_, _19014_, _19012_, _19011_, _19010_, _19009_, _19008_, _19007_, _19006_, _19005_, _19004_, _19003_, _19001_, _19000_, _18999_, _18998_, _18997_, _18996_, _18995_, _18994_, _18993_, _18992_, _19022_, _19021_, _19020_, _19019_, _19018_, _19017_, _19016_, _19013_, _19002_, _18991_ }) );
  \$mux  #( .WIDTH(32) ) _46006_ ( .A(_stream_conv2d_16_source_19_source_pat_fsm_2), .B(1), .S(_06696_), .Y({ _19047_, _19046_, _19044_, _19043_, _19042_, _19041_, _19040_, _19039_, _19038_, _19037_, _19036_, _19035_, _19033_, _19032_, _19031_, _19030_, _19029_, _19028_, _19027_, _19026_, _19025_, _19024_, _19054_, _19053_, _19052_, _19051_, _19050_, _19049_, _19048_, _19045_, _19034_, _19023_ }) );
  \$mux  #( .WIDTH(32) ) _46007_ ( .A(_24823_), .B(0), .S(RST), .Y(_02525_) );
  \$mux  #( .WIDTH(2) ) _46008_ ( .A(__tmp_1170_1), .B(2'h0), .S(RST), .Y(_01140_) );
  \$mux  #( .WIDTH(2) ) _46009_ ( .A(_stream_matmul_29_source_6_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01139_) );
  \$mux  #( .WIDTH(2) ) _46010_ ( .A(__tmp_495_1), .B(2'h0), .S(RST), .Y(_01236_) );
  \$mux  #( .WIDTH(2) ) _46011_ ( .A(_stream_conv2d_16_source_19_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01235_) );
  \$mux  #( .WIDTH(32) ) _46012_ ( .A(_stream_conv2d_16_source_8_source_pat_fsm_1), .B(2), .S(_06838_), .Y({ _19111_, _19110_, _19108_, _19107_, _19106_, _19105_, _19104_, _19103_, _19102_, _19101_, _19100_, _19099_, _19097_, _19096_, _19095_, _19094_, _19093_, _19092_, _19091_, _19090_, _19089_, _19088_, _19118_, _19117_, _19116_, _19115_, _19114_, _19113_, _19112_, _19109_, _19098_, _19087_ }) );
  \$mux  #( .WIDTH(32) ) _46013_ ( .A(_stream_conv2d_16_source_8_source_pat_fsm_1), .B(1), .S(_06691_), .Y({ _19143_, _19142_, _19140_, _19139_, _19138_, _19137_, _19136_, _19135_, _19134_, _19133_, _19132_, _19131_, _19129_, _19128_, _19127_, _19126_, _19125_, _19124_, _19123_, _19122_, _19121_, _19120_, _19150_, _19149_, _19148_, _19147_, _19146_, _19145_, _19144_, _19141_, _19130_, _19119_ }) );
  \$mux  #( .WIDTH(32) ) _46014_ ( .A(_24824_), .B(0), .S(RST), .Y(_02696_) );
  \$mux  #( .WIDTH(2) ) _46015_ ( .A(__tmp_1181_1), .B(2'h0), .S(RST), .Y(_01143_) );
  \$mux  #( .WIDTH(2) ) _46016_ ( .A(_stream_matmul_29_source_8_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01142_) );
  \$mux  #( .WIDTH(2) ) _46017_ ( .A(__tmp_475_1), .B(2'h0), .S(RST), .Y(_01233_) );
  \$mux  #( .WIDTH(2) ) _46018_ ( .A(_stream_conv2d_16_source_8_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01232_) );
  \$mux  #( .WIDTH(32) ) _46019_ ( .A(_stream_conv2d_16_source_6_source_pat_fsm_0), .B(2), .S(_06837_), .Y({ _19207_, _19206_, _19204_, _19203_, _19202_, _19201_, _19200_, _19199_, _19198_, _19197_, _19196_, _19195_, _19193_, _19192_, _19191_, _19190_, _19189_, _19188_, _19187_, _19186_, _19185_, _19184_, _19214_, _19213_, _19212_, _19211_, _19210_, _19209_, _19208_, _19205_, _19194_, _19183_ }) );
  \$mux  #( .WIDTH(32) ) _46020_ ( .A(_stream_conv2d_16_source_6_source_pat_fsm_0), .B(1), .S(_06686_), .Y({ _19239_, _19238_, _19236_, _19235_, _19234_, _19233_, _19232_, _19231_, _19230_, _19229_, _19228_, _19227_, _19225_, _19224_, _19223_, _19222_, _19221_, _19220_, _19219_, _19218_, _19217_, _19216_, _19246_, _19245_, _19244_, _19243_, _19242_, _19241_, _19240_, _19237_, _19226_, _19215_ }) );
  \$mux  #( .WIDTH(32) ) _46021_ ( .A(_24825_), .B(0), .S(RST), .Y(_02687_) );
  \$mux  #( .WIDTH(2) ) _46022_ ( .A(__tmp_1027_1), .B(2'h0), .S(RST), .Y(_01110_) );
  \$mux  #( .WIDTH(2) ) _46023_ ( .A(_stream_max_pool_serial_18_source_1_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01109_) );
  \$mux  #( .WIDTH(2) ) _46024_ ( .A(__tmp_464_1), .B(2'h0), .S(RST), .Y(_01230_) );
  \$mux  #( .WIDTH(2) ) _46025_ ( .A(_stream_conv2d_16_source_6_source_ram_raddr[1:0]), .B(2'h0), .S(RST), .Y(_01229_) );
  \$mux  #( .WIDTH(9) ) _46026_ ( .A({ conv2d_16_stream_pad_mask_2_2, conv2d_16_stream_pad_mask_2_1, conv2d_16_stream_pad_mask_2_0, conv2d_16_stream_pad_mask_1_2, conv2d_16_stream_pad_mask_1_1, conv2d_16_stream_pad_mask_1_0, conv2d_16_stream_pad_mask_0_2, conv2d_16_stream_pad_mask_0_1, conv2d_16_stream_pad_mask_0_0 }), .B(conv2d_16_stream_pad_masks), .S(_05990_), .Y(_24826_) );
  \$mux  #( .WIDTH(9) ) _46027_ ( .A(_24826_), .B(9'h000), .S(RST), .Y(_03276_) );
  \$mux  #( .WIDTH(32) ) _46028_ ( .A(conv2d_16_och_count), .B(conv2d_16_och_count_buf), .S(_05991_), .Y(_24827_) );
  \$mux  #( .WIDTH(32) ) _46029_ ( .A(_24827_), .B(0), .S(RST), .Y(_03241_) );
  \$mux  #( .WIDTH(2) ) _46030_ ( .A(conv2d_16_row_select), .B(conv2d_16_row_select_buf), .S(_05991_), .Y(_24828_) );
  \$mux  #( .WIDTH(2) ) _46031_ ( .A(_24828_), .B(2'h0), .S(RST), .Y(_03261_) );
  \$mux  #( .WIDTH(32) ) _46032_ ( .A(conv2d_16_row_count), .B(conv2d_16_row_count_buf), .S(_05991_), .Y(_24829_) );
  \$mux  #( .WIDTH(32) ) _46033_ ( .A(_24829_), .B(0), .S(RST), .Y(_03259_) );
  \$mux  #( .WIDTH(32) ) _46034_ ( .A(conv2d_16_out_page_comp_offset), .B(conv2d_16_out_page_comp_offset_buf), .S(_05991_), .Y(_24830_) );
  \$mux  #( .WIDTH(32) ) _46035_ ( .A(_24830_), .B(0), .S(RST), .Y(_03250_) );
  \$mux  #( .WIDTH(32) ) _46036_ ( .A(conv2d_16_act_page_comp_offset_2), .B(conv2d_16_act_page_comp_offset_buf_2), .S(_05991_), .Y(_24831_) );
  \$mux  #( .WIDTH(32) ) _46037_ ( .A(_24831_), .B(0), .S(RST), .Y(_03217_) );
  \$mux  #( .WIDTH(32) ) _46038_ ( .A(conv2d_16_act_page_comp_offset_1), .B(conv2d_16_act_page_comp_offset_buf_1), .S(_05991_), .Y(_24832_) );
  \$mux  #( .WIDTH(32) ) _46039_ ( .A(_24832_), .B(0), .S(RST), .Y(_03216_) );
  \$mux  #( .WIDTH(32) ) _46040_ ( .A(conv2d_16_act_page_comp_offset_0), .B(conv2d_16_act_page_comp_offset_buf_0), .S(_05991_), .Y(_24833_) );
  \$mux  #( .WIDTH(32) ) _46041_ ( .A(_24833_), .B(0), .S(RST), .Y(_03215_) );
  \$mux  #( .WIDTH(32) ) _46042_ ( .A(conv2d_16_filter_page_comp_offset), .B(conv2d_16_filter_page_comp_offset_buf), .S(_05991_), .Y(_24834_) );
  \$mux  #( .WIDTH(32) ) _46043_ ( .A(_24834_), .B(0), .S(RST), .Y(_03235_) );
  \$mux  #( .WIDTH(32) ) _46044_ ( .A(2), .B(0), .S(_06156_), .Y({ _19271_, _19270_, _19268_, _19267_, _19266_, _19265_, _19264_, _19263_, _19262_, _19261_, _19260_, _19259_, _19257_, _19256_, _19255_, _19254_, _19253_, _19252_, _19251_, _19250_, _19249_, _19248_, _19278_, _19277_, _19276_, _19275_, _19274_, _19273_, _19272_, _19269_, _19258_, _19247_ }) );
  \$mux  #( .WIDTH(32) ) _46045_ ( .A(5), .B(conv2d_16_comp_fsm), .S(_stream_conv2d_16_source_busy), .Y({ _19335_, _19334_, _19332_, _19331_, _19330_, _19329_, _19328_, _19327_, _19326_, _19325_, _19324_, _19323_, _19321_, _19320_, _19319_, _19318_, _19317_, _19316_, _19315_, _19314_, _19313_, _19312_, _19342_, _19341_, _19340_, _19339_, _19338_, _19337_, _19336_, _19333_, _19322_, _19311_ }) );
  \$mux  #( .WIDTH(32) ) _46046_ ( .A(conv2d_16_comp_fsm), .B(1), .S(_06836_), .Y({ _19367_, _19366_, _19364_, _19363_, _19362_, _19361_, _19360_, _19359_, _19358_, _19357_, _19356_, _19355_, _19353_, _19352_, _19351_, _19350_, _19349_, _19348_, _19347_, _19346_, _19345_, _19344_, _19374_, _19373_, _19372_, _19371_, _19370_, _19369_, _19368_, _19365_, _19354_, _19343_ }) );
  \$mux  #( .WIDTH(32) ) _46047_ ( .A(_24835_), .B(0), .S(RST), .Y(_03228_) );
  \$mux  #( .WIDTH(32) ) _46048_ ( .A(_24460_), .B(0), .S(_06156_), .Y({ _19399_, _19398_, _19396_, _19395_, _19394_, _19393_, _19392_, _19391_, _19390_, _19389_, _19388_, _19387_, _19385_, _19384_, _19383_, _19382_, _19381_, _19380_, _19379_, _19378_, _19377_, _19376_, _19406_, _19405_, _19404_, _19403_, _19402_, _19401_, _19400_, _19397_, _19386_, _19375_ }) );
  \$mux  #( .WIDTH(32) ) _46049_ ( .A(_24836_), .B(0), .S(RST), .Y(_03275_) );
  \$mux  #( .WIDTH(32) ) _46050_ ( .A(conv2d_16_stream_act_local_8), .B(_24459_), .S(_19439_), .Y(_24837_) );
  \$mux  #( .WIDTH(32) ) _46051_ ( .A(_24837_), .B({ cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset }), .S(_06156_), .Y({ _19464_, _19463_, _19461_, _19460_, _19459_, _19458_, _19457_, _19456_, _19455_, _19454_, _19453_, _19452_, _19450_, _19449_, _19448_, _19447_, _19446_, _19445_, _19444_, _19443_, _19442_, _19441_, _19471_, _19470_, _19469_, _19468_, _19467_, _19466_, _19465_, _19462_, _19451_, _19440_ }) );
  \$mux  #( .WIDTH(32) ) _46052_ ( .A(_24838_), .B(0), .S(RST), .Y(_03274_) );
  \$mux  #( .WIDTH(32) ) _46053_ ( .A(conv2d_16_stream_act_local_7), .B(_24458_), .S(_19504_), .Y(_24839_) );
  \$mux  #( .WIDTH(32) ) _46054_ ( .A(_24839_), .B(0), .S(_06156_), .Y({ _19529_, _19528_, _19526_, _19525_, _19524_, _19523_, _19522_, _19521_, _19520_, _19519_, _19518_, _19517_, _19515_, _19514_, _19513_, _19512_, _19511_, _19510_, _19509_, _19508_, _19507_, _19506_, _19536_, _19535_, _19534_, _19533_, _19532_, _19531_, _19530_, _19527_, _19516_, _19505_ }) );
  \$mux  #( .WIDTH(32) ) _46055_ ( .A(_24840_), .B(0), .S(RST), .Y(_03273_) );
  \$mux  #( .WIDTH(32) ) _46056_ ( .A(conv2d_16_stream_act_local_6), .B(_24457_), .S(_19569_), .Y(_24841_) );
  \$mux  #( .WIDTH(32) ) _46057_ ( .A(_24841_), .B(0), .S(_06156_), .Y({ _19594_, _19593_, _19591_, _19590_, _19589_, _19588_, _19587_, _19586_, _19585_, _19584_, _19583_, _19582_, _19580_, _19579_, _19578_, _19577_, _19576_, _19575_, _19574_, _19573_, _19572_, _19571_, _19601_, _19600_, _19599_, _19598_, _19597_, _19596_, _19595_, _19592_, _19581_, _19570_ }) );
  \$mux  #( .WIDTH(32) ) _46058_ ( .A(_24842_), .B(0), .S(RST), .Y(_03272_) );
  \$mux  #( .WIDTH(32) ) _46059_ ( .A(conv2d_16_stream_act_local_5), .B(_24456_), .S(_19439_), .Y(_24843_) );
  \$mux  #( .WIDTH(32) ) _46060_ ( .A(_24843_), .B({ cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset }), .S(_06156_), .Y({ _19658_, _19657_, _19655_, _19654_, _19653_, _19652_, _19651_, _19650_, _19649_, _19648_, _19647_, _19646_, _19644_, _19643_, _19642_, _19641_, _19640_, _19639_, _19638_, _19637_, _19636_, _19635_, _19665_, _19664_, _19663_, _19662_, _19661_, _19660_, _19659_, _19656_, _19645_, _19634_ }) );
  \$mux  #( .WIDTH(32) ) _46061_ ( .A(_24844_), .B(0), .S(RST), .Y(_03271_) );
  \$mux  #( .WIDTH(32) ) _46062_ ( .A(conv2d_16_stream_act_local_4), .B(_24455_), .S(_19504_), .Y(_24845_) );
  \$mux  #( .WIDTH(32) ) _46063_ ( .A(_24845_), .B(0), .S(_06156_), .Y({ _19722_, _19721_, _19719_, _19718_, _19717_, _19716_, _19715_, _19714_, _19713_, _19712_, _19711_, _19710_, _19708_, _19707_, _19706_, _19705_, _19704_, _19703_, _19702_, _19701_, _19700_, _19699_, _19729_, _19728_, _19727_, _19726_, _19725_, _19724_, _19723_, _19720_, _19709_, _19698_ }) );
  \$mux  #( .WIDTH(32) ) _46064_ ( .A(_24846_), .B(0), .S(RST), .Y(_03270_) );
  \$mux  #( .WIDTH(32) ) _46065_ ( .A(conv2d_16_stream_act_local_3), .B(_24454_), .S(_19569_), .Y(_24847_) );
  \$mux  #( .WIDTH(32) ) _46066_ ( .A(_24847_), .B(0), .S(_06156_), .Y({ _19786_, _19785_, _19783_, _19782_, _19781_, _19780_, _19779_, _19778_, _19777_, _19776_, _19775_, _19774_, _19772_, _19771_, _19770_, _19769_, _19768_, _19767_, _19766_, _19765_, _19764_, _19763_, _19793_, _19792_, _19791_, _19790_, _19789_, _19788_, _19787_, _19784_, _19773_, _19762_ }) );
  \$mux  #( .WIDTH(32) ) _46067_ ( .A(_24848_), .B(0), .S(RST), .Y(_03269_) );
  \$mux  #( .WIDTH(32) ) _46068_ ( .A(conv2d_16_stream_act_local_2), .B(_24453_), .S(_19439_), .Y(_24849_) );
  \$mux  #( .WIDTH(32) ) _46069_ ( .A(_24849_), .B({ cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset[6], cparam_conv2d_16_stream_act_local_large_offset }), .S(_06156_), .Y({ _19850_, _19849_, _19847_, _19846_, _19845_, _19844_, _19843_, _19842_, _19841_, _19840_, _19839_, _19838_, _19836_, _19835_, _19834_, _19833_, _19832_, _19831_, _19830_, _19829_, _19828_, _19827_, _19857_, _19856_, _19855_, _19854_, _19853_, _19852_, _19851_, _19848_, _19837_, _19826_ }) );
  \$mux  #( .WIDTH(32) ) _46070_ ( .A(_24850_), .B(0), .S(RST), .Y(_03268_) );
  \$mux  #( .WIDTH(32) ) _46071_ ( .A(conv2d_16_stream_act_local_1), .B(_24452_), .S(_19504_), .Y(_24851_) );
  \$mux  #( .WIDTH(32) ) _46072_ ( .A(_24851_), .B(0), .S(_06156_), .Y({ _19914_, _19913_, _19911_, _19910_, _19909_, _19908_, _19907_, _19906_, _19905_, _19904_, _19903_, _19902_, _19900_, _19899_, _19898_, _19897_, _19896_, _19895_, _19894_, _19893_, _19892_, _19891_, _19921_, _19920_, _19919_, _19918_, _19917_, _19916_, _19915_, _19912_, _19901_, _19890_ }) );
  \$mux  #( .WIDTH(32) ) _46073_ ( .A(_24852_), .B(0), .S(RST), .Y(_03267_) );
  \$mux  #( .WIDTH(32) ) _46074_ ( .A(conv2d_16_stream_act_local_0), .B(_24451_), .S(_19569_), .Y(_24853_) );
  \$mux  #( .WIDTH(32) ) _46075_ ( .A(_24853_), .B(0), .S(_06156_), .Y({ _19978_, _19977_, _19975_, _19974_, _19973_, _19972_, _19971_, _19970_, _19969_, _19968_, _19967_, _19966_, _19964_, _19963_, _19962_, _19961_, _19960_, _19959_, _19958_, _19957_, _19956_, _19955_, _19985_, _19984_, _19983_, _19982_, _19981_, _19980_, _19979_, _19976_, _19965_, _19954_ }) );
  \$mux  #( .WIDTH(32) ) _46076_ ( .A(_24854_), .B(0), .S(RST), .Y(_03266_) );
  \$mux  #( .WIDTH(2) ) _46077_ ( .A(_24462_), .B(_28939_), .S(_06157_), .Y(_24855_) );
  \$mux  #( .WIDTH(2) ) _46078_ ( .A(_24855_), .B(2'h2), .S(_06156_), .Y({ _20019_, _20018_ }) );
  \$mux  #( .WIDTH(2) ) _46079_ ( .A(_24856_), .B(2'h0), .S(RST), .Y(_03227_) );
  \$mux  #( .WIDTH(32) ) _46080_ ( .A(_24461_), .B(0), .S(_06156_), .Y({ _20046_, _20045_, _20043_, _20042_, _20041_, _20040_, _20039_, _20038_, _20037_, _20036_, _20035_, _20034_, _20032_, _20031_, _20030_, _20029_, _20028_, _20027_, _20026_, _20025_, _20024_, _20023_, _20053_, _20052_, _20051_, _20050_, _20049_, _20048_, _20047_, _20044_, _20033_, _20022_ }) );
  \$mux  #( .WIDTH(32) ) _46081_ ( .A(_24857_), .B(0), .S(RST), .Y(_03226_) );
  \$mux  #( .WIDTH(32) ) _46082_ ( .A(conv2d_16_sync_comp_count), .B(_24450_), .S(_stream_conv2d_16_end_flag), .Y(_24858_) );
  \$mux  #( .WIDTH(32) ) _46083_ ( .A(0), .B(_24858_), .S(_06018_), .Y(_24859_) );
  \$mux  #( .WIDTH(32) ) _46084_ ( .A(_24859_), .B(0), .S(RST), .Y(_03277_) );
  \$mux  #( .WIDTH(32) ) _46085_ ( .A({ 25'h0000000, cparam_conv2d_16_bias_num }), .B(conv2d_16_next_stream_num_ops), .S(_05991_), .Y(_24860_) );
  \$mux  #( .WIDTH(32) ) _46086_ ( .A(_24860_), .B(0), .S(RST), .Y(_03238_) );
  \$mux  #( .WIDTH(9) ) _46087_ ( .A(req_block_size_400), .B({ 5'h00, cparam_conv2d_16_inc_act_laddr_large[5:2] }), .S(set_req_401), .Y(_24861_) );
  \$mux  #( .WIDTH(9) ) _46088_ ( .A(_24861_), .B(9'h000), .S(_RESETN_inv_2), .Y(_03872_) );
  \$mux  #( .WIDTH(9) ) _46089_ ( .A(req_block_size_343), .B({ 5'h00, cparam_conv2d_16_inc_act_laddr_large[5:2] }), .S(set_req_344), .Y(_24862_) );
  \$mux  #( .WIDTH(9) ) _46090_ ( .A(_24862_), .B(9'h000), .S(_RESETN_inv_2), .Y(_03871_) );
  \$mux  #( .WIDTH(9) ) _46091_ ( .A(req_block_size_286), .B({ 5'h00, cparam_conv2d_16_inc_act_laddr_large[5:2] }), .S(set_req_287), .Y(_24863_) );
  \$mux  #( .WIDTH(9) ) _46092_ ( .A(_24863_), .B(9'h000), .S(_RESETN_inv_2), .Y(_03869_) );
  \$mux  #( .WIDTH(10) ) _46093_ ( .A(req_block_size_33), .B({ 7'h00, cparam_conv2d_16_filter_read_block[5:3] }), .S(set_req_34), .Y(_24864_) );
  \$mux  #( .WIDTH(10) ) _46094_ ( .A(_24864_), .B(10'h000), .S(_RESETN_inv_2), .Y(_03870_) );
  \$mux  #( .WIDTH(1) ) _46095_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_9_1), .S(_05995_), .Y(_24865_) );
  \$mux  #( .WIDTH(1) ) _46096_ ( .A(_24865_), .B(1'h0), .S(_RESETN_inv_2), .Y(_00689_) );
  \$mux  #( .WIDTH(1) ) _46097_ ( .A(_wvalid_1154), .B(1'h0), .S(__maxi_read_fsm_cond_3_9_1), .Y(_24866_) );
  \$mux  #( .WIDTH(1) ) _46098_ ( .A(_24866_), .B(_wvalid_1154), .S(_05993_), .Y(_24867_) );
  \$mux  #( .WIDTH(1) ) _46099_ ( .A(_24867_), .B(1'h1), .S(_06833_), .Y(_24868_) );
  \$mux  #( .WIDTH(1) ) _46100_ ( .A(_24868_), .B(_24867_), .S(_05995_), .Y(_24869_) );
  \$mux  #( .WIDTH(1) ) _46101_ ( .A(_24869_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03183_) );
  \$mux  #( .WIDTH(32) ) _46102_ ( .A(_wdata_1153), .B(maxi_rdata), .S(_06833_), .Y(_24870_) );
  \$mux  #( .WIDTH(32) ) _46103_ ( .A(_24870_), .B(_wdata_1153), .S(_05995_), .Y(_24871_) );
  \$mux  #( .WIDTH(32) ) _46104_ ( .A(_24871_), .B(0), .S(_RESETN_inv_2), .Y(_03175_) );
  \$mux  #( .WIDTH(1) ) _46105_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_8_1), .S(_05995_), .Y(_24872_) );
  \$mux  #( .WIDTH(1) ) _46106_ ( .A(_24872_), .B(1'h0), .S(_RESETN_inv_2), .Y(_00688_) );
  \$mux  #( .WIDTH(1) ) _46107_ ( .A(_wvalid_1135), .B(1'h0), .S(__maxi_read_fsm_cond_3_8_1), .Y(_24873_) );
  \$mux  #( .WIDTH(1) ) _46108_ ( .A(_24873_), .B(_wvalid_1135), .S(_05993_), .Y(_24874_) );
  \$mux  #( .WIDTH(1) ) _46109_ ( .A(_24874_), .B(1'h1), .S(_06832_), .Y(_24875_) );
  \$mux  #( .WIDTH(1) ) _46110_ ( .A(_24875_), .B(_24874_), .S(_05995_), .Y(_24876_) );
  \$mux  #( .WIDTH(1) ) _46111_ ( .A(_24876_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03182_) );
  \$mux  #( .WIDTH(32) ) _46112_ ( .A(_wdata_1134), .B(maxi_rdata), .S(_06832_), .Y(_24877_) );
  \$mux  #( .WIDTH(32) ) _46113_ ( .A(_24877_), .B(_wdata_1134), .S(_05995_), .Y(_24878_) );
  \$mux  #( .WIDTH(32) ) _46114_ ( .A(_24878_), .B(0), .S(_RESETN_inv_2), .Y(_03174_) );
  \$mux  #( .WIDTH(1) ) _46115_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_7_1), .S(_05995_), .Y(_24879_) );
  \$mux  #( .WIDTH(1) ) _46116_ ( .A(_24879_), .B(1'h0), .S(_RESETN_inv_2), .Y(_00687_) );
  \$mux  #( .WIDTH(1) ) _46117_ ( .A(_wvalid_1123), .B(1'h0), .S(__maxi_read_fsm_cond_3_7_1), .Y(_24880_) );
  \$mux  #( .WIDTH(1) ) _46118_ ( .A(_24880_), .B(_wvalid_1123), .S(_05993_), .Y(_24881_) );
  \$mux  #( .WIDTH(1) ) _46119_ ( .A(_24881_), .B(1'h1), .S(_06831_), .Y(_24882_) );
  \$mux  #( .WIDTH(1) ) _46120_ ( .A(_24882_), .B(_24881_), .S(_05995_), .Y(_24883_) );
  \$mux  #( .WIDTH(1) ) _46121_ ( .A(_24883_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03181_) );
  \$mux  #( .WIDTH(32) ) _46122_ ( .A(_wdata_1122), .B(maxi_rdata), .S(_06831_), .Y(_24884_) );
  \$mux  #( .WIDTH(32) ) _46123_ ( .A(_24884_), .B(_wdata_1122), .S(_05995_), .Y(_24885_) );
  \$mux  #( .WIDTH(32) ) _46124_ ( .A(_24885_), .B(0), .S(_RESETN_inv_2), .Y(_03173_) );
  \$mux  #( .WIDTH(1) ) _46125_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_6_1), .S(_05995_), .Y(_24886_) );
  \$mux  #( .WIDTH(1) ) _46126_ ( .A(_24886_), .B(1'h0), .S(_RESETN_inv_2), .Y(_00686_) );
  \$mux  #( .WIDTH(1) ) _46127_ ( .A(_wvalid_404), .B(1'h0), .S(__maxi_read_fsm_cond_3_6_1), .Y(_24887_) );
  \$mux  #( .WIDTH(1) ) _46128_ ( .A(_24887_), .B(_wvalid_404), .S(_05993_), .Y(_24888_) );
  \$mux  #( .WIDTH(1) ) _46129_ ( .A(_24888_), .B(1'h1), .S(_06830_), .Y(_24889_) );
  \$mux  #( .WIDTH(1) ) _46130_ ( .A(_24889_), .B(_24888_), .S(_05995_), .Y(_24890_) );
  \$mux  #( .WIDTH(1) ) _46131_ ( .A(_24890_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03189_) );
  \$mux  #( .WIDTH(32) ) _46132_ ( .A(_wdata_403), .B(maxi_rdata), .S(_06830_), .Y(_24891_) );
  \$mux  #( .WIDTH(32) ) _46133_ ( .A(_24891_), .B(_wdata_403), .S(_05995_), .Y(_24892_) );
  \$mux  #( .WIDTH(32) ) _46134_ ( .A(_24892_), .B(0), .S(_RESETN_inv_2), .Y(_03180_) );
  \$mux  #( .WIDTH(1) ) _46135_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_5_1), .S(_05995_), .Y(_24893_) );
  \$mux  #( .WIDTH(1) ) _46136_ ( .A(_24893_), .B(1'h0), .S(_RESETN_inv_2), .Y(_00685_) );
  \$mux  #( .WIDTH(1) ) _46137_ ( .A(_wvalid_347), .B(1'h0), .S(__maxi_read_fsm_cond_3_5_1), .Y(_24894_) );
  \$mux  #( .WIDTH(1) ) _46138_ ( .A(_24894_), .B(_wvalid_347), .S(_05993_), .Y(_24895_) );
  \$mux  #( .WIDTH(1) ) _46139_ ( .A(_24895_), .B(1'h1), .S(_06829_), .Y(_24896_) );
  \$mux  #( .WIDTH(1) ) _46140_ ( .A(_24896_), .B(_24895_), .S(_05995_), .Y(_24897_) );
  \$mux  #( .WIDTH(1) ) _46141_ ( .A(_24897_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03187_) );
  \$mux  #( .WIDTH(32) ) _46142_ ( .A(_wdata_346), .B(maxi_rdata), .S(_06829_), .Y(_24898_) );
  \$mux  #( .WIDTH(32) ) _46143_ ( .A(_24898_), .B(_wdata_346), .S(_05995_), .Y(_24899_) );
  \$mux  #( .WIDTH(32) ) _46144_ ( .A(_24899_), .B(0), .S(_RESETN_inv_2), .Y(_03178_) );
  \$mux  #( .WIDTH(1) ) _46145_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_4_1), .S(_05995_), .Y(_24900_) );
  \$mux  #( .WIDTH(1) ) _46146_ ( .A(_24900_), .B(1'h0), .S(_RESETN_inv_2), .Y(_00684_) );
  \$mux  #( .WIDTH(1) ) _46147_ ( .A(_wvalid_290), .B(1'h0), .S(__maxi_read_fsm_cond_3_4_1), .Y(_24901_) );
  \$mux  #( .WIDTH(1) ) _46148_ ( .A(_24901_), .B(_wvalid_290), .S(_05993_), .Y(_24902_) );
  \$mux  #( .WIDTH(1) ) _46149_ ( .A(_24902_), .B(1'h1), .S(_06828_), .Y(_24903_) );
  \$mux  #( .WIDTH(1) ) _46150_ ( .A(_24903_), .B(_24902_), .S(_05995_), .Y(_24904_) );
  \$mux  #( .WIDTH(1) ) _46151_ ( .A(_24904_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03186_) );
  \$mux  #( .WIDTH(32) ) _46152_ ( .A(_wdata_289), .B(maxi_rdata), .S(_06828_), .Y(_24905_) );
  \$mux  #( .WIDTH(32) ) _46153_ ( .A(_24905_), .B(_wdata_289), .S(_05995_), .Y(_24906_) );
  \$mux  #( .WIDTH(32) ) _46154_ ( .A(_24906_), .B(0), .S(_RESETN_inv_2), .Y(_03177_) );
  \$mux  #( .WIDTH(1) ) _46155_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_3_1), .S(_05995_), .Y(_24907_) );
  \$mux  #( .WIDTH(1) ) _46156_ ( .A(_24907_), .B(1'h0), .S(_RESETN_inv_2), .Y(_00683_) );
  \$mux  #( .WIDTH(1) ) _46157_ ( .A(_wvalid_37), .B(1'h0), .S(__maxi_read_fsm_cond_3_3_1), .Y(_24908_) );
  \$mux  #( .WIDTH(1) ) _46158_ ( .A(_24908_), .B(_wvalid_37), .S(_05993_), .Y(_24909_) );
  \$mux  #( .WIDTH(1) ) _46159_ ( .A(_24909_), .B(1'h1), .S(_06827_), .Y(_24910_) );
  \$mux  #( .WIDTH(1) ) _46160_ ( .A(_24910_), .B(_24909_), .S(_05995_), .Y(_24911_) );
  \$mux  #( .WIDTH(1) ) _46161_ ( .A(_24911_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03188_) );
  \$mux  #( .WIDTH(32) ) _46162_ ( .A(_wdata_36), .B(maxi_rdata), .S(_06827_), .Y(_24912_) );
  \$mux  #( .WIDTH(32) ) _46163_ ( .A(_24912_), .B(_wdata_36), .S(_05995_), .Y(_24913_) );
  \$mux  #( .WIDTH(32) ) _46164_ ( .A(_24913_), .B(0), .S(_RESETN_inv_2), .Y(_03179_) );
  \$mux  #( .WIDTH(1) ) _46165_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_2_1), .S(_05995_), .Y(_24914_) );
  \$mux  #( .WIDTH(1) ) _46166_ ( .A(_24914_), .B(1'h0), .S(_RESETN_inv_2), .Y(_00682_) );
  \$mux  #( .WIDTH(1) ) _46167_ ( .A(_wvalid_24), .B(1'h0), .S(__maxi_read_fsm_cond_3_2_1), .Y(_24915_) );
  \$mux  #( .WIDTH(1) ) _46168_ ( .A(_24915_), .B(_wvalid_24), .S(_05993_), .Y(_24916_) );
  \$mux  #( .WIDTH(1) ) _46169_ ( .A(_24916_), .B(1'h1), .S(_06826_), .Y(_24917_) );
  \$mux  #( .WIDTH(1) ) _46170_ ( .A(_24917_), .B(_24916_), .S(_05995_), .Y(_24918_) );
  \$mux  #( .WIDTH(1) ) _46171_ ( .A(_24918_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03185_) );
  \$mux  #( .WIDTH(32) ) _46172_ ( .A(_wdata_23), .B(maxi_rdata), .S(_06826_), .Y(_24919_) );
  \$mux  #( .WIDTH(32) ) _46173_ ( .A(_24919_), .B(_wdata_23), .S(_05995_), .Y(_24920_) );
  \$mux  #( .WIDTH(32) ) _46174_ ( .A(_24920_), .B(0), .S(_RESETN_inv_2), .Y(_03176_) );
  \$mux  #( .WIDTH(1) ) _46175_ ( .A(1'h1), .B(__maxi_read_fsm_cond_4_1_1), .S(_05994_), .Y(_24921_) );
  \$mux  #( .WIDTH(1) ) _46176_ ( .A(_24921_), .B(1'h0), .S(_RESETN_inv_2), .Y(_00690_) );
  \$mux  #( .WIDTH(1) ) _46177_ ( .A(axim_flag_21), .B(1'h0), .S(__maxi_read_fsm_cond_4_1_1), .Y(_24922_) );
  \$mux  #( .WIDTH(1) ) _46178_ ( .A(_24922_), .B(axim_flag_21), .S(_05992_), .Y(_24923_) );
  \$mux  #( .WIDTH(1) ) _46179_ ( .A(1'h1), .B(_24923_), .S(_05994_), .Y(_24924_) );
  \$mux  #( .WIDTH(1) ) _46180_ ( .A(_24924_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03199_) );
  \$mux  #( .WIDTH(1) ) _46181_ ( .A(1'h1), .B(__maxi_read_fsm_cond_3_0_1), .S(_05995_), .Y(_24925_) );
  \$mux  #( .WIDTH(1) ) _46182_ ( .A(_24925_), .B(1'h0), .S(_RESETN_inv_2), .Y(_00681_) );
  \$mux  #( .WIDTH(32) ) _46183_ ( .A(_maxi_read_fsm), .B(0), .S(_RESETN_inv_2), .Y(_01581_) );
  \$mux  #( .WIDTH(1) ) _46184_ ( .A(_wvalid_11), .B(1'h0), .S(__maxi_read_fsm_cond_3_0_1), .Y(_24926_) );
  \$mux  #( .WIDTH(1) ) _46185_ ( .A(_24926_), .B(_wvalid_11), .S(_05993_), .Y(_24927_) );
  \$mux  #( .WIDTH(1) ) _46186_ ( .A(_24927_), .B(1'h1), .S(_06824_), .Y(_24928_) );
  \$mux  #( .WIDTH(1) ) _46187_ ( .A(_24928_), .B(_24927_), .S(_05995_), .Y(_24929_) );
  \$mux  #( .WIDTH(1) ) _46188_ ( .A(_24929_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03184_) );
  \$mux  #( .WIDTH(32) ) _46189_ ( .A(_wdata_10), .B(maxi_rdata), .S(_06824_), .Y(_24930_) );
  \$mux  #( .WIDTH(32) ) _46190_ ( .A(_24930_), .B(_wdata_10), .S(_05995_), .Y(_24931_) );
  \$mux  #( .WIDTH(32) ) _46191_ ( .A(_24931_), .B(0), .S(_RESETN_inv_2), .Y(_03172_) );
  \$mux  #( .WIDTH(33) ) _46192_ ( .A(_28938_), .B(_28937_), .S(_06155_), .Y(_24932_) );
  \$mux  #( .WIDTH(33) ) _46193_ ( .A(_24932_), .B(33'h000000000), .S(_06175_), .Y(_24933_) );
  \$mux  #( .WIDTH(33) ) _46194_ ( .A(_24933_), .B(_28937_), .S(_06823_), .Y({ _20111_, _20110_, _20109_, _20107_, _20106_, _20105_, _20104_, _20103_, _20102_, _20101_, _20100_, _20099_, _20098_, _20096_, _20095_, _20094_, _20093_, _20092_, _20091_, _20090_, _20089_, _20088_, _20087_, _20118_, _20117_, _20116_, _20115_, _20114_, _20113_, _20112_, _20108_, _20097_, _20086_ }) );
  \$mux  #( .WIDTH(33) ) _46195_ ( .A(_maxi_read_rest_size), .B(_maxi_read_size), .S(_maxi_read_start), .Y({ _20177_, _20176_, _20175_, _20173_, _20172_, _20171_, _20170_, _20169_, _20168_, _20167_, _20166_, _20165_, _20164_, _20162_, _20161_, _20160_, _20159_, _20158_, _20157_, _20156_, _20155_, _20154_, _20153_, _20184_, _20183_, _20182_, _20181_, _20180_, _20179_, _20178_, _20174_, _20163_, _20152_ }) );
  \$mux  #( .WIDTH(33) ) _46196_ ( .A(_24934_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01786_) );
  \$mux  #( .WIDTH(33) ) _46197_ ( .A(33'h000000100), .B({ 2'h0, _28519_[30:0] }), .S(_06155_), .Y(_24935_) );
  \$mux  #( .WIDTH(33) ) _46198_ ( .A(_24935_), .B(_maxi_read_rest_size), .S(_06175_), .Y(_24936_) );
  \$mux  #( .WIDTH(33) ) _46199_ ( .A(_24936_), .B({ 2'h0, _28519_[30:0] }), .S(_06823_), .Y(_24937_) );
  \$mux  #( .WIDTH(33) ) _46200_ ( .A(_24937_), .B(_maxi_read_cur_size), .S(_05996_), .Y(_24938_) );
  \$mux  #( .WIDTH(33) ) _46201_ ( .A(_24938_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01779_) );
  \$mux  #( .WIDTH(32) ) _46202_ ( .A(_maxi_read_cur_global_addr), .B(_24449_[31:0]), .S(_06825_), .Y({ _20209_, _20208_, _20206_, _20205_, _20204_, _20203_, _20202_, _20201_, _20200_, _20199_, _20198_, _20197_, _20195_, _20194_, _20193_, _20192_, _20191_, _20190_, _20189_, _20188_, _20187_, _20186_, _20216_, _20215_, _20214_, _20213_, _20212_, _20211_, _20210_, _20207_, _20196_, _20185_ }) );
  \$mux  #( .WIDTH(32) ) _46203_ ( .A(_maxi_read_cur_global_addr), .B({ _24448_[31:2], 2'h0 }), .S(_maxi_read_start), .Y({ _20273_, _20272_, _20270_, _20269_, _20268_, _20267_, _20266_, _20265_, _20264_, _20263_, _20262_, _20261_, _20259_, _20258_, _20257_, _20256_, _20255_, _20254_, _20253_, _20252_, _20251_, _20250_, _20280_, _20279_, _20278_, _20277_, _20276_, _20275_, _20274_, _20271_, _20260_, _20249_ }) );
  \$mux  #( .WIDTH(32) ) _46204_ ( .A(_24939_), .B(0), .S(_RESETN_inv_2), .Y(_01778_) );
  \$mux  #( .WIDTH(32) ) _46205_ ( .A(_maxi_read_fsm), .B(1), .S(_06834_), .Y(_24941_) );
  \$mux  #( .WIDTH(32) ) _46206_ ( .A(_24941_), .B(4), .S(_06835_), .Y({ _20337_, _20336_, _20334_, _20333_, _20332_, _20331_, _20330_, _20329_, _20328_, _20327_, _20326_, _20325_, _20323_, _20322_, _20321_, _20320_, _20319_, _20318_, _20317_, _20316_, _20315_, _20314_, _20344_, _20343_, _20342_, _20341_, _20340_, _20339_, _20338_, _20335_, _20324_, _20313_ }) );
  \$mux  #( .WIDTH(32) ) _46207_ ( .A(_maxi_read_fsm), .B(3), .S(_06875_), .Y({ _20369_, _20368_, _20366_, _20365_, _20364_, _20363_, _20362_, _20361_, _20360_, _20359_, _20358_, _20357_, _20355_, _20354_, _20353_, _20352_, _20351_, _20350_, _20349_, _20348_, _20347_, _20346_, _20376_, _20375_, _20374_, _20373_, _20372_, _20371_, _20370_, _20367_, _20356_, _20345_ }) );
  \$mux  #( .WIDTH(32) ) _46208_ ( .A(_maxi_read_fsm), .B(1), .S(_06518_), .Y(_24942_) );
  \$mux  #( .WIDTH(32) ) _46209_ ( .A(_24942_), .B(1), .S(_06482_), .Y(_24943_) );
  \$mux  #( .WIDTH(32) ) _46210_ ( .A(_24943_), .B(1), .S(_06360_), .Y(_24944_) );
  \$mux  #( .WIDTH(32) ) _46211_ ( .A(_24944_), .B(1), .S(_06554_), .Y(_24945_) );
  \$mux  #( .WIDTH(32) ) _46212_ ( .A(_24945_), .B(1), .S(_06601_), .Y(_24946_) );
  \$mux  #( .WIDTH(32) ) _46213_ ( .A(_24946_), .B(1), .S(_06630_), .Y(_24947_) );
  \$mux  #( .WIDTH(32) ) _46214_ ( .A(_24947_), .B(1), .S(_06562_), .Y(_24948_) );
  \$mux  #( .WIDTH(32) ) _46215_ ( .A(_24948_), .B(1), .S(_06374_), .Y(_24949_) );
  \$mux  #( .WIDTH(32) ) _46216_ ( .A(_24949_), .B(1), .S(_06592_), .Y({ _20401_, _20400_, _20398_, _20397_, _20396_, _20395_, _20394_, _20393_, _20392_, _20391_, _20390_, _20389_, _20387_, _20386_, _20385_, _20384_, _20383_, _20382_, _20381_, _20380_, _20379_, _20378_, _20408_, _20407_, _20406_, _20405_, _20404_, _20403_, _20402_, _20399_, _20388_, _20377_ }) );
  \$mux  #( .WIDTH(32) ) _46217_ ( .A(_24940_), .B(0), .S(_RESETN_inv_2), .Y(_01780_) );
  \$mux  #( .WIDTH(1) ) _46218_ ( .A(1'h1), .B(_control_conv2d_16_cond_48_10_1), .S(_06009_), .Y(_24950_) );
  \$mux  #( .WIDTH(1) ) _46219_ ( .A(_24950_), .B(1'h0), .S(RST), .Y(_01569_) );
  \$mux  #( .WIDTH(1) ) _46220_ ( .A(axim_flag_970), .B(1'h0), .S(_control_conv2d_16_cond_48_10_1), .Y(_24951_) );
  \$mux  #( .WIDTH(1) ) _46221_ ( .A(_24951_), .B(axim_flag_970), .S(_05997_), .Y(_24952_) );
  \$mux  #( .WIDTH(1) ) _46222_ ( .A(1'h1), .B(_24952_), .S(_06009_), .Y(_24953_) );
  \$mux  #( .WIDTH(1) ) _46223_ ( .A(_24953_), .B(1'h0), .S(RST), .Y(_03205_) );
  \$mux  #( .WIDTH(1) ) _46224_ ( .A(1'h1), .B(_control_conv2d_16_cond_38_9_1), .S(_06010_), .Y(_24954_) );
  \$mux  #( .WIDTH(1) ) _46225_ ( .A(_24954_), .B(1'h0), .S(RST), .Y(_01567_) );
  \$mux  #( .WIDTH(1) ) _46226_ ( .A(axim_flag_402), .B(1'h0), .S(_control_conv2d_16_cond_38_9_1), .Y(_24955_) );
  \$mux  #( .WIDTH(1) ) _46227_ ( .A(_24955_), .B(axim_flag_402), .S(_05998_), .Y(_24956_) );
  \$mux  #( .WIDTH(1) ) _46228_ ( .A(1'h1), .B(_24956_), .S(_06010_), .Y(_24957_) );
  \$mux  #( .WIDTH(1) ) _46229_ ( .A(_24957_), .B(1'h0), .S(RST), .Y(_03204_) );
  \$mux  #( .WIDTH(1) ) _46230_ ( .A(1'h1), .B(_control_conv2d_16_cond_37_8_1), .S(_06011_), .Y(_24958_) );
  \$mux  #( .WIDTH(1) ) _46231_ ( .A(_24958_), .B(1'h0), .S(RST), .Y(_01566_) );
  \$mux  #( .WIDTH(1) ) _46232_ ( .A(set_req_401), .B(1'h0), .S(_control_conv2d_16_cond_37_8_1), .Y(_24959_) );
  \$mux  #( .WIDTH(1) ) _46233_ ( .A(_24959_), .B(set_req_401), .S(_05999_), .Y(_24960_) );
  \$mux  #( .WIDTH(1) ) _46234_ ( .A(1'h1), .B(_24960_), .S(_06011_), .Y(_24961_) );
  \$mux  #( .WIDTH(1) ) _46235_ ( .A(_24961_), .B(1'h0), .S(RST), .Y(_03879_) );
  \$mux  #( .WIDTH(1) ) _46236_ ( .A(1'h1), .B(_control_conv2d_16_cond_31_7_1), .S(_06012_), .Y(_24962_) );
  \$mux  #( .WIDTH(1) ) _46237_ ( .A(_24962_), .B(1'h0), .S(RST), .Y(_01565_) );
  \$mux  #( .WIDTH(1) ) _46238_ ( .A(axim_flag_345), .B(1'h0), .S(_control_conv2d_16_cond_31_7_1), .Y(_24963_) );
  \$mux  #( .WIDTH(1) ) _46239_ ( .A(_24963_), .B(axim_flag_345), .S(_06000_), .Y(_24964_) );
  \$mux  #( .WIDTH(1) ) _46240_ ( .A(1'h1), .B(_24964_), .S(_06012_), .Y(_24965_) );
  \$mux  #( .WIDTH(1) ) _46241_ ( .A(_24965_), .B(1'h0), .S(RST), .Y(_03202_) );
  \$mux  #( .WIDTH(1) ) _46242_ ( .A(1'h1), .B(_control_conv2d_16_cond_30_6_1), .S(_06013_), .Y(_24966_) );
  \$mux  #( .WIDTH(1) ) _46243_ ( .A(_24966_), .B(1'h0), .S(RST), .Y(_01564_) );
  \$mux  #( .WIDTH(1) ) _46244_ ( .A(set_req_344), .B(1'h0), .S(_control_conv2d_16_cond_30_6_1), .Y(_24967_) );
  \$mux  #( .WIDTH(1) ) _46245_ ( .A(_24967_), .B(set_req_344), .S(_06001_), .Y(_24968_) );
  \$mux  #( .WIDTH(1) ) _46246_ ( .A(1'h1), .B(_24968_), .S(_06013_), .Y(_24969_) );
  \$mux  #( .WIDTH(1) ) _46247_ ( .A(_24969_), .B(1'h0), .S(RST), .Y(_03877_) );
  \$mux  #( .WIDTH(1) ) _46248_ ( .A(1'h1), .B(_control_conv2d_16_cond_24_5_1), .S(_06014_), .Y(_24970_) );
  \$mux  #( .WIDTH(1) ) _46249_ ( .A(_24970_), .B(1'h0), .S(RST), .Y(_01563_) );
  \$mux  #( .WIDTH(1) ) _46250_ ( .A(axim_flag_288), .B(1'h0), .S(_control_conv2d_16_cond_24_5_1), .Y(_24971_) );
  \$mux  #( .WIDTH(1) ) _46251_ ( .A(_24971_), .B(axim_flag_288), .S(_06002_), .Y(_24972_) );
  \$mux  #( .WIDTH(1) ) _46252_ ( .A(1'h1), .B(_24972_), .S(_06014_), .Y(_24973_) );
  \$mux  #( .WIDTH(1) ) _46253_ ( .A(_24973_), .B(1'h0), .S(RST), .Y(_03201_) );
  \$mux  #( .WIDTH(1) ) _46254_ ( .A(1'h1), .B(_control_conv2d_16_cond_23_4_1), .S(_06015_), .Y(_24974_) );
  \$mux  #( .WIDTH(1) ) _46255_ ( .A(_24974_), .B(1'h0), .S(RST), .Y(_01562_) );
  \$mux  #( .WIDTH(1) ) _46256_ ( .A(set_req_287), .B(1'h0), .S(_control_conv2d_16_cond_23_4_1), .Y(_24975_) );
  \$mux  #( .WIDTH(1) ) _46257_ ( .A(_24975_), .B(set_req_287), .S(_06003_), .Y(_24976_) );
  \$mux  #( .WIDTH(1) ) _46258_ ( .A(1'h1), .B(_24976_), .S(_06015_), .Y(_24977_) );
  \$mux  #( .WIDTH(1) ) _46259_ ( .A(_24977_), .B(1'h0), .S(RST), .Y(_03876_) );
  \$mux  #( .WIDTH(1) ) _46260_ ( .A(1'h1), .B(_control_conv2d_16_cond_15_3_1), .S(_06016_), .Y(_24978_) );
  \$mux  #( .WIDTH(1) ) _46261_ ( .A(_24978_), .B(1'h0), .S(RST), .Y(_01561_) );
  \$mux  #( .WIDTH(1) ) _46262_ ( .A(axim_flag_35), .B(1'h0), .S(_control_conv2d_16_cond_15_3_1), .Y(_24979_) );
  \$mux  #( .WIDTH(1) ) _46263_ ( .A(_24979_), .B(axim_flag_35), .S(_06004_), .Y(_24980_) );
  \$mux  #( .WIDTH(1) ) _46264_ ( .A(1'h1), .B(_24980_), .S(_06016_), .Y(_24981_) );
  \$mux  #( .WIDTH(1) ) _46265_ ( .A(_24981_), .B(1'h0), .S(RST), .Y(_03203_) );
  \$mux  #( .WIDTH(1) ) _46266_ ( .A(1'h1), .B(_control_conv2d_16_cond_14_2_1), .S(_06017_), .Y(_24982_) );
  \$mux  #( .WIDTH(1) ) _46267_ ( .A(_24982_), .B(1'h0), .S(RST), .Y(_01560_) );
  \$mux  #( .WIDTH(1) ) _46268_ ( .A(set_req_34), .B(1'h0), .S(_control_conv2d_16_cond_14_2_1), .Y(_24983_) );
  \$mux  #( .WIDTH(1) ) _46269_ ( .A(_24983_), .B(set_req_34), .S(_06005_), .Y(_24984_) );
  \$mux  #( .WIDTH(1) ) _46270_ ( .A(1'h1), .B(_24984_), .S(_06017_), .Y(_24985_) );
  \$mux  #( .WIDTH(1) ) _46271_ ( .A(_24985_), .B(1'h0), .S(RST), .Y(_03878_) );
  \$mux  #( .WIDTH(1) ) _46272_ ( .A(1'h1), .B(_control_conv2d_16_cond_8_1_1), .S(_06019_), .Y(_24986_) );
  \$mux  #( .WIDTH(1) ) _46273_ ( .A(_24986_), .B(1'h0), .S(RST), .Y(_01570_) );
  \$mux  #( .WIDTH(1) ) _46274_ ( .A(axim_flag_22), .B(1'h0), .S(_control_conv2d_16_cond_8_1_1), .Y(_24987_) );
  \$mux  #( .WIDTH(1) ) _46275_ ( .A(_24987_), .B(axim_flag_22), .S(_06006_), .Y(_24988_) );
  \$mux  #( .WIDTH(1) ) _46276_ ( .A(1'h1), .B(_24988_), .S(_06019_), .Y(_24989_) );
  \$mux  #( .WIDTH(1) ) _46277_ ( .A(_24989_), .B(1'h0), .S(RST), .Y(_03200_) );
  \$mux  #( .WIDTH(1) ) _46278_ ( .A(1'h1), .B(_control_conv2d_16_cond_3_0_1), .S(_06020_), .Y(_24990_) );
  \$mux  #( .WIDTH(1) ) _46279_ ( .A(_24990_), .B(1'h0), .S(RST), .Y(_01568_) );
  \$mux  #( .WIDTH(32) ) _46280_ ( .A(control_conv2d_16), .B(0), .S(RST), .Y(_01583_) );
  \$mux  #( .WIDTH(1) ) _46281_ ( .A(axim_flag_9), .B(1'h0), .S(_control_conv2d_16_cond_3_0_1), .Y(_24991_) );
  \$mux  #( .WIDTH(1) ) _46282_ ( .A(_24991_), .B(axim_flag_9), .S(_06007_), .Y(_24992_) );
  \$mux  #( .WIDTH(1) ) _46283_ ( .A(1'h1), .B(_24992_), .S(_06020_), .Y(_24993_) );
  \$mux  #( .WIDTH(1) ) _46284_ ( .A(_24993_), .B(1'h0), .S(RST), .Y(_03206_) );
  \$mux  #( .WIDTH(1) ) _46285_ ( .A(conv2d_16_skip_write_out), .B(1'h0), .S(_06822_), .Y(_20409_) );
  \$mux  #( .WIDTH(1) ) _46286_ ( .A(_24994_), .B(1'h1), .S(RST), .Y(_03265_) );
  \$mux  #( .WIDTH(1) ) _46287_ ( .A(conv2d_16_skip_comp), .B(1'h1), .S(conv2d_16_update_filter), .Y(_20411_) );
  \$mux  #( .WIDTH(1) ) _46288_ ( .A(_24995_), .B(1'h0), .S(RST), .Y(_03262_) );
  \$mux  #( .WIDTH(1) ) _46289_ ( .A(conv2d_16_skip_read_act), .B(1'h1), .S(conv2d_16_update_filter), .Y(_20413_) );
  \$mux  #( .WIDTH(1) ) _46290_ ( .A(_24996_), .B(1'h0), .S(RST), .Y(_03263_) );
  \$mux  #( .WIDTH(1) ) _46291_ ( .A(conv2d_16_skip_read_filter), .B(1'h1), .S(conv2d_16_update_filter), .Y(_20415_) );
  \$mux  #( .WIDTH(1) ) _46292_ ( .A(_24997_), .B(1'h0), .S(RST), .Y(_03264_) );
  \$mux  #( .WIDTH(32) ) _46293_ ( .A(0), .B(conv2d_16_out_laddr_offset), .S(conv2d_16_skip_write_out), .Y({ _20441_, _20440_, _20438_, _20437_, _20436_, _20435_, _20434_, _20433_, _20432_, _20431_, _20430_, _20429_, _20427_, _20426_, _20425_, _20424_, _20423_, _20422_, _20421_, _20420_, _20419_, _20418_, _20448_, _20447_, _20446_, _20445_, _20444_, _20443_, _20442_, _20439_, _20428_, _20417_ }) );
  \$mux  #( .WIDTH(32) ) _46294_ ( .A(_24430_), .B(conv2d_16_out_laddr_offset), .S(_05722_), .Y({ _20473_, _20472_, _20470_, _20469_, _20468_, _20467_, _20466_, _20465_, _20464_, _20463_, _20462_, _20461_, _20459_, _20458_, _20457_, _20456_, _20455_, _20454_, _20453_, _20452_, _20451_, _20450_, _20480_, _20479_, _20478_, _20477_, _20476_, _20475_, _20474_, _20471_, _20460_, _20449_ }) );
  \$mux  #( .WIDTH(32) ) _46295_ ( .A(_24998_), .B(0), .S(RST), .Y(_03247_) );
  \$mux  #( .WIDTH(32) ) _46296_ ( .A(0), .B(1024), .S(conv2d_16_out_page), .Y({ _20505_, _20504_, _20502_, _20501_, _20500_, _20499_, _20498_, _20497_, _20496_, _20495_, _20494_, _20493_, _20491_, _20490_, _20489_, _20488_, _20487_, _20486_, _20485_, _20484_, _20483_, _20482_, _20512_, _20511_, _20510_, _20509_, _20508_, _20507_, _20506_, _20503_, _20492_, _20481_ }) );
  \$mux  #( .WIDTH(32) ) _46297_ ( .A(_24999_), .B(0), .S(RST), .Y(_03251_) );
  \$mux  #( .WIDTH(32) ) _46298_ ( .A(1024), .B(0), .S(conv2d_16_out_page), .Y({ _20569_, _20568_, _20566_, _20565_, _20564_, _20563_, _20562_, _20561_, _20560_, _20559_, _20558_, _20557_, _20555_, _20554_, _20553_, _20552_, _20551_, _20550_, _20549_, _20548_, _20547_, _20546_, _20576_, _20575_, _20574_, _20573_, _20572_, _20571_, _20570_, _20567_, _20556_, _20545_ }) );
  \$mux  #( .WIDTH(32) ) _46299_ ( .A(_25000_), .B(0), .S(RST), .Y(_03249_) );
  \$mux  #( .WIDTH(1) ) _46300_ ( .A(1'h1), .B(1'h0), .S(conv2d_16_out_page), .Y(_20609_) );
  \$mux  #( .WIDTH(1) ) _46301_ ( .A(_25001_), .B(1'h0), .S(RST), .Y(_03248_) );
  \$mux  #( .WIDTH(32) ) _46302_ ( .A(conv2d_16_filter_page_dma_offset), .B(_24435_), .S(conv2d_16_update_filter), .Y(_25002_) );
  \$mux  #( .WIDTH(32) ) _46303_ ( .A(_25002_), .B(0), .S(_06817_), .Y({ _20635_, _20634_, _20632_, _20631_, _20630_, _20629_, _20628_, _20627_, _20626_, _20625_, _20624_, _20623_, _20621_, _20620_, _20619_, _20618_, _20617_, _20616_, _20615_, _20614_, _20613_, _20612_, _20642_, _20641_, _20640_, _20639_, _20638_, _20637_, _20636_, _20633_, _20622_, _20611_ }) );
  \$mux  #( .WIDTH(32) ) _46304_ ( .A(_25003_), .B(0), .S(RST), .Y(_03236_) );
  \$mux  #( .WIDTH(32) ) _46305_ ( .A(conv2d_16_filter_page_comp_offset), .B(_24434_), .S(conv2d_16_update_filter), .Y(_25004_) );
  \$mux  #( .WIDTH(32) ) _46306_ ( .A(_25004_), .B(0), .S(_06817_), .Y({ _20699_, _20698_, _20696_, _20695_, _20694_, _20693_, _20692_, _20691_, _20690_, _20689_, _20688_, _20687_, _20685_, _20684_, _20683_, _20682_, _20681_, _20680_, _20679_, _20678_, _20677_, _20676_, _20706_, _20705_, _20704_, _20703_, _20702_, _20701_, _20700_, _20697_, _20686_, _20675_ }) );
  \$mux  #( .WIDTH(32) ) _46307_ ( .A(_25005_), .B(0), .S(RST), .Y(_03234_) );
  \$mux  #( .WIDTH(32) ) _46308_ ( .A(conv2d_16_act_page_dma_offset_2), .B(_24444_), .S(conv2d_16_mux_next_dma_flag_2), .Y(_25006_) );
  \$mux  #( .WIDTH(32) ) _46309_ ( .A(_25006_), .B(0), .S(_06820_), .Y(_25007_) );
  \$mux  #( .WIDTH(32) ) _46310_ ( .A(_25007_), .B(0), .S(conv2d_16_update_filter), .Y({ _20763_, _20762_, _20760_, _20759_, _20758_, _20757_, _20756_, _20755_, _20754_, _20753_, _20752_, _20751_, _20749_, _20748_, _20747_, _20746_, _20745_, _20744_, _20743_, _20742_, _20741_, _20740_, _20770_, _20769_, _20768_, _20767_, _20766_, _20765_, _20764_, _20761_, _20750_, _20739_ }) );
  \$mux  #( .WIDTH(32) ) _46311_ ( .A(_25008_), .B(0), .S(RST), .Y(_03220_) );
  \$mux  #( .WIDTH(32) ) _46312_ ( .A(conv2d_16_act_page_dma_offset_1), .B(_24442_), .S(conv2d_16_mux_next_dma_flag_1), .Y(_25009_) );
  \$mux  #( .WIDTH(32) ) _46313_ ( .A(_25009_), .B(0), .S(_06819_), .Y(_25010_) );
  \$mux  #( .WIDTH(32) ) _46314_ ( .A(_25010_), .B(0), .S(conv2d_16_update_filter), .Y({ _20827_, _20826_, _20824_, _20823_, _20822_, _20821_, _20820_, _20819_, _20818_, _20817_, _20816_, _20815_, _20813_, _20812_, _20811_, _20810_, _20809_, _20808_, _20807_, _20806_, _20805_, _20804_, _20834_, _20833_, _20832_, _20831_, _20830_, _20829_, _20828_, _20825_, _20814_, _20803_ }) );
  \$mux  #( .WIDTH(32) ) _46315_ ( .A(_25011_), .B(0), .S(RST), .Y(_03219_) );
  \$mux  #( .WIDTH(32) ) _46316_ ( .A(conv2d_16_act_page_dma_offset_0), .B(_24440_), .S(conv2d_16_mux_next_dma_flag_0), .Y(_25012_) );
  \$mux  #( .WIDTH(32) ) _46317_ ( .A(_25012_), .B(0), .S(_06818_), .Y(_25013_) );
  \$mux  #( .WIDTH(32) ) _46318_ ( .A(_25013_), .B(0), .S(conv2d_16_update_filter), .Y({ _20891_, _20890_, _20888_, _20887_, _20886_, _20885_, _20884_, _20883_, _20882_, _20881_, _20880_, _20879_, _20877_, _20876_, _20875_, _20874_, _20873_, _20872_, _20871_, _20870_, _20869_, _20868_, _20898_, _20897_, _20896_, _20895_, _20894_, _20893_, _20892_, _20889_, _20878_, _20867_ }) );
  \$mux  #( .WIDTH(32) ) _46319_ ( .A(_25014_), .B(0), .S(RST), .Y(_03218_) );
  \$mux  #( .WIDTH(32) ) _46320_ ( .A(conv2d_16_act_page_comp_offset_2), .B(_24443_), .S(conv2d_16_mux_next_dma_flag_2), .Y(_25015_) );
  \$mux  #( .WIDTH(32) ) _46321_ ( .A(_25015_), .B(0), .S(_06820_), .Y(_25016_) );
  \$mux  #( .WIDTH(32) ) _46322_ ( .A(_25016_), .B(0), .S(conv2d_16_update_filter), .Y({ _20955_, _20954_, _20952_, _20951_, _20950_, _20949_, _20948_, _20947_, _20946_, _20945_, _20944_, _20943_, _20941_, _20940_, _20939_, _20938_, _20937_, _20936_, _20935_, _20934_, _20933_, _20932_, _20962_, _20961_, _20960_, _20959_, _20958_, _20957_, _20956_, _20953_, _20942_, _20931_ }) );
  \$mux  #( .WIDTH(32) ) _46323_ ( .A(_25017_), .B(0), .S(RST), .Y(_03214_) );
  \$mux  #( .WIDTH(32) ) _46324_ ( .A(conv2d_16_act_page_comp_offset_1), .B(_24441_), .S(conv2d_16_mux_next_dma_flag_1), .Y(_25018_) );
  \$mux  #( .WIDTH(32) ) _46325_ ( .A(_25018_), .B(0), .S(_06819_), .Y(_25019_) );
  \$mux  #( .WIDTH(32) ) _46326_ ( .A(_25019_), .B(0), .S(conv2d_16_update_filter), .Y({ _21019_, _21018_, _21016_, _21015_, _21014_, _21013_, _21012_, _21011_, _21010_, _21009_, _21008_, _21007_, _21005_, _21004_, _21003_, _21002_, _21001_, _21000_, _20999_, _20998_, _20997_, _20996_, _21026_, _21025_, _21024_, _21023_, _21022_, _21021_, _21020_, _21017_, _21006_, _20995_ }) );
  \$mux  #( .WIDTH(32) ) _46327_ ( .A(_25020_), .B(0), .S(RST), .Y(_03213_) );
  \$mux  #( .WIDTH(32) ) _46328_ ( .A(conv2d_16_act_page_comp_offset_0), .B(_24439_), .S(conv2d_16_mux_next_dma_flag_0), .Y(_25021_) );
  \$mux  #( .WIDTH(32) ) _46329_ ( .A(_25021_), .B(0), .S(_06818_), .Y(_25022_) );
  \$mux  #( .WIDTH(32) ) _46330_ ( .A(_25022_), .B(0), .S(conv2d_16_update_filter), .Y({ _21083_, _21082_, _21080_, _21079_, _21078_, _21077_, _21076_, _21075_, _21074_, _21073_, _21072_, _21071_, _21069_, _21068_, _21067_, _21066_, _21065_, _21064_, _21063_, _21062_, _21061_, _21060_, _21090_, _21089_, _21088_, _21087_, _21086_, _21085_, _21084_, _21081_, _21070_, _21059_ }) );
  \$mux  #( .WIDTH(32) ) _46331_ ( .A(_25023_), .B(0), .S(RST), .Y(_03212_) );
  \$mux  #( .WIDTH(2) ) _46332_ ( .A(conv2d_16_row_select), .B(2'h0), .S(conv2d_16_update_filter), .Y({ _21124_, _21123_ }) );
  \$mux  #( .WIDTH(2) ) _46333_ ( .A(_25024_), .B(2'h0), .S(RST), .Y(_03257_) );
  \$mux  #( .WIDTH(32) ) _46334_ ( .A(_25025_), .B(0), .S(RST), .Y(_03255_) );
  \$mux  #( .WIDTH(32) ) _46335_ ( .A(_25026_), .B(0), .S(RST), .Y(_03254_) );
  \$mux  #( .WIDTH(32) ) _46336_ ( .A(_25027_), .B(0), .S(RST), .Y(_03256_) );
  \$mux  #( .WIDTH(32) ) _46337_ ( .A(0), .B(conv2d_16_out_ram_select), .S(conv2d_16_skip_write_out), .Y({ _21247_, _21246_, _21244_, _21243_, _21242_, _21241_, _21240_, _21239_, _21238_, _21237_, _21236_, _21235_, _21233_, _21232_, _21231_, _21230_, _21229_, _21228_, _21227_, _21226_, _21225_, _21224_, _21254_, _21253_, _21252_, _21251_, _21250_, _21249_, _21248_, _21245_, _21234_, _21223_ }) );
  \$mux  #( .WIDTH(32) ) _46338_ ( .A(0), .B(_24431_), .S(_05722_), .Y({ _21279_, _21278_, _21276_, _21275_, _21274_, _21273_, _21272_, _21271_, _21270_, _21269_, _21268_, _21267_, _21265_, _21264_, _21263_, _21262_, _21261_, _21260_, _21259_, _21258_, _21257_, _21256_, _21286_, _21285_, _21284_, _21283_, _21282_, _21281_, _21280_, _21277_, _21266_, _21255_ }) );
  \$mux  #( .WIDTH(32) ) _46339_ ( .A(_25028_), .B(0), .S(RST), .Y(_03252_) );
  \$mux  #( .WIDTH(32) ) _46340_ ( .A(_24446_), .B(conv2d_16_out_row_count), .S(conv2d_16_skip_write_out), .Y(_25029_) );
  \$mux  #( .WIDTH(32) ) _46341_ ( .A(_25029_), .B(0), .S(_06821_), .Y({ _21311_, _21310_, _21308_, _21307_, _21306_, _21305_, _21304_, _21303_, _21302_, _21301_, _21300_, _21299_, _21297_, _21296_, _21295_, _21294_, _21293_, _21292_, _21291_, _21290_, _21289_, _21288_, _21318_, _21317_, _21316_, _21315_, _21314_, _21313_, _21312_, _21309_, _21298_, _21287_ }) );
  \$mux  #( .WIDTH(32) ) _46342_ ( .A(_25030_), .B(0), .S(RST), .Y(_03253_) );
  \$mux  #( .WIDTH(2) ) _46343_ ( .A(_24438_), .B(_28935_[1:0]), .S(_06154_), .Y(_25031_) );
  \$mux  #( .WIDTH(2) ) _46344_ ( .A(_25031_), .B(2'h0), .S(conv2d_16_update_filter), .Y({ _21352_, _21351_ }) );
  \$mux  #( .WIDTH(2) ) _46345_ ( .A(_25032_), .B(2'h0), .S(RST), .Y(_03260_) );
  \$mux  #( .WIDTH(32) ) _46346_ ( .A(conv2d_16_och_count), .B(_24433_), .S(conv2d_16_update_filter), .Y({ _21379_, _21378_, _21376_, _21375_, _21374_, _21373_, _21372_, _21371_, _21370_, _21369_, _21368_, _21367_, _21365_, _21364_, _21363_, _21362_, _21361_, _21360_, _21359_, _21358_, _21357_, _21356_, _21386_, _21385_, _21384_, _21383_, _21382_, _21381_, _21380_, _21377_, _21366_, _21355_ }) );
  \$mux  #( .WIDTH(32) ) _46347_ ( .A(_25033_), .B(0), .S(RST), .Y(_03240_) );
  \$mux  #( .WIDTH(32) ) _46348_ ( .A(conv2d_16_bat_count), .B(0), .S(conv2d_16_update_filter), .Y({ _21443_, _21442_, _21440_, _21439_, _21438_, _21437_, _21436_, _21435_, _21434_, _21433_, _21432_, _21431_, _21429_, _21428_, _21427_, _21426_, _21425_, _21424_, _21423_, _21422_, _21421_, _21420_, _21450_, _21449_, _21448_, _21447_, _21446_, _21445_, _21444_, _21441_, _21430_, _21419_ }) );
  \$mux  #( .WIDTH(32) ) _46349_ ( .A(_25034_), .B(0), .S(RST), .Y(_03225_) );
  \$mux  #( .WIDTH(32) ) _46350_ ( .A(_24437_), .B(0), .S(conv2d_16_update_filter), .Y({ _21507_, _21506_, _21504_, _21503_, _21502_, _21501_, _21500_, _21499_, _21498_, _21497_, _21496_, _21495_, _21493_, _21492_, _21491_, _21490_, _21489_, _21488_, _21487_, _21486_, _21485_, _21484_, _21514_, _21513_, _21512_, _21511_, _21510_, _21509_, _21508_, _21505_, _21494_, _21483_ }) );
  \$mux  #( .WIDTH(32) ) _46351_ ( .A(_25035_), .B(0), .S(RST), .Y(_03258_) );
  \$mux  #( .WIDTH(32) ) _46352_ ( .A(conv2d_16_next_out_write_size), .B(512), .S(_05514_), .Y(_25036_) );
  \$mux  #( .WIDTH(32) ) _46353_ ( .A(_25036_), .B(0), .S(RST), .Y(_03237_) );
  \$mux  #( .WIDTH(32) ) _46354_ ( .A(_25037_), .B(0), .S(RST), .Y(_03278_) );
  \$mux  #( .WIDTH(1) ) _46355_ ( .A(_25038_), .B(1'h0), .S(RST), .Y(_03232_) );
  \$mux  #( .WIDTH(1) ) _46356_ ( .A(1'h0), .B(1'h1), .S(conv2d_16_update_filter), .Y(_21579_) );
  \$mux  #( .WIDTH(1) ) _46357_ ( .A(_25039_), .B(1'h0), .S(RST), .Y(_03231_) );
  \$mux  #( .WIDTH(1) ) _46358_ ( .A(conv2d_16_dma_flag_0), .B(1'h1), .S(_05514_), .Y(_25040_) );
  \$mux  #( .WIDTH(1) ) _46359_ ( .A(_25040_), .B(1'h0), .S(RST), .Y(_03230_) );
  \$mux  #( .WIDTH(32) ) _46360_ ( .A(conv2d_16_out_base_offset_och), .B(_24447_), .S(_06821_), .Y({ _21605_, _21604_, _21602_, _21601_, _21600_, _21599_, _21598_, _21597_, _21596_, _21595_, _21594_, _21593_, _21591_, _21590_, _21589_, _21588_, _21587_, _21586_, _21585_, _21584_, _21583_, _21582_, _21612_, _21611_, _21610_, _21609_, _21608_, _21607_, _21606_, _21603_, _21592_, _21581_ }) );
  \$mux  #( .WIDTH(32) ) _46361_ ( .A(_25041_), .B(0), .S(RST), .Y(_03244_) );
  \$mux  #( .WIDTH(32) ) _46362_ ( .A(conv2d_16_out_base_offset_bat), .B(0), .S(_06821_), .Y({ _21669_, _21668_, _21666_, _21665_, _21664_, _21663_, _21662_, _21661_, _21660_, _21659_, _21658_, _21657_, _21655_, _21654_, _21653_, _21652_, _21651_, _21650_, _21649_, _21648_, _21647_, _21646_, _21676_, _21675_, _21674_, _21673_, _21672_, _21671_, _21670_, _21667_, _21656_, _21645_ }) );
  \$mux  #( .WIDTH(32) ) _46363_ ( .A(_25042_), .B(0), .S(RST), .Y(_03242_) );
  \$mux  #( .WIDTH(32) ) _46364_ ( .A(_24445_), .B(conv2d_16_out_base_offset_row), .S(conv2d_16_skip_write_out), .Y(_25043_) );
  \$mux  #( .WIDTH(32) ) _46365_ ( .A(_25043_), .B(0), .S(_06821_), .Y({ _21733_, _21732_, _21730_, _21729_, _21728_, _21727_, _21726_, _21725_, _21724_, _21723_, _21722_, _21721_, _21719_, _21718_, _21717_, _21716_, _21715_, _21714_, _21713_, _21712_, _21711_, _21710_, _21740_, _21739_, _21738_, _21737_, _21736_, _21735_, _21734_, _21731_, _21720_, _21709_ }) );
  \$mux  #( .WIDTH(32) ) _46366_ ( .A(_25044_), .B(0), .S(RST), .Y(_03245_) );
  \$mux  #( .WIDTH(32) ) _46367_ ( .A(0), .B(conv2d_16_out_base_offset_col), .S(conv2d_16_skip_write_out), .Y({ _21797_, _21796_, _21794_, _21793_, _21792_, _21791_, _21790_, _21789_, _21788_, _21787_, _21786_, _21785_, _21783_, _21782_, _21781_, _21780_, _21779_, _21778_, _21777_, _21776_, _21775_, _21774_, _21804_, _21803_, _21802_, _21801_, _21800_, _21799_, _21798_, _21795_, _21784_, _21773_ }) );
  \$mux  #( .WIDTH(32) ) _46368_ ( .A(_25045_), .B(0), .S(RST), .Y(_03243_) );
  \$mux  #( .WIDTH(32) ) _46369_ ( .A(0), .B(conv2d_16_out_base_offset_val), .S(_06021_), .Y(_25046_) );
  \$mux  #( .WIDTH(32) ) _46370_ ( .A(_25046_), .B(0), .S(RST), .Y(_03246_) );
  \$mux  #( .WIDTH(32) ) _46371_ ( .A(conv2d_16_filter_base_offset), .B(_24432_), .S(conv2d_16_update_filter), .Y({ _21861_, _21860_, _21858_, _21857_, _21856_, _21855_, _21854_, _21853_, _21852_, _21851_, _21850_, _21849_, _21847_, _21846_, _21845_, _21844_, _21843_, _21842_, _21841_, _21840_, _21839_, _21838_, _21868_, _21867_, _21866_, _21865_, _21864_, _21863_, _21862_, _21859_, _21848_, _21837_ }) );
  \$mux  #( .WIDTH(32) ) _46372_ ( .A(_25047_), .B(0), .S(RST), .Y(_03233_) );
  \$mux  #( .WIDTH(32) ) _46373_ ( .A(conv2d_16_act_base_offset_bat), .B(0), .S(conv2d_16_update_filter), .Y({ _21925_, _21924_, _21922_, _21921_, _21920_, _21919_, _21918_, _21917_, _21916_, _21915_, _21914_, _21913_, _21911_, _21910_, _21909_, _21908_, _21907_, _21906_, _21905_, _21904_, _21903_, _21902_, _21932_, _21931_, _21930_, _21929_, _21928_, _21927_, _21926_, _21923_, _21912_, _21901_ }) );
  \$mux  #( .WIDTH(32) ) _46374_ ( .A(_25048_), .B(0), .S(RST), .Y(_03210_) );
  \$mux  #( .WIDTH(32) ) _46375_ ( .A(_24436_), .B(0), .S(conv2d_16_update_filter), .Y({ _21989_, _21988_, _21986_, _21985_, _21984_, _21983_, _21982_, _21981_, _21980_, _21979_, _21978_, _21977_, _21975_, _21974_, _21973_, _21972_, _21971_, _21970_, _21969_, _21968_, _21967_, _21966_, _21996_, _21995_, _21994_, _21993_, _21992_, _21991_, _21990_, _21987_, _21976_, _21965_ }) );
  \$mux  #( .WIDTH(32) ) _46376_ ( .A(_25049_), .B(0), .S(RST), .Y(_03211_) );
  \$mux  #( .WIDTH(32) ) _46377_ ( .A(0), .B(control_conv2d_16), .S(_05740_), .Y(_25050_) );
  \$mux  #( .WIDTH(32) ) _46378_ ( .A(0), .B(_25050_), .S(_05736_), .Y(_25051_) );
  \$mux  #( .WIDTH(32) ) _46379_ ( .A(0), .B(_25051_), .S(_05732_), .Y({ _22053_, _22052_, _22050_, _22049_, _22048_, _22047_, _22046_, _22045_, _22044_, _22043_, _22042_, _22041_, _22039_, _22038_, _22037_, _22036_, _22035_, _22034_, _22033_, _22032_, _22031_, _22030_, _22060_, _22059_, _22058_, _22057_, _22056_, _22055_, _22054_, _22051_, _22040_, _22029_ }) );
  \$mux  #( .WIDTH(32) ) _46380_ ( .A(control_conv2d_16), .B(55), .S(_maxi_write_idle), .Y({ _22117_, _22116_, _22114_, _22113_, _22112_, _22111_, _22110_, _22109_, _22108_, _22107_, _22106_, _22105_, _22103_, _22102_, _22101_, _22100_, _22099_, _22098_, _22097_, _22096_, _22095_, _22094_, _22124_, _22123_, _22122_, _22121_, _22120_, _22119_, _22118_, _22115_, _22104_, _22093_ }) );
  \$mux  #( .WIDTH(32) ) _46381_ ( .A(21), .B(13), .S(conv2d_16_update_filter), .Y(_25053_) );
  \$mux  #( .WIDTH(32) ) _46382_ ( .A(_25053_), .B(54), .S(_06821_), .Y({ _22149_, _22148_, _22146_, _22145_, _22144_, _22143_, _22142_, _22141_, _22140_, _22139_, _22138_, _22137_, _22135_, _22134_, _22133_, _22132_, _22131_, _22130_, _22129_, _22128_, _22127_, _22126_, _22156_, _22155_, _22154_, _22153_, _22152_, _22151_, _22150_, _22147_, _22136_, _22125_ }) );
  \$mux  #( .WIDTH(32) ) _46383_ ( .A(control_conv2d_16), .B(48), .S(_maxi_write_idle), .Y({ _22181_, _22180_, _22178_, _22177_, _22176_, _22175_, _22174_, _22173_, _22172_, _22171_, _22170_, _22169_, _22167_, _22166_, _22165_, _22164_, _22163_, _22162_, _22161_, _22160_, _22159_, _22158_, _22188_, _22187_, _22186_, _22185_, _22184_, _22183_, _22182_, _22179_, _22168_, _22157_ }) );
  \$mux  #( .WIDTH(32) ) _46384_ ( .A(47), .B(51), .S(conv2d_16_dma_out_mask_0), .Y({ _22213_, _22212_, _22210_, _22209_, _22208_, _22207_, _22206_, _22205_, _22204_, _22203_, _22202_, _22201_, _22199_, _22198_, _22197_, _22196_, _22195_, _22194_, _22193_, _22192_, _22191_, _22190_, _22220_, _22219_, _22218_, _22217_, _22216_, _22215_, _22214_, _22211_, _22200_, _22189_ }) );
  \$mux  #( .WIDTH(32) ) _46385_ ( .A(control_conv2d_16), .B(46), .S(_06153_), .Y(_25054_) );
  \$mux  #( .WIDTH(32) ) _46386_ ( .A(_25054_), .B(53), .S(conv2d_16_skip_write_out), .Y({ _22245_, _22244_, _22242_, _22241_, _22240_, _22239_, _22238_, _22237_, _22236_, _22235_, _22234_, _22233_, _22231_, _22230_, _22229_, _22228_, _22227_, _22226_, _22225_, _22224_, _22223_, _22222_, _22252_, _22251_, _22250_, _22249_, _22248_, _22247_, _22246_, _22243_, _22232_, _22221_ }) );
  \$mux  #( .WIDTH(32) ) _46387_ ( .A(45), .B(control_conv2d_16), .S(_05727_), .Y({ _22277_, _22276_, _22274_, _22273_, _22272_, _22271_, _22270_, _22269_, _22268_, _22267_, _22266_, _22265_, _22263_, _22262_, _22261_, _22260_, _22259_, _22258_, _22257_, _22256_, _22255_, _22254_, _22284_, _22283_, _22282_, _22281_, _22280_, _22279_, _22278_, _22275_, _22264_, _22253_ }) );
  \$mux  #( .WIDTH(32) ) _46388_ ( .A(control_conv2d_16), .B(42), .S(_maxi_read_idle), .Y({ _22309_, _22308_, _22306_, _22305_, _22304_, _22303_, _22302_, _22301_, _22300_, _22299_, _22298_, _22297_, _22295_, _22294_, _22293_, _22292_, _22291_, _22290_, _22289_, _22288_, _22287_, _22286_, _22316_, _22315_, _22314_, _22313_, _22312_, _22311_, _22310_, _22307_, _22296_, _22285_ }) );
  \$mux  #( .WIDTH(32) ) _46389_ ( .A(control_conv2d_16), .B(37), .S(_maxi_read_idle), .Y({ _22341_, _22340_, _22338_, _22337_, _22336_, _22335_, _22334_, _22333_, _22332_, _22331_, _22330_, _22329_, _22327_, _22326_, _22325_, _22324_, _22323_, _22322_, _22321_, _22320_, _22319_, _22318_, _22348_, _22347_, _22346_, _22345_, _22344_, _22343_, _22342_, _22339_, _22328_, _22317_ }) );
  \$mux  #( .WIDTH(32) ) _46390_ ( .A(36), .B(42), .S(_06881_), .Y({ _22373_, _22372_, _22370_, _22369_, _22368_, _22367_, _22366_, _22365_, _22364_, _22363_, _22362_, _22361_, _22359_, _22358_, _22357_, _22356_, _22355_, _22354_, _22353_, _22352_, _22351_, _22350_, _22380_, _22379_, _22378_, _22377_, _22376_, _22375_, _22374_, _22371_, _22360_, _22349_ }) );
  \$mux  #( .WIDTH(32) ) _46391_ ( .A(control_conv2d_16), .B(35), .S(_maxi_read_idle), .Y({ _22405_, _22404_, _22402_, _22401_, _22400_, _22399_, _22398_, _22397_, _22396_, _22395_, _22394_, _22393_, _22391_, _22390_, _22389_, _22388_, _22387_, _22386_, _22385_, _22384_, _22383_, _22382_, _22412_, _22411_, _22410_, _22409_, _22408_, _22407_, _22406_, _22403_, _22392_, _22381_ }) );
  \$mux  #( .WIDTH(32) ) _46392_ ( .A(control_conv2d_16), .B(30), .S(_maxi_read_idle), .Y({ _22437_, _22436_, _22434_, _22433_, _22432_, _22431_, _22430_, _22429_, _22428_, _22427_, _22426_, _22425_, _22423_, _22422_, _22421_, _22420_, _22419_, _22418_, _22417_, _22416_, _22415_, _22414_, _22444_, _22443_, _22442_, _22441_, _22440_, _22439_, _22438_, _22435_, _22424_, _22413_ }) );
  \$mux  #( .WIDTH(32) ) _46393_ ( .A(29), .B(35), .S(_06880_), .Y({ _22469_, _22468_, _22466_, _22465_, _22464_, _22463_, _22462_, _22461_, _22460_, _22459_, _22458_, _22457_, _22455_, _22454_, _22453_, _22452_, _22451_, _22450_, _22449_, _22448_, _22447_, _22446_, _22476_, _22475_, _22474_, _22473_, _22472_, _22471_, _22470_, _22467_, _22456_, _22445_ }) );
  \$mux  #( .WIDTH(32) ) _46394_ ( .A(control_conv2d_16), .B(28), .S(_maxi_read_idle), .Y({ _22501_, _22500_, _22498_, _22497_, _22496_, _22495_, _22494_, _22493_, _22492_, _22491_, _22490_, _22489_, _22487_, _22486_, _22485_, _22484_, _22483_, _22482_, _22481_, _22480_, _22479_, _22478_, _22508_, _22507_, _22506_, _22505_, _22504_, _22503_, _22502_, _22499_, _22488_, _22477_ }) );
  \$mux  #( .WIDTH(32) ) _46395_ ( .A(control_conv2d_16), .B(23), .S(_maxi_read_idle), .Y({ _22533_, _22532_, _22530_, _22529_, _22528_, _22527_, _22526_, _22525_, _22524_, _22523_, _22522_, _22521_, _22519_, _22518_, _22517_, _22516_, _22515_, _22514_, _22513_, _22512_, _22511_, _22510_, _22540_, _22539_, _22538_, _22537_, _22536_, _22535_, _22534_, _22531_, _22520_, _22509_ }) );
  \$mux  #( .WIDTH(32) ) _46396_ ( .A(22), .B(28), .S(_06879_), .Y(_25055_) );
  \$mux  #( .WIDTH(32) ) _46397_ ( .A(_25055_), .B(43), .S(conv2d_16_skip_read_act), .Y({ _22565_, _22564_, _22562_, _22561_, _22560_, _22559_, _22558_, _22557_, _22556_, _22555_, _22554_, _22553_, _22551_, _22550_, _22549_, _22548_, _22547_, _22546_, _22545_, _22544_, _22543_, _22542_, _22572_, _22571_, _22570_, _22569_, _22568_, _22567_, _22566_, _22563_, _22552_, _22541_ }) );
  \$mux  #( .WIDTH(32) ) _46398_ ( .A(control_conv2d_16), .B(19), .S(_maxi_read_idle), .Y({ _22597_, _22596_, _22594_, _22593_, _22592_, _22591_, _22590_, _22589_, _22588_, _22587_, _22586_, _22585_, _22583_, _22582_, _22581_, _22580_, _22579_, _22578_, _22577_, _22576_, _22575_, _22574_, _22604_, _22603_, _22602_, _22601_, _22600_, _22599_, _22598_, _22595_, _22584_, _22573_ }) );
  \$mux  #( .WIDTH(32) ) _46399_ ( .A(control_conv2d_16), .B(14), .S(_maxi_read_idle), .Y(_25056_) );
  \$mux  #( .WIDTH(32) ) _46400_ ( .A(_25056_), .B(20), .S(conv2d_16_skip_read_filter), .Y({ _22629_, _22628_, _22626_, _22625_, _22624_, _22623_, _22622_, _22621_, _22620_, _22619_, _22618_, _22617_, _22615_, _22614_, _22613_, _22612_, _22611_, _22610_, _22609_, _22608_, _22607_, _22606_, _22636_, _22635_, _22634_, _22633_, _22632_, _22631_, _22630_, _22627_, _22616_, _22605_ }) );
  \$mux  #( .WIDTH(32) ) _46401_ ( .A(control_conv2d_16), .B(12), .S(_maxi_read_idle), .Y({ _22661_, _22660_, _22658_, _22657_, _22656_, _22655_, _22654_, _22653_, _22652_, _22651_, _22650_, _22649_, _22647_, _22646_, _22645_, _22644_, _22643_, _22642_, _22641_, _22640_, _22639_, _22638_, _22668_, _22667_, _22666_, _22665_, _22664_, _22663_, _22662_, _22659_, _22648_, _22637_ }) );
  \$mux  #( .WIDTH(32) ) _46402_ ( .A(control_conv2d_16), .B(8), .S(_maxi_read_idle), .Y({ _22693_, _22692_, _22690_, _22689_, _22688_, _22687_, _22686_, _22685_, _22684_, _22683_, _22682_, _22681_, _22679_, _22678_, _22677_, _22676_, _22675_, _22674_, _22673_, _22672_, _22671_, _22670_, _22700_, _22699_, _22698_, _22697_, _22696_, _22695_, _22694_, _22691_, _22680_, _22669_ }) );
  \$mux  #( .WIDTH(32) ) _46403_ ( .A(control_conv2d_16), .B(7), .S(_maxi_read_idle), .Y({ _22725_, _22724_, _22722_, _22721_, _22720_, _22719_, _22718_, _22717_, _22716_, _22715_, _22714_, _22713_, _22711_, _22710_, _22709_, _22708_, _22707_, _22706_, _22705_, _22704_, _22703_, _22702_, _22732_, _22731_, _22730_, _22729_, _22728_, _22727_, _22726_, _22723_, _22712_, _22701_ }) );
  \$mux  #( .WIDTH(32) ) _46404_ ( .A(control_conv2d_16), .B(3), .S(_maxi_read_idle), .Y({ _22757_, _22756_, _22754_, _22753_, _22752_, _22751_, _22750_, _22749_, _22748_, _22747_, _22746_, _22745_, _22743_, _22742_, _22741_, _22740_, _22739_, _22738_, _22737_, _22736_, _22735_, _22734_, _22764_, _22763_, _22762_, _22761_, _22760_, _22759_, _22758_, _22755_, _22744_, _22733_ }) );
  \$mux  #( .WIDTH(32) ) _46405_ ( .A(1), .B(control_conv2d_16), .S(_05741_), .Y(_25057_) );
  \$mux  #( .WIDTH(32) ) _46406_ ( .A(1), .B(_25057_), .S(_05737_), .Y(_25058_) );
  \$mux  #( .WIDTH(32) ) _46407_ ( .A(1), .B(_25058_), .S(_05733_), .Y({ _22789_, _22788_, _22786_, _22785_, _22784_, _22783_, _22782_, _22781_, _22780_, _22779_, _22778_, _22777_, _22775_, _22774_, _22773_, _22772_, _22771_, _22770_, _22769_, _22768_, _22767_, _22766_, _22796_, _22795_, _22794_, _22793_, _22792_, _22791_, _22790_, _22787_, _22776_, _22765_ }) );
  \$mux  #( .WIDTH(32) ) _46408_ ( .A(_25052_), .B(0), .S(RST), .Y(_03207_) );
  \$mux  #( .WIDTH(32) ) _46409_ ( .A(_25059_), .B(0), .S(RST), .Y(_03288_) );
  \$mux  #( .WIDTH(32) ) _46410_ ( .A(_25060_), .B(0), .S(RST), .Y(_03287_) );
  \$mux  #( .WIDTH(32) ) _46411_ ( .A(_25061_), .B(0), .S(RST), .Y(_03286_) );
  \$mux  #( .WIDTH(32) ) _46412_ ( .A(_25062_), .B(0), .S(RST), .Y(_03285_) );
  \$mux  #( .WIDTH(32) ) _46413_ ( .A(_25063_), .B(0), .S(RST), .Y(_03301_) );
  \$mux  #( .WIDTH(32) ) _46414_ ( .A(_25064_), .B(0), .S(RST), .Y(_03339_) );
  \$mux  #( .WIDTH(32) ) _46415_ ( .A(_25065_), .B(0), .S(RST), .Y(_03345_) );
  \$mux  #( .WIDTH(32) ) _46416_ ( .A(_25066_), .B(0), .S(RST), .Y(_03224_) );
  \$mux  #( .WIDTH(32) ) _46417_ ( .A(_25067_), .B(0), .S(RST), .Y(_03223_) );
  \$mux  #( .WIDTH(32) ) _46418_ ( .A(_25068_), .B(0), .S(RST), .Y(_03222_) );
  \$mux  #( .WIDTH(32) ) _46419_ ( .A(_25069_), .B(0), .S(RST), .Y(_03221_) );
  \$mux  #( .WIDTH(32) ) _46420_ ( .A(_25070_), .B(0), .S(RST), .Y(_03239_) );
  \$mux  #( .WIDTH(32) ) _46421_ ( .A(87), .B(main_fsm), .S(_05924_), .Y({ _23237_, _23236_, _23234_, _23233_, _23232_, _23231_, _23230_, _23229_, _23228_, _23227_, _23226_, _23225_, _23223_, _23222_, _23221_, _23220_, _23219_, _23218_, _23217_, _23216_, _23215_, _23214_, _23244_, _23243_, _23242_, _23241_, _23240_, _23239_, _23238_, _23235_, _23224_, _23213_ }) );
  \$mux  #( .WIDTH(32) ) _46422_ ( .A(77), .B(main_fsm), .S(_05924_), .Y({ _23269_, _23268_, _23266_, _23265_, _23264_, _23263_, _23262_, _23261_, _23260_, _23259_, _23258_, _23257_, _23255_, _23254_, _23253_, _23252_, _23251_, _23250_, _23249_, _23248_, _23247_, _23246_, _23276_, _23275_, _23274_, _23273_, _23272_, _23271_, _23270_, _23267_, _23256_, _23245_ }) );
  \$mux  #( .WIDTH(32) ) _46423_ ( .A(67), .B(main_fsm), .S(_05924_), .Y({ _23301_, _23300_, _23298_, _23297_, _23296_, _23295_, _23294_, _23293_, _23292_, _23291_, _23290_, _23289_, _23287_, _23286_, _23285_, _23284_, _23283_, _23282_, _23281_, _23280_, _23279_, _23278_, _23308_, _23307_, _23306_, _23305_, _23304_, _23303_, _23302_, _23299_, _23288_, _23277_ }) );
  \$mux  #( .WIDTH(32) ) _46424_ ( .A(55), .B(main_fsm), .S(_05942_), .Y({ _23333_, _23332_, _23330_, _23329_, _23328_, _23327_, _23326_, _23325_, _23324_, _23323_, _23322_, _23321_, _23319_, _23318_, _23317_, _23316_, _23315_, _23314_, _23313_, _23312_, _23311_, _23310_, _23340_, _23339_, _23338_, _23337_, _23336_, _23335_, _23334_, _23331_, _23320_, _23309_ }) );
  \$mux  #( .WIDTH(32) ) _46425_ ( .A(48), .B(main_fsm), .S(_06008_), .Y({ _23365_, _23364_, _23362_, _23361_, _23360_, _23359_, _23358_, _23357_, _23356_, _23355_, _23354_, _23353_, _23351_, _23350_, _23349_, _23348_, _23347_, _23346_, _23345_, _23344_, _23343_, _23342_, _23372_, _23371_, _23370_, _23369_, _23368_, _23367_, _23366_, _23363_, _23352_, _23341_ }) );
  \$mux  #( .WIDTH(32) ) _46426_ ( .A(38), .B(main_fsm), .S(_05942_), .Y({ _23397_, _23396_, _23394_, _23393_, _23392_, _23391_, _23390_, _23389_, _23388_, _23387_, _23386_, _23385_, _23383_, _23382_, _23381_, _23380_, _23379_, _23378_, _23377_, _23376_, _23375_, _23374_, _23404_, _23403_, _23402_, _23401_, _23400_, _23399_, _23398_, _23395_, _23384_, _23373_ }) );
  \$mux  #( .WIDTH(32) ) _46427_ ( .A(31), .B(main_fsm), .S(_06008_), .Y({ _23429_, _23428_, _23426_, _23425_, _23424_, _23423_, _23422_, _23421_, _23420_, _23419_, _23418_, _23417_, _23415_, _23414_, _23413_, _23412_, _23411_, _23410_, _23409_, _23408_, _23407_, _23406_, _23436_, _23435_, _23434_, _23433_, _23432_, _23431_, _23430_, _23427_, _23416_, _23405_ }) );
  \$mux  #( .WIDTH(32) ) _46428_ ( .A(21), .B(main_fsm), .S(_05942_), .Y({ _23461_, _23460_, _23458_, _23457_, _23456_, _23455_, _23454_, _23453_, _23452_, _23451_, _23450_, _23449_, _23447_, _23446_, _23445_, _23444_, _23443_, _23442_, _23441_, _23440_, _23439_, _23438_, _23468_, _23467_, _23466_, _23465_, _23464_, _23463_, _23462_, _23459_, _23448_, _23437_ }) );
  \$mux  #( .WIDTH(32) ) _46429_ ( .A(14), .B(main_fsm), .S(_06008_), .Y({ _23493_, _23492_, _23490_, _23489_, _23488_, _23487_, _23486_, _23485_, _23484_, _23483_, _23482_, _23481_, _23479_, _23478_, _23477_, _23476_, _23475_, _23474_, _23473_, _23472_, _23471_, _23470_, _23500_, _23499_, _23498_, _23497_, _23496_, _23495_, _23494_, _23491_, _23480_, _23469_ }) );
  \$mux  #( .WIDTH(32) ) _46430_ ( .A(main_fsm), .B(1), .S(_06885_), .Y({ _23525_, _23524_, _23522_, _23521_, _23520_, _23519_, _23518_, _23517_, _23516_, _23515_, _23514_, _23513_, _23511_, _23510_, _23509_, _23508_, _23507_, _23506_, _23505_, _23504_, _23503_, _23502_, _23532_, _23531_, _23530_, _23529_, _23528_, _23527_, _23526_, _23523_, _23512_, _23501_ }) );
  \$mux  #( .WIDTH(32) ) _46431_ ( .A(_25071_), .B(0), .S(RST), .Y(_03279_) );
  \$mux  #( .WIDTH(2) ) _46432_ ( .A(_25072_), .B(2'h0), .S(RST), .Y(_03293_) );
  \$mux  #( .WIDTH(2) ) _46433_ ( .A(_25073_), .B(2'h0), .S(RST), .Y(_03344_) );
  \$mux  #( .WIDTH(2) ) _46434_ ( .A(_25074_), .B(2'h0), .S(RST), .Y(_03229_) );
  \$mux  #( .WIDTH(1) ) _46435_ ( .A(_stream_matmul_29_source_busy), .B(1'h1), .S(_stream_matmul_29_start_flag), .Y(_23534_) );
  \$mux  #( .WIDTH(1) ) _46436_ ( .A(_25075_), .B(1'h0), .S(RST), .Y(_02767_) );
  \$mux  #( .WIDTH(1) ) _46437_ ( .A(1'h0), .B(1'h1), .S(__tmp_1307_38), .Y(_25076_) );
  \$mux  #( .WIDTH(1) ) _46438_ ( .A(_25076_), .B(1'h0), .S(RST), .Y(_02769_) );
  \$mux  #( .WIDTH(1) ) _46439_ ( .A(1'h0), .B(1'h1), .S(__tmp_1305_42), .Y(_25077_) );
  \$mux  #( .WIDTH(1) ) _46440_ ( .A(_25077_), .B(1'h0), .S(RST), .Y(_02712_) );
  \$mux  #( .WIDTH(1) ) _46441_ ( .A(1'h0), .B(1'h1), .S(_stream_matmul_29_start_flag), .Y(_25078_) );
  \$mux  #( .WIDTH(1) ) _46442_ ( .A(_25078_), .B(1'h0), .S(_05685_), .Y(_25079_) );
  \$mux  #( .WIDTH(1) ) _46443_ ( .A(_25079_), .B(1'h0), .S(RST), .Y(_02768_) );
  \$mux  #( .WIDTH(32) ) _46444_ ( .A(_stream_matmul_29_fsm), .B(3), .S(_stream_matmul_29_done), .Y({ _23591_, _23590_, _23588_, _23587_, _23586_, _23585_, _23584_, _23583_, _23582_, _23581_, _23580_, _23579_, _23577_, _23576_, _23575_, _23574_, _23573_, _23572_, _23571_, _23570_, _23569_, _23568_, _23598_, _23597_, _23596_, _23595_, _23594_, _23593_, _23592_, _23589_, _23578_, _23567_ }) );
  \$mux  #( .WIDTH(32) ) _46445_ ( .A(_stream_matmul_29_fsm), .B(1), .S(_stream_matmul_29_start_flag), .Y({ _23623_, _23622_, _23620_, _23619_, _23618_, _23617_, _23616_, _23615_, _23614_, _23613_, _23612_, _23611_, _23609_, _23608_, _23607_, _23606_, _23605_, _23604_, _23603_, _23602_, _23601_, _23600_, _23630_, _23629_, _23628_, _23627_, _23626_, _23625_, _23624_, _23621_, _23610_, _23599_ }) );
  \$mux  #( .WIDTH(32) ) _46446_ ( .A(_25080_), .B(0), .S(RST), .Y(_02713_) );
  \$mux  #( .WIDTH(1) ) _46447_ ( .A(__tmp_1305_41), .B(1'h0), .S(RST), .Y(_01220_) );
  \$mux  #( .WIDTH(1) ) _46448_ ( .A(__tmp_1305_40), .B(1'h0), .S(RST), .Y(_01219_) );
  \$mux  #( .WIDTH(1) ) _46449_ ( .A(__tmp_1305_39), .B(1'h0), .S(RST), .Y(_01218_) );
  \$mux  #( .WIDTH(1) ) _46450_ ( .A(__tmp_1307_38), .B(1'h0), .S(RST), .Y(_01217_) );
  \$mux  #( .WIDTH(1) ) _46451_ ( .A(__tmp_1307_37), .B(1'h0), .S(RST), .Y(_01216_) );
  \$mux  #( .WIDTH(1) ) _46452_ ( .A(__tmp_1307_36), .B(1'h0), .S(RST), .Y(_01215_) );
  \$mux  #( .WIDTH(1) ) _46453_ ( .A(__tmp_1307_35), .B(1'h0), .S(RST), .Y(_01214_) );
  \$mux  #( .WIDTH(1) ) _46454_ ( .A(__tmp_1307_34), .B(1'h0), .S(RST), .Y(_01213_) );
  \$mux  #( .WIDTH(1) ) _46455_ ( .A(__tmp_1307_33), .B(1'h0), .S(RST), .Y(_01212_) );
  \$mux  #( .WIDTH(1) ) _46456_ ( .A(__tmp_1307_32), .B(1'h0), .S(RST), .Y(_01211_) );
  \$mux  #( .WIDTH(1) ) _46457_ ( .A(__tmp_1307_31), .B(1'h0), .S(RST), .Y(_01210_) );
  \$mux  #( .WIDTH(1) ) _46458_ ( .A(__tmp_1307_30), .B(1'h0), .S(RST), .Y(_01209_) );
  \$mux  #( .WIDTH(1) ) _46459_ ( .A(__tmp_1307_29), .B(1'h0), .S(RST), .Y(_01208_) );
  \$mux  #( .WIDTH(1) ) _46460_ ( .A(__tmp_1307_28), .B(1'h0), .S(RST), .Y(_01207_) );
  \$mux  #( .WIDTH(1) ) _46461_ ( .A(__tmp_1307_27), .B(1'h0), .S(RST), .Y(_01206_) );
  \$mux  #( .WIDTH(1) ) _46462_ ( .A(__tmp_1307_26), .B(1'h0), .S(RST), .Y(_01205_) );
  \$mux  #( .WIDTH(1) ) _46463_ ( .A(__tmp_1291_25), .B(1'h0), .S(RST), .Y(_01204_) );
  \$mux  #( .WIDTH(1) ) _46464_ ( .A(__tmp_1291_24), .B(1'h0), .S(RST), .Y(_01203_) );
  \$mux  #( .WIDTH(1) ) _46465_ ( .A(__tmp_1291_23), .B(1'h0), .S(RST), .Y(_01202_) );
  \$mux  #( .WIDTH(1) ) _46466_ ( .A(__tmp_1291_22), .B(1'h0), .S(RST), .Y(_01201_) );
  \$mux  #( .WIDTH(1) ) _46467_ ( .A(__tmp_1291_21), .B(1'h0), .S(RST), .Y(_01200_) );
  \$mux  #( .WIDTH(1) ) _46468_ ( .A(__tmp_1291_20), .B(1'h0), .S(RST), .Y(_01199_) );
  \$mux  #( .WIDTH(1) ) _46469_ ( .A(__tmp_1299_19), .B(1'h0), .S(RST), .Y(_01198_) );
  \$mux  #( .WIDTH(1) ) _46470_ ( .A(__tmp_1299_18), .B(1'h0), .S(RST), .Y(_01197_) );
  \$mux  #( .WIDTH(1) ) _46471_ ( .A(__tmp_1299_17), .B(1'h0), .S(RST), .Y(_01196_) );
  \$mux  #( .WIDTH(1) ) _46472_ ( .A(__tmp_1299_16), .B(1'h0), .S(RST), .Y(_01195_) );
  \$mux  #( .WIDTH(1) ) _46473_ ( .A(__tmp_1299_15), .B(1'h0), .S(RST), .Y(_01194_) );
  \$mux  #( .WIDTH(1) ) _46474_ ( .A(__tmp_1299_14), .B(1'h0), .S(RST), .Y(_01193_) );
  \$mux  #( .WIDTH(1) ) _46475_ ( .A(__tmp_1299_13), .B(1'h0), .S(RST), .Y(_01192_) );
  \$mux  #( .WIDTH(1) ) _46476_ ( .A(__tmp_1299_12), .B(1'h0), .S(RST), .Y(_01191_) );
  \$mux  #( .WIDTH(1) ) _46477_ ( .A(__tmp_1249_27), .B(1'h0), .S(RST), .Y(_01178_) );
  \$mux  #( .WIDTH(1) ) _46478_ ( .A(__tmp_1249_26), .B(1'h0), .S(RST), .Y(_01177_) );
  \$mux  #( .WIDTH(1) ) _46479_ ( .A(__tmp_1249_25), .B(1'h0), .S(RST), .Y(_01176_) );
  \$mux  #( .WIDTH(1) ) _46480_ ( .A(__tmp_1249_24), .B(1'h0), .S(RST), .Y(_01175_) );
  \$mux  #( .WIDTH(1) ) _46481_ ( .A(__tmp_1249_23), .B(1'h0), .S(RST), .Y(_01174_) );
  \$mux  #( .WIDTH(1) ) _46482_ ( .A(__tmp_1249_22), .B(1'h0), .S(RST), .Y(_01173_) );
  \$mux  #( .WIDTH(1) ) _46483_ ( .A(__tmp_1249_21), .B(1'h0), .S(RST), .Y(_01172_) );
  \$mux  #( .WIDTH(1) ) _46484_ ( .A(__tmp_1249_20), .B(1'h0), .S(RST), .Y(_01171_) );
  \$mux  #( .WIDTH(1) ) _46485_ ( .A(__tmp_1249_19), .B(1'h0), .S(RST), .Y(_01170_) );
  \$mux  #( .WIDTH(1) ) _46486_ ( .A(__tmp_1249_18), .B(1'h0), .S(RST), .Y(_01169_) );
  \$mux  #( .WIDTH(1) ) _46487_ ( .A(__tmp_1249_17), .B(1'h0), .S(RST), .Y(_01167_) );
  \$mux  #( .WIDTH(1) ) _46488_ ( .A(__tmp_1249_16), .B(1'h0), .S(RST), .Y(_01166_) );
  \$mux  #( .WIDTH(1) ) _46489_ ( .A(__tmp_1249_15), .B(1'h0), .S(RST), .Y(_01165_) );
  \$mux  #( .WIDTH(1) ) _46490_ ( .A(__tmp_1249_14), .B(1'h0), .S(RST), .Y(_01164_) );
  \$mux  #( .WIDTH(1) ) _46491_ ( .A(__tmp_1249_13), .B(1'h0), .S(RST), .Y(_01163_) );
  \$mux  #( .WIDTH(1) ) _46492_ ( .A(__tmp_1249_12), .B(1'h0), .S(RST), .Y(_01162_) );
  \$mux  #( .WIDTH(1) ) _46493_ ( .A(__tmp_1249_11), .B(1'h0), .S(RST), .Y(_01161_) );
  \$mux  #( .WIDTH(1) ) _46494_ ( .A(__tmp_1249_10), .B(1'h0), .S(RST), .Y(_01160_) );
  \$mux  #( .WIDTH(1) ) _46495_ ( .A(__tmp_1249_9), .B(1'h0), .S(RST), .Y(_01159_) );
  \$mux  #( .WIDTH(1) ) _46496_ ( .A(__tmp_1249_8), .B(1'h0), .S(RST), .Y(_01168_) );
  \$mux  #( .WIDTH(1) ) _46497_ ( .A(__tmp_1249_7), .B(1'h0), .S(RST), .Y(_01158_) );
  \$mux  #( .WIDTH(1) ) _46498_ ( .A(__tmp_1249_6), .B(1'h0), .S(RST), .Y(_01157_) );
  \$mux  #( .WIDTH(1) ) _46499_ ( .A(__tmp_1249_5), .B(1'h0), .S(RST), .Y(_01156_) );
  \$mux  #( .WIDTH(1) ) _46500_ ( .A(__tmp_1249_4), .B(1'h0), .S(RST), .Y(_01155_) );
  \$mux  #( .WIDTH(1) ) _46501_ ( .A(__tmp_1249_3), .B(1'h0), .S(RST), .Y(_01154_) );
  \$mux  #( .WIDTH(1) ) _46502_ ( .A(__tmp_1249_2), .B(1'h0), .S(RST), .Y(_01153_) );
  \$mux  #( .WIDTH(1) ) _46503_ ( .A(__tmp_1249_1), .B(1'h0), .S(RST), .Y(_01152_) );
  \$mux  #( .WIDTH(1) ) _46504_ ( .A(_tmp_1227), .B(1'h0), .S(RST), .Y(_01151_) );
  \$mux  #( .WIDTH(1) ) _46505_ ( .A(__stream_matmul_29_start_41), .B(1'h0), .S(RST), .Y(_01054_) );
  \$mux  #( .WIDTH(1) ) _46506_ ( .A(__stream_matmul_29_start_40), .B(1'h0), .S(RST), .Y(_01053_) );
  \$mux  #( .WIDTH(1) ) _46507_ ( .A(__stream_matmul_29_start_39), .B(1'h0), .S(RST), .Y(_01052_) );
  \$mux  #( .WIDTH(1) ) _46508_ ( .A(__stream_matmul_29_start_38), .B(1'h0), .S(RST), .Y(_01050_) );
  \$mux  #( .WIDTH(1) ) _46509_ ( .A(__stream_matmul_29_start_37), .B(1'h0), .S(RST), .Y(_01049_) );
  \$mux  #( .WIDTH(1) ) _46510_ ( .A(__stream_matmul_29_start_36), .B(1'h0), .S(RST), .Y(_01048_) );
  \$mux  #( .WIDTH(1) ) _46511_ ( .A(__stream_matmul_29_start_35), .B(1'h0), .S(RST), .Y(_01047_) );
  \$mux  #( .WIDTH(1) ) _46512_ ( .A(__stream_matmul_29_start_34), .B(1'h0), .S(RST), .Y(_01046_) );
  \$mux  #( .WIDTH(1) ) _46513_ ( .A(__stream_matmul_29_start_33), .B(1'h0), .S(RST), .Y(_01045_) );
  \$mux  #( .WIDTH(1) ) _46514_ ( .A(__stream_matmul_29_start_32), .B(1'h0), .S(RST), .Y(_01044_) );
  \$mux  #( .WIDTH(1) ) _46515_ ( .A(__stream_matmul_29_start_31), .B(1'h0), .S(RST), .Y(_01043_) );
  \$mux  #( .WIDTH(1) ) _46516_ ( .A(__stream_matmul_29_start_30), .B(1'h0), .S(RST), .Y(_01042_) );
  \$mux  #( .WIDTH(1) ) _46517_ ( .A(__stream_matmul_29_start_29), .B(1'h0), .S(RST), .Y(_01041_) );
  \$mux  #( .WIDTH(1) ) _46518_ ( .A(__stream_matmul_29_start_28), .B(1'h0), .S(RST), .Y(_01039_) );
  \$mux  #( .WIDTH(1) ) _46519_ ( .A(__stream_matmul_29_start_27), .B(1'h0), .S(RST), .Y(_01038_) );
  \$mux  #( .WIDTH(1) ) _46520_ ( .A(__stream_matmul_29_start_26), .B(1'h0), .S(RST), .Y(_01037_) );
  \$mux  #( .WIDTH(1) ) _46521_ ( .A(__stream_matmul_29_start_25), .B(1'h0), .S(RST), .Y(_01036_) );
  \$mux  #( .WIDTH(1) ) _46522_ ( .A(__stream_matmul_29_start_24), .B(1'h0), .S(RST), .Y(_01035_) );
  \$mux  #( .WIDTH(1) ) _46523_ ( .A(__stream_matmul_29_start_23), .B(1'h0), .S(RST), .Y(_01034_) );
  \$mux  #( .WIDTH(1) ) _46524_ ( .A(__stream_matmul_29_start_22), .B(1'h0), .S(RST), .Y(_01033_) );
  \$mux  #( .WIDTH(1) ) _46525_ ( .A(__stream_matmul_29_start_21), .B(1'h0), .S(RST), .Y(_01032_) );
  \$mux  #( .WIDTH(1) ) _46526_ ( .A(__stream_matmul_29_start_20), .B(1'h0), .S(RST), .Y(_01031_) );
  \$mux  #( .WIDTH(1) ) _46527_ ( .A(__stream_matmul_29_start_19), .B(1'h0), .S(RST), .Y(_01030_) );
  \$mux  #( .WIDTH(1) ) _46528_ ( .A(__stream_matmul_29_start_18), .B(1'h0), .S(RST), .Y(_01028_) );
  \$mux  #( .WIDTH(1) ) _46529_ ( .A(__stream_matmul_29_start_17), .B(1'h0), .S(RST), .Y(_01027_) );
  \$mux  #( .WIDTH(1) ) _46530_ ( .A(__stream_matmul_29_start_16), .B(1'h0), .S(RST), .Y(_01026_) );
  \$mux  #( .WIDTH(1) ) _46531_ ( .A(__stream_matmul_29_start_15), .B(1'h0), .S(RST), .Y(_01025_) );
  \$mux  #( .WIDTH(1) ) _46532_ ( .A(__stream_matmul_29_start_14), .B(1'h0), .S(RST), .Y(_01024_) );
  \$mux  #( .WIDTH(1) ) _46533_ ( .A(__stream_matmul_29_start_13), .B(1'h0), .S(RST), .Y(_01023_) );
  \$mux  #( .WIDTH(1) ) _46534_ ( .A(__stream_matmul_29_start_12), .B(1'h0), .S(RST), .Y(_01022_) );
  \$mux  #( .WIDTH(1) ) _46535_ ( .A(__stream_matmul_29_start_11), .B(1'h0), .S(RST), .Y(_01021_) );
  \$mux  #( .WIDTH(1) ) _46536_ ( .A(__stream_matmul_29_start_10), .B(1'h0), .S(RST), .Y(_01020_) );
  \$mux  #( .WIDTH(1) ) _46537_ ( .A(__stream_matmul_29_start_9), .B(1'h0), .S(RST), .Y(_01019_) );
  \$mux  #( .WIDTH(1) ) _46538_ ( .A(__stream_matmul_29_start_8), .B(1'h0), .S(RST), .Y(_01060_) );
  \$mux  #( .WIDTH(1) ) _46539_ ( .A(__stream_matmul_29_start_7), .B(1'h0), .S(RST), .Y(_01059_) );
  \$mux  #( .WIDTH(1) ) _46540_ ( .A(__stream_matmul_29_start_6), .B(1'h0), .S(RST), .Y(_01058_) );
  \$mux  #( .WIDTH(1) ) _46541_ ( .A(__stream_matmul_29_start_5), .B(1'h0), .S(RST), .Y(_01057_) );
  \$mux  #( .WIDTH(1) ) _46542_ ( .A(__stream_matmul_29_start_4), .B(1'h0), .S(RST), .Y(_01056_) );
  \$mux  #( .WIDTH(1) ) _46543_ ( .A(__stream_matmul_29_start_3), .B(1'h0), .S(RST), .Y(_01055_) );
  \$mux  #( .WIDTH(1) ) _46544_ ( .A(__stream_matmul_29_start_2), .B(1'h0), .S(RST), .Y(_01051_) );
  \$mux  #( .WIDTH(1) ) _46545_ ( .A(__stream_matmul_29_start_1), .B(1'h0), .S(RST), .Y(_01040_) );
  \$mux  #( .WIDTH(1) ) _46546_ ( .A(_stream_matmul_29_start), .B(1'h0), .S(RST), .Y(_01029_) );
  \$mux  #( .WIDTH(1) ) _46547_ ( .A(__set_flag_1224_40), .B(1'h0), .S(RST), .Y(_00749_) );
  \$mux  #( .WIDTH(1) ) _46548_ ( .A(__set_flag_1224_39), .B(1'h0), .S(RST), .Y(_00748_) );
  \$mux  #( .WIDTH(1) ) _46549_ ( .A(__set_flag_1224_38), .B(1'h0), .S(RST), .Y(_00746_) );
  \$mux  #( .WIDTH(1) ) _46550_ ( .A(__set_flag_1224_37), .B(1'h0), .S(RST), .Y(_00745_) );
  \$mux  #( .WIDTH(1) ) _46551_ ( .A(__set_flag_1224_36), .B(1'h0), .S(RST), .Y(_00744_) );
  \$mux  #( .WIDTH(1) ) _46552_ ( .A(__set_flag_1224_35), .B(1'h0), .S(RST), .Y(_00743_) );
  \$mux  #( .WIDTH(1) ) _46553_ ( .A(__set_flag_1224_34), .B(1'h0), .S(RST), .Y(_00742_) );
  \$mux  #( .WIDTH(1) ) _46554_ ( .A(__set_flag_1224_33), .B(1'h0), .S(RST), .Y(_00741_) );
  \$mux  #( .WIDTH(1) ) _46555_ ( .A(__set_flag_1224_32), .B(1'h0), .S(RST), .Y(_00740_) );
  \$mux  #( .WIDTH(1) ) _46556_ ( .A(__set_flag_1224_31), .B(1'h0), .S(RST), .Y(_00739_) );
  \$mux  #( .WIDTH(1) ) _46557_ ( .A(__set_flag_1224_30), .B(1'h0), .S(RST), .Y(_00738_) );
  \$mux  #( .WIDTH(1) ) _46558_ ( .A(__set_flag_1224_29), .B(1'h0), .S(RST), .Y(_00737_) );
  \$mux  #( .WIDTH(1) ) _46559_ ( .A(__set_flag_1224_28), .B(1'h0), .S(RST), .Y(_00735_) );
  \$mux  #( .WIDTH(1) ) _46560_ ( .A(__set_flag_1224_27), .B(1'h0), .S(RST), .Y(_00734_) );
  \$mux  #( .WIDTH(1) ) _46561_ ( .A(__set_flag_1224_26), .B(1'h0), .S(RST), .Y(_00733_) );
  \$mux  #( .WIDTH(1) ) _46562_ ( .A(__set_flag_1224_25), .B(1'h0), .S(RST), .Y(_00732_) );
  \$mux  #( .WIDTH(1) ) _46563_ ( .A(__set_flag_1224_24), .B(1'h0), .S(RST), .Y(_00731_) );
  \$mux  #( .WIDTH(1) ) _46564_ ( .A(__set_flag_1224_23), .B(1'h0), .S(RST), .Y(_00730_) );
  \$mux  #( .WIDTH(1) ) _46565_ ( .A(__set_flag_1224_22), .B(1'h0), .S(RST), .Y(_00729_) );
  \$mux  #( .WIDTH(1) ) _46566_ ( .A(__set_flag_1224_21), .B(1'h0), .S(RST), .Y(_00728_) );
  \$mux  #( .WIDTH(1) ) _46567_ ( .A(__set_flag_1224_20), .B(1'h0), .S(RST), .Y(_00727_) );
  \$mux  #( .WIDTH(1) ) _46568_ ( .A(__set_flag_1224_19), .B(1'h0), .S(RST), .Y(_00726_) );
  \$mux  #( .WIDTH(1) ) _46569_ ( .A(__set_flag_1224_18), .B(1'h0), .S(RST), .Y(_00724_) );
  \$mux  #( .WIDTH(1) ) _46570_ ( .A(__set_flag_1224_17), .B(1'h0), .S(RST), .Y(_00723_) );
  \$mux  #( .WIDTH(1) ) _46571_ ( .A(__set_flag_1224_16), .B(1'h0), .S(RST), .Y(_00722_) );
  \$mux  #( .WIDTH(1) ) _46572_ ( .A(__set_flag_1224_15), .B(1'h0), .S(RST), .Y(_00721_) );
  \$mux  #( .WIDTH(1) ) _46573_ ( .A(__set_flag_1224_14), .B(1'h0), .S(RST), .Y(_00720_) );
  \$mux  #( .WIDTH(1) ) _46574_ ( .A(__set_flag_1224_13), .B(1'h0), .S(RST), .Y(_00719_) );
  \$mux  #( .WIDTH(1) ) _46575_ ( .A(__set_flag_1224_12), .B(1'h0), .S(RST), .Y(_00718_) );
  \$mux  #( .WIDTH(1) ) _46576_ ( .A(__set_flag_1224_11), .B(1'h0), .S(RST), .Y(_00717_) );
  \$mux  #( .WIDTH(1) ) _46577_ ( .A(__set_flag_1224_10), .B(1'h0), .S(RST), .Y(_00716_) );
  \$mux  #( .WIDTH(1) ) _46578_ ( .A(__set_flag_1224_9), .B(1'h0), .S(RST), .Y(_00715_) );
  \$mux  #( .WIDTH(1) ) _46579_ ( .A(__set_flag_1224_8), .B(1'h0), .S(RST), .Y(_00755_) );
  \$mux  #( .WIDTH(1) ) _46580_ ( .A(__set_flag_1224_7), .B(1'h0), .S(RST), .Y(_00754_) );
  \$mux  #( .WIDTH(1) ) _46581_ ( .A(__set_flag_1224_6), .B(1'h0), .S(RST), .Y(_00753_) );
  \$mux  #( .WIDTH(1) ) _46582_ ( .A(__set_flag_1224_5), .B(1'h0), .S(RST), .Y(_00752_) );
  \$mux  #( .WIDTH(1) ) _46583_ ( .A(__set_flag_1224_4), .B(1'h0), .S(RST), .Y(_00751_) );
  \$mux  #( .WIDTH(1) ) _46584_ ( .A(__set_flag_1224_3), .B(1'h0), .S(RST), .Y(_00750_) );
  \$mux  #( .WIDTH(1) ) _46585_ ( .A(__set_flag_1224_2), .B(1'h0), .S(RST), .Y(_00747_) );
  \$mux  #( .WIDTH(1) ) _46586_ ( .A(__set_flag_1224_1), .B(1'h0), .S(RST), .Y(_00736_) );
  \$mux  #( .WIDTH(1) ) _46587_ ( .A(_set_flag_1224), .B(1'h0), .S(RST), .Y(_00725_) );
  \$mux  #( .WIDTH(33) ) _46588_ ( .A(__stream_matmul_29_sink_21_sink_size_1_40), .B(33'h000000000), .S(RST), .Y(_01012_) );
  \$mux  #( .WIDTH(33) ) _46589_ ( .A(__stream_matmul_29_sink_21_sink_size_1_39), .B(33'h000000000), .S(RST), .Y(_01011_) );
  \$mux  #( .WIDTH(33) ) _46590_ ( .A(__stream_matmul_29_sink_21_sink_size_1_38), .B(33'h000000000), .S(RST), .Y(_01009_) );
  \$mux  #( .WIDTH(33) ) _46591_ ( .A(__stream_matmul_29_sink_21_sink_size_1_37), .B(33'h000000000), .S(RST), .Y(_01008_) );
  \$mux  #( .WIDTH(33) ) _46592_ ( .A(__stream_matmul_29_sink_21_sink_size_1_36), .B(33'h000000000), .S(RST), .Y(_01007_) );
  \$mux  #( .WIDTH(33) ) _46593_ ( .A(__stream_matmul_29_sink_21_sink_size_1_35), .B(33'h000000000), .S(RST), .Y(_01006_) );
  \$mux  #( .WIDTH(33) ) _46594_ ( .A(__stream_matmul_29_sink_21_sink_size_1_34), .B(33'h000000000), .S(RST), .Y(_01005_) );
  \$mux  #( .WIDTH(33) ) _46595_ ( .A(__stream_matmul_29_sink_21_sink_size_1_33), .B(33'h000000000), .S(RST), .Y(_01004_) );
  \$mux  #( .WIDTH(33) ) _46596_ ( .A(__stream_matmul_29_sink_21_sink_size_1_32), .B(33'h000000000), .S(RST), .Y(_01003_) );
  \$mux  #( .WIDTH(33) ) _46597_ ( .A(__stream_matmul_29_sink_21_sink_size_1_31), .B(33'h000000000), .S(RST), .Y(_01002_) );
  \$mux  #( .WIDTH(33) ) _46598_ ( .A(__stream_matmul_29_sink_21_sink_size_1_30), .B(33'h000000000), .S(RST), .Y(_01001_) );
  \$mux  #( .WIDTH(33) ) _46599_ ( .A(__stream_matmul_29_sink_21_sink_size_1_29), .B(33'h000000000), .S(RST), .Y(_01000_) );
  \$mux  #( .WIDTH(33) ) _46600_ ( .A(__stream_matmul_29_sink_21_sink_size_1_28), .B(33'h000000000), .S(RST), .Y(_00998_) );
  \$mux  #( .WIDTH(33) ) _46601_ ( .A(__stream_matmul_29_sink_21_sink_size_1_27), .B(33'h000000000), .S(RST), .Y(_00997_) );
  \$mux  #( .WIDTH(33) ) _46602_ ( .A(__stream_matmul_29_sink_21_sink_size_1_26), .B(33'h000000000), .S(RST), .Y(_00996_) );
  \$mux  #( .WIDTH(33) ) _46603_ ( .A(__stream_matmul_29_sink_21_sink_size_1_25), .B(33'h000000000), .S(RST), .Y(_00995_) );
  \$mux  #( .WIDTH(33) ) _46604_ ( .A(__stream_matmul_29_sink_21_sink_size_1_24), .B(33'h000000000), .S(RST), .Y(_00994_) );
  \$mux  #( .WIDTH(33) ) _46605_ ( .A(__stream_matmul_29_sink_21_sink_size_1_23), .B(33'h000000000), .S(RST), .Y(_00993_) );
  \$mux  #( .WIDTH(33) ) _46606_ ( .A(__stream_matmul_29_sink_21_sink_size_1_22), .B(33'h000000000), .S(RST), .Y(_00992_) );
  \$mux  #( .WIDTH(33) ) _46607_ ( .A(__stream_matmul_29_sink_21_sink_size_1_21), .B(33'h000000000), .S(RST), .Y(_00991_) );
  \$mux  #( .WIDTH(33) ) _46608_ ( .A(__stream_matmul_29_sink_21_sink_size_1_20), .B(33'h000000000), .S(RST), .Y(_00990_) );
  \$mux  #( .WIDTH(33) ) _46609_ ( .A(__stream_matmul_29_sink_21_sink_size_1_19), .B(33'h000000000), .S(RST), .Y(_00989_) );
  \$mux  #( .WIDTH(33) ) _46610_ ( .A(__stream_matmul_29_sink_21_sink_size_1_18), .B(33'h000000000), .S(RST), .Y(_00987_) );
  \$mux  #( .WIDTH(33) ) _46611_ ( .A(__stream_matmul_29_sink_21_sink_size_1_17), .B(33'h000000000), .S(RST), .Y(_00986_) );
  \$mux  #( .WIDTH(33) ) _46612_ ( .A(__stream_matmul_29_sink_21_sink_size_1_16), .B(33'h000000000), .S(RST), .Y(_00985_) );
  \$mux  #( .WIDTH(33) ) _46613_ ( .A(__stream_matmul_29_sink_21_sink_size_1_15), .B(33'h000000000), .S(RST), .Y(_00984_) );
  \$mux  #( .WIDTH(33) ) _46614_ ( .A(__stream_matmul_29_sink_21_sink_size_1_14), .B(33'h000000000), .S(RST), .Y(_00983_) );
  \$mux  #( .WIDTH(33) ) _46615_ ( .A(__stream_matmul_29_sink_21_sink_size_1_13), .B(33'h000000000), .S(RST), .Y(_00982_) );
  \$mux  #( .WIDTH(33) ) _46616_ ( .A(__stream_matmul_29_sink_21_sink_size_1_12), .B(33'h000000000), .S(RST), .Y(_00981_) );
  \$mux  #( .WIDTH(33) ) _46617_ ( .A(__stream_matmul_29_sink_21_sink_size_1_11), .B(33'h000000000), .S(RST), .Y(_00980_) );
  \$mux  #( .WIDTH(33) ) _46618_ ( .A(__stream_matmul_29_sink_21_sink_size_1_10), .B(33'h000000000), .S(RST), .Y(_00979_) );
  \$mux  #( .WIDTH(33) ) _46619_ ( .A(__stream_matmul_29_sink_21_sink_size_1_9), .B(33'h000000000), .S(RST), .Y(_00978_) );
  \$mux  #( .WIDTH(33) ) _46620_ ( .A(__stream_matmul_29_sink_21_sink_size_1_8), .B(33'h000000000), .S(RST), .Y(_01018_) );
  \$mux  #( .WIDTH(33) ) _46621_ ( .A(__stream_matmul_29_sink_21_sink_size_1_7), .B(33'h000000000), .S(RST), .Y(_01017_) );
  \$mux  #( .WIDTH(33) ) _46622_ ( .A(__stream_matmul_29_sink_21_sink_size_1_6), .B(33'h000000000), .S(RST), .Y(_01016_) );
  \$mux  #( .WIDTH(33) ) _46623_ ( .A(__stream_matmul_29_sink_21_sink_size_1_5), .B(33'h000000000), .S(RST), .Y(_01015_) );
  \$mux  #( .WIDTH(33) ) _46624_ ( .A(__stream_matmul_29_sink_21_sink_size_1_4), .B(33'h000000000), .S(RST), .Y(_01014_) );
  \$mux  #( .WIDTH(33) ) _46625_ ( .A(__stream_matmul_29_sink_21_sink_size_1_3), .B(33'h000000000), .S(RST), .Y(_01013_) );
  \$mux  #( .WIDTH(33) ) _46626_ ( .A(__stream_matmul_29_sink_21_sink_size_1_2), .B(33'h000000000), .S(RST), .Y(_01010_) );
  \$mux  #( .WIDTH(33) ) _46627_ ( .A(__stream_matmul_29_sink_21_sink_size_1_1), .B(33'h000000000), .S(RST), .Y(_00999_) );
  \$mux  #( .WIDTH(33) ) _46628_ ( .A({ 1'h0, matmul_29_next_stream_num_ops }), .B(33'h000000000), .S(RST), .Y(_00988_) );
  \$mux  #( .WIDTH(32) ) _46629_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_40), .B(0), .S(RST), .Y(_00971_) );
  \$mux  #( .WIDTH(32) ) _46630_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_39), .B(0), .S(RST), .Y(_00970_) );
  \$mux  #( .WIDTH(32) ) _46631_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_38), .B(0), .S(RST), .Y(_00968_) );
  \$mux  #( .WIDTH(32) ) _46632_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_37), .B(0), .S(RST), .Y(_00967_) );
  \$mux  #( .WIDTH(32) ) _46633_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_36), .B(0), .S(RST), .Y(_00966_) );
  \$mux  #( .WIDTH(32) ) _46634_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_35), .B(0), .S(RST), .Y(_00965_) );
  \$mux  #( .WIDTH(32) ) _46635_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_34), .B(0), .S(RST), .Y(_00964_) );
  \$mux  #( .WIDTH(32) ) _46636_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_33), .B(0), .S(RST), .Y(_00963_) );
  \$mux  #( .WIDTH(32) ) _46637_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_32), .B(0), .S(RST), .Y(_00962_) );
  \$mux  #( .WIDTH(32) ) _46638_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_31), .B(0), .S(RST), .Y(_00961_) );
  \$mux  #( .WIDTH(32) ) _46639_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_30), .B(0), .S(RST), .Y(_00960_) );
  \$mux  #( .WIDTH(32) ) _46640_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_29), .B(0), .S(RST), .Y(_00959_) );
  \$mux  #( .WIDTH(32) ) _46641_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_28), .B(0), .S(RST), .Y(_00957_) );
  \$mux  #( .WIDTH(32) ) _46642_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_27), .B(0), .S(RST), .Y(_00956_) );
  \$mux  #( .WIDTH(32) ) _46643_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_26), .B(0), .S(RST), .Y(_00955_) );
  \$mux  #( .WIDTH(32) ) _46644_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_25), .B(0), .S(RST), .Y(_00954_) );
  \$mux  #( .WIDTH(32) ) _46645_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_24), .B(0), .S(RST), .Y(_00953_) );
  \$mux  #( .WIDTH(32) ) _46646_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_23), .B(0), .S(RST), .Y(_00952_) );
  \$mux  #( .WIDTH(32) ) _46647_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_22), .B(0), .S(RST), .Y(_00951_) );
  \$mux  #( .WIDTH(32) ) _46648_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_21), .B(0), .S(RST), .Y(_00950_) );
  \$mux  #( .WIDTH(32) ) _46649_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_20), .B(0), .S(RST), .Y(_00949_) );
  \$mux  #( .WIDTH(32) ) _46650_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_19), .B(0), .S(RST), .Y(_00948_) );
  \$mux  #( .WIDTH(32) ) _46651_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_18), .B(0), .S(RST), .Y(_00946_) );
  \$mux  #( .WIDTH(32) ) _46652_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_17), .B(0), .S(RST), .Y(_00945_) );
  \$mux  #( .WIDTH(32) ) _46653_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_16), .B(0), .S(RST), .Y(_00944_) );
  \$mux  #( .WIDTH(32) ) _46654_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_15), .B(0), .S(RST), .Y(_00943_) );
  \$mux  #( .WIDTH(32) ) _46655_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_14), .B(0), .S(RST), .Y(_00942_) );
  \$mux  #( .WIDTH(32) ) _46656_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_13), .B(0), .S(RST), .Y(_00941_) );
  \$mux  #( .WIDTH(32) ) _46657_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_12), .B(0), .S(RST), .Y(_00940_) );
  \$mux  #( .WIDTH(32) ) _46658_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_11), .B(0), .S(RST), .Y(_00939_) );
  \$mux  #( .WIDTH(32) ) _46659_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_10), .B(0), .S(RST), .Y(_00938_) );
  \$mux  #( .WIDTH(32) ) _46660_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_9), .B(0), .S(RST), .Y(_00937_) );
  \$mux  #( .WIDTH(32) ) _46661_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_8), .B(0), .S(RST), .Y(_00977_) );
  \$mux  #( .WIDTH(32) ) _46662_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_7), .B(0), .S(RST), .Y(_00976_) );
  \$mux  #( .WIDTH(32) ) _46663_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_6), .B(0), .S(RST), .Y(_00975_) );
  \$mux  #( .WIDTH(32) ) _46664_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_5), .B(0), .S(RST), .Y(_00974_) );
  \$mux  #( .WIDTH(32) ) _46665_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_4), .B(0), .S(RST), .Y(_00973_) );
  \$mux  #( .WIDTH(32) ) _46666_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_3), .B(0), .S(RST), .Y(_00972_) );
  \$mux  #( .WIDTH(32) ) _46667_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_2), .B(0), .S(RST), .Y(_00969_) );
  \$mux  #( .WIDTH(32) ) _46668_ ( .A(__stream_matmul_29_sink_21_sink_offset_0_1), .B(0), .S(RST), .Y(_00958_) );
  \$mux  #( .WIDTH(32) ) _46669_ ( .A(_24428_), .B(0), .S(RST), .Y(_00947_) );
  \$mux  #( .WIDTH(4) ) _46670_ ( .A(__variable_wdata_864), .B(_stream_matmul_29_source_20_source_ram_rdata), .S(_stream_matmul_29_source_20_source_ram_rvalid), .Y(_25082_) );
  \$mux  #( .WIDTH(4) ) _46671_ ( .A(_25082_), .B(4'h0), .S(RST), .Y(_01462_) );
  \$mux  #( .WIDTH(1) ) _46672_ ( .A(_tmp_1223), .B(1'h0), .S(RST), .Y(_01150_) );
  \$mux  #( .WIDTH(32) ) _46673_ ( .A(_source_stream_matmul_29_source_20_pat_stride_buf_3), .B(_source_stream_matmul_29_source_20_pat_stride_3), .S(_06810_), .Y(_25083_) );
  \$mux  #( .WIDTH(32) ) _46674_ ( .A(_25083_), .B(0), .S(RST), .Y(_02411_) );
  \$mux  #( .WIDTH(32) ) _46675_ ( .A(_source_stream_matmul_29_source_20_pat_stride_buf_2), .B(_source_stream_matmul_29_source_20_pat_stride_2), .S(_06810_), .Y(_25084_) );
  \$mux  #( .WIDTH(32) ) _46676_ ( .A(_25084_), .B(0), .S(RST), .Y(_02410_) );
  \$mux  #( .WIDTH(32) ) _46677_ ( .A(_source_stream_matmul_29_source_20_pat_stride_buf_1), .B(_source_stream_matmul_29_source_20_pat_stride_1), .S(_06810_), .Y(_25085_) );
  \$mux  #( .WIDTH(32) ) _46678_ ( .A(_25085_), .B(0), .S(RST), .Y(_02409_) );
  \$mux  #( .WIDTH(32) ) _46679_ ( .A(_source_stream_matmul_29_source_20_pat_stride_buf_0), .B(_source_stream_matmul_29_source_20_pat_stride_0), .S(_06810_), .Y(_25086_) );
  \$mux  #( .WIDTH(32) ) _46680_ ( .A(_25086_), .B(0), .S(RST), .Y(_02408_) );
  \$mux  #( .WIDTH(33) ) _46681_ ( .A(_source_stream_matmul_29_source_20_pat_size_buf_3), .B(_source_stream_matmul_29_source_20_pat_size_3), .S(_06810_), .Y(_25087_) );
  \$mux  #( .WIDTH(33) ) _46682_ ( .A(_25087_), .B(33'h000000000), .S(RST), .Y(_02403_) );
  \$mux  #( .WIDTH(33) ) _46683_ ( .A(_source_stream_matmul_29_source_20_pat_size_buf_2), .B(_source_stream_matmul_29_source_20_pat_size_2), .S(_06810_), .Y(_25088_) );
  \$mux  #( .WIDTH(33) ) _46684_ ( .A(_25088_), .B(33'h000000000), .S(RST), .Y(_02402_) );
  \$mux  #( .WIDTH(33) ) _46685_ ( .A(_source_stream_matmul_29_source_20_pat_size_buf_1), .B(_source_stream_matmul_29_source_20_pat_size_1), .S(_06810_), .Y(_25089_) );
  \$mux  #( .WIDTH(33) ) _46686_ ( .A(_25089_), .B(33'h000000000), .S(RST), .Y(_02401_) );
  \$mux  #( .WIDTH(33) ) _46687_ ( .A(_source_stream_matmul_29_source_20_pat_size_buf_0), .B(_source_stream_matmul_29_source_20_pat_size_0), .S(_06810_), .Y(_25090_) );
  \$mux  #( .WIDTH(33) ) _46688_ ( .A(_25090_), .B(33'h000000000), .S(RST), .Y(_02400_) );
  \$mux  #( .WIDTH(33) ) _46689_ ( .A(_source_stream_matmul_29_source_20_pat_count_3), .B(_28924_), .S(_06810_), .Y(_25091_) );
  \$mux  #( .WIDTH(33) ) _46690_ ( .A(_25091_), .B(_28931_), .S(_06813_), .Y(_25092_) );
  \$mux  #( .WIDTH(33) ) _46691_ ( .A(_25092_), .B(_28932_), .S(_06814_), .Y(_25093_) );
  \$mux  #( .WIDTH(33) ) _46692_ ( .A(_25093_), .B(33'h000000000), .S(RST), .Y(_02391_) );
  \$mux  #( .WIDTH(33) ) _46693_ ( .A(_source_stream_matmul_29_source_20_pat_count_2), .B(_28923_), .S(_06810_), .Y(_25094_) );
  \$mux  #( .WIDTH(33) ) _46694_ ( .A(_25094_), .B(_28929_), .S(_06812_), .Y(_25095_) );
  \$mux  #( .WIDTH(33) ) _46695_ ( .A(_25095_), .B(_28930_), .S(_06813_), .Y(_25096_) );
  \$mux  #( .WIDTH(33) ) _46696_ ( .A(_25096_), .B(33'h000000000), .S(RST), .Y(_02390_) );
  \$mux  #( .WIDTH(33) ) _46697_ ( .A(_source_stream_matmul_29_source_20_pat_count_1), .B(_28922_), .S(_06810_), .Y(_25097_) );
  \$mux  #( .WIDTH(33) ) _46698_ ( .A(_25097_), .B(_28927_), .S(_06811_), .Y(_25098_) );
  \$mux  #( .WIDTH(33) ) _46699_ ( .A(_25098_), .B(_28928_), .S(_06812_), .Y(_25099_) );
  \$mux  #( .WIDTH(33) ) _46700_ ( .A(_25099_), .B(33'h000000000), .S(RST), .Y(_02389_) );
  \$mux  #( .WIDTH(33) ) _46701_ ( .A(_source_stream_matmul_29_source_20_pat_count_0), .B(_28921_), .S(_06810_), .Y(_25100_) );
  \$mux  #( .WIDTH(33) ) _46702_ ( .A(_28925_), .B(_25100_), .S(_05909_), .Y(_25101_) );
  \$mux  #( .WIDTH(33) ) _46703_ ( .A(_25101_), .B(_28926_), .S(_06811_), .Y(_25102_) );
  \$mux  #( .WIDTH(33) ) _46704_ ( .A(_25102_), .B(33'h000000000), .S(RST), .Y(_02388_) );
  \$mux  #( .WIDTH(32) ) _46705_ ( .A(_source_stream_matmul_29_source_20_pat_stride_3), .B(0), .S(_set_flag_1224), .Y(_25103_) );
  \$mux  #( .WIDTH(32) ) _46706_ ( .A(_25103_), .B(0), .S(RST), .Y(_02407_) );
  \$mux  #( .WIDTH(32) ) _46707_ ( .A(_source_stream_matmul_29_source_20_pat_stride_2), .B(0), .S(_set_flag_1224), .Y(_25104_) );
  \$mux  #( .WIDTH(32) ) _46708_ ( .A(_25104_), .B(0), .S(RST), .Y(_02406_) );
  \$mux  #( .WIDTH(32) ) _46709_ ( .A(_source_stream_matmul_29_source_20_pat_stride_1), .B({ 21'h000000, cparam_matmul_29_act_bat_step }), .S(_set_flag_1224), .Y(_25105_) );
  \$mux  #( .WIDTH(32) ) _46710_ ( .A(_25105_), .B(0), .S(RST), .Y(_02405_) );
  \$mux  #( .WIDTH(32) ) _46711_ ( .A(_source_stream_matmul_29_source_20_pat_stride_0), .B(1), .S(_set_flag_1224), .Y(_25106_) );
  \$mux  #( .WIDTH(32) ) _46712_ ( .A(_25106_), .B(0), .S(RST), .Y(_02404_) );
  \$mux  #( .WIDTH(33) ) _46713_ ( .A(_source_stream_matmul_29_source_20_pat_size_3), .B(33'h000000001), .S(_set_flag_1224), .Y(_25107_) );
  \$mux  #( .WIDTH(33) ) _46714_ ( .A(_25107_), .B(33'h000000000), .S(RST), .Y(_02399_) );
  \$mux  #( .WIDTH(33) ) _46715_ ( .A(_source_stream_matmul_29_source_20_pat_size_2), .B(33'h000000001), .S(_set_flag_1224), .Y(_25108_) );
  \$mux  #( .WIDTH(33) ) _46716_ ( .A(_25108_), .B(33'h000000000), .S(RST), .Y(_02398_) );
  \$mux  #( .WIDTH(33) ) _46717_ ( .A(_source_stream_matmul_29_source_20_pat_size_1), .B({ 1'h0, matmul_29_next_stream_num_ops }), .S(_set_flag_1224), .Y(_25109_) );
  \$mux  #( .WIDTH(33) ) _46718_ ( .A(_25109_), .B(33'h000000000), .S(RST), .Y(_02397_) );
  \$mux  #( .WIDTH(33) ) _46719_ ( .A(_source_stream_matmul_29_source_20_pat_size_0), .B({ 22'h000000, cparam_matmul_29_act_bat_step }), .S(_set_flag_1224), .Y(_25110_) );
  \$mux  #( .WIDTH(33) ) _46720_ ( .A(_25110_), .B(33'h000000000), .S(RST), .Y(_02396_) );
  \$mux  #( .WIDTH(32) ) _46721_ ( .A(_source_stream_matmul_29_source_20_pat_cur_offset_3), .B(0), .S(_06810_), .Y(_25111_) );
  \$mux  #( .WIDTH(32) ) _46722_ ( .A(_25111_), .B(_24427_), .S(_06813_), .Y(_25112_) );
  \$mux  #( .WIDTH(32) ) _46723_ ( .A(_25112_), .B(0), .S(_06814_), .Y(_25113_) );
  \$mux  #( .WIDTH(32) ) _46724_ ( .A(_25113_), .B(0), .S(RST), .Y(_02395_) );
  \$mux  #( .WIDTH(32) ) _46725_ ( .A(_source_stream_matmul_29_source_20_pat_cur_offset_2), .B(0), .S(_06810_), .Y(_25114_) );
  \$mux  #( .WIDTH(32) ) _46726_ ( .A(_25114_), .B(_24426_), .S(_06812_), .Y(_25115_) );
  \$mux  #( .WIDTH(32) ) _46727_ ( .A(_25115_), .B(0), .S(_06813_), .Y(_25116_) );
  \$mux  #( .WIDTH(32) ) _46728_ ( .A(_25116_), .B(0), .S(RST), .Y(_02394_) );
  \$mux  #( .WIDTH(32) ) _46729_ ( .A(_source_stream_matmul_29_source_20_pat_cur_offset_1), .B(0), .S(_06810_), .Y(_25117_) );
  \$mux  #( .WIDTH(32) ) _46730_ ( .A(_25117_), .B(_24425_), .S(_06811_), .Y(_25118_) );
  \$mux  #( .WIDTH(32) ) _46731_ ( .A(_25118_), .B(0), .S(_06812_), .Y(_25119_) );
  \$mux  #( .WIDTH(32) ) _46732_ ( .A(_25119_), .B(0), .S(RST), .Y(_02393_) );
  \$mux  #( .WIDTH(32) ) _46733_ ( .A(_source_stream_matmul_29_source_20_pat_cur_offset_0), .B(0), .S(_06810_), .Y(_25120_) );
  \$mux  #( .WIDTH(32) ) _46734_ ( .A(_24424_), .B(_25120_), .S(_05909_), .Y(_25121_) );
  \$mux  #( .WIDTH(32) ) _46735_ ( .A(_25121_), .B(0), .S(_06811_), .Y(_25122_) );
  \$mux  #( .WIDTH(32) ) _46736_ ( .A(_25122_), .B(0), .S(RST), .Y(_02392_) );
  \$mux  #( .WIDTH(8) ) _46737_ ( .A(__variable_wdata_850), .B(_stream_matmul_29_source_19_source_ram_rdata), .S(_stream_matmul_29_source_19_source_ram_rvalid), .Y(_25123_) );
  \$mux  #( .WIDTH(8) ) _46738_ ( .A(_25123_), .B(8'h00), .S(RST), .Y(_01461_) );
  \$mux  #( .WIDTH(32) ) _46739_ ( .A(_source_stream_matmul_29_source_19_pat_stride_buf_3), .B(_source_stream_matmul_29_source_19_pat_stride_3), .S(_06805_), .Y(_25124_) );
  \$mux  #( .WIDTH(32) ) _46740_ ( .A(_25124_), .B(0), .S(RST), .Y(_02387_) );
  \$mux  #( .WIDTH(32) ) _46741_ ( .A(_source_stream_matmul_29_source_19_pat_stride_buf_2), .B(_source_stream_matmul_29_source_19_pat_stride_2), .S(_06805_), .Y(_25125_) );
  \$mux  #( .WIDTH(32) ) _46742_ ( .A(_25125_), .B(0), .S(RST), .Y(_02386_) );
  \$mux  #( .WIDTH(32) ) _46743_ ( .A(_source_stream_matmul_29_source_19_pat_stride_buf_1), .B(_source_stream_matmul_29_source_19_pat_stride_1), .S(_06805_), .Y(_25126_) );
  \$mux  #( .WIDTH(32) ) _46744_ ( .A(_25126_), .B(0), .S(RST), .Y(_02385_) );
  \$mux  #( .WIDTH(32) ) _46745_ ( .A(_source_stream_matmul_29_source_19_pat_stride_buf_0), .B(_source_stream_matmul_29_source_19_pat_stride_0), .S(_06805_), .Y(_25127_) );
  \$mux  #( .WIDTH(32) ) _46746_ ( .A(_25127_), .B(0), .S(RST), .Y(_02384_) );
  \$mux  #( .WIDTH(33) ) _46747_ ( .A(_source_stream_matmul_29_source_19_pat_size_buf_3), .B(_source_stream_matmul_29_source_19_pat_size_3), .S(_06805_), .Y(_25128_) );
  \$mux  #( .WIDTH(33) ) _46748_ ( .A(_25128_), .B(33'h000000000), .S(RST), .Y(_02379_) );
  \$mux  #( .WIDTH(33) ) _46749_ ( .A(_source_stream_matmul_29_source_19_pat_size_buf_2), .B(_source_stream_matmul_29_source_19_pat_size_2), .S(_06805_), .Y(_25129_) );
  \$mux  #( .WIDTH(33) ) _46750_ ( .A(_25129_), .B(33'h000000000), .S(RST), .Y(_02378_) );
  \$mux  #( .WIDTH(33) ) _46751_ ( .A(_source_stream_matmul_29_source_19_pat_size_buf_1), .B(_source_stream_matmul_29_source_19_pat_size_1), .S(_06805_), .Y(_25130_) );
  \$mux  #( .WIDTH(33) ) _46752_ ( .A(_25130_), .B(33'h000000000), .S(RST), .Y(_02377_) );
  \$mux  #( .WIDTH(33) ) _46753_ ( .A(_source_stream_matmul_29_source_19_pat_size_buf_0), .B(_source_stream_matmul_29_source_19_pat_size_0), .S(_06805_), .Y(_25131_) );
  \$mux  #( .WIDTH(33) ) _46754_ ( .A(_25131_), .B(33'h000000000), .S(RST), .Y(_02376_) );
  \$mux  #( .WIDTH(33) ) _46755_ ( .A(_source_stream_matmul_29_source_19_pat_count_3), .B(_28912_), .S(_06805_), .Y(_25132_) );
  \$mux  #( .WIDTH(33) ) _46756_ ( .A(_25132_), .B(_28919_), .S(_06808_), .Y(_25133_) );
  \$mux  #( .WIDTH(33) ) _46757_ ( .A(_25133_), .B(_28920_), .S(_06809_), .Y(_25134_) );
  \$mux  #( .WIDTH(33) ) _46758_ ( .A(_25134_), .B(33'h000000000), .S(RST), .Y(_02367_) );
  \$mux  #( .WIDTH(33) ) _46759_ ( .A(_source_stream_matmul_29_source_19_pat_count_2), .B(_28911_), .S(_06805_), .Y(_25135_) );
  \$mux  #( .WIDTH(33) ) _46760_ ( .A(_25135_), .B(_28917_), .S(_06807_), .Y(_25136_) );
  \$mux  #( .WIDTH(33) ) _46761_ ( .A(_25136_), .B(_28918_), .S(_06808_), .Y(_25137_) );
  \$mux  #( .WIDTH(33) ) _46762_ ( .A(_25137_), .B(33'h000000000), .S(RST), .Y(_02366_) );
  \$mux  #( .WIDTH(33) ) _46763_ ( .A(_source_stream_matmul_29_source_19_pat_count_1), .B(_28910_), .S(_06805_), .Y(_25138_) );
  \$mux  #( .WIDTH(33) ) _46764_ ( .A(_25138_), .B(_28915_), .S(_06806_), .Y(_25139_) );
  \$mux  #( .WIDTH(33) ) _46765_ ( .A(_25139_), .B(_28916_), .S(_06807_), .Y(_25140_) );
  \$mux  #( .WIDTH(33) ) _46766_ ( .A(_25140_), .B(33'h000000000), .S(RST), .Y(_02365_) );
  \$mux  #( .WIDTH(33) ) _46767_ ( .A(_source_stream_matmul_29_source_19_pat_count_0), .B(_28909_), .S(_06805_), .Y(_25141_) );
  \$mux  #( .WIDTH(33) ) _46768_ ( .A(_28913_), .B(_25141_), .S(_05913_), .Y(_25142_) );
  \$mux  #( .WIDTH(33) ) _46769_ ( .A(_25142_), .B(_28914_), .S(_06806_), .Y(_25143_) );
  \$mux  #( .WIDTH(33) ) _46770_ ( .A(_25143_), .B(33'h000000000), .S(RST), .Y(_02364_) );
  \$mux  #( .WIDTH(32) ) _46771_ ( .A(_source_stream_matmul_29_source_19_pat_stride_3), .B(0), .S(_set_flag_1224), .Y(_25144_) );
  \$mux  #( .WIDTH(32) ) _46772_ ( .A(_25144_), .B(0), .S(RST), .Y(_02383_) );
  \$mux  #( .WIDTH(32) ) _46773_ ( .A(_source_stream_matmul_29_source_19_pat_stride_2), .B(0), .S(_set_flag_1224), .Y(_25145_) );
  \$mux  #( .WIDTH(32) ) _46774_ ( .A(_25145_), .B(0), .S(RST), .Y(_02382_) );
  \$mux  #( .WIDTH(32) ) _46775_ ( .A(_source_stream_matmul_29_source_19_pat_stride_1), .B(0), .S(_set_flag_1224), .Y(_25146_) );
  \$mux  #( .WIDTH(32) ) _46776_ ( .A(_25146_), .B(0), .S(RST), .Y(_02381_) );
  \$mux  #( .WIDTH(32) ) _46777_ ( .A(_source_stream_matmul_29_source_19_pat_stride_0), .B(1), .S(_set_flag_1224), .Y(_25147_) );
  \$mux  #( .WIDTH(32) ) _46778_ ( .A(_25147_), .B(0), .S(RST), .Y(_02380_) );
  \$mux  #( .WIDTH(33) ) _46779_ ( .A(_source_stream_matmul_29_source_19_pat_size_3), .B(33'h000000001), .S(_set_flag_1224), .Y(_25148_) );
  \$mux  #( .WIDTH(33) ) _46780_ ( .A(_25148_), .B(33'h000000000), .S(RST), .Y(_02375_) );
  \$mux  #( .WIDTH(33) ) _46781_ ( .A(_source_stream_matmul_29_source_19_pat_size_2), .B(33'h000000001), .S(_set_flag_1224), .Y(_25149_) );
  \$mux  #( .WIDTH(33) ) _46782_ ( .A(_25149_), .B(33'h000000000), .S(RST), .Y(_02374_) );
  \$mux  #( .WIDTH(33) ) _46783_ ( .A(_source_stream_matmul_29_source_19_pat_size_1), .B({ 1'h0, matmul_29_next_stream_num_ops }), .S(_set_flag_1224), .Y(_25150_) );
  \$mux  #( .WIDTH(33) ) _46784_ ( .A(_25150_), .B(33'h000000000), .S(RST), .Y(_02373_) );
  \$mux  #( .WIDTH(33) ) _46785_ ( .A(_source_stream_matmul_29_source_19_pat_size_0), .B({ 22'h000000, cparam_matmul_29_act_bat_step }), .S(_set_flag_1224), .Y(_25151_) );
  \$mux  #( .WIDTH(33) ) _46786_ ( .A(_25151_), .B(33'h000000000), .S(RST), .Y(_02372_) );
  \$mux  #( .WIDTH(32) ) _46787_ ( .A(_source_stream_matmul_29_source_19_pat_cur_offset_3), .B(0), .S(_06805_), .Y(_25152_) );
  \$mux  #( .WIDTH(32) ) _46788_ ( .A(_25152_), .B(_24423_), .S(_06808_), .Y(_25153_) );
  \$mux  #( .WIDTH(32) ) _46789_ ( .A(_25153_), .B(0), .S(_06809_), .Y(_25154_) );
  \$mux  #( .WIDTH(32) ) _46790_ ( .A(_25154_), .B(0), .S(RST), .Y(_02371_) );
  \$mux  #( .WIDTH(32) ) _46791_ ( .A(_source_stream_matmul_29_source_19_pat_cur_offset_2), .B(0), .S(_06805_), .Y(_25155_) );
  \$mux  #( .WIDTH(32) ) _46792_ ( .A(_25155_), .B(_24422_), .S(_06807_), .Y(_25156_) );
  \$mux  #( .WIDTH(32) ) _46793_ ( .A(_25156_), .B(0), .S(_06808_), .Y(_25157_) );
  \$mux  #( .WIDTH(32) ) _46794_ ( .A(_25157_), .B(0), .S(RST), .Y(_02370_) );
  \$mux  #( .WIDTH(32) ) _46795_ ( .A(_source_stream_matmul_29_source_19_pat_cur_offset_1), .B(0), .S(_06805_), .Y(_25158_) );
  \$mux  #( .WIDTH(32) ) _46796_ ( .A(_25158_), .B(_24421_), .S(_06806_), .Y(_25159_) );
  \$mux  #( .WIDTH(32) ) _46797_ ( .A(_25159_), .B(0), .S(_06807_), .Y(_25160_) );
  \$mux  #( .WIDTH(32) ) _46798_ ( .A(_25160_), .B(0), .S(RST), .Y(_02369_) );
  \$mux  #( .WIDTH(32) ) _46799_ ( .A(_source_stream_matmul_29_source_19_pat_cur_offset_0), .B(0), .S(_06805_), .Y(_25161_) );
  \$mux  #( .WIDTH(32) ) _46800_ ( .A(_24420_), .B(_25161_), .S(_05913_), .Y(_25162_) );
  \$mux  #( .WIDTH(32) ) _46801_ ( .A(_25162_), .B(0), .S(_06806_), .Y(_25163_) );
  \$mux  #( .WIDTH(32) ) _46802_ ( .A(_25163_), .B(0), .S(RST), .Y(_02368_) );
  \$mux  #( .WIDTH(2) ) _46803_ ( .A(__variable_wdata_849), .B(_stream_matmul_29_constant_18_next_constant_data), .S(_stream_matmul_29_start), .Y(_25164_) );
  \$mux  #( .WIDTH(2) ) _46804_ ( .A(_25164_), .B(2'h0), .S(RST), .Y(_01460_) );
  \$mux  #( .WIDTH(4) ) _46805_ ( .A(__variable_wdata_848), .B(_stream_matmul_29_constant_17_next_constant_data), .S(_stream_matmul_29_start), .Y(_25165_) );
  \$mux  #( .WIDTH(4) ) _46806_ ( .A(_25165_), .B(4'h0), .S(RST), .Y(_01459_) );
  \$mux  #( .WIDTH(1) ) _46807_ ( .A(__variable_wdata_847), .B(_stream_matmul_29_constant_16_next_constant_data), .S(_stream_matmul_29_start), .Y(_25166_) );
  \$mux  #( .WIDTH(1) ) _46808_ ( .A(_25166_), .B(1'h0), .S(RST), .Y(_01458_) );
  \$mux  #( .WIDTH(1) ) _46809_ ( .A(__variable_wdata_846), .B(_stream_matmul_29_constant_15_next_constant_data), .S(_stream_matmul_29_start), .Y(_25167_) );
  \$mux  #( .WIDTH(1) ) _46810_ ( .A(_25167_), .B(1'h0), .S(RST), .Y(_01457_) );
  \$mux  #( .WIDTH(8) ) _46811_ ( .A(__variable_wdata_840), .B(_stream_matmul_29_source_14_source_empty_data), .S(_stream_matmul_29_start), .Y(_25168_) );
  \$mux  #( .WIDTH(8) ) _46812_ ( .A(_25168_), .B(8'h00), .S(RST), .Y(_01456_) );
  \$mux  #( .WIDTH(8) ) _46813_ ( .A(__variable_wdata_833), .B(_stream_matmul_29_source_12_source_empty_data), .S(_stream_matmul_29_start), .Y(_25169_) );
  \$mux  #( .WIDTH(8) ) _46814_ ( .A(_25169_), .B(8'h00), .S(RST), .Y(_01455_) );
  \$mux  #( .WIDTH(8) ) _46815_ ( .A(__variable_wdata_826), .B(_stream_matmul_29_source_10_source_empty_data), .S(_stream_matmul_29_start), .Y(_25170_) );
  \$mux  #( .WIDTH(8) ) _46816_ ( .A(_25170_), .B(8'h00), .S(RST), .Y(_01454_) );
  \$mux  #( .WIDTH(8) ) _46817_ ( .A(__variable_wdata_819), .B(_stream_matmul_29_source_8_source_ram_rdata), .S(_stream_matmul_29_source_8_source_ram_rvalid), .Y(_25171_) );
  \$mux  #( .WIDTH(8) ) _46818_ ( .A(_25171_), .B(8'h00), .S(RST), .Y(_01453_) );
  \$mux  #( .WIDTH(32) ) _46819_ ( .A(_source_stream_matmul_29_source_8_pat_stride_buf_3), .B(_source_stream_matmul_29_source_8_pat_stride_3), .S(_06800_), .Y(_25172_) );
  \$mux  #( .WIDTH(32) ) _46820_ ( .A(_25172_), .B(0), .S(RST), .Y(_02459_) );
  \$mux  #( .WIDTH(32) ) _46821_ ( .A(_source_stream_matmul_29_source_8_pat_stride_buf_2), .B(_source_stream_matmul_29_source_8_pat_stride_2), .S(_06800_), .Y(_25173_) );
  \$mux  #( .WIDTH(32) ) _46822_ ( .A(_25173_), .B(0), .S(RST), .Y(_02458_) );
  \$mux  #( .WIDTH(32) ) _46823_ ( .A(_source_stream_matmul_29_source_8_pat_stride_buf_1), .B(_source_stream_matmul_29_source_8_pat_stride_1), .S(_06800_), .Y(_25174_) );
  \$mux  #( .WIDTH(32) ) _46824_ ( .A(_25174_), .B(0), .S(RST), .Y(_02457_) );
  \$mux  #( .WIDTH(32) ) _46825_ ( .A(_source_stream_matmul_29_source_8_pat_stride_buf_0), .B(_source_stream_matmul_29_source_8_pat_stride_0), .S(_06800_), .Y(_25175_) );
  \$mux  #( .WIDTH(32) ) _46826_ ( .A(_25175_), .B(0), .S(RST), .Y(_02456_) );
  \$mux  #( .WIDTH(33) ) _46827_ ( .A(_source_stream_matmul_29_source_8_pat_size_buf_3), .B(_source_stream_matmul_29_source_8_pat_size_3), .S(_06800_), .Y(_25176_) );
  \$mux  #( .WIDTH(33) ) _46828_ ( .A(_25176_), .B(33'h000000000), .S(RST), .Y(_02451_) );
  \$mux  #( .WIDTH(33) ) _46829_ ( .A(_source_stream_matmul_29_source_8_pat_size_buf_2), .B(_source_stream_matmul_29_source_8_pat_size_2), .S(_06800_), .Y(_25177_) );
  \$mux  #( .WIDTH(33) ) _46830_ ( .A(_25177_), .B(33'h000000000), .S(RST), .Y(_02450_) );
  \$mux  #( .WIDTH(33) ) _46831_ ( .A(_source_stream_matmul_29_source_8_pat_size_buf_1), .B(_source_stream_matmul_29_source_8_pat_size_1), .S(_06800_), .Y(_25178_) );
  \$mux  #( .WIDTH(33) ) _46832_ ( .A(_25178_), .B(33'h000000000), .S(RST), .Y(_02449_) );
  \$mux  #( .WIDTH(33) ) _46833_ ( .A(_source_stream_matmul_29_source_8_pat_size_buf_0), .B(_source_stream_matmul_29_source_8_pat_size_0), .S(_06800_), .Y(_25179_) );
  \$mux  #( .WIDTH(33) ) _46834_ ( .A(_25179_), .B(33'h000000000), .S(RST), .Y(_02448_) );
  \$mux  #( .WIDTH(33) ) _46835_ ( .A(_source_stream_matmul_29_source_8_pat_count_3), .B(_28900_), .S(_06800_), .Y(_25180_) );
  \$mux  #( .WIDTH(33) ) _46836_ ( .A(_25180_), .B(_28907_), .S(_06803_), .Y(_25181_) );
  \$mux  #( .WIDTH(33) ) _46837_ ( .A(_25181_), .B(_28908_), .S(_06804_), .Y(_25182_) );
  \$mux  #( .WIDTH(33) ) _46838_ ( .A(_25182_), .B(33'h000000000), .S(RST), .Y(_02439_) );
  \$mux  #( .WIDTH(33) ) _46839_ ( .A(_source_stream_matmul_29_source_8_pat_count_2), .B(_28899_), .S(_06800_), .Y(_25183_) );
  \$mux  #( .WIDTH(33) ) _46840_ ( .A(_25183_), .B(_28905_), .S(_06802_), .Y(_25184_) );
  \$mux  #( .WIDTH(33) ) _46841_ ( .A(_25184_), .B(_28906_), .S(_06803_), .Y(_25185_) );
  \$mux  #( .WIDTH(33) ) _46842_ ( .A(_25185_), .B(33'h000000000), .S(RST), .Y(_02438_) );
  \$mux  #( .WIDTH(33) ) _46843_ ( .A(_source_stream_matmul_29_source_8_pat_count_1), .B(_28898_), .S(_06800_), .Y(_25186_) );
  \$mux  #( .WIDTH(33) ) _46844_ ( .A(_25186_), .B(_28903_), .S(_06801_), .Y(_25187_) );
  \$mux  #( .WIDTH(33) ) _46845_ ( .A(_25187_), .B(_28904_), .S(_06802_), .Y(_25188_) );
  \$mux  #( .WIDTH(33) ) _46846_ ( .A(_25188_), .B(33'h000000000), .S(RST), .Y(_02437_) );
  \$mux  #( .WIDTH(33) ) _46847_ ( .A(_source_stream_matmul_29_source_8_pat_count_0), .B(_28897_), .S(_06800_), .Y(_25189_) );
  \$mux  #( .WIDTH(33) ) _46848_ ( .A(_28901_), .B(_25189_), .S(_05911_), .Y(_25190_) );
  \$mux  #( .WIDTH(33) ) _46849_ ( .A(_25190_), .B(_28902_), .S(_06801_), .Y(_25191_) );
  \$mux  #( .WIDTH(33) ) _46850_ ( .A(_25191_), .B(33'h000000000), .S(RST), .Y(_02436_) );
  \$mux  #( .WIDTH(32) ) _46851_ ( .A(_source_stream_matmul_29_source_8_pat_stride_3), .B(0), .S(_set_flag_1224), .Y(_25192_) );
  \$mux  #( .WIDTH(32) ) _46852_ ( .A(_25192_), .B(0), .S(RST), .Y(_02455_) );
  \$mux  #( .WIDTH(32) ) _46853_ ( .A(_source_stream_matmul_29_source_8_pat_stride_2), .B(0), .S(_set_flag_1224), .Y(_25193_) );
  \$mux  #( .WIDTH(32) ) _46854_ ( .A(_25193_), .B(0), .S(RST), .Y(_02454_) );
  \$mux  #( .WIDTH(32) ) _46855_ ( .A(_source_stream_matmul_29_source_8_pat_stride_1), .B(0), .S(_set_flag_1224), .Y(_25194_) );
  \$mux  #( .WIDTH(32) ) _46856_ ( .A(_25194_), .B(0), .S(RST), .Y(_02453_) );
  \$mux  #( .WIDTH(32) ) _46857_ ( .A(_source_stream_matmul_29_source_8_pat_stride_0), .B(0), .S(_set_flag_1224), .Y(_25195_) );
  \$mux  #( .WIDTH(32) ) _46858_ ( .A(_25195_), .B(0), .S(RST), .Y(_02452_) );
  \$mux  #( .WIDTH(33) ) _46859_ ( .A(_source_stream_matmul_29_source_8_pat_size_3), .B(33'h000000001), .S(_set_flag_1224), .Y(_25196_) );
  \$mux  #( .WIDTH(33) ) _46860_ ( .A(_25196_), .B(33'h000000000), .S(RST), .Y(_02447_) );
  \$mux  #( .WIDTH(33) ) _46861_ ( .A(_source_stream_matmul_29_source_8_pat_size_2), .B(33'h000000001), .S(_set_flag_1224), .Y(_25197_) );
  \$mux  #( .WIDTH(33) ) _46862_ ( .A(_25197_), .B(33'h000000000), .S(RST), .Y(_02446_) );
  \$mux  #( .WIDTH(33) ) _46863_ ( .A(_source_stream_matmul_29_source_8_pat_size_1), .B({ 1'h0, matmul_29_next_stream_num_ops }), .S(_set_flag_1224), .Y(_25198_) );
  \$mux  #( .WIDTH(33) ) _46864_ ( .A(_25198_), .B(33'h000000000), .S(RST), .Y(_02445_) );
  \$mux  #( .WIDTH(33) ) _46865_ ( .A(_source_stream_matmul_29_source_8_pat_size_0), .B({ 22'h000000, cparam_matmul_29_act_bat_step }), .S(_set_flag_1224), .Y(_25199_) );
  \$mux  #( .WIDTH(33) ) _46866_ ( .A(_25199_), .B(33'h000000000), .S(RST), .Y(_02444_) );
  \$mux  #( .WIDTH(32) ) _46867_ ( .A(_source_stream_matmul_29_source_8_pat_cur_offset_3), .B(0), .S(_06800_), .Y(_25200_) );
  \$mux  #( .WIDTH(32) ) _46868_ ( .A(_25200_), .B(_24418_), .S(_06803_), .Y(_25201_) );
  \$mux  #( .WIDTH(32) ) _46869_ ( .A(_25201_), .B(0), .S(_06804_), .Y(_25202_) );
  \$mux  #( .WIDTH(32) ) _46870_ ( .A(_25202_), .B(0), .S(RST), .Y(_02443_) );
  \$mux  #( .WIDTH(32) ) _46871_ ( .A(_source_stream_matmul_29_source_8_pat_cur_offset_2), .B(0), .S(_06800_), .Y(_25203_) );
  \$mux  #( .WIDTH(32) ) _46872_ ( .A(_25203_), .B(_24417_), .S(_06802_), .Y(_25204_) );
  \$mux  #( .WIDTH(32) ) _46873_ ( .A(_25204_), .B(0), .S(_06803_), .Y(_25205_) );
  \$mux  #( .WIDTH(32) ) _46874_ ( .A(_25205_), .B(0), .S(RST), .Y(_02442_) );
  \$mux  #( .WIDTH(32) ) _46875_ ( .A(_source_stream_matmul_29_source_8_pat_cur_offset_1), .B(0), .S(_06800_), .Y(_25206_) );
  \$mux  #( .WIDTH(32) ) _46876_ ( .A(_25206_), .B(_24416_), .S(_06801_), .Y(_25207_) );
  \$mux  #( .WIDTH(32) ) _46877_ ( .A(_25207_), .B(0), .S(_06802_), .Y(_25208_) );
  \$mux  #( .WIDTH(32) ) _46878_ ( .A(_25208_), .B(0), .S(RST), .Y(_02441_) );
  \$mux  #( .WIDTH(32) ) _46879_ ( .A(_source_stream_matmul_29_source_8_pat_cur_offset_0), .B(0), .S(_06800_), .Y(_25209_) );
  \$mux  #( .WIDTH(32) ) _46880_ ( .A(_24415_), .B(_25209_), .S(_05911_), .Y(_25210_) );
  \$mux  #( .WIDTH(32) ) _46881_ ( .A(_25210_), .B(0), .S(_06801_), .Y(_25211_) );
  \$mux  #( .WIDTH(32) ) _46882_ ( .A(_25211_), .B(0), .S(RST), .Y(_02440_) );
  \$mux  #( .WIDTH(8) ) _46883_ ( .A(__variable_wdata_812), .B(_stream_matmul_29_source_6_source_ram_rdata), .S(_stream_matmul_29_source_6_source_ram_rvalid), .Y(_25212_) );
  \$mux  #( .WIDTH(8) ) _46884_ ( .A(_25212_), .B(8'h00), .S(RST), .Y(_01452_) );
  \$mux  #( .WIDTH(32) ) _46885_ ( .A(_source_stream_matmul_29_source_6_pat_stride_buf_3), .B(_source_stream_matmul_29_source_6_pat_stride_3), .S(_06795_), .Y(_25213_) );
  \$mux  #( .WIDTH(32) ) _46886_ ( .A(_25213_), .B(0), .S(RST), .Y(_02435_) );
  \$mux  #( .WIDTH(32) ) _46887_ ( .A(_source_stream_matmul_29_source_6_pat_stride_buf_2), .B(_source_stream_matmul_29_source_6_pat_stride_2), .S(_06795_), .Y(_25214_) );
  \$mux  #( .WIDTH(32) ) _46888_ ( .A(_25214_), .B(0), .S(RST), .Y(_02434_) );
  \$mux  #( .WIDTH(32) ) _46889_ ( .A(_source_stream_matmul_29_source_6_pat_stride_buf_1), .B(_source_stream_matmul_29_source_6_pat_stride_1), .S(_06795_), .Y(_25215_) );
  \$mux  #( .WIDTH(32) ) _46890_ ( .A(_25215_), .B(0), .S(RST), .Y(_02433_) );
  \$mux  #( .WIDTH(32) ) _46891_ ( .A(_source_stream_matmul_29_source_6_pat_stride_buf_0), .B(_source_stream_matmul_29_source_6_pat_stride_0), .S(_06795_), .Y(_25216_) );
  \$mux  #( .WIDTH(32) ) _46892_ ( .A(_25216_), .B(0), .S(RST), .Y(_02432_) );
  \$mux  #( .WIDTH(33) ) _46893_ ( .A(_source_stream_matmul_29_source_6_pat_size_buf_3), .B(_source_stream_matmul_29_source_6_pat_size_3), .S(_06795_), .Y(_25217_) );
  \$mux  #( .WIDTH(33) ) _46894_ ( .A(_25217_), .B(33'h000000000), .S(RST), .Y(_02427_) );
  \$mux  #( .WIDTH(33) ) _46895_ ( .A(_source_stream_matmul_29_source_6_pat_size_buf_2), .B(_source_stream_matmul_29_source_6_pat_size_2), .S(_06795_), .Y(_25218_) );
  \$mux  #( .WIDTH(33) ) _46896_ ( .A(_25218_), .B(33'h000000000), .S(RST), .Y(_02426_) );
  \$mux  #( .WIDTH(33) ) _46897_ ( .A(_source_stream_matmul_29_source_6_pat_size_buf_1), .B(_source_stream_matmul_29_source_6_pat_size_1), .S(_06795_), .Y(_25219_) );
  \$mux  #( .WIDTH(33) ) _46898_ ( .A(_25219_), .B(33'h000000000), .S(RST), .Y(_02425_) );
  \$mux  #( .WIDTH(33) ) _46899_ ( .A(_source_stream_matmul_29_source_6_pat_size_buf_0), .B(_source_stream_matmul_29_source_6_pat_size_0), .S(_06795_), .Y(_25220_) );
  \$mux  #( .WIDTH(33) ) _46900_ ( .A(_25220_), .B(33'h000000000), .S(RST), .Y(_02424_) );
  \$mux  #( .WIDTH(33) ) _46901_ ( .A(_source_stream_matmul_29_source_6_pat_count_3), .B(_28888_), .S(_06795_), .Y(_25221_) );
  \$mux  #( .WIDTH(33) ) _46902_ ( .A(_25221_), .B(_28895_), .S(_06798_), .Y(_25222_) );
  \$mux  #( .WIDTH(33) ) _46903_ ( .A(_25222_), .B(_28896_), .S(_06799_), .Y(_25223_) );
  \$mux  #( .WIDTH(33) ) _46904_ ( .A(_25223_), .B(33'h000000000), .S(RST), .Y(_02415_) );
  \$mux  #( .WIDTH(33) ) _46905_ ( .A(_source_stream_matmul_29_source_6_pat_count_2), .B(_28887_), .S(_06795_), .Y(_25224_) );
  \$mux  #( .WIDTH(33) ) _46906_ ( .A(_25224_), .B(_28893_), .S(_06797_), .Y(_25225_) );
  \$mux  #( .WIDTH(33) ) _46907_ ( .A(_25225_), .B(_28894_), .S(_06798_), .Y(_25226_) );
  \$mux  #( .WIDTH(33) ) _46908_ ( .A(_25226_), .B(33'h000000000), .S(RST), .Y(_02414_) );
  \$mux  #( .WIDTH(33) ) _46909_ ( .A(_source_stream_matmul_29_source_6_pat_count_1), .B(_28886_), .S(_06795_), .Y(_25227_) );
  \$mux  #( .WIDTH(33) ) _46910_ ( .A(_25227_), .B(_28891_), .S(_06796_), .Y(_25228_) );
  \$mux  #( .WIDTH(33) ) _46911_ ( .A(_25228_), .B(_28892_), .S(_06797_), .Y(_25229_) );
  \$mux  #( .WIDTH(33) ) _46912_ ( .A(_25229_), .B(33'h000000000), .S(RST), .Y(_02413_) );
  \$mux  #( .WIDTH(33) ) _46913_ ( .A(_source_stream_matmul_29_source_6_pat_count_0), .B(_28885_), .S(_06795_), .Y(_25230_) );
  \$mux  #( .WIDTH(33) ) _46914_ ( .A(_28889_), .B(_25230_), .S(_05912_), .Y(_25231_) );
  \$mux  #( .WIDTH(33) ) _46915_ ( .A(_25231_), .B(_28890_), .S(_06796_), .Y(_25232_) );
  \$mux  #( .WIDTH(33) ) _46916_ ( .A(_25232_), .B(33'h000000000), .S(RST), .Y(_02412_) );
  \$mux  #( .WIDTH(32) ) _46917_ ( .A(_source_stream_matmul_29_source_6_pat_stride_3), .B(0), .S(_set_flag_1224), .Y(_25233_) );
  \$mux  #( .WIDTH(32) ) _46918_ ( .A(_25233_), .B(0), .S(RST), .Y(_02431_) );
  \$mux  #( .WIDTH(32) ) _46919_ ( .A(_source_stream_matmul_29_source_6_pat_stride_2), .B(0), .S(_set_flag_1224), .Y(_25234_) );
  \$mux  #( .WIDTH(32) ) _46920_ ( .A(_25234_), .B(0), .S(RST), .Y(_02430_) );
  \$mux  #( .WIDTH(32) ) _46921_ ( .A(_source_stream_matmul_29_source_6_pat_stride_1), .B(_29294_), .S(_set_flag_1224), .Y(_25235_) );
  \$mux  #( .WIDTH(32) ) _46922_ ( .A(_25235_), .B(0), .S(RST), .Y(_02429_) );
  \$mux  #( .WIDTH(32) ) _46923_ ( .A(_source_stream_matmul_29_source_6_pat_stride_0), .B(0), .S(_set_flag_1224), .Y(_25236_) );
  \$mux  #( .WIDTH(32) ) _46924_ ( .A(_25236_), .B(0), .S(RST), .Y(_02428_) );
  \$mux  #( .WIDTH(33) ) _46925_ ( .A(_source_stream_matmul_29_source_6_pat_size_3), .B(33'h000000001), .S(_set_flag_1224), .Y(_25237_) );
  \$mux  #( .WIDTH(33) ) _46926_ ( .A(_25237_), .B(33'h000000000), .S(RST), .Y(_02423_) );
  \$mux  #( .WIDTH(33) ) _46927_ ( .A(_source_stream_matmul_29_source_6_pat_size_2), .B(33'h000000001), .S(_set_flag_1224), .Y(_25238_) );
  \$mux  #( .WIDTH(33) ) _46928_ ( .A(_25238_), .B(33'h000000000), .S(RST), .Y(_02422_) );
  \$mux  #( .WIDTH(33) ) _46929_ ( .A(_source_stream_matmul_29_source_6_pat_size_1), .B({ 1'h0, matmul_29_next_stream_num_ops }), .S(_set_flag_1224), .Y(_25239_) );
  \$mux  #( .WIDTH(33) ) _46930_ ( .A(_25239_), .B(33'h000000000), .S(RST), .Y(_02421_) );
  \$mux  #( .WIDTH(33) ) _46931_ ( .A(_source_stream_matmul_29_source_6_pat_size_0), .B({ 22'h000000, cparam_matmul_29_act_bat_step }), .S(_set_flag_1224), .Y(_25240_) );
  \$mux  #( .WIDTH(33) ) _46932_ ( .A(_25240_), .B(33'h000000000), .S(RST), .Y(_02420_) );
  \$mux  #( .WIDTH(32) ) _46933_ ( .A(_source_stream_matmul_29_source_6_pat_cur_offset_3), .B(0), .S(_06795_), .Y(_25241_) );
  \$mux  #( .WIDTH(32) ) _46934_ ( .A(_25241_), .B(_24414_), .S(_06798_), .Y(_25242_) );
  \$mux  #( .WIDTH(32) ) _46935_ ( .A(_25242_), .B(0), .S(_06799_), .Y(_25243_) );
  \$mux  #( .WIDTH(32) ) _46936_ ( .A(_25243_), .B(0), .S(RST), .Y(_02419_) );
  \$mux  #( .WIDTH(32) ) _46937_ ( .A(_source_stream_matmul_29_source_6_pat_cur_offset_2), .B(0), .S(_06795_), .Y(_25244_) );
  \$mux  #( .WIDTH(32) ) _46938_ ( .A(_25244_), .B(_24413_), .S(_06797_), .Y(_25245_) );
  \$mux  #( .WIDTH(32) ) _46939_ ( .A(_25245_), .B(0), .S(_06798_), .Y(_25246_) );
  \$mux  #( .WIDTH(32) ) _46940_ ( .A(_25246_), .B(0), .S(RST), .Y(_02418_) );
  \$mux  #( .WIDTH(32) ) _46941_ ( .A(_source_stream_matmul_29_source_6_pat_cur_offset_1), .B(0), .S(_06795_), .Y(_25247_) );
  \$mux  #( .WIDTH(32) ) _46942_ ( .A(_25247_), .B(_24412_), .S(_06796_), .Y(_25248_) );
  \$mux  #( .WIDTH(32) ) _46943_ ( .A(_25248_), .B(0), .S(_06797_), .Y(_25249_) );
  \$mux  #( .WIDTH(32) ) _46944_ ( .A(_25249_), .B(0), .S(RST), .Y(_02417_) );
  \$mux  #( .WIDTH(32) ) _46945_ ( .A(_source_stream_matmul_29_source_6_pat_cur_offset_0), .B(0), .S(_06795_), .Y(_25250_) );
  \$mux  #( .WIDTH(32) ) _46946_ ( .A(_24411_), .B(_25250_), .S(_05912_), .Y(_25251_) );
  \$mux  #( .WIDTH(32) ) _46947_ ( .A(_25251_), .B(0), .S(_06796_), .Y(_25252_) );
  \$mux  #( .WIDTH(32) ) _46948_ ( .A(_25252_), .B(0), .S(RST), .Y(_02416_) );
  \$mux  #( .WIDTH(1) ) _46949_ ( .A(__variable_wdata_799), .B(_stream_matmul_29_constant_3_next_constant_data), .S(_stream_matmul_29_start), .Y(_25253_) );
  \$mux  #( .WIDTH(1) ) _46950_ ( .A(_25253_), .B(1'h0), .S(RST), .Y(_01451_) );
  \$mux  #( .WIDTH(1) ) _46951_ ( .A(__variable_wdata_798), .B(_stream_matmul_29_constant_2_next_constant_data), .S(_stream_matmul_29_start), .Y(_25254_) );
  \$mux  #( .WIDTH(1) ) _46952_ ( .A(_25254_), .B(1'h0), .S(RST), .Y(_01450_) );
  \$mux  #( .WIDTH(1) ) _46953_ ( .A(__variable_wdata_797), .B(_stream_matmul_29_constant_1_next_constant_data), .S(_stream_matmul_29_start), .Y(_25255_) );
  \$mux  #( .WIDTH(1) ) _46954_ ( .A(_25255_), .B(1'h0), .S(RST), .Y(_01449_) );
  \$mux  #( .WIDTH(11) ) _46955_ ( .A(__variable_wdata_796), .B(_stream_matmul_29_constant_0_next_constant_data), .S(_stream_matmul_29_start), .Y(_25256_) );
  \$mux  #( .WIDTH(11) ) _46956_ ( .A(_25256_), .B(11'h000), .S(RST), .Y(_01448_) );
  \$mux  #( .WIDTH(1) ) _46957_ ( .A(1'h1), .B(1'h0), .S(_05917_), .Y(_25081_) );
  \$mux  #( .WIDTH(1) ) _46958_ ( .A(_25081_), .B(1'h0), .S(RST), .Y(_01872_) );
  \$mux  #( .WIDTH(1) ) _46959_ ( .A(__delay_data_1615), .B(1'h0), .S(RST), .Y(_00483_) );
  \$mux  #( .WIDTH(8) ) _46960_ ( .A(_29292_), .B(8'h00), .S(RST), .Y(_01559_) );
  \$mux  #( .WIDTH(1) ) _46961_ ( .A(__delay_data_1614), .B(1'h0), .S(RST), .Y(_00482_) );
  \$mux  #( .WIDTH(8) ) _46962_ ( .A(__delay_data_1564), .B(8'h00), .S(RST), .Y(_00481_) );
  \$mux  #( .WIDTH(1) ) _46963_ ( .A(__delay_data_1599), .B(1'h0), .S(RST), .Y(_00480_) );
  \$mux  #( .WIDTH(8) ) _46964_ ( .A(_29291_), .B(8'h00), .S(RST), .Y(_01558_) );
  \$mux  #( .WIDTH(1) ) _46965_ ( .A(__delay_data_1598), .B(1'h0), .S(RST), .Y(_00479_) );
  \$mux  #( .WIDTH(8) ) _46966_ ( .A(__delay_data_1528), .B(8'h00), .S(RST), .Y(_00444_) );
  \$mux  #( .WIDTH(1) ) _46967_ ( .A(__delay_data_1562), .B(1'h0), .S(RST), .Y(_00443_) );
  \$mux  #( .WIDTH(1) ) _46968_ ( .A(__delay_data_1597), .B(1'h0), .S(RST), .Y(_00478_) );
  \$mux  #( .WIDTH(1) ) _46969_ ( .A(__delay_data_1561), .B(1'h0), .S(RST), .Y(_00442_) );
  \$mux  #( .WIDTH(1) ) _46970_ ( .A(__delay_data_1596), .B(1'h0), .S(RST), .Y(_00477_) );
  \$mux  #( .WIDTH(1) ) _46971_ ( .A(__delay_data_1560), .B(1'h0), .S(RST), .Y(_00441_) );
  \$mux  #( .WIDTH(1) ) _46972_ ( .A(__delay_data_1595), .B(1'h0), .S(RST), .Y(_00476_) );
  \$mux  #( .WIDTH(1) ) _46973_ ( .A(__delay_data_1559), .B(1'h0), .S(RST), .Y(_00440_) );
  \$mux  #( .WIDTH(1) ) _46974_ ( .A(__delay_data_1594), .B(1'h0), .S(RST), .Y(_00475_) );
  \$mux  #( .WIDTH(1) ) _46975_ ( .A(__delay_data_1558), .B(1'h0), .S(RST), .Y(_00439_) );
  \$mux  #( .WIDTH(1) ) _46976_ ( .A(__delay_data_1593), .B(1'h0), .S(RST), .Y(_00474_) );
  \$mux  #( .WIDTH(1) ) _46977_ ( .A(__delay_data_1557), .B(1'h0), .S(RST), .Y(_00438_) );
  \$mux  #( .WIDTH(1) ) _46978_ ( .A(__delay_data_1592), .B(1'h0), .S(RST), .Y(_00473_) );
  \$mux  #( .WIDTH(1) ) _46979_ ( .A(__delay_data_1556), .B(1'h0), .S(RST), .Y(_00437_) );
  \$mux  #( .WIDTH(1) ) _46980_ ( .A(__delay_data_1591), .B(1'h0), .S(RST), .Y(_00472_) );
  \$mux  #( .WIDTH(1) ) _46981_ ( .A(__delay_data_1555), .B(1'h0), .S(RST), .Y(_00436_) );
  \$mux  #( .WIDTH(1) ) _46982_ ( .A(__delay_data_1590), .B(1'h0), .S(RST), .Y(_00471_) );
  \$mux  #( .WIDTH(1) ) _46983_ ( .A(__delay_data_1554), .B(1'h0), .S(RST), .Y(_00435_) );
  \$mux  #( .WIDTH(1) ) _46984_ ( .A(__delay_data_1589), .B(1'h0), .S(RST), .Y(_00470_) );
  \$mux  #( .WIDTH(1) ) _46985_ ( .A(__delay_data_1553), .B(1'h0), .S(RST), .Y(_00434_) );
  \$mux  #( .WIDTH(1) ) _46986_ ( .A(__delay_data_1588), .B(1'h0), .S(RST), .Y(_00469_) );
  \$mux  #( .WIDTH(1) ) _46987_ ( .A(__delay_data_1552), .B(1'h0), .S(RST), .Y(_00433_) );
  \$mux  #( .WIDTH(1) ) _46988_ ( .A(__delay_data_1587), .B(1'h0), .S(RST), .Y(_00468_) );
  \$mux  #( .WIDTH(1) ) _46989_ ( .A(__delay_data_1551), .B(1'h0), .S(RST), .Y(_00432_) );
  \$mux  #( .WIDTH(1) ) _46990_ ( .A(__delay_data_1586), .B(1'h0), .S(RST), .Y(_00467_) );
  \$mux  #( .WIDTH(1) ) _46991_ ( .A(__delay_data_1550), .B(1'h0), .S(RST), .Y(_00431_) );
  \$mux  #( .WIDTH(8) ) _46992_ ( .A(__delay_data_1526), .B(8'h00), .S(RST), .Y(_00408_) );
  \$mux  #( .WIDTH(8) ) _46993_ ( .A(__delay_data_1504), .B(8'h00), .S(RST), .Y(_00386_) );
  \$mux  #( .WIDTH(32) ) _46994_ ( .A(_24410_), .B(0), .S(RST), .Y(_01817_) );
  \$mux  #( .WIDTH(1) ) _46995_ ( .A(__delay_data_1585), .B(1'h0), .S(RST), .Y(_00466_) );
  \$mux  #( .WIDTH(1) ) _46996_ ( .A(__delay_data_1549), .B(1'h0), .S(RST), .Y(_00430_) );
  \$mux  #( .WIDTH(8) ) _46997_ ( .A(__delay_data_1525), .B(8'h00), .S(RST), .Y(_00407_) );
  \$mux  #( .WIDTH(8) ) _46998_ ( .A(__delay_data_1503), .B(8'h00), .S(RST), .Y(_00385_) );
  \$mux  #( .WIDTH(8) ) _46999_ ( .A(__delay_data_1480), .B(8'h00), .S(RST), .Y(_00362_) );
  \$mux  #( .WIDTH(1) ) _47000_ ( .A(__delay_data_1584), .B(1'h0), .S(RST), .Y(_00465_) );
  \$mux  #( .WIDTH(1) ) _47001_ ( .A(__delay_data_1548), .B(1'h0), .S(RST), .Y(_00429_) );
  \$mux  #( .WIDTH(8) ) _47002_ ( .A(__delay_data_1524), .B(8'h00), .S(RST), .Y(_00406_) );
  \$mux  #( .WIDTH(8) ) _47003_ ( .A(__delay_data_1502), .B(8'h00), .S(RST), .Y(_00384_) );
  \$mux  #( .WIDTH(8) ) _47004_ ( .A(__delay_data_1479), .B(8'h00), .S(RST), .Y(_00361_) );
  \$mux  #( .WIDTH(1) ) _47005_ ( .A(__delay_data_1583), .B(1'h0), .S(RST), .Y(_00464_) );
  \$mux  #( .WIDTH(1) ) _47006_ ( .A(__delay_data_1547), .B(1'h0), .S(RST), .Y(_00428_) );
  \$mux  #( .WIDTH(8) ) _47007_ ( .A(__delay_data_1523), .B(8'h00), .S(RST), .Y(_00405_) );
  \$mux  #( .WIDTH(8) ) _47008_ ( .A(__delay_data_1501), .B(8'h00), .S(RST), .Y(_00383_) );
  \$mux  #( .WIDTH(8) ) _47009_ ( .A(__delay_data_1478), .B(8'h00), .S(RST), .Y(_00360_) );
  \$mux  #( .WIDTH(1) ) _47010_ ( .A(__delay_data_1582), .B(1'h0), .S(RST), .Y(_00463_) );
  \$mux  #( .WIDTH(1) ) _47011_ ( .A(__delay_data_1546), .B(1'h0), .S(RST), .Y(_00427_) );
  \$mux  #( .WIDTH(8) ) _47012_ ( .A(__delay_data_1522), .B(8'h00), .S(RST), .Y(_00404_) );
  \$mux  #( .WIDTH(8) ) _47013_ ( .A(__delay_data_1500), .B(8'h00), .S(RST), .Y(_00382_) );
  \$mux  #( .WIDTH(8) ) _47014_ ( .A(__delay_data_1477), .B(8'h00), .S(RST), .Y(_00359_) );
  \$mux  #( .WIDTH(1) ) _47015_ ( .A(__delay_data_1581), .B(1'h0), .S(RST), .Y(_00462_) );
  \$mux  #( .WIDTH(1) ) _47016_ ( .A(__delay_data_1545), .B(1'h0), .S(RST), .Y(_00426_) );
  \$mux  #( .WIDTH(8) ) _47017_ ( .A(__delay_data_1521), .B(8'h00), .S(RST), .Y(_00403_) );
  \$mux  #( .WIDTH(8) ) _47018_ ( .A(__delay_data_1499), .B(8'h00), .S(RST), .Y(_00381_) );
  \$mux  #( .WIDTH(8) ) _47019_ ( .A(__delay_data_1476), .B(8'h00), .S(RST), .Y(_00358_) );
  \$mux  #( .WIDTH(1) ) _47020_ ( .A(__delay_data_1580), .B(1'h0), .S(RST), .Y(_00461_) );
  \$mux  #( .WIDTH(1) ) _47021_ ( .A(__delay_data_1544), .B(1'h0), .S(RST), .Y(_00425_) );
  \$mux  #( .WIDTH(8) ) _47022_ ( .A(__delay_data_1520), .B(8'h00), .S(RST), .Y(_00402_) );
  \$mux  #( .WIDTH(8) ) _47023_ ( .A(__delay_data_1498), .B(8'h00), .S(RST), .Y(_00380_) );
  \$mux  #( .WIDTH(8) ) _47024_ ( .A(__delay_data_1475), .B(8'h00), .S(RST), .Y(_00357_) );
  \$mux  #( .WIDTH(1) ) _47025_ ( .A(__delay_data_1579), .B(1'h0), .S(RST), .Y(_00460_) );
  \$mux  #( .WIDTH(1) ) _47026_ ( .A(__delay_data_1543), .B(1'h0), .S(RST), .Y(_00424_) );
  \$mux  #( .WIDTH(8) ) _47027_ ( .A(__delay_data_1519), .B(8'h00), .S(RST), .Y(_00401_) );
  \$mux  #( .WIDTH(8) ) _47028_ ( .A(__delay_data_1497), .B(8'h00), .S(RST), .Y(_00379_) );
  \$mux  #( .WIDTH(8) ) _47029_ ( .A(__delay_data_1474), .B(8'h00), .S(RST), .Y(_00356_) );
  \$mux  #( .WIDTH(1) ) _47030_ ( .A(__delay_data_1578), .B(1'h0), .S(RST), .Y(_00459_) );
  \$mux  #( .WIDTH(1) ) _47031_ ( .A(__delay_data_1542), .B(1'h0), .S(RST), .Y(_00423_) );
  \$mux  #( .WIDTH(8) ) _47032_ ( .A(__delay_data_1518), .B(8'h00), .S(RST), .Y(_00400_) );
  \$mux  #( .WIDTH(8) ) _47033_ ( .A(__delay_data_1496), .B(8'h00), .S(RST), .Y(_00378_) );
  \$mux  #( .WIDTH(8) ) _47034_ ( .A(__delay_data_1473), .B(8'h00), .S(RST), .Y(_00355_) );
  \$mux  #( .WIDTH(11) ) _47035_ ( .A(__delay_data_1458), .B(11'h000), .S(RST), .Y(_00340_) );
  \$mux  #( .WIDTH(8) ) _47036_ ( .A(__delay_data_1442), .B(8'h00), .S(RST), .Y(_00324_) );
  \$mux  #( .WIDTH(32) ) _47037_ ( .A(__variable_wdata_22), .B(0), .S(RST), .Y(_01104_) );
  \$mux  #( .WIDTH(1) ) _47038_ ( .A(__delay_data_1577), .B(1'h0), .S(RST), .Y(_00458_) );
  \$mux  #( .WIDTH(1) ) _47039_ ( .A(__delay_data_1541), .B(1'h0), .S(RST), .Y(_00422_) );
  \$mux  #( .WIDTH(8) ) _47040_ ( .A(__delay_data_1517), .B(8'h00), .S(RST), .Y(_00399_) );
  \$mux  #( .WIDTH(8) ) _47041_ ( .A(__delay_data_1495), .B(8'h00), .S(RST), .Y(_00377_) );
  \$mux  #( .WIDTH(8) ) _47042_ ( .A(__delay_data_1472), .B(8'h00), .S(RST), .Y(_00354_) );
  \$mux  #( .WIDTH(11) ) _47043_ ( .A(__delay_data_1457), .B(11'h000), .S(RST), .Y(_00339_) );
  \$mux  #( .WIDTH(8) ) _47044_ ( .A(__delay_data_1441), .B(8'h00), .S(RST), .Y(_00323_) );
  \$mux  #( .WIDTH(1) ) _47045_ ( .A(__delay_data_1576), .B(1'h0), .S(RST), .Y(_00457_) );
  \$mux  #( .WIDTH(1) ) _47046_ ( .A(__delay_data_1540), .B(1'h0), .S(RST), .Y(_00421_) );
  \$mux  #( .WIDTH(8) ) _47047_ ( .A(__delay_data_1516), .B(8'h00), .S(RST), .Y(_00398_) );
  \$mux  #( .WIDTH(8) ) _47048_ ( .A(__delay_data_1494), .B(8'h00), .S(RST), .Y(_00376_) );
  \$mux  #( .WIDTH(8) ) _47049_ ( .A(__delay_data_1471), .B(8'h00), .S(RST), .Y(_00353_) );
  \$mux  #( .WIDTH(11) ) _47050_ ( .A(__delay_data_1456), .B(11'h000), .S(RST), .Y(_00338_) );
  \$mux  #( .WIDTH(8) ) _47051_ ( .A(__delay_data_1440), .B(8'h00), .S(RST), .Y(_00322_) );
  \$mux  #( .WIDTH(1) ) _47052_ ( .A(__delay_data_1575), .B(1'h0), .S(RST), .Y(_00456_) );
  \$mux  #( .WIDTH(1) ) _47053_ ( .A(__delay_data_1539), .B(1'h0), .S(RST), .Y(_00420_) );
  \$mux  #( .WIDTH(8) ) _47054_ ( .A(__delay_data_1515), .B(8'h00), .S(RST), .Y(_00397_) );
  \$mux  #( .WIDTH(8) ) _47055_ ( .A(__delay_data_1493), .B(8'h00), .S(RST), .Y(_00375_) );
  \$mux  #( .WIDTH(8) ) _47056_ ( .A(__delay_data_1470), .B(8'h00), .S(RST), .Y(_00352_) );
  \$mux  #( .WIDTH(11) ) _47057_ ( .A(__delay_data_1455), .B(11'h000), .S(RST), .Y(_00337_) );
  \$mux  #( .WIDTH(8) ) _47058_ ( .A(__delay_data_1439), .B(8'h00), .S(RST), .Y(_00321_) );
  \$mux  #( .WIDTH(1) ) _47059_ ( .A(__delay_data_1574), .B(1'h0), .S(RST), .Y(_00455_) );
  \$mux  #( .WIDTH(1) ) _47060_ ( .A(__delay_data_1538), .B(1'h0), .S(RST), .Y(_00419_) );
  \$mux  #( .WIDTH(8) ) _47061_ ( .A(__delay_data_1514), .B(8'h00), .S(RST), .Y(_00396_) );
  \$mux  #( .WIDTH(8) ) _47062_ ( .A(__delay_data_1492), .B(8'h00), .S(RST), .Y(_00374_) );
  \$mux  #( .WIDTH(8) ) _47063_ ( .A(__delay_data_1469), .B(8'h00), .S(RST), .Y(_00351_) );
  \$mux  #( .WIDTH(11) ) _47064_ ( .A(__delay_data_1454), .B(11'h000), .S(RST), .Y(_00336_) );
  \$mux  #( .WIDTH(8) ) _47065_ ( .A(__delay_data_1438), .B(8'h00), .S(RST), .Y(_00320_) );
  \$mux  #( .WIDTH(1) ) _47066_ ( .A(__delay_data_1573), .B(1'h0), .S(RST), .Y(_00454_) );
  \$mux  #( .WIDTH(1) ) _47067_ ( .A(__delay_data_1537), .B(1'h0), .S(RST), .Y(_00418_) );
  \$mux  #( .WIDTH(8) ) _47068_ ( .A(__delay_data_1513), .B(8'h00), .S(RST), .Y(_00395_) );
  \$mux  #( .WIDTH(8) ) _47069_ ( .A(__delay_data_1491), .B(8'h00), .S(RST), .Y(_00373_) );
  \$mux  #( .WIDTH(8) ) _47070_ ( .A(__delay_data_1468), .B(8'h00), .S(RST), .Y(_00350_) );
  \$mux  #( .WIDTH(11) ) _47071_ ( .A(__delay_data_1453), .B(11'h000), .S(RST), .Y(_00335_) );
  \$mux  #( .WIDTH(8) ) _47072_ ( .A(__delay_data_1437), .B(8'h00), .S(RST), .Y(_00319_) );
  \$mux  #( .WIDTH(1) ) _47073_ ( .A(__delay_data_1572), .B(1'h0), .S(RST), .Y(_00453_) );
  \$mux  #( .WIDTH(1) ) _47074_ ( .A(__delay_data_1536), .B(1'h0), .S(RST), .Y(_00417_) );
  \$mux  #( .WIDTH(8) ) _47075_ ( .A(__delay_data_1512), .B(8'h00), .S(RST), .Y(_00394_) );
  \$mux  #( .WIDTH(8) ) _47076_ ( .A(__delay_data_1490), .B(8'h00), .S(RST), .Y(_00372_) );
  \$mux  #( .WIDTH(8) ) _47077_ ( .A(__delay_data_1467), .B(8'h00), .S(RST), .Y(_00349_) );
  \$mux  #( .WIDTH(11) ) _47078_ ( .A(__delay_data_1452), .B(11'h000), .S(RST), .Y(_00334_) );
  \$mux  #( .WIDTH(8) ) _47079_ ( .A(__delay_data_1436), .B(8'h00), .S(RST), .Y(_00318_) );
  \$mux  #( .WIDTH(1) ) _47080_ ( .A(__delay_data_1571), .B(1'h0), .S(RST), .Y(_00452_) );
  \$mux  #( .WIDTH(1) ) _47081_ ( .A(__delay_data_1535), .B(1'h0), .S(RST), .Y(_00416_) );
  \$mux  #( .WIDTH(8) ) _47082_ ( .A(__delay_data_1511), .B(8'h00), .S(RST), .Y(_00393_) );
  \$mux  #( .WIDTH(8) ) _47083_ ( .A(__delay_data_1489), .B(8'h00), .S(RST), .Y(_00371_) );
  \$mux  #( .WIDTH(8) ) _47084_ ( .A(__delay_data_1466), .B(8'h00), .S(RST), .Y(_00348_) );
  \$mux  #( .WIDTH(11) ) _47085_ ( .A(__delay_data_1451), .B(11'h000), .S(RST), .Y(_00333_) );
  \$mux  #( .WIDTH(8) ) _47086_ ( .A(__delay_data_1435), .B(8'h00), .S(RST), .Y(_00317_) );
  \$mux  #( .WIDTH(1) ) _47087_ ( .A(__delay_data_1570), .B(1'h0), .S(RST), .Y(_00451_) );
  \$mux  #( .WIDTH(1) ) _47088_ ( .A(__delay_data_1534), .B(1'h0), .S(RST), .Y(_00415_) );
  \$mux  #( .WIDTH(8) ) _47089_ ( .A(__delay_data_1510), .B(8'h00), .S(RST), .Y(_00392_) );
  \$mux  #( .WIDTH(8) ) _47090_ ( .A(__delay_data_1488), .B(8'h00), .S(RST), .Y(_00370_) );
  \$mux  #( .WIDTH(8) ) _47091_ ( .A(__delay_data_1465), .B(8'h00), .S(RST), .Y(_00347_) );
  \$mux  #( .WIDTH(11) ) _47092_ ( .A(__delay_data_1450), .B(11'h000), .S(RST), .Y(_00332_) );
  \$mux  #( .WIDTH(8) ) _47093_ ( .A(__delay_data_1434), .B(8'h00), .S(RST), .Y(_00316_) );
  \$mux  #( .WIDTH(1) ) _47094_ ( .A(__delay_data_1569), .B(1'h0), .S(RST), .Y(_00450_) );
  \$mux  #( .WIDTH(1) ) _47095_ ( .A(__delay_data_1533), .B(1'h0), .S(RST), .Y(_00414_) );
  \$mux  #( .WIDTH(8) ) _47096_ ( .A(__delay_data_1509), .B(8'h00), .S(RST), .Y(_00391_) );
  \$mux  #( .WIDTH(8) ) _47097_ ( .A(__delay_data_1487), .B(8'h00), .S(RST), .Y(_00369_) );
  \$mux  #( .WIDTH(8) ) _47098_ ( .A(__delay_data_1464), .B(8'h00), .S(RST), .Y(_00346_) );
  \$mux  #( .WIDTH(11) ) _47099_ ( .A(__delay_data_1449), .B(11'h000), .S(RST), .Y(_00331_) );
  \$mux  #( .WIDTH(8) ) _47100_ ( .A(__delay_data_1433), .B(8'h00), .S(RST), .Y(_00315_) );
  \$mux  #( .WIDTH(1) ) _47101_ ( .A(__delay_data_1568), .B(1'h0), .S(RST), .Y(_00449_) );
  \$mux  #( .WIDTH(1) ) _47102_ ( .A(__delay_data_1532), .B(1'h0), .S(RST), .Y(_00413_) );
  \$mux  #( .WIDTH(8) ) _47103_ ( .A(__delay_data_1508), .B(8'h00), .S(RST), .Y(_00390_) );
  \$mux  #( .WIDTH(8) ) _47104_ ( .A(__delay_data_1486), .B(8'h00), .S(RST), .Y(_00368_) );
  \$mux  #( .WIDTH(8) ) _47105_ ( .A(__delay_data_1463), .B(8'h00), .S(RST), .Y(_00345_) );
  \$mux  #( .WIDTH(11) ) _47106_ ( .A(__delay_data_1448), .B(11'h000), .S(RST), .Y(_00330_) );
  \$mux  #( .WIDTH(8) ) _47107_ ( .A(__delay_data_1432), .B(8'h00), .S(RST), .Y(_00314_) );
  \$mux  #( .WIDTH(1) ) _47108_ ( .A(__delay_data_1567), .B(1'h0), .S(RST), .Y(_00448_) );
  \$mux  #( .WIDTH(1) ) _47109_ ( .A(__delay_data_1531), .B(1'h0), .S(RST), .Y(_00412_) );
  \$mux  #( .WIDTH(8) ) _47110_ ( .A(__delay_data_1507), .B(8'h00), .S(RST), .Y(_00389_) );
  \$mux  #( .WIDTH(8) ) _47111_ ( .A(__delay_data_1485), .B(8'h00), .S(RST), .Y(_00367_) );
  \$mux  #( .WIDTH(8) ) _47112_ ( .A(__delay_data_1462), .B(8'h00), .S(RST), .Y(_00344_) );
  \$mux  #( .WIDTH(11) ) _47113_ ( .A(__delay_data_1447), .B(11'h000), .S(RST), .Y(_00329_) );
  \$mux  #( .WIDTH(8) ) _47114_ ( .A(__delay_data_1431), .B(8'h00), .S(RST), .Y(_00313_) );
  \$mux  #( .WIDTH(1) ) _47115_ ( .A(__delay_data_1566), .B(1'h0), .S(RST), .Y(_00447_) );
  \$mux  #( .WIDTH(1) ) _47116_ ( .A(__delay_data_1530), .B(1'h0), .S(RST), .Y(_00411_) );
  \$mux  #( .WIDTH(8) ) _47117_ ( .A(__delay_data_1506), .B(8'h00), .S(RST), .Y(_00388_) );
  \$mux  #( .WIDTH(8) ) _47118_ ( .A(__delay_data_1484), .B(8'h00), .S(RST), .Y(_00366_) );
  \$mux  #( .WIDTH(8) ) _47119_ ( .A(__delay_data_1461), .B(8'h00), .S(RST), .Y(_00343_) );
  \$mux  #( .WIDTH(11) ) _47120_ ( .A(__delay_data_1446), .B(11'h000), .S(RST), .Y(_00328_) );
  \$mux  #( .WIDTH(8) ) _47121_ ( .A(__delay_data_1430), .B(8'h00), .S(RST), .Y(_00312_) );
  \$mux  #( .WIDTH(8) ) _47122_ ( .A(__delay_data_1427), .B(8'h00), .S(RST), .Y(_00309_) );
  \$mux  #( .WIDTH(4) ) _47123_ ( .A(__delay_data_1425), .B(4'h0), .S(RST), .Y(_00307_) );
  \$mux  #( .WIDTH(8) ) _47124_ ( .A(_29290_), .B(8'h00), .S(RST), .Y(_01557_) );
  \$mux  #( .WIDTH(1) ) _47125_ ( .A(__delay_data_1565), .B(1'h0), .S(RST), .Y(_00446_) );
  \$mux  #( .WIDTH(1) ) _47126_ ( .A(__delay_data_1529), .B(1'h0), .S(RST), .Y(_00410_) );
  \$mux  #( .WIDTH(8) ) _47127_ ( .A(_plus_data_885), .B(8'h00), .S(RST), .Y(_00387_) );
  \$mux  #( .WIDTH(8) ) _47128_ ( .A(__delay_data_1483), .B(8'h00), .S(RST), .Y(_00365_) );
  \$mux  #( .WIDTH(8) ) _47129_ ( .A(__delay_data_1460), .B(8'h00), .S(RST), .Y(_00342_) );
  \$mux  #( .WIDTH(11) ) _47130_ ( .A(__delay_data_1445), .B(11'h000), .S(RST), .Y(_00327_) );
  \$mux  #( .WIDTH(8) ) _47131_ ( .A(_plus_data_880), .B(8'h00), .S(RST), .Y(_00311_) );
  \$mux  #( .WIDTH(8) ) _47132_ ( .A(_plus_data_875), .B(8'h00), .S(RST), .Y(_00308_) );
  \$mux  #( .WIDTH(4) ) _47133_ ( .A(__delay_data_1424), .B(4'h0), .S(RST), .Y(_00306_) );
  \$mux  #( .WIDTH(1) ) _47134_ ( .A(__delay_data_1420), .B(1'h0), .S(RST), .Y(_00302_) );
  \$mux  #( .WIDTH(8) ) _47135_ ( .A(_29289_), .B(8'h00), .S(RST), .Y(_01556_) );
  \$mux  #( .WIDTH(1) ) _47136_ ( .A(_eq_data_894), .B(1'h0), .S(RST), .Y(_00445_) );
  \$mux  #( .WIDTH(1) ) _47137_ ( .A(_eq_data_891), .B(1'h0), .S(RST), .Y(_00409_) );
  \$mux  #( .WIDTH(8) ) _47138_ ( .A(_cond_data_824), .B(8'h00), .S(RST), .Y(_00364_) );
  \$mux  #( .WIDTH(8) ) _47139_ ( .A(_cond_data_817), .B(8'h00), .S(RST), .Y(_00341_) );
  \$mux  #( .WIDTH(11) ) _47140_ ( .A(__delay_data_1444), .B(11'h000), .S(RST), .Y(_00326_) );
  \$mux  #( .WIDTH(4) ) _47141_ ( .A(__delay_data_1423), .B(4'h0), .S(RST), .Y(_00305_) );
  \$mux  #( .WIDTH(1) ) _47142_ ( .A(__delay_data_1419), .B(1'h0), .S(RST), .Y(_00301_) );
  \$mux  #( .WIDTH(1) ) _47143_ ( .A(_eq_data_855), .B(1'h0), .S(RST), .Y(_00299_) );
  \$mux  #( .WIDTH(8) ) _47144_ ( .A(_24409_), .B(8'h00), .S(RST), .Y(_01818_) );
  \$mux  #( .WIDTH(8) ) _47145_ ( .A(_24408_), .B(8'h00), .S(RST), .Y(_01816_) );
  \$mux  #( .WIDTH(8) ) _47146_ ( .A(_24407_), .B(8'h00), .S(RST), .Y(_01815_) );
  \$mux  #( .WIDTH(8) ) _47147_ ( .A(_29288_), .B(8'h00), .S(RST), .Y(_01555_) );
  \$mux  #( .WIDTH(4) ) _47148_ ( .A(__variable_wdata_848), .B(4'h0), .S(RST), .Y(_00363_) );
  \$mux  #( .WIDTH(11) ) _47149_ ( .A(__variable_wdata_796), .B(11'h000), .S(RST), .Y(_00325_) );
  \$mux  #( .WIDTH(1) ) _47150_ ( .A(__variable_wdata_847), .B(1'h0), .S(RST), .Y(_00310_) );
  \$mux  #( .WIDTH(4) ) _47151_ ( .A(__variable_wdata_864), .B(4'h0), .S(RST), .Y(_00304_) );
  \$mux  #( .WIDTH(1) ) _47152_ ( .A(__variable_wdata_846), .B(1'h0), .S(RST), .Y(_00303_) );
  \$mux  #( .WIDTH(1) ) _47153_ ( .A(__variable_wdata_799), .B(1'h0), .S(RST), .Y(_00300_) );
  \$mux  #( .WIDTH(8) ) _47154_ ( .A(__variable_wdata_850), .B(8'h00), .S(RST), .Y(_00298_) );
  \$mux  #( .WIDTH(1) ) _47155_ ( .A(_06145_), .B(1'h0), .S(RST), .Y(_01689_) );
  \$mux  #( .WIDTH(1) ) _47156_ ( .A(_06144_), .B(1'h0), .S(RST), .Y(_01688_) );
  \$mux  #( .WIDTH(1) ) _47157_ ( .A(_06143_), .B(1'h0), .S(RST), .Y(_01687_) );
  \$mux  #( .WIDTH(1) ) _47158_ ( .A(_06142_), .B(1'h0), .S(RST), .Y(_01686_) );
  \$mux  #( .WIDTH(8) ) _47159_ ( .A(__variable_wdata_840), .B(8'h00), .S(RST), .Y(_01553_) );
  \$mux  #( .WIDTH(8) ) _47160_ ( .A(__variable_wdata_833), .B(8'h00), .S(RST), .Y(_01552_) );
  \$mux  #( .WIDTH(8) ) _47161_ ( .A(__variable_wdata_826), .B(8'h00), .S(RST), .Y(_01551_) );
  \$mux  #( .WIDTH(8) ) _47162_ ( .A(__variable_wdata_819), .B(8'h00), .S(RST), .Y(_01550_) );
  \$mux  #( .WIDTH(8) ) _47163_ ( .A(__variable_wdata_812), .B(8'h00), .S(RST), .Y(_01549_) );
  \$mux  #( .WIDTH(8) ) _47164_ ( .A(_stream_matmul_29_sink_21_sink_wdata), .B(_cond_data_896), .S(_06816_), .Y(_25257_) );
  \$mux  #( .WIDTH(8) ) _47165_ ( .A(_25257_), .B(8'h00), .S(RST), .Y(_02723_) );
  \$mux  #( .WIDTH(1) ) _47166_ ( .A(1'h0), .B(1'h1), .S(_06816_), .Y(_25258_) );
  \$mux  #( .WIDTH(1) ) _47167_ ( .A(_25258_), .B(1'h0), .S(RST), .Y(_02724_) );
  \$mux  #( .WIDTH(32) ) _47168_ ( .A(_stream_matmul_29_sink_21_sink_waddr), .B(_28933_), .S(_06815_), .Y(_25259_) );
  \$mux  #( .WIDTH(32) ) _47169_ ( .A(_25259_), .B(_24429_), .S(_06816_), .Y(_25260_) );
  \$mux  #( .WIDTH(32) ) _47170_ ( .A(_25260_), .B(0), .S(RST), .Y(_02722_) );
  \$mux  #( .WIDTH(8) ) _47171_ ( .A(_stream_matmul_29_sink_21_sink_ram_sel), .B(8'h05), .S(__set_flag_1224_41), .Y(_25261_) );
  \$mux  #( .WIDTH(8) ) _47172_ ( .A(_25261_), .B(8'h00), .S(RST), .Y(_02718_) );
  \$mux  #( .WIDTH(32) ) _47173_ ( .A(_stream_matmul_29_sink_21_sink_stride_buf), .B(_stream_matmul_29_sink_21_sink_stride), .S(_06815_), .Y(_25262_) );
  \$mux  #( .WIDTH(32) ) _47174_ ( .A(_25262_), .B(0), .S(RST), .Y(_02721_) );
  \$mux  #( .WIDTH(33) ) _47175_ ( .A(_stream_matmul_29_sink_21_sink_count), .B(_stream_matmul_29_sink_21_sink_size), .S(_06815_), .Y(_25263_) );
  \$mux  #( .WIDTH(33) ) _47176_ ( .A(_25263_), .B(_28934_), .S(_06816_), .Y(_25264_) );
  \$mux  #( .WIDTH(33) ) _47177_ ( .A(_25264_), .B(33'h000000000), .S(RST), .Y(_02714_) );
  \$mux  #( .WIDTH(32) ) _47178_ ( .A(_stream_matmul_29_sink_21_sink_stride), .B(1), .S(__set_flag_1224_41), .Y(_25265_) );
  \$mux  #( .WIDTH(32) ) _47179_ ( .A(_25265_), .B(0), .S(RST), .Y(_02720_) );
  \$mux  #( .WIDTH(33) ) _47180_ ( .A(_stream_matmul_29_sink_21_sink_size), .B(__stream_matmul_29_sink_21_sink_size_1_41), .S(__set_flag_1224_41), .Y(_25266_) );
  \$mux  #( .WIDTH(33) ) _47181_ ( .A(_25266_), .B(33'h000000000), .S(RST), .Y(_02719_) );
  \$mux  #( .WIDTH(32) ) _47182_ ( .A(_stream_matmul_29_sink_21_sink_offset), .B(__stream_matmul_29_sink_21_sink_offset_0_41), .S(__set_flag_1224_41), .Y(_25267_) );
  \$mux  #( .WIDTH(32) ) _47183_ ( .A(_25267_), .B(0), .S(RST), .Y(_02717_) );
  \$mux  #( .WIDTH(3) ) _47184_ ( .A(_stream_matmul_29_sink_21_sink_mode), .B(3'h1), .S(__set_flag_1224_41), .Y(_25268_) );
  \$mux  #( .WIDTH(3) ) _47185_ ( .A(_25268_), .B(3'h0), .S(RST), .Y(_02716_) );
  \$mux  #( .WIDTH(1) ) _47186_ ( .A(1'h0), .B(1'h1), .S(__tmp_1223_1), .Y(_25269_) );
  \$mux  #( .WIDTH(1) ) _47187_ ( .A(_25269_), .B(1'h0), .S(RST), .Y(_02747_) );
  \$mux  #( .WIDTH(1) ) _47188_ ( .A(1'h1), .B(_stream_matmul_29_source_20_source_ram_renable), .S(_05909_), .Y(_25270_) );
  \$mux  #( .WIDTH(1) ) _47189_ ( .A(1'h0), .B(_25270_), .S(_05908_), .Y(_25271_) );
  \$mux  #( .WIDTH(1) ) _47190_ ( .A(_25271_), .B(1'h0), .S(RST), .Y(_02746_) );
  \$mux  #( .WIDTH(32) ) _47191_ ( .A(_stream_matmul_29_source_20_source_pat_all_offset), .B(_stream_matmul_29_source_20_source_ram_raddr), .S(_05909_), .Y(_25272_) );
  \$mux  #( .WIDTH(32) ) _47192_ ( .A(_25272_), .B(0), .S(RST), .Y(_02745_) );
  \$mux  #( .WIDTH(8) ) _47193_ ( .A(_stream_matmul_29_source_20_source_ram_sel), .B(8'h04), .S(_set_flag_1224), .Y(_25273_) );
  \$mux  #( .WIDTH(8) ) _47194_ ( .A(_25273_), .B(8'h00), .S(RST), .Y(_02748_) );
  \$mux  #( .WIDTH(32) ) _47195_ ( .A(_stream_matmul_29_source_20_source_offset_buf), .B(_stream_matmul_29_source_20_source_offset), .S(_06810_), .Y(_25274_) );
  \$mux  #( .WIDTH(32) ) _47196_ ( .A(_25274_), .B(0), .S(RST), .Y(_02743_) );
  \$mux  #( .WIDTH(32) ) _47197_ ( .A(_stream_matmul_29_source_20_source_offset), .B(matmul_29_filter_page_comp_offset_buf), .S(_set_flag_1224), .Y(_25275_) );
  \$mux  #( .WIDTH(32) ) _47198_ ( .A(_25275_), .B(0), .S(RST), .Y(_02742_) );
  \$mux  #( .WIDTH(3) ) _47199_ ( .A(_stream_matmul_29_source_20_source_mode), .B(3'h2), .S(_set_flag_1224), .Y(_25276_) );
  \$mux  #( .WIDTH(3) ) _47200_ ( .A(_25276_), .B(3'h0), .S(RST), .Y(_02741_) );
  \$mux  #( .WIDTH(1) ) _47201_ ( .A(_stream_matmul_29_source_20_idle), .B(1'h0), .S(_06810_), .Y(_25277_) );
  \$mux  #( .WIDTH(1) ) _47202_ ( .A(1'h1), .B(_25277_), .S(_05908_), .Y(_25278_) );
  \$mux  #( .WIDTH(1) ) _47203_ ( .A(_25278_), .B(1'h1), .S(RST), .Y(_02740_) );
  \$mux  #( .WIDTH(1) ) _47204_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id3_0_cond_5_1), .Y(_25279_) );
  \$mux  #( .WIDTH(1) ) _47205_ ( .A(_25279_), .B(1'h0), .S(RST), .Y(_02738_) );
  \$mux  #( .WIDTH(1) ) _47206_ ( .A(1'h1), .B(_stream_matmul_29_source_19_source_ram_renable), .S(_05913_), .Y(_25280_) );
  \$mux  #( .WIDTH(1) ) _47207_ ( .A(1'h0), .B(_25280_), .S(_05910_), .Y(_25281_) );
  \$mux  #( .WIDTH(1) ) _47208_ ( .A(_25281_), .B(1'h0), .S(RST), .Y(_02737_) );
  \$mux  #( .WIDTH(32) ) _47209_ ( .A(_stream_matmul_29_source_19_source_pat_all_offset), .B(_stream_matmul_29_source_19_source_ram_raddr), .S(_05913_), .Y(_25282_) );
  \$mux  #( .WIDTH(32) ) _47210_ ( .A(_25282_), .B(0), .S(RST), .Y(_02736_) );
  \$mux  #( .WIDTH(8) ) _47211_ ( .A(_stream_matmul_29_source_19_source_ram_sel), .B(8'h03), .S(_set_flag_1224), .Y(_25283_) );
  \$mux  #( .WIDTH(8) ) _47212_ ( .A(_25283_), .B(8'h00), .S(RST), .Y(_02739_) );
  \$mux  #( .WIDTH(32) ) _47213_ ( .A(_stream_matmul_29_source_19_source_offset_buf), .B(_stream_matmul_29_source_19_source_offset), .S(_06805_), .Y(_25284_) );
  \$mux  #( .WIDTH(32) ) _47214_ ( .A(_25284_), .B(0), .S(RST), .Y(_02734_) );
  \$mux  #( .WIDTH(32) ) _47215_ ( .A(_stream_matmul_29_source_19_source_offset), .B(_24419_), .S(_set_flag_1224), .Y(_25285_) );
  \$mux  #( .WIDTH(32) ) _47216_ ( .A(_25285_), .B(0), .S(RST), .Y(_02733_) );
  \$mux  #( .WIDTH(3) ) _47217_ ( .A(_stream_matmul_29_source_19_source_mode), .B(3'h2), .S(_set_flag_1224), .Y(_25286_) );
  \$mux  #( .WIDTH(3) ) _47218_ ( .A(_25286_), .B(3'h0), .S(RST), .Y(_02732_) );
  \$mux  #( .WIDTH(1) ) _47219_ ( .A(_stream_matmul_29_source_19_idle), .B(1'h0), .S(_06805_), .Y(_25287_) );
  \$mux  #( .WIDTH(1) ) _47220_ ( .A(1'h1), .B(_25287_), .S(_05910_), .Y(_25288_) );
  \$mux  #( .WIDTH(1) ) _47221_ ( .A(_25288_), .B(1'h1), .S(RST), .Y(_02731_) );
  \$mux  #( .WIDTH(2) ) _47222_ ( .A(_stream_matmul_29_constant_18_next_constant_data), .B({ 1'h0, cparam_matmul_29_keep_filter }), .S(_set_flag_1224), .Y(_25289_) );
  \$mux  #( .WIDTH(2) ) _47223_ ( .A(_25289_), .B(2'h0), .S(RST), .Y(_02708_) );
  \$mux  #( .WIDTH(4) ) _47224_ ( .A(_stream_matmul_29_constant_17_next_constant_data), .B(cparam_matmul_29_cshamt_out_value), .S(_set_flag_1224), .Y(_25290_) );
  \$mux  #( .WIDTH(4) ) _47225_ ( .A(_25290_), .B(4'h0), .S(RST), .Y(_02707_) );
  \$mux  #( .WIDTH(1) ) _47226_ ( .A(_stream_matmul_29_constant_16_next_constant_data), .B(1'h0), .S(_set_flag_1224), .Y(_25291_) );
  \$mux  #( .WIDTH(1) ) _47227_ ( .A(_25291_), .B(1'h0), .S(RST), .Y(_02706_) );
  \$mux  #( .WIDTH(1) ) _47228_ ( .A(_stream_matmul_29_constant_15_next_constant_data), .B(1'h0), .S(_set_flag_1224), .Y(_25292_) );
  \$mux  #( .WIDTH(1) ) _47229_ ( .A(_25292_), .B(1'h0), .S(RST), .Y(_02705_) );
  \$mux  #( .WIDTH(8) ) _47230_ ( .A(_stream_matmul_29_source_14_source_empty_data), .B(8'h00), .S(_set_flag_1224), .Y(_25293_) );
  \$mux  #( .WIDTH(8) ) _47231_ ( .A(_25293_), .B(8'h00), .S(RST), .Y(_02730_) );
  \$mux  #( .WIDTH(1) ) _47232_ ( .A(_stream_matmul_29_source_14_idle), .B(1'h1), .S(_stream_matmul_29_start), .Y(_25294_) );
  \$mux  #( .WIDTH(1) ) _47233_ ( .A(_25294_), .B(1'h1), .S(RST), .Y(_02729_) );
  \$mux  #( .WIDTH(8) ) _47234_ ( .A(_stream_matmul_29_source_12_source_empty_data), .B(8'h00), .S(_set_flag_1224), .Y(_25295_) );
  \$mux  #( .WIDTH(8) ) _47235_ ( .A(_25295_), .B(8'h00), .S(RST), .Y(_02728_) );
  \$mux  #( .WIDTH(1) ) _47236_ ( .A(_stream_matmul_29_source_12_idle), .B(1'h1), .S(_stream_matmul_29_start), .Y(_25296_) );
  \$mux  #( .WIDTH(1) ) _47237_ ( .A(_25296_), .B(1'h1), .S(RST), .Y(_02727_) );
  \$mux  #( .WIDTH(8) ) _47238_ ( .A(_stream_matmul_29_source_10_source_empty_data), .B(8'h00), .S(_set_flag_1224), .Y(_25297_) );
  \$mux  #( .WIDTH(8) ) _47239_ ( .A(_25297_), .B(8'h00), .S(RST), .Y(_02726_) );
  \$mux  #( .WIDTH(1) ) _47240_ ( .A(_stream_matmul_29_source_10_idle), .B(1'h1), .S(_stream_matmul_29_start), .Y(_25298_) );
  \$mux  #( .WIDTH(1) ) _47241_ ( .A(_25298_), .B(1'h1), .S(RST), .Y(_02725_) );
  \$mux  #( .WIDTH(1) ) _47242_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id0_3_cond_5_1), .Y(_25299_) );
  \$mux  #( .WIDTH(1) ) _47243_ ( .A(_25299_), .B(1'h0), .S(RST), .Y(_02765_) );
  \$mux  #( .WIDTH(1) ) _47244_ ( .A(1'h1), .B(_stream_matmul_29_source_8_source_ram_renable), .S(_05911_), .Y(_25300_) );
  \$mux  #( .WIDTH(1) ) _47245_ ( .A(1'h0), .B(_25300_), .S(_05914_), .Y(_25301_) );
  \$mux  #( .WIDTH(1) ) _47246_ ( .A(_25301_), .B(1'h0), .S(RST), .Y(_02764_) );
  \$mux  #( .WIDTH(32) ) _47247_ ( .A(_stream_matmul_29_source_8_source_pat_all_offset), .B(_stream_matmul_29_source_8_source_ram_raddr), .S(_05911_), .Y(_25302_) );
  \$mux  #( .WIDTH(32) ) _47248_ ( .A(_25302_), .B(0), .S(RST), .Y(_02763_) );
  \$mux  #( .WIDTH(8) ) _47249_ ( .A(_stream_matmul_29_source_8_source_ram_sel), .B(8'h02), .S(_set_flag_1224), .Y(_25303_) );
  \$mux  #( .WIDTH(8) ) _47250_ ( .A(_25303_), .B(8'h00), .S(RST), .Y(_02766_) );
  \$mux  #( .WIDTH(32) ) _47251_ ( .A(_stream_matmul_29_source_8_source_offset_buf), .B(_stream_matmul_29_source_8_source_offset), .S(_06800_), .Y(_25304_) );
  \$mux  #( .WIDTH(32) ) _47252_ ( .A(_25304_), .B(0), .S(RST), .Y(_02761_) );
  \$mux  #( .WIDTH(32) ) _47253_ ( .A(_stream_matmul_29_source_8_source_offset), .B(0), .S(_set_flag_1224), .Y(_25305_) );
  \$mux  #( .WIDTH(32) ) _47254_ ( .A(_25305_), .B(0), .S(RST), .Y(_02760_) );
  \$mux  #( .WIDTH(3) ) _47255_ ( .A(_stream_matmul_29_source_8_source_mode), .B(3'h2), .S(_set_flag_1224), .Y(_25306_) );
  \$mux  #( .WIDTH(3) ) _47256_ ( .A(_25306_), .B(3'h0), .S(RST), .Y(_02759_) );
  \$mux  #( .WIDTH(1) ) _47257_ ( .A(_stream_matmul_29_source_8_idle), .B(1'h0), .S(_06800_), .Y(_25307_) );
  \$mux  #( .WIDTH(1) ) _47258_ ( .A(1'h1), .B(_25307_), .S(_05914_), .Y(_25308_) );
  \$mux  #( .WIDTH(1) ) _47259_ ( .A(_25308_), .B(1'h1), .S(RST), .Y(_02758_) );
  \$mux  #( .WIDTH(1) ) _47260_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id2_0_cond_6_1), .Y(_25309_) );
  \$mux  #( .WIDTH(1) ) _47261_ ( .A(_25309_), .B(1'h0), .S(RST), .Y(_02756_) );
  \$mux  #( .WIDTH(1) ) _47262_ ( .A(1'h1), .B(_stream_matmul_29_source_6_source_ram_renable), .S(_05912_), .Y(_25310_) );
  \$mux  #( .WIDTH(1) ) _47263_ ( .A(1'h0), .B(_25310_), .S(_05915_), .Y(_25311_) );
  \$mux  #( .WIDTH(1) ) _47264_ ( .A(_25311_), .B(1'h0), .S(RST), .Y(_02755_) );
  \$mux  #( .WIDTH(32) ) _47265_ ( .A(_stream_matmul_29_source_6_source_pat_all_offset), .B(_stream_matmul_29_source_6_source_ram_raddr), .S(_05912_), .Y(_25312_) );
  \$mux  #( .WIDTH(32) ) _47266_ ( .A(_25312_), .B(0), .S(RST), .Y(_02754_) );
  \$mux  #( .WIDTH(8) ) _47267_ ( .A(_stream_matmul_29_source_6_source_ram_sel), .B(8'h01), .S(_set_flag_1224), .Y(_25313_) );
  \$mux  #( .WIDTH(8) ) _47268_ ( .A(_25313_), .B(8'h00), .S(RST), .Y(_02757_) );
  \$mux  #( .WIDTH(32) ) _47269_ ( .A(_stream_matmul_29_source_6_source_offset_buf), .B(_stream_matmul_29_source_6_source_offset), .S(_06795_), .Y(_25314_) );
  \$mux  #( .WIDTH(32) ) _47270_ ( .A(_25314_), .B(0), .S(RST), .Y(_02752_) );
  \$mux  #( .WIDTH(32) ) _47271_ ( .A(_stream_matmul_29_source_6_source_offset), .B(_29293_), .S(_set_flag_1224), .Y(_25315_) );
  \$mux  #( .WIDTH(32) ) _47272_ ( .A(_25315_), .B(0), .S(RST), .Y(_02751_) );
  \$mux  #( .WIDTH(3) ) _47273_ ( .A(_stream_matmul_29_source_6_source_mode), .B(3'h2), .S(_set_flag_1224), .Y(_25316_) );
  \$mux  #( .WIDTH(3) ) _47274_ ( .A(_25316_), .B(3'h0), .S(RST), .Y(_02750_) );
  \$mux  #( .WIDTH(1) ) _47275_ ( .A(_stream_matmul_29_source_6_idle), .B(1'h0), .S(_06795_), .Y(_25317_) );
  \$mux  #( .WIDTH(1) ) _47276_ ( .A(1'h1), .B(_25317_), .S(_05915_), .Y(_25318_) );
  \$mux  #( .WIDTH(1) ) _47277_ ( .A(_25318_), .B(1'h1), .S(RST), .Y(_02749_) );
  \$mux  #( .WIDTH(1) ) _47278_ ( .A(_stream_matmul_29_constant_3_next_constant_data), .B(matmul_29_stream_pad_masks), .S(_set_flag_1224), .Y(_25319_) );
  \$mux  #( .WIDTH(1) ) _47279_ ( .A(_25319_), .B(1'h0), .S(RST), .Y(_02711_) );
  \$mux  #( .WIDTH(1) ) _47280_ ( .A(_stream_matmul_29_constant_2_next_constant_data), .B(matmul_29_row_select_buf), .S(_set_flag_1224), .Y(_25320_) );
  \$mux  #( .WIDTH(1) ) _47281_ ( .A(_25320_), .B(1'h0), .S(RST), .Y(_02710_) );
  \$mux  #( .WIDTH(1) ) _47282_ ( .A(_stream_matmul_29_constant_1_next_constant_data), .B(matmul_29_col_select), .S(_set_flag_1224), .Y(_25321_) );
  \$mux  #( .WIDTH(1) ) _47283_ ( .A(_25321_), .B(1'h0), .S(RST), .Y(_02709_) );
  \$mux  #( .WIDTH(11) ) _47284_ ( .A(_stream_matmul_29_constant_0_next_constant_data), .B(cparam_matmul_29_act_bat_step), .S(_set_flag_1224), .Y(_25322_) );
  \$mux  #( .WIDTH(11) ) _47285_ ( .A(_25322_), .B(11'h000), .S(RST), .Y(_02704_) );
  \$mux  #( .WIDTH(1) ) _47286_ ( .A(_stream_max_pool_serial_18_reduce_reset), .B(1'h0), .S(__tmp_1046_5), .Y(_25323_) );
  \$mux  #( .WIDTH(1) ) _47287_ ( .A(_25323_), .B(1'h1), .S(__tmp_1060_1), .Y(_25324_) );
  \$mux  #( .WIDTH(1) ) _47288_ ( .A(_25324_), .B(1'h1), .S(RST), .Y(_02774_) );
  \$mux  #( .WIDTH(1) ) _47289_ ( .A(_stream_max_pool_serial_18_source_busy), .B(1'h1), .S(_stream_max_pool_serial_18_start_flag), .Y(_23632_) );
  \$mux  #( .WIDTH(1) ) _47290_ ( .A(_25325_), .B(1'h0), .S(RST), .Y(_02795_) );
  \$mux  #( .WIDTH(1) ) _47291_ ( .A(1'h0), .B(1'h1), .S(__tmp_1070_6), .Y(_25326_) );
  \$mux  #( .WIDTH(1) ) _47292_ ( .A(_25326_), .B(1'h0), .S(RST), .Y(_02797_) );
  \$mux  #( .WIDTH(1) ) _47293_ ( .A(1'h0), .B(1'h1), .S(__tmp_1068_10), .Y(_25327_) );
  \$mux  #( .WIDTH(1) ) _47294_ ( .A(_25327_), .B(1'h0), .S(RST), .Y(_02772_) );
  \$mux  #( .WIDTH(1) ) _47295_ ( .A(1'h0), .B(1'h1), .S(_stream_max_pool_serial_18_start_flag), .Y(_25328_) );
  \$mux  #( .WIDTH(1) ) _47296_ ( .A(_25328_), .B(1'h0), .S(_05686_), .Y(_25329_) );
  \$mux  #( .WIDTH(1) ) _47297_ ( .A(_25329_), .B(1'h0), .S(RST), .Y(_02796_) );
  \$mux  #( .WIDTH(32) ) _47298_ ( .A(_stream_max_pool_serial_18_fsm), .B(3), .S(_stream_max_pool_serial_18_source_1_idle), .Y({ _23689_, _23688_, _23686_, _23685_, _23684_, _23683_, _23682_, _23681_, _23680_, _23679_, _23678_, _23677_, _23675_, _23674_, _23673_, _23672_, _23671_, _23670_, _23669_, _23668_, _23667_, _23666_, _23696_, _23695_, _23694_, _23693_, _23692_, _23691_, _23690_, _23687_, _23676_, _23665_ }) );
  \$mux  #( .WIDTH(32) ) _47299_ ( .A(_stream_max_pool_serial_18_fsm), .B(1), .S(_stream_max_pool_serial_18_start_flag), .Y({ _23721_, _23720_, _23718_, _23717_, _23716_, _23715_, _23714_, _23713_, _23712_, _23711_, _23710_, _23709_, _23707_, _23706_, _23705_, _23704_, _23703_, _23702_, _23701_, _23700_, _23699_, _23698_, _23728_, _23727_, _23726_, _23725_, _23724_, _23723_, _23722_, _23719_, _23708_, _23697_ }) );
  \$mux  #( .WIDTH(32) ) _47300_ ( .A(_25330_), .B(0), .S(RST), .Y(_02773_) );
  \$mux  #( .WIDTH(1) ) _47301_ ( .A(__tmp_1068_9), .B(1'h0), .S(RST), .Y(_01126_) );
  \$mux  #( .WIDTH(1) ) _47302_ ( .A(__tmp_1068_8), .B(1'h0), .S(RST), .Y(_01130_) );
  \$mux  #( .WIDTH(1) ) _47303_ ( .A(__tmp_1068_7), .B(1'h0), .S(RST), .Y(_01129_) );
  \$mux  #( .WIDTH(1) ) _47304_ ( .A(__tmp_1070_6), .B(1'h0), .S(RST), .Y(_01128_) );
  \$mux  #( .WIDTH(1) ) _47305_ ( .A(__tmp_1060_5), .B(1'h0), .S(RST), .Y(_01127_) );
  \$mux  #( .WIDTH(1) ) _47306_ ( .A(__tmp_1042_8), .B(1'h0), .S(RST), .Y(_01120_) );
  \$mux  #( .WIDTH(1) ) _47307_ ( .A(__tmp_1046_7), .B(1'h0), .S(RST), .Y(_01119_) );
  \$mux  #( .WIDTH(1) ) _47308_ ( .A(__tmp_1046_6), .B(1'h0), .S(RST), .Y(_01118_) );
  \$mux  #( .WIDTH(1) ) _47309_ ( .A(__tmp_1046_5), .B(1'h0), .S(RST), .Y(_01117_) );
  \$mux  #( .WIDTH(1) ) _47310_ ( .A(__tmp_1046_4), .B(1'h0), .S(RST), .Y(_01116_) );
  \$mux  #( .WIDTH(1) ) _47311_ ( .A(__tmp_1046_3), .B(1'h0), .S(RST), .Y(_01115_) );
  \$mux  #( .WIDTH(1) ) _47312_ ( .A(__tmp_1046_2), .B(1'h0), .S(RST), .Y(_01114_) );
  \$mux  #( .WIDTH(1) ) _47313_ ( .A(__tmp_1046_1), .B(1'h0), .S(RST), .Y(_01113_) );
  \$mux  #( .WIDTH(1) ) _47314_ ( .A(_tmp_1040), .B(1'h0), .S(RST), .Y(_01112_) );
  \$mux  #( .WIDTH(1) ) _47315_ ( .A(1'h1), .B(1'h0), .S(_05936_), .Y(_25331_) );
  \$mux  #( .WIDTH(1) ) _47316_ ( .A(_25331_), .B(1'h0), .S(RST), .Y(_01871_) );
  \$mux  #( .WIDTH(1) ) _47317_ ( .A(__stream_max_pool_serial_18_start_9), .B(1'h0), .S(RST), .Y(_01079_) );
  \$mux  #( .WIDTH(1) ) _47318_ ( .A(__stream_max_pool_serial_18_start_8), .B(1'h0), .S(RST), .Y(_01088_) );
  \$mux  #( .WIDTH(1) ) _47319_ ( .A(__stream_max_pool_serial_18_start_7), .B(1'h0), .S(RST), .Y(_01087_) );
  \$mux  #( .WIDTH(1) ) _47320_ ( .A(__stream_max_pool_serial_18_start_6), .B(1'h0), .S(RST), .Y(_01086_) );
  \$mux  #( .WIDTH(1) ) _47321_ ( .A(__stream_max_pool_serial_18_start_5), .B(1'h0), .S(RST), .Y(_01085_) );
  \$mux  #( .WIDTH(1) ) _47322_ ( .A(__stream_max_pool_serial_18_start_4), .B(1'h0), .S(RST), .Y(_01084_) );
  \$mux  #( .WIDTH(1) ) _47323_ ( .A(__stream_max_pool_serial_18_start_3), .B(1'h0), .S(RST), .Y(_01083_) );
  \$mux  #( .WIDTH(1) ) _47324_ ( .A(__stream_max_pool_serial_18_start_2), .B(1'h0), .S(RST), .Y(_01082_) );
  \$mux  #( .WIDTH(1) ) _47325_ ( .A(__stream_max_pool_serial_18_start_1), .B(1'h0), .S(RST), .Y(_01081_) );
  \$mux  #( .WIDTH(1) ) _47326_ ( .A(_stream_max_pool_serial_18_start), .B(1'h0), .S(RST), .Y(_01080_) );
  \$mux  #( .WIDTH(1) ) _47327_ ( .A(__set_flag_1036_8), .B(1'h0), .S(RST), .Y(_00714_) );
  \$mux  #( .WIDTH(1) ) _47328_ ( .A(__set_flag_1036_7), .B(1'h0), .S(RST), .Y(_00713_) );
  \$mux  #( .WIDTH(1) ) _47329_ ( .A(__set_flag_1036_6), .B(1'h0), .S(RST), .Y(_00712_) );
  \$mux  #( .WIDTH(1) ) _47330_ ( .A(__set_flag_1036_5), .B(1'h0), .S(RST), .Y(_00711_) );
  \$mux  #( .WIDTH(1) ) _47331_ ( .A(__set_flag_1036_4), .B(1'h0), .S(RST), .Y(_00710_) );
  \$mux  #( .WIDTH(1) ) _47332_ ( .A(__set_flag_1036_3), .B(1'h0), .S(RST), .Y(_00709_) );
  \$mux  #( .WIDTH(1) ) _47333_ ( .A(__set_flag_1036_2), .B(1'h0), .S(RST), .Y(_00708_) );
  \$mux  #( .WIDTH(1) ) _47334_ ( .A(__set_flag_1036_1), .B(1'h0), .S(RST), .Y(_00707_) );
  \$mux  #( .WIDTH(1) ) _47335_ ( .A(_set_flag_1036), .B(1'h0), .S(RST), .Y(_00706_) );
  \$mux  #( .WIDTH(33) ) _47336_ ( .A(__stream_max_pool_serial_18_sink_3_sink_size_1_8), .B(33'h000000000), .S(RST), .Y(_01078_) );
  \$mux  #( .WIDTH(33) ) _47337_ ( .A(__stream_max_pool_serial_18_sink_3_sink_size_1_7), .B(33'h000000000), .S(RST), .Y(_01077_) );
  \$mux  #( .WIDTH(33) ) _47338_ ( .A(__stream_max_pool_serial_18_sink_3_sink_size_1_6), .B(33'h000000000), .S(RST), .Y(_01076_) );
  \$mux  #( .WIDTH(33) ) _47339_ ( .A(__stream_max_pool_serial_18_sink_3_sink_size_1_5), .B(33'h000000000), .S(RST), .Y(_01075_) );
  \$mux  #( .WIDTH(33) ) _47340_ ( .A(__stream_max_pool_serial_18_sink_3_sink_size_1_4), .B(33'h000000000), .S(RST), .Y(_01074_) );
  \$mux  #( .WIDTH(33) ) _47341_ ( .A(__stream_max_pool_serial_18_sink_3_sink_size_1_3), .B(33'h000000000), .S(RST), .Y(_01073_) );
  \$mux  #( .WIDTH(33) ) _47342_ ( .A(__stream_max_pool_serial_18_sink_3_sink_size_1_2), .B(33'h000000000), .S(RST), .Y(_01072_) );
  \$mux  #( .WIDTH(33) ) _47343_ ( .A(__stream_max_pool_serial_18_sink_3_sink_size_1_1), .B(33'h000000000), .S(RST), .Y(_01071_) );
  \$mux  #( .WIDTH(33) ) _47344_ ( .A({ 26'h0000000, cparam_max_pool_serial_18_inc_out_laddr }), .B(33'h000000000), .S(RST), .Y(_01070_) );
  \$mux  #( .WIDTH(32) ) _47345_ ( .A(__stream_max_pool_serial_18_sink_3_sink_offset_0_8), .B(0), .S(RST), .Y(_01069_) );
  \$mux  #( .WIDTH(32) ) _47346_ ( .A(__stream_max_pool_serial_18_sink_3_sink_offset_0_7), .B(0), .S(RST), .Y(_01068_) );
  \$mux  #( .WIDTH(32) ) _47347_ ( .A(__stream_max_pool_serial_18_sink_3_sink_offset_0_6), .B(0), .S(RST), .Y(_01067_) );
  \$mux  #( .WIDTH(32) ) _47348_ ( .A(__stream_max_pool_serial_18_sink_3_sink_offset_0_5), .B(0), .S(RST), .Y(_01066_) );
  \$mux  #( .WIDTH(32) ) _47349_ ( .A(__stream_max_pool_serial_18_sink_3_sink_offset_0_4), .B(0), .S(RST), .Y(_01065_) );
  \$mux  #( .WIDTH(32) ) _47350_ ( .A(__stream_max_pool_serial_18_sink_3_sink_offset_0_3), .B(0), .S(RST), .Y(_01064_) );
  \$mux  #( .WIDTH(32) ) _47351_ ( .A(__stream_max_pool_serial_18_sink_3_sink_offset_0_2), .B(0), .S(RST), .Y(_01063_) );
  \$mux  #( .WIDTH(32) ) _47352_ ( .A(__stream_max_pool_serial_18_sink_3_sink_offset_0_1), .B(0), .S(RST), .Y(_01062_) );
  \$mux  #( .WIDTH(32) ) _47353_ ( .A(_24405_), .B(0), .S(RST), .Y(_01061_) );
  \$mux  #( .WIDTH(8) ) _47354_ ( .A(__variable_wdata_778), .B(_stream_max_pool_serial_18_source_1_source_ram_rdata), .S(_stream_max_pool_serial_18_source_1_source_ram_rvalid), .Y(_25333_) );
  \$mux  #( .WIDTH(8) ) _47355_ ( .A(_25333_), .B(8'h00), .S(RST), .Y(_01446_) );
  \$mux  #( .WIDTH(32) ) _47356_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_stride_buf_3), .B(_source_stream_max_pool_serial_18_source_1_pat_stride_3), .S(_06788_), .Y(_25334_) );
  \$mux  #( .WIDTH(32) ) _47357_ ( .A(_25334_), .B(0), .S(RST), .Y(_02483_) );
  \$mux  #( .WIDTH(32) ) _47358_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_stride_buf_2), .B(_source_stream_max_pool_serial_18_source_1_pat_stride_2), .S(_06788_), .Y(_25335_) );
  \$mux  #( .WIDTH(32) ) _47359_ ( .A(_25335_), .B(0), .S(RST), .Y(_02482_) );
  \$mux  #( .WIDTH(32) ) _47360_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_stride_buf_1), .B(_source_stream_max_pool_serial_18_source_1_pat_stride_1), .S(_06788_), .Y(_25336_) );
  \$mux  #( .WIDTH(32) ) _47361_ ( .A(_25336_), .B(0), .S(RST), .Y(_02481_) );
  \$mux  #( .WIDTH(32) ) _47362_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_stride_buf_0), .B(_source_stream_max_pool_serial_18_source_1_pat_stride_0), .S(_06788_), .Y(_25337_) );
  \$mux  #( .WIDTH(32) ) _47363_ ( .A(_25337_), .B(0), .S(RST), .Y(_02480_) );
  \$mux  #( .WIDTH(33) ) _47364_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_buf_3), .B(_source_stream_max_pool_serial_18_source_1_pat_size_3), .S(_06788_), .Y(_25338_) );
  \$mux  #( .WIDTH(33) ) _47365_ ( .A(_25338_), .B(33'h000000000), .S(RST), .Y(_02475_) );
  \$mux  #( .WIDTH(33) ) _47366_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_buf_2), .B(_source_stream_max_pool_serial_18_source_1_pat_size_2), .S(_06788_), .Y(_25339_) );
  \$mux  #( .WIDTH(33) ) _47367_ ( .A(_25339_), .B(33'h000000000), .S(RST), .Y(_02474_) );
  \$mux  #( .WIDTH(33) ) _47368_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_buf_1), .B(_source_stream_max_pool_serial_18_source_1_pat_size_1), .S(_06788_), .Y(_25340_) );
  \$mux  #( .WIDTH(33) ) _47369_ ( .A(_25340_), .B(33'h000000000), .S(RST), .Y(_02473_) );
  \$mux  #( .WIDTH(33) ) _47370_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_buf_0), .B(_source_stream_max_pool_serial_18_source_1_pat_size_0), .S(_06788_), .Y(_25341_) );
  \$mux  #( .WIDTH(33) ) _47371_ ( .A(_25341_), .B(33'h000000000), .S(RST), .Y(_02472_) );
  \$mux  #( .WIDTH(33) ) _47372_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_3), .B(_28874_), .S(_06788_), .Y(_25342_) );
  \$mux  #( .WIDTH(33) ) _47373_ ( .A(_25342_), .B(_28881_), .S(_06791_), .Y(_25343_) );
  \$mux  #( .WIDTH(33) ) _47374_ ( .A(_25343_), .B(_28882_), .S(_06792_), .Y(_25344_) );
  \$mux  #( .WIDTH(33) ) _47375_ ( .A(_25344_), .B(33'h000000000), .S(RST), .Y(_02463_) );
  \$mux  #( .WIDTH(33) ) _47376_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_2), .B(_28873_), .S(_06788_), .Y(_25345_) );
  \$mux  #( .WIDTH(33) ) _47377_ ( .A(_25345_), .B(_28879_), .S(_06790_), .Y(_25346_) );
  \$mux  #( .WIDTH(33) ) _47378_ ( .A(_25346_), .B(_28880_), .S(_06791_), .Y(_25347_) );
  \$mux  #( .WIDTH(33) ) _47379_ ( .A(_25347_), .B(33'h000000000), .S(RST), .Y(_02462_) );
  \$mux  #( .WIDTH(33) ) _47380_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_1), .B(_28872_), .S(_06788_), .Y(_25348_) );
  \$mux  #( .WIDTH(33) ) _47381_ ( .A(_25348_), .B(_28877_), .S(_06789_), .Y(_25349_) );
  \$mux  #( .WIDTH(33) ) _47382_ ( .A(_25349_), .B(_28878_), .S(_06790_), .Y(_25350_) );
  \$mux  #( .WIDTH(33) ) _47383_ ( .A(_25350_), .B(33'h000000000), .S(RST), .Y(_02461_) );
  \$mux  #( .WIDTH(33) ) _47384_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_count_0), .B(_28871_), .S(_06788_), .Y(_25351_) );
  \$mux  #( .WIDTH(33) ) _47385_ ( .A(_28875_), .B(_25351_), .S(_05932_), .Y(_25352_) );
  \$mux  #( .WIDTH(33) ) _47386_ ( .A(_25352_), .B(_28876_), .S(_06789_), .Y(_25353_) );
  \$mux  #( .WIDTH(33) ) _47387_ ( .A(_25353_), .B(33'h000000000), .S(RST), .Y(_02460_) );
  \$mux  #( .WIDTH(32) ) _47388_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_stride_3), .B(0), .S(_set_flag_1036), .Y(_25354_) );
  \$mux  #( .WIDTH(32) ) _47389_ ( .A(_25354_), .B(0), .S(RST), .Y(_02479_) );
  \$mux  #( .WIDTH(32) ) _47390_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_stride_2), .B(1), .S(_set_flag_1036), .Y(_25355_) );
  \$mux  #( .WIDTH(32) ) _47391_ ( .A(_25355_), .B(0), .S(RST), .Y(_02478_) );
  \$mux  #( .WIDTH(32) ) _47392_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_stride_1), .B(512), .S(_set_flag_1036), .Y(_25356_) );
  \$mux  #( .WIDTH(32) ) _47393_ ( .A(_25356_), .B(0), .S(RST), .Y(_02477_) );
  \$mux  #( .WIDTH(32) ) _47394_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_stride_0), .B({ 25'h0000000, cparam_max_pool_serial_18_inc_out_laddr }), .S(_set_flag_1036), .Y(_25357_) );
  \$mux  #( .WIDTH(32) ) _47395_ ( .A(_25357_), .B(0), .S(RST), .Y(_02476_) );
  \$mux  #( .WIDTH(33) ) _47396_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_3), .B(33'h000000001), .S(_set_flag_1036), .Y(_25358_) );
  \$mux  #( .WIDTH(33) ) _47397_ ( .A(_25358_), .B(33'h000000000), .S(RST), .Y(_02471_) );
  \$mux  #( .WIDTH(33) ) _47398_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_2), .B({ 26'h0000000, cparam_max_pool_serial_18_inc_out_laddr }), .S(_set_flag_1036), .Y(_25359_) );
  \$mux  #( .WIDTH(33) ) _47399_ ( .A(_25359_), .B(33'h000000000), .S(RST), .Y(_02470_) );
  \$mux  #( .WIDTH(33) ) _47400_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_1), .B(33'h000000002), .S(_set_flag_1036), .Y(_25360_) );
  \$mux  #( .WIDTH(33) ) _47401_ ( .A(_25360_), .B(33'h000000000), .S(RST), .Y(_02469_) );
  \$mux  #( .WIDTH(33) ) _47402_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_size_0), .B(33'h000000002), .S(_set_flag_1036), .Y(_25361_) );
  \$mux  #( .WIDTH(33) ) _47403_ ( .A(_25361_), .B(33'h000000000), .S(RST), .Y(_02468_) );
  \$mux  #( .WIDTH(32) ) _47404_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_3), .B(0), .S(_06788_), .Y(_25362_) );
  \$mux  #( .WIDTH(32) ) _47405_ ( .A(_25362_), .B(_24404_), .S(_06791_), .Y(_25363_) );
  \$mux  #( .WIDTH(32) ) _47406_ ( .A(_25363_), .B(0), .S(_06792_), .Y(_25364_) );
  \$mux  #( .WIDTH(32) ) _47407_ ( .A(_25364_), .B(0), .S(RST), .Y(_02467_) );
  \$mux  #( .WIDTH(32) ) _47408_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_2), .B(0), .S(_06788_), .Y(_25365_) );
  \$mux  #( .WIDTH(32) ) _47409_ ( .A(_25365_), .B(_24403_), .S(_06790_), .Y(_25366_) );
  \$mux  #( .WIDTH(32) ) _47410_ ( .A(_25366_), .B(0), .S(_06791_), .Y(_25367_) );
  \$mux  #( .WIDTH(32) ) _47411_ ( .A(_25367_), .B(0), .S(RST), .Y(_02466_) );
  \$mux  #( .WIDTH(32) ) _47412_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_1), .B(0), .S(_06788_), .Y(_25368_) );
  \$mux  #( .WIDTH(32) ) _47413_ ( .A(_25368_), .B(_24402_), .S(_06789_), .Y(_25369_) );
  \$mux  #( .WIDTH(32) ) _47414_ ( .A(_25369_), .B(0), .S(_06790_), .Y(_25370_) );
  \$mux  #( .WIDTH(32) ) _47415_ ( .A(_25370_), .B(0), .S(RST), .Y(_02465_) );
  \$mux  #( .WIDTH(32) ) _47416_ ( .A(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_0), .B(0), .S(_06788_), .Y(_25371_) );
  \$mux  #( .WIDTH(32) ) _47417_ ( .A(_24401_), .B(_25371_), .S(_05932_), .Y(_25372_) );
  \$mux  #( .WIDTH(32) ) _47418_ ( .A(_25372_), .B(0), .S(_06789_), .Y(_25373_) );
  \$mux  #( .WIDTH(32) ) _47419_ ( .A(_25373_), .B(0), .S(RST), .Y(_02464_) );
  \$mux  #( .WIDTH(4) ) _47420_ ( .A(__variable_wdata_779), .B(_stream_max_pool_serial_18_constant_2_next_constant_data), .S(_stream_max_pool_serial_18_start), .Y(_25374_) );
  \$mux  #( .WIDTH(4) ) _47421_ ( .A(_25374_), .B(4'h0), .S(RST), .Y(_01447_) );
  \$mux  #( .WIDTH(3) ) _47422_ ( .A(__variable_wdata_777), .B(_stream_max_pool_serial_18_constant_0_next_constant_data), .S(_stream_max_pool_serial_18_start), .Y(_25375_) );
  \$mux  #( .WIDTH(3) ) _47423_ ( .A(_25375_), .B(3'h0), .S(RST), .Y(_01445_) );
  \$mux  #( .WIDTH(1) ) _47424_ ( .A(1'h1), .B(1'h0), .S(_05935_), .Y(_25332_) );
  \$mux  #( .WIDTH(1) ) _47425_ ( .A(_25332_), .B(1'h0), .S(RST), .Y(_01870_) );
  \$mux  #( .WIDTH(1) ) _47426_ ( .A(_pulse_data_213), .B(1'h0), .S(RST), .Y(_01103_) );
  \$mux  #( .WIDTH(8) ) _47427_ ( .A(_reducemax_data_211), .B(8'h00), .S(RST), .Y(_01102_) );
  \$mux  #( .WIDTH(3) ) _47428_ ( .A(__delay_data_1415), .B(3'h0), .S(RST), .Y(_00297_) );
  \$mux  #( .WIDTH(9) ) _47429_ ( .A(_29281_), .B(9'h000), .S(RST), .Y(_01548_) );
  \$mux  #( .WIDTH(3) ) _47430_ ( .A(__delay_data_1414), .B(3'h0), .S(RST), .Y(_00296_) );
  \$mux  #( .WIDTH(8) ) _47431_ ( .A(__delay_data_1412), .B(8'h00), .S(RST), .Y(_00294_) );
  \$mux  #( .WIDTH(1) ) _47432_ ( .A(_28508_[0]), .B(1'h0), .S(RST), .Y(_01819_) );
  \$mux  #( .WIDTH(3) ) _47433_ ( .A(__variable_wdata_777), .B(3'h0), .S(RST), .Y(_00295_) );
  \$mux  #( .WIDTH(8) ) _47434_ ( .A(__variable_wdata_778), .B(8'h00), .S(RST), .Y(_00293_) );
  \$mux  #( .WIDTH(4) ) _47435_ ( .A(__variable_wdata_779), .B(4'h0), .S(RST), .Y(_00292_) );
  \$mux  #( .WIDTH(32) ) _47436_ ( .A(_29280_), .B(0), .S(_stream_max_pool_serial_18_reduce_reset), .Y(_25376_) );
  \$mux  #( .WIDTH(32) ) _47437_ ( .A(_25376_), .B(0), .S(RST), .Y(_01579_) );
  \$mux  #( .WIDTH(32) ) _47438_ ( .A(_counter_count_782), .B(0), .S(_stream_max_pool_serial_18_reduce_reset), .Y(_25377_) );
  \$mux  #( .WIDTH(32) ) _47439_ ( .A(_25377_), .B(0), .S(RST), .Y(_01580_) );
  \$mux  #( .WIDTH(8) ) _47440_ ( .A(_stream_max_pool_serial_18_sink_3_sink_wdata), .B(__substreamoutput_data_793), .S(_06794_), .Y(_25378_) );
  \$mux  #( .WIDTH(8) ) _47441_ ( .A(_25378_), .B(8'h00), .S(RST), .Y(_02784_) );
  \$mux  #( .WIDTH(1) ) _47442_ ( .A(1'h0), .B(1'h1), .S(_06794_), .Y(_25379_) );
  \$mux  #( .WIDTH(1) ) _47443_ ( .A(_25379_), .B(1'h0), .S(RST), .Y(_02785_) );
  \$mux  #( .WIDTH(32) ) _47444_ ( .A(_stream_max_pool_serial_18_sink_3_sink_waddr), .B(_28883_), .S(_06793_), .Y(_25380_) );
  \$mux  #( .WIDTH(32) ) _47445_ ( .A(_25380_), .B(_24406_), .S(_06794_), .Y(_25381_) );
  \$mux  #( .WIDTH(32) ) _47446_ ( .A(_25381_), .B(0), .S(RST), .Y(_02783_) );
  \$mux  #( .WIDTH(8) ) _47447_ ( .A(_stream_max_pool_serial_18_sink_3_sink_ram_sel), .B(8'h02), .S(__set_flag_1036_9), .Y(_25382_) );
  \$mux  #( .WIDTH(8) ) _47448_ ( .A(_25382_), .B(8'h00), .S(RST), .Y(_02779_) );
  \$mux  #( .WIDTH(32) ) _47449_ ( .A(_stream_max_pool_serial_18_sink_3_sink_stride_buf), .B(_stream_max_pool_serial_18_sink_3_sink_stride), .S(_06793_), .Y(_25383_) );
  \$mux  #( .WIDTH(32) ) _47450_ ( .A(_25383_), .B(0), .S(RST), .Y(_02782_) );
  \$mux  #( .WIDTH(33) ) _47451_ ( .A(_stream_max_pool_serial_18_sink_3_sink_count), .B(_stream_max_pool_serial_18_sink_3_sink_size), .S(_06793_), .Y(_25384_) );
  \$mux  #( .WIDTH(33) ) _47452_ ( .A(_25384_), .B(_28884_), .S(_06794_), .Y(_25385_) );
  \$mux  #( .WIDTH(33) ) _47453_ ( .A(_25385_), .B(33'h000000000), .S(RST), .Y(_02775_) );
  \$mux  #( .WIDTH(32) ) _47454_ ( .A(_stream_max_pool_serial_18_sink_3_sink_stride), .B(1), .S(__set_flag_1036_9), .Y(_25386_) );
  \$mux  #( .WIDTH(32) ) _47455_ ( .A(_25386_), .B(0), .S(RST), .Y(_02781_) );
  \$mux  #( .WIDTH(33) ) _47456_ ( .A(_stream_max_pool_serial_18_sink_3_sink_size), .B(__stream_max_pool_serial_18_sink_3_sink_size_1_9), .S(__set_flag_1036_9), .Y(_25387_) );
  \$mux  #( .WIDTH(33) ) _47457_ ( .A(_25387_), .B(33'h000000000), .S(RST), .Y(_02780_) );
  \$mux  #( .WIDTH(32) ) _47458_ ( .A(_stream_max_pool_serial_18_sink_3_sink_offset), .B(__stream_max_pool_serial_18_sink_3_sink_offset_0_9), .S(__set_flag_1036_9), .Y(_25388_) );
  \$mux  #( .WIDTH(32) ) _47459_ ( .A(_25388_), .B(0), .S(RST), .Y(_02778_) );
  \$mux  #( .WIDTH(3) ) _47460_ ( .A(_stream_max_pool_serial_18_sink_3_sink_mode), .B(3'h1), .S(__set_flag_1036_9), .Y(_25389_) );
  \$mux  #( .WIDTH(3) ) _47461_ ( .A(_25389_), .B(3'h0), .S(RST), .Y(_02777_) );
  \$mux  #( .WIDTH(4) ) _47462_ ( .A(_stream_max_pool_serial_18_constant_2_next_constant_data), .B(max_pool_serial_18_stream_pad_masks), .S(_set_flag_1036), .Y(_25390_) );
  \$mux  #( .WIDTH(4) ) _47463_ ( .A(_25390_), .B(4'h0), .S(RST), .Y(_02771_) );
  \$mux  #( .WIDTH(1) ) _47464_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id1_0_cond_4_1), .Y(_25391_) );
  \$mux  #( .WIDTH(1) ) _47465_ ( .A(_25391_), .B(1'h0), .S(RST), .Y(_02793_) );
  \$mux  #( .WIDTH(1) ) _47466_ ( .A(1'h1), .B(_stream_max_pool_serial_18_source_1_source_ram_renable), .S(_05932_), .Y(_25392_) );
  \$mux  #( .WIDTH(1) ) _47467_ ( .A(1'h0), .B(_25392_), .S(_05933_), .Y(_25393_) );
  \$mux  #( .WIDTH(1) ) _47468_ ( .A(_25393_), .B(1'h0), .S(RST), .Y(_02792_) );
  \$mux  #( .WIDTH(32) ) _47469_ ( .A(_stream_max_pool_serial_18_source_1_source_pat_all_offset), .B(_stream_max_pool_serial_18_source_1_source_ram_raddr), .S(_05932_), .Y(_25394_) );
  \$mux  #( .WIDTH(32) ) _47470_ ( .A(_25394_), .B(0), .S(RST), .Y(_02791_) );
  \$mux  #( .WIDTH(8) ) _47471_ ( .A(_stream_max_pool_serial_18_source_1_source_ram_sel), .B(8'h01), .S(_set_flag_1036), .Y(_25395_) );
  \$mux  #( .WIDTH(8) ) _47472_ ( .A(_25395_), .B(8'h00), .S(RST), .Y(_02794_) );
  \$mux  #( .WIDTH(32) ) _47473_ ( .A(_stream_max_pool_serial_18_source_1_source_offset_buf), .B(_stream_max_pool_serial_18_source_1_source_offset), .S(_06788_), .Y(_25396_) );
  \$mux  #( .WIDTH(32) ) _47474_ ( .A(_25396_), .B(0), .S(RST), .Y(_02789_) );
  \$mux  #( .WIDTH(32) ) _47475_ ( .A(_stream_max_pool_serial_18_source_1_source_offset), .B(_24400_), .S(_set_flag_1036), .Y(_25397_) );
  \$mux  #( .WIDTH(32) ) _47476_ ( .A(_25397_), .B(0), .S(RST), .Y(_02788_) );
  \$mux  #( .WIDTH(3) ) _47477_ ( .A(_stream_max_pool_serial_18_source_1_source_mode), .B(3'h2), .S(_set_flag_1036), .Y(_25398_) );
  \$mux  #( .WIDTH(3) ) _47478_ ( .A(_25398_), .B(3'h0), .S(RST), .Y(_02787_) );
  \$mux  #( .WIDTH(1) ) _47479_ ( .A(_stream_max_pool_serial_18_source_1_idle), .B(1'h0), .S(_06788_), .Y(_25399_) );
  \$mux  #( .WIDTH(1) ) _47480_ ( .A(1'h1), .B(_25399_), .S(_05933_), .Y(_25400_) );
  \$mux  #( .WIDTH(1) ) _47481_ ( .A(_25400_), .B(1'h1), .S(RST), .Y(_02786_) );
  \$mux  #( .WIDTH(3) ) _47482_ ( .A(_stream_max_pool_serial_18_constant_0_next_constant_data), .B(3'h4), .S(_set_flag_1036), .Y(_25401_) );
  \$mux  #( .WIDTH(3) ) _47483_ ( .A(_25401_), .B(3'h0), .S(RST), .Y(_02770_) );
  \$mux  #( .WIDTH(1) ) _47484_ ( .A(_stream_conv2d_16_source_busy), .B(1'h1), .S(_stream_conv2d_16_start_flag), .Y(_23730_) );
  \$mux  #( .WIDTH(1) ) _47485_ ( .A(_25402_), .B(1'h0), .S(RST), .Y(_02701_) );
  \$mux  #( .WIDTH(1) ) _47486_ ( .A(1'h0), .B(1'h1), .S(__tmp_969_42), .Y(_25403_) );
  \$mux  #( .WIDTH(1) ) _47487_ ( .A(_25403_), .B(1'h0), .S(RST), .Y(_02703_) );
  \$mux  #( .WIDTH(1) ) _47488_ ( .A(1'h0), .B(1'h1), .S(__tmp_967_46), .Y(_25404_) );
  \$mux  #( .WIDTH(1) ) _47489_ ( .A(_25404_), .B(1'h0), .S(RST), .Y(_02502_) );
  \$mux  #( .WIDTH(1) ) _47490_ ( .A(1'h0), .B(1'h1), .S(_stream_conv2d_16_start_flag), .Y(_25405_) );
  \$mux  #( .WIDTH(1) ) _47491_ ( .A(_25405_), .B(1'h0), .S(_05687_), .Y(_25406_) );
  \$mux  #( .WIDTH(1) ) _47492_ ( .A(_25406_), .B(1'h0), .S(RST), .Y(_02702_) );
  \$mux  #( .WIDTH(32) ) _47493_ ( .A(_stream_conv2d_16_fsm), .B(3), .S(_stream_conv2d_16_done), .Y({ _23787_, _23786_, _23784_, _23783_, _23782_, _23781_, _23780_, _23779_, _23778_, _23777_, _23776_, _23775_, _23773_, _23772_, _23771_, _23770_, _23769_, _23768_, _23767_, _23766_, _23765_, _23764_, _23794_, _23793_, _23792_, _23791_, _23790_, _23789_, _23788_, _23785_, _23774_, _23763_ }) );
  \$mux  #( .WIDTH(32) ) _47494_ ( .A(_stream_conv2d_16_fsm), .B(1), .S(_stream_conv2d_16_start_flag), .Y({ _23819_, _23818_, _23816_, _23815_, _23814_, _23813_, _23812_, _23811_, _23810_, _23809_, _23808_, _23807_, _23805_, _23804_, _23803_, _23802_, _23801_, _23800_, _23799_, _23798_, _23797_, _23796_, _23826_, _23825_, _23824_, _23823_, _23822_, _23821_, _23820_, _23817_, _23806_, _23795_ }) );
  \$mux  #( .WIDTH(32) ) _47495_ ( .A(_25407_), .B(0), .S(RST), .Y(_02503_) );
  \$mux  #( .WIDTH(1) ) _47496_ ( .A(__tmp_967_45), .B(1'h0), .S(RST), .Y(_01368_) );
  \$mux  #( .WIDTH(1) ) _47497_ ( .A(__tmp_967_44), .B(1'h0), .S(RST), .Y(_01367_) );
  \$mux  #( .WIDTH(1) ) _47498_ ( .A(__tmp_967_43), .B(1'h0), .S(RST), .Y(_01366_) );
  \$mux  #( .WIDTH(1) ) _47499_ ( .A(__tmp_969_42), .B(1'h0), .S(RST), .Y(_01365_) );
  \$mux  #( .WIDTH(1) ) _47500_ ( .A(__tmp_969_41), .B(1'h0), .S(RST), .Y(_01364_) );
  \$mux  #( .WIDTH(1) ) _47501_ ( .A(__tmp_969_40), .B(1'h0), .S(RST), .Y(_01363_) );
  \$mux  #( .WIDTH(1) ) _47502_ ( .A(__tmp_969_39), .B(1'h0), .S(RST), .Y(_01362_) );
  \$mux  #( .WIDTH(1) ) _47503_ ( .A(__tmp_969_38), .B(1'h0), .S(RST), .Y(_01361_) );
  \$mux  #( .WIDTH(1) ) _47504_ ( .A(__tmp_969_37), .B(1'h0), .S(RST), .Y(_01360_) );
  \$mux  #( .WIDTH(1) ) _47505_ ( .A(__tmp_969_36), .B(1'h0), .S(RST), .Y(_01359_) );
  \$mux  #( .WIDTH(1) ) _47506_ ( .A(__tmp_969_35), .B(1'h0), .S(RST), .Y(_01358_) );
  \$mux  #( .WIDTH(1) ) _47507_ ( .A(__tmp_969_34), .B(1'h0), .S(RST), .Y(_01357_) );
  \$mux  #( .WIDTH(1) ) _47508_ ( .A(__tmp_969_33), .B(1'h0), .S(RST), .Y(_01356_) );
  \$mux  #( .WIDTH(1) ) _47509_ ( .A(__tmp_969_32), .B(1'h0), .S(RST), .Y(_01355_) );
  \$mux  #( .WIDTH(1) ) _47510_ ( .A(__tmp_969_31), .B(1'h0), .S(RST), .Y(_01354_) );
  \$mux  #( .WIDTH(1) ) _47511_ ( .A(__tmp_969_30), .B(1'h0), .S(RST), .Y(_01353_) );
  \$mux  #( .WIDTH(1) ) _47512_ ( .A(__tmp_969_29), .B(1'h0), .S(RST), .Y(_01352_) );
  \$mux  #( .WIDTH(1) ) _47513_ ( .A(__tmp_969_28), .B(1'h0), .S(RST), .Y(_01351_) );
  \$mux  #( .WIDTH(1) ) _47514_ ( .A(__tmp_969_27), .B(1'h0), .S(RST), .Y(_01350_) );
  \$mux  #( .WIDTH(1) ) _47515_ ( .A(__tmp_969_26), .B(1'h0), .S(RST), .Y(_01349_) );
  \$mux  #( .WIDTH(1) ) _47516_ ( .A(__tmp_969_25), .B(1'h0), .S(RST), .Y(_01348_) );
  \$mux  #( .WIDTH(1) ) _47517_ ( .A(__tmp_969_24), .B(1'h0), .S(RST), .Y(_01347_) );
  \$mux  #( .WIDTH(1) ) _47518_ ( .A(__tmp_969_23), .B(1'h0), .S(RST), .Y(_01346_) );
  \$mux  #( .WIDTH(1) ) _47519_ ( .A(__tmp_969_22), .B(1'h0), .S(RST), .Y(_01345_) );
  \$mux  #( .WIDTH(1) ) _47520_ ( .A(__tmp_969_21), .B(1'h0), .S(RST), .Y(_01344_) );
  \$mux  #( .WIDTH(1) ) _47521_ ( .A(__tmp_969_20), .B(1'h0), .S(RST), .Y(_01343_) );
  \$mux  #( .WIDTH(1) ) _47522_ ( .A(__tmp_969_19), .B(1'h0), .S(RST), .Y(_01342_) );
  \$mux  #( .WIDTH(1) ) _47523_ ( .A(__tmp_969_18), .B(1'h0), .S(RST), .Y(_01341_) );
  \$mux  #( .WIDTH(1) ) _47524_ ( .A(__tmp_969_17), .B(1'h0), .S(RST), .Y(_01340_) );
  \$mux  #( .WIDTH(1) ) _47525_ ( .A(__tmp_969_16), .B(1'h0), .S(RST), .Y(_01339_) );
  \$mux  #( .WIDTH(1) ) _47526_ ( .A(__tmp_969_15), .B(1'h0), .S(RST), .Y(_01338_) );
  \$mux  #( .WIDTH(1) ) _47527_ ( .A(__tmp_969_14), .B(1'h0), .S(RST), .Y(_01337_) );
  \$mux  #( .WIDTH(1) ) _47528_ ( .A(__tmp_969_13), .B(1'h0), .S(RST), .Y(_01336_) );
  \$mux  #( .WIDTH(1) ) _47529_ ( .A(__tmp_959_12), .B(1'h0), .S(RST), .Y(_01335_) );
  \$mux  #( .WIDTH(1) ) _47530_ ( .A(__tmp_799_32), .B(1'h0), .S(RST), .Y(_01321_) );
  \$mux  #( .WIDTH(1) ) _47531_ ( .A(__tmp_799_31), .B(1'h0), .S(RST), .Y(_01320_) );
  \$mux  #( .WIDTH(1) ) _47532_ ( .A(__tmp_799_33), .B(1'h0), .S(RST), .Y(_01322_) );
  \$mux  #( .WIDTH(1) ) _47533_ ( .A(__tmp_799_30), .B(1'h0), .S(RST), .Y(_01319_) );
  \$mux  #( .WIDTH(1) ) _47534_ ( .A(__tmp_799_29), .B(1'h0), .S(RST), .Y(_01318_) );
  \$mux  #( .WIDTH(1) ) _47535_ ( .A(__tmp_799_28), .B(1'h0), .S(RST), .Y(_01317_) );
  \$mux  #( .WIDTH(1) ) _47536_ ( .A(__tmp_799_27), .B(1'h0), .S(RST), .Y(_01316_) );
  \$mux  #( .WIDTH(1) ) _47537_ ( .A(__tmp_799_26), .B(1'h0), .S(RST), .Y(_01315_) );
  \$mux  #( .WIDTH(1) ) _47538_ ( .A(__tmp_799_25), .B(1'h0), .S(RST), .Y(_01314_) );
  \$mux  #( .WIDTH(1) ) _47539_ ( .A(__tmp_799_24), .B(1'h0), .S(RST), .Y(_01313_) );
  \$mux  #( .WIDTH(1) ) _47540_ ( .A(__tmp_799_23), .B(1'h0), .S(RST), .Y(_01312_) );
  \$mux  #( .WIDTH(1) ) _47541_ ( .A(__tmp_799_22), .B(1'h0), .S(RST), .Y(_01311_) );
  \$mux  #( .WIDTH(1) ) _47542_ ( .A(__tmp_799_21), .B(1'h0), .S(RST), .Y(_01310_) );
  \$mux  #( .WIDTH(1) ) _47543_ ( .A(__tmp_799_20), .B(1'h0), .S(RST), .Y(_01309_) );
  \$mux  #( .WIDTH(1) ) _47544_ ( .A(__tmp_799_19), .B(1'h0), .S(RST), .Y(_01308_) );
  \$mux  #( .WIDTH(1) ) _47545_ ( .A(__tmp_799_18), .B(1'h0), .S(RST), .Y(_01307_) );
  \$mux  #( .WIDTH(1) ) _47546_ ( .A(__tmp_799_17), .B(1'h0), .S(RST), .Y(_01306_) );
  \$mux  #( .WIDTH(1) ) _47547_ ( .A(__tmp_799_16), .B(1'h0), .S(RST), .Y(_01305_) );
  \$mux  #( .WIDTH(1) ) _47548_ ( .A(__tmp_799_15), .B(1'h0), .S(RST), .Y(_01304_) );
  \$mux  #( .WIDTH(1) ) _47549_ ( .A(__tmp_799_14), .B(1'h0), .S(RST), .Y(_01303_) );
  \$mux  #( .WIDTH(1) ) _47550_ ( .A(__tmp_799_13), .B(1'h0), .S(RST), .Y(_01302_) );
  \$mux  #( .WIDTH(1) ) _47551_ ( .A(__tmp_799_12), .B(1'h0), .S(RST), .Y(_01301_) );
  \$mux  #( .WIDTH(1) ) _47552_ ( .A(__tmp_799_11), .B(1'h0), .S(RST), .Y(_01296_) );
  \$mux  #( .WIDTH(1) ) _47553_ ( .A(__tmp_799_10), .B(1'h0), .S(RST), .Y(_01295_) );
  \$mux  #( .WIDTH(1) ) _47554_ ( .A(__tmp_799_9), .B(1'h0), .S(RST), .Y(_01294_) );
  \$mux  #( .WIDTH(1) ) _47555_ ( .A(__tmp_799_8), .B(1'h0), .S(RST), .Y(_01300_) );
  \$mux  #( .WIDTH(1) ) _47556_ ( .A(__tmp_799_7), .B(1'h0), .S(RST), .Y(_01299_) );
  \$mux  #( .WIDTH(1) ) _47557_ ( .A(__tmp_799_6), .B(1'h0), .S(RST), .Y(_01298_) );
  \$mux  #( .WIDTH(1) ) _47558_ ( .A(__tmp_799_5), .B(1'h0), .S(RST), .Y(_01297_) );
  \$mux  #( .WIDTH(1) ) _47559_ ( .A(__tmp_799_4), .B(1'h0), .S(RST), .Y(_01293_) );
  \$mux  #( .WIDTH(1) ) _47560_ ( .A(__tmp_799_3), .B(1'h0), .S(RST), .Y(_01292_) );
  \$mux  #( .WIDTH(1) ) _47561_ ( .A(__tmp_799_2), .B(1'h0), .S(RST), .Y(_01291_) );
  \$mux  #( .WIDTH(1) ) _47562_ ( .A(__tmp_799_1), .B(1'h0), .S(RST), .Y(_01290_) );
  \$mux  #( .WIDTH(1) ) _47563_ ( .A(_tmp_713), .B(1'h0), .S(RST), .Y(_01289_) );
  \$mux  #( .WIDTH(1) ) _47564_ ( .A(__stream_conv2d_16_start_45), .B(1'h0), .S(RST), .Y(_00930_) );
  \$mux  #( .WIDTH(1) ) _47565_ ( .A(__stream_conv2d_16_start_44), .B(1'h0), .S(RST), .Y(_00929_) );
  \$mux  #( .WIDTH(1) ) _47566_ ( .A(__stream_conv2d_16_start_43), .B(1'h0), .S(RST), .Y(_00928_) );
  \$mux  #( .WIDTH(1) ) _47567_ ( .A(__stream_conv2d_16_start_42), .B(1'h0), .S(RST), .Y(_00927_) );
  \$mux  #( .WIDTH(1) ) _47568_ ( .A(__stream_conv2d_16_start_41), .B(1'h0), .S(RST), .Y(_00926_) );
  \$mux  #( .WIDTH(1) ) _47569_ ( .A(__stream_conv2d_16_start_40), .B(1'h0), .S(RST), .Y(_00925_) );
  \$mux  #( .WIDTH(1) ) _47570_ ( .A(__stream_conv2d_16_start_39), .B(1'h0), .S(RST), .Y(_00924_) );
  \$mux  #( .WIDTH(1) ) _47571_ ( .A(__stream_conv2d_16_start_38), .B(1'h0), .S(RST), .Y(_00922_) );
  \$mux  #( .WIDTH(1) ) _47572_ ( .A(__stream_conv2d_16_start_37), .B(1'h0), .S(RST), .Y(_00921_) );
  \$mux  #( .WIDTH(1) ) _47573_ ( .A(__stream_conv2d_16_start_36), .B(1'h0), .S(RST), .Y(_00920_) );
  \$mux  #( .WIDTH(1) ) _47574_ ( .A(__stream_conv2d_16_start_35), .B(1'h0), .S(RST), .Y(_00919_) );
  \$mux  #( .WIDTH(1) ) _47575_ ( .A(__stream_conv2d_16_start_34), .B(1'h0), .S(RST), .Y(_00918_) );
  \$mux  #( .WIDTH(1) ) _47576_ ( .A(__stream_conv2d_16_start_33), .B(1'h0), .S(RST), .Y(_00917_) );
  \$mux  #( .WIDTH(1) ) _47577_ ( .A(__stream_conv2d_16_start_32), .B(1'h0), .S(RST), .Y(_00916_) );
  \$mux  #( .WIDTH(1) ) _47578_ ( .A(__stream_conv2d_16_start_31), .B(1'h0), .S(RST), .Y(_00915_) );
  \$mux  #( .WIDTH(1) ) _47579_ ( .A(__stream_conv2d_16_start_30), .B(1'h0), .S(RST), .Y(_00914_) );
  \$mux  #( .WIDTH(1) ) _47580_ ( .A(__stream_conv2d_16_start_29), .B(1'h0), .S(RST), .Y(_00913_) );
  \$mux  #( .WIDTH(1) ) _47581_ ( .A(__stream_conv2d_16_start_28), .B(1'h0), .S(RST), .Y(_00911_) );
  \$mux  #( .WIDTH(1) ) _47582_ ( .A(__stream_conv2d_16_start_27), .B(1'h0), .S(RST), .Y(_00910_) );
  \$mux  #( .WIDTH(1) ) _47583_ ( .A(__stream_conv2d_16_start_26), .B(1'h0), .S(RST), .Y(_00909_) );
  \$mux  #( .WIDTH(1) ) _47584_ ( .A(__stream_conv2d_16_start_25), .B(1'h0), .S(RST), .Y(_00908_) );
  \$mux  #( .WIDTH(1) ) _47585_ ( .A(__stream_conv2d_16_start_24), .B(1'h0), .S(RST), .Y(_00907_) );
  \$mux  #( .WIDTH(1) ) _47586_ ( .A(__stream_conv2d_16_start_23), .B(1'h0), .S(RST), .Y(_00906_) );
  \$mux  #( .WIDTH(1) ) _47587_ ( .A(__stream_conv2d_16_start_22), .B(1'h0), .S(RST), .Y(_00905_) );
  \$mux  #( .WIDTH(1) ) _47588_ ( .A(__stream_conv2d_16_start_21), .B(1'h0), .S(RST), .Y(_00904_) );
  \$mux  #( .WIDTH(1) ) _47589_ ( .A(__stream_conv2d_16_start_20), .B(1'h0), .S(RST), .Y(_00903_) );
  \$mux  #( .WIDTH(1) ) _47590_ ( .A(__stream_conv2d_16_start_19), .B(1'h0), .S(RST), .Y(_00902_) );
  \$mux  #( .WIDTH(1) ) _47591_ ( .A(__stream_conv2d_16_start_18), .B(1'h0), .S(RST), .Y(_00900_) );
  \$mux  #( .WIDTH(1) ) _47592_ ( .A(__stream_conv2d_16_start_17), .B(1'h0), .S(RST), .Y(_00899_) );
  \$mux  #( .WIDTH(1) ) _47593_ ( .A(__stream_conv2d_16_start_16), .B(1'h0), .S(RST), .Y(_00898_) );
  \$mux  #( .WIDTH(1) ) _47594_ ( .A(__stream_conv2d_16_start_15), .B(1'h0), .S(RST), .Y(_00897_) );
  \$mux  #( .WIDTH(1) ) _47595_ ( .A(__stream_conv2d_16_start_14), .B(1'h0), .S(RST), .Y(_00896_) );
  \$mux  #( .WIDTH(1) ) _47596_ ( .A(__stream_conv2d_16_start_13), .B(1'h0), .S(RST), .Y(_00895_) );
  \$mux  #( .WIDTH(1) ) _47597_ ( .A(__stream_conv2d_16_start_12), .B(1'h0), .S(RST), .Y(_00894_) );
  \$mux  #( .WIDTH(1) ) _47598_ ( .A(__stream_conv2d_16_start_11), .B(1'h0), .S(RST), .Y(_00893_) );
  \$mux  #( .WIDTH(1) ) _47599_ ( .A(__stream_conv2d_16_start_10), .B(1'h0), .S(RST), .Y(_00892_) );
  \$mux  #( .WIDTH(1) ) _47600_ ( .A(__stream_conv2d_16_start_9), .B(1'h0), .S(RST), .Y(_00891_) );
  \$mux  #( .WIDTH(1) ) _47601_ ( .A(__stream_conv2d_16_start_8), .B(1'h0), .S(RST), .Y(_00936_) );
  \$mux  #( .WIDTH(1) ) _47602_ ( .A(__stream_conv2d_16_start_7), .B(1'h0), .S(RST), .Y(_00935_) );
  \$mux  #( .WIDTH(1) ) _47603_ ( .A(__stream_conv2d_16_start_6), .B(1'h0), .S(RST), .Y(_00934_) );
  \$mux  #( .WIDTH(1) ) _47604_ ( .A(__stream_conv2d_16_start_5), .B(1'h0), .S(RST), .Y(_00933_) );
  \$mux  #( .WIDTH(1) ) _47605_ ( .A(__stream_conv2d_16_start_4), .B(1'h0), .S(RST), .Y(_00932_) );
  \$mux  #( .WIDTH(1) ) _47606_ ( .A(__stream_conv2d_16_start_3), .B(1'h0), .S(RST), .Y(_00931_) );
  \$mux  #( .WIDTH(1) ) _47607_ ( .A(__stream_conv2d_16_start_2), .B(1'h0), .S(RST), .Y(_00923_) );
  \$mux  #( .WIDTH(1) ) _47608_ ( .A(__stream_conv2d_16_start_1), .B(1'h0), .S(RST), .Y(_00912_) );
  \$mux  #( .WIDTH(1) ) _47609_ ( .A(_stream_conv2d_16_start), .B(1'h0), .S(RST), .Y(_00901_) );
  \$mux  #( .WIDTH(1) ) _47610_ ( .A(__set_flag_710_42), .B(1'h0), .S(RST), .Y(_00792_) );
  \$mux  #( .WIDTH(1) ) _47611_ ( .A(__set_flag_710_41), .B(1'h0), .S(RST), .Y(_00791_) );
  \$mux  #( .WIDTH(1) ) _47612_ ( .A(__set_flag_710_40), .B(1'h0), .S(RST), .Y(_00790_) );
  \$mux  #( .WIDTH(1) ) _47613_ ( .A(__set_flag_710_39), .B(1'h0), .S(RST), .Y(_00789_) );
  \$mux  #( .WIDTH(1) ) _47614_ ( .A(__set_flag_710_36), .B(1'h0), .S(RST), .Y(_00785_) );
  \$mux  #( .WIDTH(1) ) _47615_ ( .A(__set_flag_710_34), .B(1'h0), .S(RST), .Y(_00783_) );
  \$mux  #( .WIDTH(1) ) _47616_ ( .A(__set_flag_710_32), .B(1'h0), .S(RST), .Y(_00781_) );
  \$mux  #( .WIDTH(1) ) _47617_ ( .A(__set_flag_710_31), .B(1'h0), .S(RST), .Y(_00780_) );
  \$mux  #( .WIDTH(1) ) _47618_ ( .A(__set_flag_710_30), .B(1'h0), .S(RST), .Y(_00779_) );
  \$mux  #( .WIDTH(1) ) _47619_ ( .A(__set_flag_710_29), .B(1'h0), .S(RST), .Y(_00778_) );
  \$mux  #( .WIDTH(1) ) _47620_ ( .A(__set_flag_710_28), .B(1'h0), .S(RST), .Y(_00776_) );
  \$mux  #( .WIDTH(1) ) _47621_ ( .A(__set_flag_710_27), .B(1'h0), .S(RST), .Y(_00775_) );
  \$mux  #( .WIDTH(1) ) _47622_ ( .A(__set_flag_710_26), .B(1'h0), .S(RST), .Y(_00774_) );
  \$mux  #( .WIDTH(1) ) _47623_ ( .A(__set_flag_710_25), .B(1'h0), .S(RST), .Y(_00773_) );
  \$mux  #( .WIDTH(1) ) _47624_ ( .A(__set_flag_710_24), .B(1'h0), .S(RST), .Y(_00772_) );
  \$mux  #( .WIDTH(1) ) _47625_ ( .A(__set_flag_710_23), .B(1'h0), .S(RST), .Y(_00771_) );
  \$mux  #( .WIDTH(1) ) _47626_ ( .A(__set_flag_710_22), .B(1'h0), .S(RST), .Y(_00770_) );
  \$mux  #( .WIDTH(1) ) _47627_ ( .A(__set_flag_710_21), .B(1'h0), .S(RST), .Y(_00769_) );
  \$mux  #( .WIDTH(1) ) _47628_ ( .A(__set_flag_710_20), .B(1'h0), .S(RST), .Y(_00768_) );
  \$mux  #( .WIDTH(1) ) _47629_ ( .A(__set_flag_710_19), .B(1'h0), .S(RST), .Y(_00767_) );
  \$mux  #( .WIDTH(1) ) _47630_ ( .A(__set_flag_710_18), .B(1'h0), .S(RST), .Y(_00765_) );
  \$mux  #( .WIDTH(1) ) _47631_ ( .A(__set_flag_710_17), .B(1'h0), .S(RST), .Y(_00764_) );
  \$mux  #( .WIDTH(1) ) _47632_ ( .A(__set_flag_710_44), .B(1'h0), .S(RST), .Y(_00794_) );
  \$mux  #( .WIDTH(1) ) _47633_ ( .A(__set_flag_710_43), .B(1'h0), .S(RST), .Y(_00793_) );
  \$mux  #( .WIDTH(1) ) _47634_ ( .A(__set_flag_710_38), .B(1'h0), .S(RST), .Y(_00787_) );
  \$mux  #( .WIDTH(1) ) _47635_ ( .A(__set_flag_710_37), .B(1'h0), .S(RST), .Y(_00786_) );
  \$mux  #( .WIDTH(1) ) _47636_ ( .A(__set_flag_710_35), .B(1'h0), .S(RST), .Y(_00784_) );
  \$mux  #( .WIDTH(1) ) _47637_ ( .A(__set_flag_710_33), .B(1'h0), .S(RST), .Y(_00782_) );
  \$mux  #( .WIDTH(1) ) _47638_ ( .A(__set_flag_710_16), .B(1'h0), .S(RST), .Y(_00763_) );
  \$mux  #( .WIDTH(1) ) _47639_ ( .A(__set_flag_710_15), .B(1'h0), .S(RST), .Y(_00762_) );
  \$mux  #( .WIDTH(1) ) _47640_ ( .A(__set_flag_710_14), .B(1'h0), .S(RST), .Y(_00761_) );
  \$mux  #( .WIDTH(1) ) _47641_ ( .A(__set_flag_710_13), .B(1'h0), .S(RST), .Y(_00760_) );
  \$mux  #( .WIDTH(1) ) _47642_ ( .A(__set_flag_710_12), .B(1'h0), .S(RST), .Y(_00759_) );
  \$mux  #( .WIDTH(1) ) _47643_ ( .A(__set_flag_710_11), .B(1'h0), .S(RST), .Y(_00758_) );
  \$mux  #( .WIDTH(1) ) _47644_ ( .A(__set_flag_710_10), .B(1'h0), .S(RST), .Y(_00757_) );
  \$mux  #( .WIDTH(1) ) _47645_ ( .A(__set_flag_710_9), .B(1'h0), .S(RST), .Y(_00756_) );
  \$mux  #( .WIDTH(1) ) _47646_ ( .A(__set_flag_710_8), .B(1'h0), .S(RST), .Y(_00800_) );
  \$mux  #( .WIDTH(1) ) _47647_ ( .A(__set_flag_710_7), .B(1'h0), .S(RST), .Y(_00799_) );
  \$mux  #( .WIDTH(1) ) _47648_ ( .A(__set_flag_710_6), .B(1'h0), .S(RST), .Y(_00798_) );
  \$mux  #( .WIDTH(1) ) _47649_ ( .A(__set_flag_710_5), .B(1'h0), .S(RST), .Y(_00797_) );
  \$mux  #( .WIDTH(1) ) _47650_ ( .A(__set_flag_710_4), .B(1'h0), .S(RST), .Y(_00796_) );
  \$mux  #( .WIDTH(1) ) _47651_ ( .A(__set_flag_710_3), .B(1'h0), .S(RST), .Y(_00795_) );
  \$mux  #( .WIDTH(1) ) _47652_ ( .A(__set_flag_710_2), .B(1'h0), .S(RST), .Y(_00788_) );
  \$mux  #( .WIDTH(1) ) _47653_ ( .A(__set_flag_710_1), .B(1'h0), .S(RST), .Y(_00777_) );
  \$mux  #( .WIDTH(1) ) _47654_ ( .A(_set_flag_710), .B(1'h0), .S(RST), .Y(_00766_) );
  \$mux  #( .WIDTH(33) ) _47655_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_44), .B(33'h000000000), .S(RST), .Y(_00884_) );
  \$mux  #( .WIDTH(33) ) _47656_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_43), .B(33'h000000000), .S(RST), .Y(_00883_) );
  \$mux  #( .WIDTH(33) ) _47657_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_42), .B(33'h000000000), .S(RST), .Y(_00882_) );
  \$mux  #( .WIDTH(33) ) _47658_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_41), .B(33'h000000000), .S(RST), .Y(_00881_) );
  \$mux  #( .WIDTH(33) ) _47659_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_40), .B(33'h000000000), .S(RST), .Y(_00880_) );
  \$mux  #( .WIDTH(33) ) _47660_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_39), .B(33'h000000000), .S(RST), .Y(_00879_) );
  \$mux  #( .WIDTH(33) ) _47661_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_38), .B(33'h000000000), .S(RST), .Y(_00877_) );
  \$mux  #( .WIDTH(33) ) _47662_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_37), .B(33'h000000000), .S(RST), .Y(_00876_) );
  \$mux  #( .WIDTH(33) ) _47663_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_36), .B(33'h000000000), .S(RST), .Y(_00875_) );
  \$mux  #( .WIDTH(33) ) _47664_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_35), .B(33'h000000000), .S(RST), .Y(_00874_) );
  \$mux  #( .WIDTH(33) ) _47665_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_34), .B(33'h000000000), .S(RST), .Y(_00873_) );
  \$mux  #( .WIDTH(33) ) _47666_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_33), .B(33'h000000000), .S(RST), .Y(_00872_) );
  \$mux  #( .WIDTH(33) ) _47667_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_32), .B(33'h000000000), .S(RST), .Y(_00871_) );
  \$mux  #( .WIDTH(33) ) _47668_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_31), .B(33'h000000000), .S(RST), .Y(_00870_) );
  \$mux  #( .WIDTH(33) ) _47669_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_30), .B(33'h000000000), .S(RST), .Y(_00869_) );
  \$mux  #( .WIDTH(33) ) _47670_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_29), .B(33'h000000000), .S(RST), .Y(_00868_) );
  \$mux  #( .WIDTH(33) ) _47671_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_28), .B(33'h000000000), .S(RST), .Y(_00866_) );
  \$mux  #( .WIDTH(33) ) _47672_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_27), .B(33'h000000000), .S(RST), .Y(_00865_) );
  \$mux  #( .WIDTH(33) ) _47673_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_26), .B(33'h000000000), .S(RST), .Y(_00864_) );
  \$mux  #( .WIDTH(33) ) _47674_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_25), .B(33'h000000000), .S(RST), .Y(_00863_) );
  \$mux  #( .WIDTH(33) ) _47675_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_24), .B(33'h000000000), .S(RST), .Y(_00862_) );
  \$mux  #( .WIDTH(33) ) _47676_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_23), .B(33'h000000000), .S(RST), .Y(_00861_) );
  \$mux  #( .WIDTH(33) ) _47677_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_22), .B(33'h000000000), .S(RST), .Y(_00860_) );
  \$mux  #( .WIDTH(33) ) _47678_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_21), .B(33'h000000000), .S(RST), .Y(_00859_) );
  \$mux  #( .WIDTH(33) ) _47679_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_20), .B(33'h000000000), .S(RST), .Y(_00858_) );
  \$mux  #( .WIDTH(33) ) _47680_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_19), .B(33'h000000000), .S(RST), .Y(_00857_) );
  \$mux  #( .WIDTH(33) ) _47681_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_18), .B(33'h000000000), .S(RST), .Y(_00855_) );
  \$mux  #( .WIDTH(33) ) _47682_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_17), .B(33'h000000000), .S(RST), .Y(_00854_) );
  \$mux  #( .WIDTH(33) ) _47683_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_16), .B(33'h000000000), .S(RST), .Y(_00853_) );
  \$mux  #( .WIDTH(33) ) _47684_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_15), .B(33'h000000000), .S(RST), .Y(_00852_) );
  \$mux  #( .WIDTH(33) ) _47685_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_14), .B(33'h000000000), .S(RST), .Y(_00851_) );
  \$mux  #( .WIDTH(33) ) _47686_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_13), .B(33'h000000000), .S(RST), .Y(_00850_) );
  \$mux  #( .WIDTH(33) ) _47687_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_12), .B(33'h000000000), .S(RST), .Y(_00849_) );
  \$mux  #( .WIDTH(33) ) _47688_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_11), .B(33'h000000000), .S(RST), .Y(_00848_) );
  \$mux  #( .WIDTH(33) ) _47689_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_10), .B(33'h000000000), .S(RST), .Y(_00847_) );
  \$mux  #( .WIDTH(33) ) _47690_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_9), .B(33'h000000000), .S(RST), .Y(_00846_) );
  \$mux  #( .WIDTH(33) ) _47691_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_8), .B(33'h000000000), .S(RST), .Y(_00890_) );
  \$mux  #( .WIDTH(33) ) _47692_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_7), .B(33'h000000000), .S(RST), .Y(_00889_) );
  \$mux  #( .WIDTH(33) ) _47693_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_6), .B(33'h000000000), .S(RST), .Y(_00888_) );
  \$mux  #( .WIDTH(33) ) _47694_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_5), .B(33'h000000000), .S(RST), .Y(_00887_) );
  \$mux  #( .WIDTH(33) ) _47695_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_4), .B(33'h000000000), .S(RST), .Y(_00886_) );
  \$mux  #( .WIDTH(33) ) _47696_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_3), .B(33'h000000000), .S(RST), .Y(_00885_) );
  \$mux  #( .WIDTH(33) ) _47697_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_2), .B(33'h000000000), .S(RST), .Y(_00878_) );
  \$mux  #( .WIDTH(33) ) _47698_ ( .A(__stream_conv2d_16_sink_37_sink_size_1_1), .B(33'h000000000), .S(RST), .Y(_00867_) );
  \$mux  #( .WIDTH(33) ) _47699_ ( .A({ 1'h0, conv2d_16_next_stream_num_ops }), .B(33'h000000000), .S(RST), .Y(_00856_) );
  \$mux  #( .WIDTH(32) ) _47700_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_44), .B(0), .S(RST), .Y(_00839_) );
  \$mux  #( .WIDTH(32) ) _47701_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_43), .B(0), .S(RST), .Y(_00838_) );
  \$mux  #( .WIDTH(32) ) _47702_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_42), .B(0), .S(RST), .Y(_00837_) );
  \$mux  #( .WIDTH(32) ) _47703_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_41), .B(0), .S(RST), .Y(_00836_) );
  \$mux  #( .WIDTH(32) ) _47704_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_40), .B(0), .S(RST), .Y(_00835_) );
  \$mux  #( .WIDTH(32) ) _47705_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_39), .B(0), .S(RST), .Y(_00834_) );
  \$mux  #( .WIDTH(32) ) _47706_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_38), .B(0), .S(RST), .Y(_00832_) );
  \$mux  #( .WIDTH(32) ) _47707_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_37), .B(0), .S(RST), .Y(_00831_) );
  \$mux  #( .WIDTH(32) ) _47708_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_36), .B(0), .S(RST), .Y(_00830_) );
  \$mux  #( .WIDTH(32) ) _47709_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_35), .B(0), .S(RST), .Y(_00829_) );
  \$mux  #( .WIDTH(32) ) _47710_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_34), .B(0), .S(RST), .Y(_00828_) );
  \$mux  #( .WIDTH(32) ) _47711_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_33), .B(0), .S(RST), .Y(_00827_) );
  \$mux  #( .WIDTH(32) ) _47712_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_32), .B(0), .S(RST), .Y(_00826_) );
  \$mux  #( .WIDTH(32) ) _47713_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_31), .B(0), .S(RST), .Y(_00825_) );
  \$mux  #( .WIDTH(32) ) _47714_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_30), .B(0), .S(RST), .Y(_00824_) );
  \$mux  #( .WIDTH(32) ) _47715_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_29), .B(0), .S(RST), .Y(_00823_) );
  \$mux  #( .WIDTH(32) ) _47716_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_28), .B(0), .S(RST), .Y(_00821_) );
  \$mux  #( .WIDTH(32) ) _47717_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_27), .B(0), .S(RST), .Y(_00820_) );
  \$mux  #( .WIDTH(32) ) _47718_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_26), .B(0), .S(RST), .Y(_00819_) );
  \$mux  #( .WIDTH(32) ) _47719_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_25), .B(0), .S(RST), .Y(_00818_) );
  \$mux  #( .WIDTH(32) ) _47720_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_24), .B(0), .S(RST), .Y(_00817_) );
  \$mux  #( .WIDTH(32) ) _47721_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_23), .B(0), .S(RST), .Y(_00816_) );
  \$mux  #( .WIDTH(32) ) _47722_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_22), .B(0), .S(RST), .Y(_00815_) );
  \$mux  #( .WIDTH(32) ) _47723_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_21), .B(0), .S(RST), .Y(_00814_) );
  \$mux  #( .WIDTH(32) ) _47724_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_20), .B(0), .S(RST), .Y(_00813_) );
  \$mux  #( .WIDTH(32) ) _47725_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_19), .B(0), .S(RST), .Y(_00812_) );
  \$mux  #( .WIDTH(32) ) _47726_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_18), .B(0), .S(RST), .Y(_00810_) );
  \$mux  #( .WIDTH(32) ) _47727_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_17), .B(0), .S(RST), .Y(_00809_) );
  \$mux  #( .WIDTH(32) ) _47728_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_16), .B(0), .S(RST), .Y(_00808_) );
  \$mux  #( .WIDTH(32) ) _47729_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_15), .B(0), .S(RST), .Y(_00807_) );
  \$mux  #( .WIDTH(32) ) _47730_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_14), .B(0), .S(RST), .Y(_00806_) );
  \$mux  #( .WIDTH(32) ) _47731_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_13), .B(0), .S(RST), .Y(_00805_) );
  \$mux  #( .WIDTH(32) ) _47732_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_12), .B(0), .S(RST), .Y(_00804_) );
  \$mux  #( .WIDTH(32) ) _47733_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_11), .B(0), .S(RST), .Y(_00803_) );
  \$mux  #( .WIDTH(32) ) _47734_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_10), .B(0), .S(RST), .Y(_00802_) );
  \$mux  #( .WIDTH(32) ) _47735_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_9), .B(0), .S(RST), .Y(_00801_) );
  \$mux  #( .WIDTH(32) ) _47736_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_8), .B(0), .S(RST), .Y(_00845_) );
  \$mux  #( .WIDTH(32) ) _47737_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_7), .B(0), .S(RST), .Y(_00844_) );
  \$mux  #( .WIDTH(32) ) _47738_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_6), .B(0), .S(RST), .Y(_00843_) );
  \$mux  #( .WIDTH(32) ) _47739_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_5), .B(0), .S(RST), .Y(_00842_) );
  \$mux  #( .WIDTH(32) ) _47740_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_4), .B(0), .S(RST), .Y(_00841_) );
  \$mux  #( .WIDTH(32) ) _47741_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_3), .B(0), .S(RST), .Y(_00840_) );
  \$mux  #( .WIDTH(32) ) _47742_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_2), .B(0), .S(RST), .Y(_00833_) );
  \$mux  #( .WIDTH(32) ) _47743_ ( .A(__stream_conv2d_16_sink_37_sink_offset_0_1), .B(0), .S(RST), .Y(_00822_) );
  \$mux  #( .WIDTH(32) ) _47744_ ( .A(_24397_), .B(0), .S(RST), .Y(_00811_) );
  \$mux  #( .WIDTH(4) ) _47745_ ( .A(__variable_wdata_510), .B(_stream_conv2d_16_source_36_source_ram_rdata), .S(_stream_conv2d_16_source_36_source_ram_rvalid), .Y(_25409_) );
  \$mux  #( .WIDTH(4) ) _47746_ ( .A(_25409_), .B(4'h0), .S(RST), .Y(_01438_) );
  \$mux  #( .WIDTH(32) ) _47747_ ( .A(_source_stream_conv2d_16_source_36_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_36_pat_stride_3), .S(_06781_), .Y(_25410_) );
  \$mux  #( .WIDTH(32) ) _47748_ ( .A(_25410_), .B(0), .S(RST), .Y(_02315_) );
  \$mux  #( .WIDTH(32) ) _47749_ ( .A(_source_stream_conv2d_16_source_36_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_36_pat_stride_2), .S(_06781_), .Y(_25411_) );
  \$mux  #( .WIDTH(32) ) _47750_ ( .A(_25411_), .B(0), .S(RST), .Y(_02314_) );
  \$mux  #( .WIDTH(32) ) _47751_ ( .A(_source_stream_conv2d_16_source_36_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_36_pat_stride_1), .S(_06781_), .Y(_25412_) );
  \$mux  #( .WIDTH(32) ) _47752_ ( .A(_25412_), .B(0), .S(RST), .Y(_02313_) );
  \$mux  #( .WIDTH(32) ) _47753_ ( .A(_source_stream_conv2d_16_source_36_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_36_pat_stride_0), .S(_06781_), .Y(_25413_) );
  \$mux  #( .WIDTH(32) ) _47754_ ( .A(_25413_), .B(0), .S(RST), .Y(_02312_) );
  \$mux  #( .WIDTH(33) ) _47755_ ( .A(_source_stream_conv2d_16_source_36_pat_size_buf_3), .B(_source_stream_conv2d_16_source_36_pat_size_3), .S(_06781_), .Y(_25414_) );
  \$mux  #( .WIDTH(33) ) _47756_ ( .A(_25414_), .B(33'h000000000), .S(RST), .Y(_02307_) );
  \$mux  #( .WIDTH(33) ) _47757_ ( .A(_source_stream_conv2d_16_source_36_pat_size_buf_2), .B(_source_stream_conv2d_16_source_36_pat_size_2), .S(_06781_), .Y(_25415_) );
  \$mux  #( .WIDTH(33) ) _47758_ ( .A(_25415_), .B(33'h000000000), .S(RST), .Y(_02306_) );
  \$mux  #( .WIDTH(33) ) _47759_ ( .A(_source_stream_conv2d_16_source_36_pat_size_buf_1), .B(_source_stream_conv2d_16_source_36_pat_size_1), .S(_06781_), .Y(_25416_) );
  \$mux  #( .WIDTH(33) ) _47760_ ( .A(_25416_), .B(33'h000000000), .S(RST), .Y(_02305_) );
  \$mux  #( .WIDTH(33) ) _47761_ ( .A(_source_stream_conv2d_16_source_36_pat_size_buf_0), .B(_source_stream_conv2d_16_source_36_pat_size_0), .S(_06781_), .Y(_25417_) );
  \$mux  #( .WIDTH(33) ) _47762_ ( .A(_25417_), .B(33'h000000000), .S(RST), .Y(_02304_) );
  \$mux  #( .WIDTH(33) ) _47763_ ( .A(_source_stream_conv2d_16_source_36_pat_count_3), .B(_28859_), .S(_06781_), .Y(_25418_) );
  \$mux  #( .WIDTH(33) ) _47764_ ( .A(_25418_), .B(_28866_), .S(_06784_), .Y(_25419_) );
  \$mux  #( .WIDTH(33) ) _47765_ ( .A(_25419_), .B(_28867_), .S(_06785_), .Y(_25420_) );
  \$mux  #( .WIDTH(33) ) _47766_ ( .A(_25420_), .B(33'h000000000), .S(RST), .Y(_02295_) );
  \$mux  #( .WIDTH(33) ) _47767_ ( .A(_source_stream_conv2d_16_source_36_pat_count_2), .B(_28858_), .S(_06781_), .Y(_25421_) );
  \$mux  #( .WIDTH(33) ) _47768_ ( .A(_25421_), .B(_28864_), .S(_06783_), .Y(_25422_) );
  \$mux  #( .WIDTH(33) ) _47769_ ( .A(_25422_), .B(_28865_), .S(_06784_), .Y(_25423_) );
  \$mux  #( .WIDTH(33) ) _47770_ ( .A(_25423_), .B(33'h000000000), .S(RST), .Y(_02294_) );
  \$mux  #( .WIDTH(33) ) _47771_ ( .A(_source_stream_conv2d_16_source_36_pat_count_1), .B(_28857_), .S(_06781_), .Y(_25424_) );
  \$mux  #( .WIDTH(33) ) _47772_ ( .A(_25424_), .B(_28862_), .S(_06782_), .Y(_25425_) );
  \$mux  #( .WIDTH(33) ) _47773_ ( .A(_25425_), .B(_28863_), .S(_06783_), .Y(_25426_) );
  \$mux  #( .WIDTH(33) ) _47774_ ( .A(_25426_), .B(33'h000000000), .S(RST), .Y(_02293_) );
  \$mux  #( .WIDTH(33) ) _47775_ ( .A(_source_stream_conv2d_16_source_36_pat_count_0), .B(_28856_), .S(_06781_), .Y(_25427_) );
  \$mux  #( .WIDTH(33) ) _47776_ ( .A(_28860_), .B(_25427_), .S(_05949_), .Y(_25428_) );
  \$mux  #( .WIDTH(33) ) _47777_ ( .A(_25428_), .B(_28861_), .S(_06782_), .Y(_25429_) );
  \$mux  #( .WIDTH(33) ) _47778_ ( .A(_25429_), .B(33'h000000000), .S(RST), .Y(_02292_) );
  \$mux  #( .WIDTH(32) ) _47779_ ( .A(_source_stream_conv2d_16_source_36_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25430_) );
  \$mux  #( .WIDTH(32) ) _47780_ ( .A(_25430_), .B(0), .S(RST), .Y(_02311_) );
  \$mux  #( .WIDTH(32) ) _47781_ ( .A(_source_stream_conv2d_16_source_36_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25431_) );
  \$mux  #( .WIDTH(32) ) _47782_ ( .A(_25431_), .B(0), .S(RST), .Y(_02310_) );
  \$mux  #( .WIDTH(32) ) _47783_ ( .A(_source_stream_conv2d_16_source_36_pat_stride_1), .B({ 26'h0000000, cparam_conv2d_16_filter_read_block }), .S(_set_flag_710), .Y(_25432_) );
  \$mux  #( .WIDTH(32) ) _47784_ ( .A(_25432_), .B(0), .S(RST), .Y(_02309_) );
  \$mux  #( .WIDTH(32) ) _47785_ ( .A(_source_stream_conv2d_16_source_36_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25433_) );
  \$mux  #( .WIDTH(32) ) _47786_ ( .A(_25433_), .B(0), .S(RST), .Y(_02308_) );
  \$mux  #( .WIDTH(33) ) _47787_ ( .A(_source_stream_conv2d_16_source_36_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25434_) );
  \$mux  #( .WIDTH(33) ) _47788_ ( .A(_25434_), .B(33'h000000000), .S(RST), .Y(_02303_) );
  \$mux  #( .WIDTH(33) ) _47789_ ( .A(_source_stream_conv2d_16_source_36_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25435_) );
  \$mux  #( .WIDTH(33) ) _47790_ ( .A(_25435_), .B(33'h000000000), .S(RST), .Y(_02302_) );
  \$mux  #( .WIDTH(33) ) _47791_ ( .A(_source_stream_conv2d_16_source_36_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25436_) );
  \$mux  #( .WIDTH(33) ) _47792_ ( .A(_25436_), .B(33'h000000000), .S(RST), .Y(_02301_) );
  \$mux  #( .WIDTH(33) ) _47793_ ( .A(_source_stream_conv2d_16_source_36_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25437_) );
  \$mux  #( .WIDTH(33) ) _47794_ ( .A(_25437_), .B(33'h000000000), .S(RST), .Y(_02300_) );
  \$mux  #( .WIDTH(32) ) _47795_ ( .A(_source_stream_conv2d_16_source_36_pat_cur_offset_3), .B(0), .S(_06781_), .Y(_25438_) );
  \$mux  #( .WIDTH(32) ) _47796_ ( .A(_25438_), .B(_24396_), .S(_06784_), .Y(_25439_) );
  \$mux  #( .WIDTH(32) ) _47797_ ( .A(_25439_), .B(0), .S(_06785_), .Y(_25440_) );
  \$mux  #( .WIDTH(32) ) _47798_ ( .A(_25440_), .B(0), .S(RST), .Y(_02299_) );
  \$mux  #( .WIDTH(32) ) _47799_ ( .A(_source_stream_conv2d_16_source_36_pat_cur_offset_2), .B(0), .S(_06781_), .Y(_25441_) );
  \$mux  #( .WIDTH(32) ) _47800_ ( .A(_25441_), .B(_24395_), .S(_06783_), .Y(_25442_) );
  \$mux  #( .WIDTH(32) ) _47801_ ( .A(_25442_), .B(0), .S(_06784_), .Y(_25443_) );
  \$mux  #( .WIDTH(32) ) _47802_ ( .A(_25443_), .B(0), .S(RST), .Y(_02298_) );
  \$mux  #( .WIDTH(32) ) _47803_ ( .A(_source_stream_conv2d_16_source_36_pat_cur_offset_1), .B(0), .S(_06781_), .Y(_25444_) );
  \$mux  #( .WIDTH(32) ) _47804_ ( .A(_25444_), .B(_24394_), .S(_06782_), .Y(_25445_) );
  \$mux  #( .WIDTH(32) ) _47805_ ( .A(_25445_), .B(0), .S(_06783_), .Y(_25446_) );
  \$mux  #( .WIDTH(32) ) _47806_ ( .A(_25446_), .B(0), .S(RST), .Y(_02297_) );
  \$mux  #( .WIDTH(32) ) _47807_ ( .A(_source_stream_conv2d_16_source_36_pat_cur_offset_0), .B(0), .S(_06781_), .Y(_25447_) );
  \$mux  #( .WIDTH(32) ) _47808_ ( .A(_24393_), .B(_25447_), .S(_05949_), .Y(_25448_) );
  \$mux  #( .WIDTH(32) ) _47809_ ( .A(_25448_), .B(0), .S(_06782_), .Y(_25449_) );
  \$mux  #( .WIDTH(32) ) _47810_ ( .A(_25449_), .B(0), .S(RST), .Y(_02296_) );
  \$mux  #( .WIDTH(4) ) _47811_ ( .A(__variable_wdata_509), .B(_stream_conv2d_16_source_35_source_ram_rdata), .S(_stream_conv2d_16_source_35_source_ram_rvalid), .Y(_25450_) );
  \$mux  #( .WIDTH(4) ) _47812_ ( .A(_25450_), .B(4'h0), .S(RST), .Y(_01437_) );
  \$mux  #( .WIDTH(32) ) _47813_ ( .A(_source_stream_conv2d_16_source_35_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_35_pat_stride_3), .S(_06776_), .Y(_25451_) );
  \$mux  #( .WIDTH(32) ) _47814_ ( .A(_25451_), .B(0), .S(RST), .Y(_02291_) );
  \$mux  #( .WIDTH(32) ) _47815_ ( .A(_source_stream_conv2d_16_source_35_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_35_pat_stride_2), .S(_06776_), .Y(_25452_) );
  \$mux  #( .WIDTH(32) ) _47816_ ( .A(_25452_), .B(0), .S(RST), .Y(_02290_) );
  \$mux  #( .WIDTH(32) ) _47817_ ( .A(_source_stream_conv2d_16_source_35_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_35_pat_stride_1), .S(_06776_), .Y(_25453_) );
  \$mux  #( .WIDTH(32) ) _47818_ ( .A(_25453_), .B(0), .S(RST), .Y(_02289_) );
  \$mux  #( .WIDTH(32) ) _47819_ ( .A(_source_stream_conv2d_16_source_35_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_35_pat_stride_0), .S(_06776_), .Y(_25454_) );
  \$mux  #( .WIDTH(32) ) _47820_ ( .A(_25454_), .B(0), .S(RST), .Y(_02288_) );
  \$mux  #( .WIDTH(33) ) _47821_ ( .A(_source_stream_conv2d_16_source_35_pat_size_buf_3), .B(_source_stream_conv2d_16_source_35_pat_size_3), .S(_06776_), .Y(_25455_) );
  \$mux  #( .WIDTH(33) ) _47822_ ( .A(_25455_), .B(33'h000000000), .S(RST), .Y(_02283_) );
  \$mux  #( .WIDTH(33) ) _47823_ ( .A(_source_stream_conv2d_16_source_35_pat_size_buf_2), .B(_source_stream_conv2d_16_source_35_pat_size_2), .S(_06776_), .Y(_25456_) );
  \$mux  #( .WIDTH(33) ) _47824_ ( .A(_25456_), .B(33'h000000000), .S(RST), .Y(_02282_) );
  \$mux  #( .WIDTH(33) ) _47825_ ( .A(_source_stream_conv2d_16_source_35_pat_size_buf_1), .B(_source_stream_conv2d_16_source_35_pat_size_1), .S(_06776_), .Y(_25457_) );
  \$mux  #( .WIDTH(33) ) _47826_ ( .A(_25457_), .B(33'h000000000), .S(RST), .Y(_02281_) );
  \$mux  #( .WIDTH(33) ) _47827_ ( .A(_source_stream_conv2d_16_source_35_pat_size_buf_0), .B(_source_stream_conv2d_16_source_35_pat_size_0), .S(_06776_), .Y(_25458_) );
  \$mux  #( .WIDTH(33) ) _47828_ ( .A(_25458_), .B(33'h000000000), .S(RST), .Y(_02280_) );
  \$mux  #( .WIDTH(33) ) _47829_ ( .A(_source_stream_conv2d_16_source_35_pat_count_3), .B(_28847_), .S(_06776_), .Y(_25459_) );
  \$mux  #( .WIDTH(33) ) _47830_ ( .A(_25459_), .B(_28854_), .S(_06779_), .Y(_25460_) );
  \$mux  #( .WIDTH(33) ) _47831_ ( .A(_25460_), .B(_28855_), .S(_06780_), .Y(_25461_) );
  \$mux  #( .WIDTH(33) ) _47832_ ( .A(_25461_), .B(33'h000000000), .S(RST), .Y(_02271_) );
  \$mux  #( .WIDTH(33) ) _47833_ ( .A(_source_stream_conv2d_16_source_35_pat_count_2), .B(_28846_), .S(_06776_), .Y(_25462_) );
  \$mux  #( .WIDTH(33) ) _47834_ ( .A(_25462_), .B(_28852_), .S(_06778_), .Y(_25463_) );
  \$mux  #( .WIDTH(33) ) _47835_ ( .A(_25463_), .B(_28853_), .S(_06779_), .Y(_25464_) );
  \$mux  #( .WIDTH(33) ) _47836_ ( .A(_25464_), .B(33'h000000000), .S(RST), .Y(_02270_) );
  \$mux  #( .WIDTH(33) ) _47837_ ( .A(_source_stream_conv2d_16_source_35_pat_count_1), .B(_28845_), .S(_06776_), .Y(_25465_) );
  \$mux  #( .WIDTH(33) ) _47838_ ( .A(_25465_), .B(_28850_), .S(_06777_), .Y(_25466_) );
  \$mux  #( .WIDTH(33) ) _47839_ ( .A(_25466_), .B(_28851_), .S(_06778_), .Y(_25467_) );
  \$mux  #( .WIDTH(33) ) _47840_ ( .A(_25467_), .B(33'h000000000), .S(RST), .Y(_02269_) );
  \$mux  #( .WIDTH(33) ) _47841_ ( .A(_source_stream_conv2d_16_source_35_pat_count_0), .B(_28844_), .S(_06776_), .Y(_25468_) );
  \$mux  #( .WIDTH(33) ) _47842_ ( .A(_28848_), .B(_25468_), .S(_05952_), .Y(_25469_) );
  \$mux  #( .WIDTH(33) ) _47843_ ( .A(_25469_), .B(_28849_), .S(_06777_), .Y(_25470_) );
  \$mux  #( .WIDTH(33) ) _47844_ ( .A(_25470_), .B(33'h000000000), .S(RST), .Y(_02268_) );
  \$mux  #( .WIDTH(32) ) _47845_ ( .A(_source_stream_conv2d_16_source_35_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25471_) );
  \$mux  #( .WIDTH(32) ) _47846_ ( .A(_25471_), .B(0), .S(RST), .Y(_02287_) );
  \$mux  #( .WIDTH(32) ) _47847_ ( .A(_source_stream_conv2d_16_source_35_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25472_) );
  \$mux  #( .WIDTH(32) ) _47848_ ( .A(_25472_), .B(0), .S(RST), .Y(_02286_) );
  \$mux  #( .WIDTH(32) ) _47849_ ( .A(_source_stream_conv2d_16_source_35_pat_stride_1), .B({ 26'h0000000, cparam_conv2d_16_filter_read_block }), .S(_set_flag_710), .Y(_25473_) );
  \$mux  #( .WIDTH(32) ) _47850_ ( .A(_25473_), .B(0), .S(RST), .Y(_02285_) );
  \$mux  #( .WIDTH(32) ) _47851_ ( .A(_source_stream_conv2d_16_source_35_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25474_) );
  \$mux  #( .WIDTH(32) ) _47852_ ( .A(_25474_), .B(0), .S(RST), .Y(_02284_) );
  \$mux  #( .WIDTH(33) ) _47853_ ( .A(_source_stream_conv2d_16_source_35_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25475_) );
  \$mux  #( .WIDTH(33) ) _47854_ ( .A(_25475_), .B(33'h000000000), .S(RST), .Y(_02279_) );
  \$mux  #( .WIDTH(33) ) _47855_ ( .A(_source_stream_conv2d_16_source_35_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25476_) );
  \$mux  #( .WIDTH(33) ) _47856_ ( .A(_25476_), .B(33'h000000000), .S(RST), .Y(_02278_) );
  \$mux  #( .WIDTH(33) ) _47857_ ( .A(_source_stream_conv2d_16_source_35_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25477_) );
  \$mux  #( .WIDTH(33) ) _47858_ ( .A(_25477_), .B(33'h000000000), .S(RST), .Y(_02277_) );
  \$mux  #( .WIDTH(33) ) _47859_ ( .A(_source_stream_conv2d_16_source_35_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25478_) );
  \$mux  #( .WIDTH(33) ) _47860_ ( .A(_25478_), .B(33'h000000000), .S(RST), .Y(_02276_) );
  \$mux  #( .WIDTH(32) ) _47861_ ( .A(_source_stream_conv2d_16_source_35_pat_cur_offset_3), .B(0), .S(_06776_), .Y(_25479_) );
  \$mux  #( .WIDTH(32) ) _47862_ ( .A(_25479_), .B(_24392_), .S(_06779_), .Y(_25480_) );
  \$mux  #( .WIDTH(32) ) _47863_ ( .A(_25480_), .B(0), .S(_06780_), .Y(_25481_) );
  \$mux  #( .WIDTH(32) ) _47864_ ( .A(_25481_), .B(0), .S(RST), .Y(_02275_) );
  \$mux  #( .WIDTH(32) ) _47865_ ( .A(_source_stream_conv2d_16_source_35_pat_cur_offset_2), .B(0), .S(_06776_), .Y(_25482_) );
  \$mux  #( .WIDTH(32) ) _47866_ ( .A(_25482_), .B(_24391_), .S(_06778_), .Y(_25483_) );
  \$mux  #( .WIDTH(32) ) _47867_ ( .A(_25483_), .B(0), .S(_06779_), .Y(_25484_) );
  \$mux  #( .WIDTH(32) ) _47868_ ( .A(_25484_), .B(0), .S(RST), .Y(_02274_) );
  \$mux  #( .WIDTH(32) ) _47869_ ( .A(_source_stream_conv2d_16_source_35_pat_cur_offset_1), .B(0), .S(_06776_), .Y(_25485_) );
  \$mux  #( .WIDTH(32) ) _47870_ ( .A(_25485_), .B(_24390_), .S(_06777_), .Y(_25486_) );
  \$mux  #( .WIDTH(32) ) _47871_ ( .A(_25486_), .B(0), .S(_06778_), .Y(_25487_) );
  \$mux  #( .WIDTH(32) ) _47872_ ( .A(_25487_), .B(0), .S(RST), .Y(_02273_) );
  \$mux  #( .WIDTH(32) ) _47873_ ( .A(_source_stream_conv2d_16_source_35_pat_cur_offset_0), .B(0), .S(_06776_), .Y(_25488_) );
  \$mux  #( .WIDTH(32) ) _47874_ ( .A(_24389_), .B(_25488_), .S(_05952_), .Y(_25489_) );
  \$mux  #( .WIDTH(32) ) _47875_ ( .A(_25489_), .B(0), .S(_06777_), .Y(_25490_) );
  \$mux  #( .WIDTH(32) ) _47876_ ( .A(_25490_), .B(0), .S(RST), .Y(_02272_) );
  \$mux  #( .WIDTH(4) ) _47877_ ( .A(__variable_wdata_508), .B(_stream_conv2d_16_source_34_source_ram_rdata), .S(_stream_conv2d_16_source_34_source_ram_rvalid), .Y(_25491_) );
  \$mux  #( .WIDTH(4) ) _47878_ ( .A(_25491_), .B(4'h0), .S(RST), .Y(_01436_) );
  \$mux  #( .WIDTH(32) ) _47879_ ( .A(_source_stream_conv2d_16_source_34_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_34_pat_stride_3), .S(_06771_), .Y(_25492_) );
  \$mux  #( .WIDTH(32) ) _47880_ ( .A(_25492_), .B(0), .S(RST), .Y(_02267_) );
  \$mux  #( .WIDTH(32) ) _47881_ ( .A(_source_stream_conv2d_16_source_34_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_34_pat_stride_2), .S(_06771_), .Y(_25493_) );
  \$mux  #( .WIDTH(32) ) _47882_ ( .A(_25493_), .B(0), .S(RST), .Y(_02266_) );
  \$mux  #( .WIDTH(32) ) _47883_ ( .A(_source_stream_conv2d_16_source_34_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_34_pat_stride_1), .S(_06771_), .Y(_25494_) );
  \$mux  #( .WIDTH(32) ) _47884_ ( .A(_25494_), .B(0), .S(RST), .Y(_02265_) );
  \$mux  #( .WIDTH(32) ) _47885_ ( .A(_source_stream_conv2d_16_source_34_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_34_pat_stride_0), .S(_06771_), .Y(_25495_) );
  \$mux  #( .WIDTH(32) ) _47886_ ( .A(_25495_), .B(0), .S(RST), .Y(_02264_) );
  \$mux  #( .WIDTH(33) ) _47887_ ( .A(_source_stream_conv2d_16_source_34_pat_size_buf_3), .B(_source_stream_conv2d_16_source_34_pat_size_3), .S(_06771_), .Y(_25496_) );
  \$mux  #( .WIDTH(33) ) _47888_ ( .A(_25496_), .B(33'h000000000), .S(RST), .Y(_02259_) );
  \$mux  #( .WIDTH(33) ) _47889_ ( .A(_source_stream_conv2d_16_source_34_pat_size_buf_2), .B(_source_stream_conv2d_16_source_34_pat_size_2), .S(_06771_), .Y(_25497_) );
  \$mux  #( .WIDTH(33) ) _47890_ ( .A(_25497_), .B(33'h000000000), .S(RST), .Y(_02258_) );
  \$mux  #( .WIDTH(33) ) _47891_ ( .A(_source_stream_conv2d_16_source_34_pat_size_buf_1), .B(_source_stream_conv2d_16_source_34_pat_size_1), .S(_06771_), .Y(_25498_) );
  \$mux  #( .WIDTH(33) ) _47892_ ( .A(_25498_), .B(33'h000000000), .S(RST), .Y(_02257_) );
  \$mux  #( .WIDTH(33) ) _47893_ ( .A(_source_stream_conv2d_16_source_34_pat_size_buf_0), .B(_source_stream_conv2d_16_source_34_pat_size_0), .S(_06771_), .Y(_25499_) );
  \$mux  #( .WIDTH(33) ) _47894_ ( .A(_25499_), .B(33'h000000000), .S(RST), .Y(_02256_) );
  \$mux  #( .WIDTH(33) ) _47895_ ( .A(_source_stream_conv2d_16_source_34_pat_count_3), .B(_28835_), .S(_06771_), .Y(_25500_) );
  \$mux  #( .WIDTH(33) ) _47896_ ( .A(_25500_), .B(_28842_), .S(_06774_), .Y(_25501_) );
  \$mux  #( .WIDTH(33) ) _47897_ ( .A(_25501_), .B(_28843_), .S(_06775_), .Y(_25502_) );
  \$mux  #( .WIDTH(33) ) _47898_ ( .A(_25502_), .B(33'h000000000), .S(RST), .Y(_02247_) );
  \$mux  #( .WIDTH(33) ) _47899_ ( .A(_source_stream_conv2d_16_source_34_pat_count_2), .B(_28834_), .S(_06771_), .Y(_25503_) );
  \$mux  #( .WIDTH(33) ) _47900_ ( .A(_25503_), .B(_28840_), .S(_06773_), .Y(_25504_) );
  \$mux  #( .WIDTH(33) ) _47901_ ( .A(_25504_), .B(_28841_), .S(_06774_), .Y(_25505_) );
  \$mux  #( .WIDTH(33) ) _47902_ ( .A(_25505_), .B(33'h000000000), .S(RST), .Y(_02246_) );
  \$mux  #( .WIDTH(33) ) _47903_ ( .A(_source_stream_conv2d_16_source_34_pat_count_1), .B(_28833_), .S(_06771_), .Y(_25506_) );
  \$mux  #( .WIDTH(33) ) _47904_ ( .A(_25506_), .B(_28838_), .S(_06772_), .Y(_25507_) );
  \$mux  #( .WIDTH(33) ) _47905_ ( .A(_25507_), .B(_28839_), .S(_06773_), .Y(_25508_) );
  \$mux  #( .WIDTH(33) ) _47906_ ( .A(_25508_), .B(33'h000000000), .S(RST), .Y(_02245_) );
  \$mux  #( .WIDTH(33) ) _47907_ ( .A(_source_stream_conv2d_16_source_34_pat_count_0), .B(_28832_), .S(_06771_), .Y(_25509_) );
  \$mux  #( .WIDTH(33) ) _47908_ ( .A(_28836_), .B(_25509_), .S(_05954_), .Y(_25510_) );
  \$mux  #( .WIDTH(33) ) _47909_ ( .A(_25510_), .B(_28837_), .S(_06772_), .Y(_25511_) );
  \$mux  #( .WIDTH(33) ) _47910_ ( .A(_25511_), .B(33'h000000000), .S(RST), .Y(_02244_) );
  \$mux  #( .WIDTH(32) ) _47911_ ( .A(_source_stream_conv2d_16_source_34_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25512_) );
  \$mux  #( .WIDTH(32) ) _47912_ ( .A(_25512_), .B(0), .S(RST), .Y(_02263_) );
  \$mux  #( .WIDTH(32) ) _47913_ ( .A(_source_stream_conv2d_16_source_34_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25513_) );
  \$mux  #( .WIDTH(32) ) _47914_ ( .A(_25513_), .B(0), .S(RST), .Y(_02262_) );
  \$mux  #( .WIDTH(32) ) _47915_ ( .A(_source_stream_conv2d_16_source_34_pat_stride_1), .B({ 26'h0000000, cparam_conv2d_16_filter_read_block }), .S(_set_flag_710), .Y(_25514_) );
  \$mux  #( .WIDTH(32) ) _47916_ ( .A(_25514_), .B(0), .S(RST), .Y(_02261_) );
  \$mux  #( .WIDTH(32) ) _47917_ ( .A(_source_stream_conv2d_16_source_34_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25515_) );
  \$mux  #( .WIDTH(32) ) _47918_ ( .A(_25515_), .B(0), .S(RST), .Y(_02260_) );
  \$mux  #( .WIDTH(33) ) _47919_ ( .A(_source_stream_conv2d_16_source_34_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25516_) );
  \$mux  #( .WIDTH(33) ) _47920_ ( .A(_25516_), .B(33'h000000000), .S(RST), .Y(_02255_) );
  \$mux  #( .WIDTH(33) ) _47921_ ( .A(_source_stream_conv2d_16_source_34_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25517_) );
  \$mux  #( .WIDTH(33) ) _47922_ ( .A(_25517_), .B(33'h000000000), .S(RST), .Y(_02254_) );
  \$mux  #( .WIDTH(33) ) _47923_ ( .A(_source_stream_conv2d_16_source_34_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25518_) );
  \$mux  #( .WIDTH(33) ) _47924_ ( .A(_25518_), .B(33'h000000000), .S(RST), .Y(_02253_) );
  \$mux  #( .WIDTH(33) ) _47925_ ( .A(_source_stream_conv2d_16_source_34_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25519_) );
  \$mux  #( .WIDTH(33) ) _47926_ ( .A(_25519_), .B(33'h000000000), .S(RST), .Y(_02252_) );
  \$mux  #( .WIDTH(32) ) _47927_ ( .A(_source_stream_conv2d_16_source_34_pat_cur_offset_3), .B(0), .S(_06771_), .Y(_25520_) );
  \$mux  #( .WIDTH(32) ) _47928_ ( .A(_25520_), .B(_24388_), .S(_06774_), .Y(_25521_) );
  \$mux  #( .WIDTH(32) ) _47929_ ( .A(_25521_), .B(0), .S(_06775_), .Y(_25522_) );
  \$mux  #( .WIDTH(32) ) _47930_ ( .A(_25522_), .B(0), .S(RST), .Y(_02251_) );
  \$mux  #( .WIDTH(32) ) _47931_ ( .A(_source_stream_conv2d_16_source_34_pat_cur_offset_2), .B(0), .S(_06771_), .Y(_25523_) );
  \$mux  #( .WIDTH(32) ) _47932_ ( .A(_25523_), .B(_24387_), .S(_06773_), .Y(_25524_) );
  \$mux  #( .WIDTH(32) ) _47933_ ( .A(_25524_), .B(0), .S(_06774_), .Y(_25525_) );
  \$mux  #( .WIDTH(32) ) _47934_ ( .A(_25525_), .B(0), .S(RST), .Y(_02250_) );
  \$mux  #( .WIDTH(32) ) _47935_ ( .A(_source_stream_conv2d_16_source_34_pat_cur_offset_1), .B(0), .S(_06771_), .Y(_25526_) );
  \$mux  #( .WIDTH(32) ) _47936_ ( .A(_25526_), .B(_24386_), .S(_06772_), .Y(_25527_) );
  \$mux  #( .WIDTH(32) ) _47937_ ( .A(_25527_), .B(0), .S(_06773_), .Y(_25528_) );
  \$mux  #( .WIDTH(32) ) _47938_ ( .A(_25528_), .B(0), .S(RST), .Y(_02249_) );
  \$mux  #( .WIDTH(32) ) _47939_ ( .A(_source_stream_conv2d_16_source_34_pat_cur_offset_0), .B(0), .S(_06771_), .Y(_25529_) );
  \$mux  #( .WIDTH(32) ) _47940_ ( .A(_24385_), .B(_25529_), .S(_05954_), .Y(_25530_) );
  \$mux  #( .WIDTH(32) ) _47941_ ( .A(_25530_), .B(0), .S(_06772_), .Y(_25531_) );
  \$mux  #( .WIDTH(32) ) _47942_ ( .A(_25531_), .B(0), .S(RST), .Y(_02248_) );
  \$mux  #( .WIDTH(4) ) _47943_ ( .A(__variable_wdata_507), .B(_stream_conv2d_16_source_33_source_ram_rdata), .S(_stream_conv2d_16_source_33_source_ram_rvalid), .Y(_25532_) );
  \$mux  #( .WIDTH(4) ) _47944_ ( .A(_25532_), .B(4'h0), .S(RST), .Y(_01435_) );
  \$mux  #( .WIDTH(32) ) _47945_ ( .A(_source_stream_conv2d_16_source_33_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_33_pat_stride_3), .S(_06766_), .Y(_25533_) );
  \$mux  #( .WIDTH(32) ) _47946_ ( .A(_25533_), .B(0), .S(RST), .Y(_02243_) );
  \$mux  #( .WIDTH(32) ) _47947_ ( .A(_source_stream_conv2d_16_source_33_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_33_pat_stride_2), .S(_06766_), .Y(_25534_) );
  \$mux  #( .WIDTH(32) ) _47948_ ( .A(_25534_), .B(0), .S(RST), .Y(_02242_) );
  \$mux  #( .WIDTH(32) ) _47949_ ( .A(_source_stream_conv2d_16_source_33_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_33_pat_stride_1), .S(_06766_), .Y(_25535_) );
  \$mux  #( .WIDTH(32) ) _47950_ ( .A(_25535_), .B(0), .S(RST), .Y(_02241_) );
  \$mux  #( .WIDTH(32) ) _47951_ ( .A(_source_stream_conv2d_16_source_33_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_33_pat_stride_0), .S(_06766_), .Y(_25536_) );
  \$mux  #( .WIDTH(32) ) _47952_ ( .A(_25536_), .B(0), .S(RST), .Y(_02240_) );
  \$mux  #( .WIDTH(33) ) _47953_ ( .A(_source_stream_conv2d_16_source_33_pat_size_buf_3), .B(_source_stream_conv2d_16_source_33_pat_size_3), .S(_06766_), .Y(_25537_) );
  \$mux  #( .WIDTH(33) ) _47954_ ( .A(_25537_), .B(33'h000000000), .S(RST), .Y(_02235_) );
  \$mux  #( .WIDTH(33) ) _47955_ ( .A(_source_stream_conv2d_16_source_33_pat_size_buf_2), .B(_source_stream_conv2d_16_source_33_pat_size_2), .S(_06766_), .Y(_25538_) );
  \$mux  #( .WIDTH(33) ) _47956_ ( .A(_25538_), .B(33'h000000000), .S(RST), .Y(_02234_) );
  \$mux  #( .WIDTH(33) ) _47957_ ( .A(_source_stream_conv2d_16_source_33_pat_size_buf_1), .B(_source_stream_conv2d_16_source_33_pat_size_1), .S(_06766_), .Y(_25539_) );
  \$mux  #( .WIDTH(33) ) _47958_ ( .A(_25539_), .B(33'h000000000), .S(RST), .Y(_02233_) );
  \$mux  #( .WIDTH(33) ) _47959_ ( .A(_source_stream_conv2d_16_source_33_pat_size_buf_0), .B(_source_stream_conv2d_16_source_33_pat_size_0), .S(_06766_), .Y(_25540_) );
  \$mux  #( .WIDTH(33) ) _47960_ ( .A(_25540_), .B(33'h000000000), .S(RST), .Y(_02232_) );
  \$mux  #( .WIDTH(33) ) _47961_ ( .A(_source_stream_conv2d_16_source_33_pat_count_3), .B(_28823_), .S(_06766_), .Y(_25541_) );
  \$mux  #( .WIDTH(33) ) _47962_ ( .A(_25541_), .B(_28830_), .S(_06769_), .Y(_25542_) );
  \$mux  #( .WIDTH(33) ) _47963_ ( .A(_25542_), .B(_28831_), .S(_06770_), .Y(_25543_) );
  \$mux  #( .WIDTH(33) ) _47964_ ( .A(_25543_), .B(33'h000000000), .S(RST), .Y(_02223_) );
  \$mux  #( .WIDTH(33) ) _47965_ ( .A(_source_stream_conv2d_16_source_33_pat_count_2), .B(_28822_), .S(_06766_), .Y(_25544_) );
  \$mux  #( .WIDTH(33) ) _47966_ ( .A(_25544_), .B(_28828_), .S(_06768_), .Y(_25545_) );
  \$mux  #( .WIDTH(33) ) _47967_ ( .A(_25545_), .B(_28829_), .S(_06769_), .Y(_25546_) );
  \$mux  #( .WIDTH(33) ) _47968_ ( .A(_25546_), .B(33'h000000000), .S(RST), .Y(_02222_) );
  \$mux  #( .WIDTH(33) ) _47969_ ( .A(_source_stream_conv2d_16_source_33_pat_count_1), .B(_28821_), .S(_06766_), .Y(_25547_) );
  \$mux  #( .WIDTH(33) ) _47970_ ( .A(_25547_), .B(_28826_), .S(_06767_), .Y(_25548_) );
  \$mux  #( .WIDTH(33) ) _47971_ ( .A(_25548_), .B(_28827_), .S(_06768_), .Y(_25549_) );
  \$mux  #( .WIDTH(33) ) _47972_ ( .A(_25549_), .B(33'h000000000), .S(RST), .Y(_02221_) );
  \$mux  #( .WIDTH(33) ) _47973_ ( .A(_source_stream_conv2d_16_source_33_pat_count_0), .B(_28820_), .S(_06766_), .Y(_25550_) );
  \$mux  #( .WIDTH(33) ) _47974_ ( .A(_28824_), .B(_25550_), .S(_05956_), .Y(_25551_) );
  \$mux  #( .WIDTH(33) ) _47975_ ( .A(_25551_), .B(_28825_), .S(_06767_), .Y(_25552_) );
  \$mux  #( .WIDTH(33) ) _47976_ ( .A(_25552_), .B(33'h000000000), .S(RST), .Y(_02220_) );
  \$mux  #( .WIDTH(32) ) _47977_ ( .A(_source_stream_conv2d_16_source_33_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25553_) );
  \$mux  #( .WIDTH(32) ) _47978_ ( .A(_25553_), .B(0), .S(RST), .Y(_02239_) );
  \$mux  #( .WIDTH(32) ) _47979_ ( .A(_source_stream_conv2d_16_source_33_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25554_) );
  \$mux  #( .WIDTH(32) ) _47980_ ( .A(_25554_), .B(0), .S(RST), .Y(_02238_) );
  \$mux  #( .WIDTH(32) ) _47981_ ( .A(_source_stream_conv2d_16_source_33_pat_stride_1), .B({ 26'h0000000, cparam_conv2d_16_filter_read_block }), .S(_set_flag_710), .Y(_25555_) );
  \$mux  #( .WIDTH(32) ) _47982_ ( .A(_25555_), .B(0), .S(RST), .Y(_02237_) );
  \$mux  #( .WIDTH(32) ) _47983_ ( .A(_source_stream_conv2d_16_source_33_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25556_) );
  \$mux  #( .WIDTH(32) ) _47984_ ( .A(_25556_), .B(0), .S(RST), .Y(_02236_) );
  \$mux  #( .WIDTH(33) ) _47985_ ( .A(_source_stream_conv2d_16_source_33_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25557_) );
  \$mux  #( .WIDTH(33) ) _47986_ ( .A(_25557_), .B(33'h000000000), .S(RST), .Y(_02231_) );
  \$mux  #( .WIDTH(33) ) _47987_ ( .A(_source_stream_conv2d_16_source_33_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25558_) );
  \$mux  #( .WIDTH(33) ) _47988_ ( .A(_25558_), .B(33'h000000000), .S(RST), .Y(_02230_) );
  \$mux  #( .WIDTH(33) ) _47989_ ( .A(_source_stream_conv2d_16_source_33_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25559_) );
  \$mux  #( .WIDTH(33) ) _47990_ ( .A(_25559_), .B(33'h000000000), .S(RST), .Y(_02229_) );
  \$mux  #( .WIDTH(33) ) _47991_ ( .A(_source_stream_conv2d_16_source_33_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25560_) );
  \$mux  #( .WIDTH(33) ) _47992_ ( .A(_25560_), .B(33'h000000000), .S(RST), .Y(_02228_) );
  \$mux  #( .WIDTH(32) ) _47993_ ( .A(_source_stream_conv2d_16_source_33_pat_cur_offset_3), .B(0), .S(_06766_), .Y(_25561_) );
  \$mux  #( .WIDTH(32) ) _47994_ ( .A(_25561_), .B(_24384_), .S(_06769_), .Y(_25562_) );
  \$mux  #( .WIDTH(32) ) _47995_ ( .A(_25562_), .B(0), .S(_06770_), .Y(_25563_) );
  \$mux  #( .WIDTH(32) ) _47996_ ( .A(_25563_), .B(0), .S(RST), .Y(_02227_) );
  \$mux  #( .WIDTH(32) ) _47997_ ( .A(_source_stream_conv2d_16_source_33_pat_cur_offset_2), .B(0), .S(_06766_), .Y(_25564_) );
  \$mux  #( .WIDTH(32) ) _47998_ ( .A(_25564_), .B(_24383_), .S(_06768_), .Y(_25565_) );
  \$mux  #( .WIDTH(32) ) _47999_ ( .A(_25565_), .B(0), .S(_06769_), .Y(_25566_) );
  \$mux  #( .WIDTH(32) ) _48000_ ( .A(_25566_), .B(0), .S(RST), .Y(_02226_) );
  \$mux  #( .WIDTH(32) ) _48001_ ( .A(_source_stream_conv2d_16_source_33_pat_cur_offset_1), .B(0), .S(_06766_), .Y(_25567_) );
  \$mux  #( .WIDTH(32) ) _48002_ ( .A(_25567_), .B(_24382_), .S(_06767_), .Y(_25568_) );
  \$mux  #( .WIDTH(32) ) _48003_ ( .A(_25568_), .B(0), .S(_06768_), .Y(_25569_) );
  \$mux  #( .WIDTH(32) ) _48004_ ( .A(_25569_), .B(0), .S(RST), .Y(_02225_) );
  \$mux  #( .WIDTH(32) ) _48005_ ( .A(_source_stream_conv2d_16_source_33_pat_cur_offset_0), .B(0), .S(_06766_), .Y(_25570_) );
  \$mux  #( .WIDTH(32) ) _48006_ ( .A(_24381_), .B(_25570_), .S(_05956_), .Y(_25571_) );
  \$mux  #( .WIDTH(32) ) _48007_ ( .A(_25571_), .B(0), .S(_06767_), .Y(_25572_) );
  \$mux  #( .WIDTH(32) ) _48008_ ( .A(_25572_), .B(0), .S(RST), .Y(_02224_) );
  \$mux  #( .WIDTH(4) ) _48009_ ( .A(__variable_wdata_506), .B(_stream_conv2d_16_source_32_source_ram_rdata), .S(_stream_conv2d_16_source_32_source_ram_rvalid), .Y(_25573_) );
  \$mux  #( .WIDTH(4) ) _48010_ ( .A(_25573_), .B(4'h0), .S(RST), .Y(_01434_) );
  \$mux  #( .WIDTH(32) ) _48011_ ( .A(_source_stream_conv2d_16_source_32_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_32_pat_stride_3), .S(_06761_), .Y(_25574_) );
  \$mux  #( .WIDTH(32) ) _48012_ ( .A(_25574_), .B(0), .S(RST), .Y(_02219_) );
  \$mux  #( .WIDTH(32) ) _48013_ ( .A(_source_stream_conv2d_16_source_32_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_32_pat_stride_2), .S(_06761_), .Y(_25575_) );
  \$mux  #( .WIDTH(32) ) _48014_ ( .A(_25575_), .B(0), .S(RST), .Y(_02218_) );
  \$mux  #( .WIDTH(32) ) _48015_ ( .A(_source_stream_conv2d_16_source_32_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_32_pat_stride_1), .S(_06761_), .Y(_25576_) );
  \$mux  #( .WIDTH(32) ) _48016_ ( .A(_25576_), .B(0), .S(RST), .Y(_02217_) );
  \$mux  #( .WIDTH(32) ) _48017_ ( .A(_source_stream_conv2d_16_source_32_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_32_pat_stride_0), .S(_06761_), .Y(_25577_) );
  \$mux  #( .WIDTH(32) ) _48018_ ( .A(_25577_), .B(0), .S(RST), .Y(_02216_) );
  \$mux  #( .WIDTH(33) ) _48019_ ( .A(_source_stream_conv2d_16_source_32_pat_size_buf_3), .B(_source_stream_conv2d_16_source_32_pat_size_3), .S(_06761_), .Y(_25578_) );
  \$mux  #( .WIDTH(33) ) _48020_ ( .A(_25578_), .B(33'h000000000), .S(RST), .Y(_02211_) );
  \$mux  #( .WIDTH(33) ) _48021_ ( .A(_source_stream_conv2d_16_source_32_pat_size_buf_2), .B(_source_stream_conv2d_16_source_32_pat_size_2), .S(_06761_), .Y(_25579_) );
  \$mux  #( .WIDTH(33) ) _48022_ ( .A(_25579_), .B(33'h000000000), .S(RST), .Y(_02210_) );
  \$mux  #( .WIDTH(33) ) _48023_ ( .A(_source_stream_conv2d_16_source_32_pat_size_buf_1), .B(_source_stream_conv2d_16_source_32_pat_size_1), .S(_06761_), .Y(_25580_) );
  \$mux  #( .WIDTH(33) ) _48024_ ( .A(_25580_), .B(33'h000000000), .S(RST), .Y(_02209_) );
  \$mux  #( .WIDTH(33) ) _48025_ ( .A(_source_stream_conv2d_16_source_32_pat_size_buf_0), .B(_source_stream_conv2d_16_source_32_pat_size_0), .S(_06761_), .Y(_25581_) );
  \$mux  #( .WIDTH(33) ) _48026_ ( .A(_25581_), .B(33'h000000000), .S(RST), .Y(_02208_) );
  \$mux  #( .WIDTH(33) ) _48027_ ( .A(_source_stream_conv2d_16_source_32_pat_count_3), .B(_28811_), .S(_06761_), .Y(_25582_) );
  \$mux  #( .WIDTH(33) ) _48028_ ( .A(_25582_), .B(_28818_), .S(_06764_), .Y(_25583_) );
  \$mux  #( .WIDTH(33) ) _48029_ ( .A(_25583_), .B(_28819_), .S(_06765_), .Y(_25584_) );
  \$mux  #( .WIDTH(33) ) _48030_ ( .A(_25584_), .B(33'h000000000), .S(RST), .Y(_02199_) );
  \$mux  #( .WIDTH(33) ) _48031_ ( .A(_source_stream_conv2d_16_source_32_pat_count_2), .B(_28810_), .S(_06761_), .Y(_25585_) );
  \$mux  #( .WIDTH(33) ) _48032_ ( .A(_25585_), .B(_28816_), .S(_06763_), .Y(_25586_) );
  \$mux  #( .WIDTH(33) ) _48033_ ( .A(_25586_), .B(_28817_), .S(_06764_), .Y(_25587_) );
  \$mux  #( .WIDTH(33) ) _48034_ ( .A(_25587_), .B(33'h000000000), .S(RST), .Y(_02198_) );
  \$mux  #( .WIDTH(33) ) _48035_ ( .A(_source_stream_conv2d_16_source_32_pat_count_1), .B(_28809_), .S(_06761_), .Y(_25588_) );
  \$mux  #( .WIDTH(33) ) _48036_ ( .A(_25588_), .B(_28814_), .S(_06762_), .Y(_25589_) );
  \$mux  #( .WIDTH(33) ) _48037_ ( .A(_25589_), .B(_28815_), .S(_06763_), .Y(_25590_) );
  \$mux  #( .WIDTH(33) ) _48038_ ( .A(_25590_), .B(33'h000000000), .S(RST), .Y(_02197_) );
  \$mux  #( .WIDTH(33) ) _48039_ ( .A(_source_stream_conv2d_16_source_32_pat_count_0), .B(_28808_), .S(_06761_), .Y(_25591_) );
  \$mux  #( .WIDTH(33) ) _48040_ ( .A(_28812_), .B(_25591_), .S(_05959_), .Y(_25592_) );
  \$mux  #( .WIDTH(33) ) _48041_ ( .A(_25592_), .B(_28813_), .S(_06762_), .Y(_25593_) );
  \$mux  #( .WIDTH(33) ) _48042_ ( .A(_25593_), .B(33'h000000000), .S(RST), .Y(_02196_) );
  \$mux  #( .WIDTH(32) ) _48043_ ( .A(_source_stream_conv2d_16_source_32_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25594_) );
  \$mux  #( .WIDTH(32) ) _48044_ ( .A(_25594_), .B(0), .S(RST), .Y(_02215_) );
  \$mux  #( .WIDTH(32) ) _48045_ ( .A(_source_stream_conv2d_16_source_32_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25595_) );
  \$mux  #( .WIDTH(32) ) _48046_ ( .A(_25595_), .B(0), .S(RST), .Y(_02214_) );
  \$mux  #( .WIDTH(32) ) _48047_ ( .A(_source_stream_conv2d_16_source_32_pat_stride_1), .B({ 26'h0000000, cparam_conv2d_16_filter_read_block }), .S(_set_flag_710), .Y(_25596_) );
  \$mux  #( .WIDTH(32) ) _48048_ ( .A(_25596_), .B(0), .S(RST), .Y(_02213_) );
  \$mux  #( .WIDTH(32) ) _48049_ ( .A(_source_stream_conv2d_16_source_32_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25597_) );
  \$mux  #( .WIDTH(32) ) _48050_ ( .A(_25597_), .B(0), .S(RST), .Y(_02212_) );
  \$mux  #( .WIDTH(33) ) _48051_ ( .A(_source_stream_conv2d_16_source_32_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25598_) );
  \$mux  #( .WIDTH(33) ) _48052_ ( .A(_25598_), .B(33'h000000000), .S(RST), .Y(_02207_) );
  \$mux  #( .WIDTH(33) ) _48053_ ( .A(_source_stream_conv2d_16_source_32_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25599_) );
  \$mux  #( .WIDTH(33) ) _48054_ ( .A(_25599_), .B(33'h000000000), .S(RST), .Y(_02206_) );
  \$mux  #( .WIDTH(33) ) _48055_ ( .A(_source_stream_conv2d_16_source_32_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25600_) );
  \$mux  #( .WIDTH(33) ) _48056_ ( .A(_25600_), .B(33'h000000000), .S(RST), .Y(_02205_) );
  \$mux  #( .WIDTH(33) ) _48057_ ( .A(_source_stream_conv2d_16_source_32_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25601_) );
  \$mux  #( .WIDTH(33) ) _48058_ ( .A(_25601_), .B(33'h000000000), .S(RST), .Y(_02204_) );
  \$mux  #( .WIDTH(32) ) _48059_ ( .A(_source_stream_conv2d_16_source_32_pat_cur_offset_3), .B(0), .S(_06761_), .Y(_25602_) );
  \$mux  #( .WIDTH(32) ) _48060_ ( .A(_25602_), .B(_24380_), .S(_06764_), .Y(_25603_) );
  \$mux  #( .WIDTH(32) ) _48061_ ( .A(_25603_), .B(0), .S(_06765_), .Y(_25604_) );
  \$mux  #( .WIDTH(32) ) _48062_ ( .A(_25604_), .B(0), .S(RST), .Y(_02203_) );
  \$mux  #( .WIDTH(32) ) _48063_ ( .A(_source_stream_conv2d_16_source_32_pat_cur_offset_2), .B(0), .S(_06761_), .Y(_25605_) );
  \$mux  #( .WIDTH(32) ) _48064_ ( .A(_25605_), .B(_24379_), .S(_06763_), .Y(_25606_) );
  \$mux  #( .WIDTH(32) ) _48065_ ( .A(_25606_), .B(0), .S(_06764_), .Y(_25607_) );
  \$mux  #( .WIDTH(32) ) _48066_ ( .A(_25607_), .B(0), .S(RST), .Y(_02202_) );
  \$mux  #( .WIDTH(32) ) _48067_ ( .A(_source_stream_conv2d_16_source_32_pat_cur_offset_1), .B(0), .S(_06761_), .Y(_25608_) );
  \$mux  #( .WIDTH(32) ) _48068_ ( .A(_25608_), .B(_24378_), .S(_06762_), .Y(_25609_) );
  \$mux  #( .WIDTH(32) ) _48069_ ( .A(_25609_), .B(0), .S(_06763_), .Y(_25610_) );
  \$mux  #( .WIDTH(32) ) _48070_ ( .A(_25610_), .B(0), .S(RST), .Y(_02201_) );
  \$mux  #( .WIDTH(32) ) _48071_ ( .A(_source_stream_conv2d_16_source_32_pat_cur_offset_0), .B(0), .S(_06761_), .Y(_25611_) );
  \$mux  #( .WIDTH(32) ) _48072_ ( .A(_24377_), .B(_25611_), .S(_05959_), .Y(_25612_) );
  \$mux  #( .WIDTH(32) ) _48073_ ( .A(_25612_), .B(0), .S(_06762_), .Y(_25613_) );
  \$mux  #( .WIDTH(32) ) _48074_ ( .A(_25613_), .B(0), .S(RST), .Y(_02200_) );
  \$mux  #( .WIDTH(4) ) _48075_ ( .A(__variable_wdata_505), .B(_stream_conv2d_16_source_31_source_ram_rdata), .S(_stream_conv2d_16_source_31_source_ram_rvalid), .Y(_25614_) );
  \$mux  #( .WIDTH(4) ) _48076_ ( .A(_25614_), .B(4'h0), .S(RST), .Y(_01433_) );
  \$mux  #( .WIDTH(32) ) _48077_ ( .A(_source_stream_conv2d_16_source_31_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_31_pat_stride_3), .S(_06756_), .Y(_25615_) );
  \$mux  #( .WIDTH(32) ) _48078_ ( .A(_25615_), .B(0), .S(RST), .Y(_02195_) );
  \$mux  #( .WIDTH(32) ) _48079_ ( .A(_source_stream_conv2d_16_source_31_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_31_pat_stride_2), .S(_06756_), .Y(_25616_) );
  \$mux  #( .WIDTH(32) ) _48080_ ( .A(_25616_), .B(0), .S(RST), .Y(_02194_) );
  \$mux  #( .WIDTH(32) ) _48081_ ( .A(_source_stream_conv2d_16_source_31_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_31_pat_stride_1), .S(_06756_), .Y(_25617_) );
  \$mux  #( .WIDTH(32) ) _48082_ ( .A(_25617_), .B(0), .S(RST), .Y(_02193_) );
  \$mux  #( .WIDTH(32) ) _48083_ ( .A(_source_stream_conv2d_16_source_31_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_31_pat_stride_0), .S(_06756_), .Y(_25618_) );
  \$mux  #( .WIDTH(32) ) _48084_ ( .A(_25618_), .B(0), .S(RST), .Y(_02192_) );
  \$mux  #( .WIDTH(33) ) _48085_ ( .A(_source_stream_conv2d_16_source_31_pat_size_buf_3), .B(_source_stream_conv2d_16_source_31_pat_size_3), .S(_06756_), .Y(_25619_) );
  \$mux  #( .WIDTH(33) ) _48086_ ( .A(_25619_), .B(33'h000000000), .S(RST), .Y(_02187_) );
  \$mux  #( .WIDTH(33) ) _48087_ ( .A(_source_stream_conv2d_16_source_31_pat_size_buf_2), .B(_source_stream_conv2d_16_source_31_pat_size_2), .S(_06756_), .Y(_25620_) );
  \$mux  #( .WIDTH(33) ) _48088_ ( .A(_25620_), .B(33'h000000000), .S(RST), .Y(_02186_) );
  \$mux  #( .WIDTH(33) ) _48089_ ( .A(_source_stream_conv2d_16_source_31_pat_size_buf_1), .B(_source_stream_conv2d_16_source_31_pat_size_1), .S(_06756_), .Y(_25621_) );
  \$mux  #( .WIDTH(33) ) _48090_ ( .A(_25621_), .B(33'h000000000), .S(RST), .Y(_02185_) );
  \$mux  #( .WIDTH(33) ) _48091_ ( .A(_source_stream_conv2d_16_source_31_pat_size_buf_0), .B(_source_stream_conv2d_16_source_31_pat_size_0), .S(_06756_), .Y(_25622_) );
  \$mux  #( .WIDTH(33) ) _48092_ ( .A(_25622_), .B(33'h000000000), .S(RST), .Y(_02184_) );
  \$mux  #( .WIDTH(33) ) _48093_ ( .A(_source_stream_conv2d_16_source_31_pat_count_3), .B(_28799_), .S(_06756_), .Y(_25623_) );
  \$mux  #( .WIDTH(33) ) _48094_ ( .A(_25623_), .B(_28806_), .S(_06759_), .Y(_25624_) );
  \$mux  #( .WIDTH(33) ) _48095_ ( .A(_25624_), .B(_28807_), .S(_06760_), .Y(_25625_) );
  \$mux  #( .WIDTH(33) ) _48096_ ( .A(_25625_), .B(33'h000000000), .S(RST), .Y(_02175_) );
  \$mux  #( .WIDTH(33) ) _48097_ ( .A(_source_stream_conv2d_16_source_31_pat_count_2), .B(_28798_), .S(_06756_), .Y(_25626_) );
  \$mux  #( .WIDTH(33) ) _48098_ ( .A(_25626_), .B(_28804_), .S(_06758_), .Y(_25627_) );
  \$mux  #( .WIDTH(33) ) _48099_ ( .A(_25627_), .B(_28805_), .S(_06759_), .Y(_25628_) );
  \$mux  #( .WIDTH(33) ) _48100_ ( .A(_25628_), .B(33'h000000000), .S(RST), .Y(_02174_) );
  \$mux  #( .WIDTH(33) ) _48101_ ( .A(_source_stream_conv2d_16_source_31_pat_count_1), .B(_28797_), .S(_06756_), .Y(_25629_) );
  \$mux  #( .WIDTH(33) ) _48102_ ( .A(_25629_), .B(_28802_), .S(_06757_), .Y(_25630_) );
  \$mux  #( .WIDTH(33) ) _48103_ ( .A(_25630_), .B(_28803_), .S(_06758_), .Y(_25631_) );
  \$mux  #( .WIDTH(33) ) _48104_ ( .A(_25631_), .B(33'h000000000), .S(RST), .Y(_02173_) );
  \$mux  #( .WIDTH(33) ) _48105_ ( .A(_source_stream_conv2d_16_source_31_pat_count_0), .B(_28796_), .S(_06756_), .Y(_25632_) );
  \$mux  #( .WIDTH(33) ) _48106_ ( .A(_28800_), .B(_25632_), .S(_05962_), .Y(_25633_) );
  \$mux  #( .WIDTH(33) ) _48107_ ( .A(_25633_), .B(_28801_), .S(_06757_), .Y(_25634_) );
  \$mux  #( .WIDTH(33) ) _48108_ ( .A(_25634_), .B(33'h000000000), .S(RST), .Y(_02172_) );
  \$mux  #( .WIDTH(32) ) _48109_ ( .A(_source_stream_conv2d_16_source_31_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25635_) );
  \$mux  #( .WIDTH(32) ) _48110_ ( .A(_25635_), .B(0), .S(RST), .Y(_02191_) );
  \$mux  #( .WIDTH(32) ) _48111_ ( .A(_source_stream_conv2d_16_source_31_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25636_) );
  \$mux  #( .WIDTH(32) ) _48112_ ( .A(_25636_), .B(0), .S(RST), .Y(_02190_) );
  \$mux  #( .WIDTH(32) ) _48113_ ( .A(_source_stream_conv2d_16_source_31_pat_stride_1), .B({ 26'h0000000, cparam_conv2d_16_filter_read_block }), .S(_set_flag_710), .Y(_25637_) );
  \$mux  #( .WIDTH(32) ) _48114_ ( .A(_25637_), .B(0), .S(RST), .Y(_02189_) );
  \$mux  #( .WIDTH(32) ) _48115_ ( .A(_source_stream_conv2d_16_source_31_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25638_) );
  \$mux  #( .WIDTH(32) ) _48116_ ( .A(_25638_), .B(0), .S(RST), .Y(_02188_) );
  \$mux  #( .WIDTH(33) ) _48117_ ( .A(_source_stream_conv2d_16_source_31_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25639_) );
  \$mux  #( .WIDTH(33) ) _48118_ ( .A(_25639_), .B(33'h000000000), .S(RST), .Y(_02183_) );
  \$mux  #( .WIDTH(33) ) _48119_ ( .A(_source_stream_conv2d_16_source_31_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25640_) );
  \$mux  #( .WIDTH(33) ) _48120_ ( .A(_25640_), .B(33'h000000000), .S(RST), .Y(_02182_) );
  \$mux  #( .WIDTH(33) ) _48121_ ( .A(_source_stream_conv2d_16_source_31_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25641_) );
  \$mux  #( .WIDTH(33) ) _48122_ ( .A(_25641_), .B(33'h000000000), .S(RST), .Y(_02181_) );
  \$mux  #( .WIDTH(33) ) _48123_ ( .A(_source_stream_conv2d_16_source_31_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25642_) );
  \$mux  #( .WIDTH(33) ) _48124_ ( .A(_25642_), .B(33'h000000000), .S(RST), .Y(_02180_) );
  \$mux  #( .WIDTH(32) ) _48125_ ( .A(_source_stream_conv2d_16_source_31_pat_cur_offset_3), .B(0), .S(_06756_), .Y(_25643_) );
  \$mux  #( .WIDTH(32) ) _48126_ ( .A(_25643_), .B(_24376_), .S(_06759_), .Y(_25644_) );
  \$mux  #( .WIDTH(32) ) _48127_ ( .A(_25644_), .B(0), .S(_06760_), .Y(_25645_) );
  \$mux  #( .WIDTH(32) ) _48128_ ( .A(_25645_), .B(0), .S(RST), .Y(_02179_) );
  \$mux  #( .WIDTH(32) ) _48129_ ( .A(_source_stream_conv2d_16_source_31_pat_cur_offset_2), .B(0), .S(_06756_), .Y(_25646_) );
  \$mux  #( .WIDTH(32) ) _48130_ ( .A(_25646_), .B(_24375_), .S(_06758_), .Y(_25647_) );
  \$mux  #( .WIDTH(32) ) _48131_ ( .A(_25647_), .B(0), .S(_06759_), .Y(_25648_) );
  \$mux  #( .WIDTH(32) ) _48132_ ( .A(_25648_), .B(0), .S(RST), .Y(_02178_) );
  \$mux  #( .WIDTH(32) ) _48133_ ( .A(_source_stream_conv2d_16_source_31_pat_cur_offset_1), .B(0), .S(_06756_), .Y(_25649_) );
  \$mux  #( .WIDTH(32) ) _48134_ ( .A(_25649_), .B(_24374_), .S(_06757_), .Y(_25650_) );
  \$mux  #( .WIDTH(32) ) _48135_ ( .A(_25650_), .B(0), .S(_06758_), .Y(_25651_) );
  \$mux  #( .WIDTH(32) ) _48136_ ( .A(_25651_), .B(0), .S(RST), .Y(_02177_) );
  \$mux  #( .WIDTH(32) ) _48137_ ( .A(_source_stream_conv2d_16_source_31_pat_cur_offset_0), .B(0), .S(_06756_), .Y(_25652_) );
  \$mux  #( .WIDTH(32) ) _48138_ ( .A(_24373_), .B(_25652_), .S(_05962_), .Y(_25653_) );
  \$mux  #( .WIDTH(32) ) _48139_ ( .A(_25653_), .B(0), .S(_06757_), .Y(_25654_) );
  \$mux  #( .WIDTH(32) ) _48140_ ( .A(_25654_), .B(0), .S(RST), .Y(_02176_) );
  \$mux  #( .WIDTH(4) ) _48141_ ( .A(__variable_wdata_504), .B(_stream_conv2d_16_source_30_source_ram_rdata), .S(_stream_conv2d_16_source_30_source_ram_rvalid), .Y(_25655_) );
  \$mux  #( .WIDTH(4) ) _48142_ ( .A(_25655_), .B(4'h0), .S(RST), .Y(_01432_) );
  \$mux  #( .WIDTH(1) ) _48143_ ( .A(_tmp_625), .B(1'h0), .S(RST), .Y(_01270_) );
  \$mux  #( .WIDTH(32) ) _48144_ ( .A(_source_stream_conv2d_16_source_30_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_30_pat_stride_3), .S(_06751_), .Y(_25656_) );
  \$mux  #( .WIDTH(32) ) _48145_ ( .A(_25656_), .B(0), .S(RST), .Y(_02171_) );
  \$mux  #( .WIDTH(32) ) _48146_ ( .A(_source_stream_conv2d_16_source_30_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_30_pat_stride_2), .S(_06751_), .Y(_25657_) );
  \$mux  #( .WIDTH(32) ) _48147_ ( .A(_25657_), .B(0), .S(RST), .Y(_02170_) );
  \$mux  #( .WIDTH(32) ) _48148_ ( .A(_source_stream_conv2d_16_source_30_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_30_pat_stride_1), .S(_06751_), .Y(_25658_) );
  \$mux  #( .WIDTH(32) ) _48149_ ( .A(_25658_), .B(0), .S(RST), .Y(_02169_) );
  \$mux  #( .WIDTH(32) ) _48150_ ( .A(_source_stream_conv2d_16_source_30_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_30_pat_stride_0), .S(_06751_), .Y(_25659_) );
  \$mux  #( .WIDTH(32) ) _48151_ ( .A(_25659_), .B(0), .S(RST), .Y(_02168_) );
  \$mux  #( .WIDTH(33) ) _48152_ ( .A(_source_stream_conv2d_16_source_30_pat_size_buf_3), .B(_source_stream_conv2d_16_source_30_pat_size_3), .S(_06751_), .Y(_25660_) );
  \$mux  #( .WIDTH(33) ) _48153_ ( .A(_25660_), .B(33'h000000000), .S(RST), .Y(_02163_) );
  \$mux  #( .WIDTH(33) ) _48154_ ( .A(_source_stream_conv2d_16_source_30_pat_size_buf_2), .B(_source_stream_conv2d_16_source_30_pat_size_2), .S(_06751_), .Y(_25661_) );
  \$mux  #( .WIDTH(33) ) _48155_ ( .A(_25661_), .B(33'h000000000), .S(RST), .Y(_02162_) );
  \$mux  #( .WIDTH(33) ) _48156_ ( .A(_source_stream_conv2d_16_source_30_pat_size_buf_1), .B(_source_stream_conv2d_16_source_30_pat_size_1), .S(_06751_), .Y(_25662_) );
  \$mux  #( .WIDTH(33) ) _48157_ ( .A(_25662_), .B(33'h000000000), .S(RST), .Y(_02161_) );
  \$mux  #( .WIDTH(33) ) _48158_ ( .A(_source_stream_conv2d_16_source_30_pat_size_buf_0), .B(_source_stream_conv2d_16_source_30_pat_size_0), .S(_06751_), .Y(_25663_) );
  \$mux  #( .WIDTH(33) ) _48159_ ( .A(_25663_), .B(33'h000000000), .S(RST), .Y(_02160_) );
  \$mux  #( .WIDTH(33) ) _48160_ ( .A(_source_stream_conv2d_16_source_30_pat_count_3), .B(_28787_), .S(_06751_), .Y(_25664_) );
  \$mux  #( .WIDTH(33) ) _48161_ ( .A(_25664_), .B(_28794_), .S(_06754_), .Y(_25665_) );
  \$mux  #( .WIDTH(33) ) _48162_ ( .A(_25665_), .B(_28795_), .S(_06755_), .Y(_25666_) );
  \$mux  #( .WIDTH(33) ) _48163_ ( .A(_25666_), .B(33'h000000000), .S(RST), .Y(_02151_) );
  \$mux  #( .WIDTH(33) ) _48164_ ( .A(_source_stream_conv2d_16_source_30_pat_count_2), .B(_28786_), .S(_06751_), .Y(_25667_) );
  \$mux  #( .WIDTH(33) ) _48165_ ( .A(_25667_), .B(_28792_), .S(_06753_), .Y(_25668_) );
  \$mux  #( .WIDTH(33) ) _48166_ ( .A(_25668_), .B(_28793_), .S(_06754_), .Y(_25669_) );
  \$mux  #( .WIDTH(33) ) _48167_ ( .A(_25669_), .B(33'h000000000), .S(RST), .Y(_02150_) );
  \$mux  #( .WIDTH(33) ) _48168_ ( .A(_source_stream_conv2d_16_source_30_pat_count_1), .B(_28785_), .S(_06751_), .Y(_25670_) );
  \$mux  #( .WIDTH(33) ) _48169_ ( .A(_25670_), .B(_28790_), .S(_06752_), .Y(_25671_) );
  \$mux  #( .WIDTH(33) ) _48170_ ( .A(_25671_), .B(_28791_), .S(_06753_), .Y(_25672_) );
  \$mux  #( .WIDTH(33) ) _48171_ ( .A(_25672_), .B(33'h000000000), .S(RST), .Y(_02149_) );
  \$mux  #( .WIDTH(33) ) _48172_ ( .A(_source_stream_conv2d_16_source_30_pat_count_0), .B(_28784_), .S(_06751_), .Y(_25673_) );
  \$mux  #( .WIDTH(33) ) _48173_ ( .A(_28788_), .B(_25673_), .S(_05960_), .Y(_25674_) );
  \$mux  #( .WIDTH(33) ) _48174_ ( .A(_25674_), .B(_28789_), .S(_06752_), .Y(_25675_) );
  \$mux  #( .WIDTH(33) ) _48175_ ( .A(_25675_), .B(33'h000000000), .S(RST), .Y(_02148_) );
  \$mux  #( .WIDTH(32) ) _48176_ ( .A(_source_stream_conv2d_16_source_30_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25676_) );
  \$mux  #( .WIDTH(32) ) _48177_ ( .A(_25676_), .B(0), .S(RST), .Y(_02167_) );
  \$mux  #( .WIDTH(32) ) _48178_ ( .A(_source_stream_conv2d_16_source_30_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25677_) );
  \$mux  #( .WIDTH(32) ) _48179_ ( .A(_25677_), .B(0), .S(RST), .Y(_02166_) );
  \$mux  #( .WIDTH(32) ) _48180_ ( .A(_source_stream_conv2d_16_source_30_pat_stride_1), .B({ 26'h0000000, cparam_conv2d_16_filter_read_block }), .S(_set_flag_710), .Y(_25678_) );
  \$mux  #( .WIDTH(32) ) _48181_ ( .A(_25678_), .B(0), .S(RST), .Y(_02165_) );
  \$mux  #( .WIDTH(32) ) _48182_ ( .A(_source_stream_conv2d_16_source_30_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25679_) );
  \$mux  #( .WIDTH(32) ) _48183_ ( .A(_25679_), .B(0), .S(RST), .Y(_02164_) );
  \$mux  #( .WIDTH(33) ) _48184_ ( .A(_source_stream_conv2d_16_source_30_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25680_) );
  \$mux  #( .WIDTH(33) ) _48185_ ( .A(_25680_), .B(33'h000000000), .S(RST), .Y(_02159_) );
  \$mux  #( .WIDTH(33) ) _48186_ ( .A(_source_stream_conv2d_16_source_30_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25681_) );
  \$mux  #( .WIDTH(33) ) _48187_ ( .A(_25681_), .B(33'h000000000), .S(RST), .Y(_02158_) );
  \$mux  #( .WIDTH(33) ) _48188_ ( .A(_source_stream_conv2d_16_source_30_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25682_) );
  \$mux  #( .WIDTH(33) ) _48189_ ( .A(_25682_), .B(33'h000000000), .S(RST), .Y(_02157_) );
  \$mux  #( .WIDTH(33) ) _48190_ ( .A(_source_stream_conv2d_16_source_30_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25683_) );
  \$mux  #( .WIDTH(33) ) _48191_ ( .A(_25683_), .B(33'h000000000), .S(RST), .Y(_02156_) );
  \$mux  #( .WIDTH(32) ) _48192_ ( .A(_source_stream_conv2d_16_source_30_pat_cur_offset_3), .B(0), .S(_06751_), .Y(_25684_) );
  \$mux  #( .WIDTH(32) ) _48193_ ( .A(_25684_), .B(_24372_), .S(_06754_), .Y(_25685_) );
  \$mux  #( .WIDTH(32) ) _48194_ ( .A(_25685_), .B(0), .S(_06755_), .Y(_25686_) );
  \$mux  #( .WIDTH(32) ) _48195_ ( .A(_25686_), .B(0), .S(RST), .Y(_02155_) );
  \$mux  #( .WIDTH(32) ) _48196_ ( .A(_source_stream_conv2d_16_source_30_pat_cur_offset_2), .B(0), .S(_06751_), .Y(_25687_) );
  \$mux  #( .WIDTH(32) ) _48197_ ( .A(_25687_), .B(_24371_), .S(_06753_), .Y(_25688_) );
  \$mux  #( .WIDTH(32) ) _48198_ ( .A(_25688_), .B(0), .S(_06754_), .Y(_25689_) );
  \$mux  #( .WIDTH(32) ) _48199_ ( .A(_25689_), .B(0), .S(RST), .Y(_02154_) );
  \$mux  #( .WIDTH(32) ) _48200_ ( .A(_source_stream_conv2d_16_source_30_pat_cur_offset_1), .B(0), .S(_06751_), .Y(_25690_) );
  \$mux  #( .WIDTH(32) ) _48201_ ( .A(_25690_), .B(_24370_), .S(_06752_), .Y(_25691_) );
  \$mux  #( .WIDTH(32) ) _48202_ ( .A(_25691_), .B(0), .S(_06753_), .Y(_25692_) );
  \$mux  #( .WIDTH(32) ) _48203_ ( .A(_25692_), .B(0), .S(RST), .Y(_02153_) );
  \$mux  #( .WIDTH(32) ) _48204_ ( .A(_source_stream_conv2d_16_source_30_pat_cur_offset_0), .B(0), .S(_06751_), .Y(_25693_) );
  \$mux  #( .WIDTH(32) ) _48205_ ( .A(_24369_), .B(_25693_), .S(_05960_), .Y(_25694_) );
  \$mux  #( .WIDTH(32) ) _48206_ ( .A(_25694_), .B(0), .S(_06752_), .Y(_25695_) );
  \$mux  #( .WIDTH(32) ) _48207_ ( .A(_25695_), .B(0), .S(RST), .Y(_02152_) );
  \$mux  #( .WIDTH(4) ) _48208_ ( .A(__variable_wdata_503), .B(_stream_conv2d_16_source_29_source_ram_rdata), .S(_stream_conv2d_16_source_29_source_ram_rvalid), .Y(_25696_) );
  \$mux  #( .WIDTH(4) ) _48209_ ( .A(_25696_), .B(4'h0), .S(RST), .Y(_01431_) );
  \$mux  #( .WIDTH(1) ) _48210_ ( .A(_tmp_611), .B(1'h0), .S(RST), .Y(_01267_) );
  \$mux  #( .WIDTH(32) ) _48211_ ( .A(_source_stream_conv2d_16_source_29_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_29_pat_stride_3), .S(_06746_), .Y(_25697_) );
  \$mux  #( .WIDTH(32) ) _48212_ ( .A(_25697_), .B(0), .S(RST), .Y(_02147_) );
  \$mux  #( .WIDTH(32) ) _48213_ ( .A(_source_stream_conv2d_16_source_29_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_29_pat_stride_2), .S(_06746_), .Y(_25698_) );
  \$mux  #( .WIDTH(32) ) _48214_ ( .A(_25698_), .B(0), .S(RST), .Y(_02146_) );
  \$mux  #( .WIDTH(32) ) _48215_ ( .A(_source_stream_conv2d_16_source_29_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_29_pat_stride_1), .S(_06746_), .Y(_25699_) );
  \$mux  #( .WIDTH(32) ) _48216_ ( .A(_25699_), .B(0), .S(RST), .Y(_02145_) );
  \$mux  #( .WIDTH(32) ) _48217_ ( .A(_source_stream_conv2d_16_source_29_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_29_pat_stride_0), .S(_06746_), .Y(_25700_) );
  \$mux  #( .WIDTH(32) ) _48218_ ( .A(_25700_), .B(0), .S(RST), .Y(_02144_) );
  \$mux  #( .WIDTH(33) ) _48219_ ( .A(_source_stream_conv2d_16_source_29_pat_size_buf_3), .B(_source_stream_conv2d_16_source_29_pat_size_3), .S(_06746_), .Y(_25701_) );
  \$mux  #( .WIDTH(33) ) _48220_ ( .A(_25701_), .B(33'h000000000), .S(RST), .Y(_02139_) );
  \$mux  #( .WIDTH(33) ) _48221_ ( .A(_source_stream_conv2d_16_source_29_pat_size_buf_2), .B(_source_stream_conv2d_16_source_29_pat_size_2), .S(_06746_), .Y(_25702_) );
  \$mux  #( .WIDTH(33) ) _48222_ ( .A(_25702_), .B(33'h000000000), .S(RST), .Y(_02138_) );
  \$mux  #( .WIDTH(33) ) _48223_ ( .A(_source_stream_conv2d_16_source_29_pat_size_buf_1), .B(_source_stream_conv2d_16_source_29_pat_size_1), .S(_06746_), .Y(_25703_) );
  \$mux  #( .WIDTH(33) ) _48224_ ( .A(_25703_), .B(33'h000000000), .S(RST), .Y(_02137_) );
  \$mux  #( .WIDTH(33) ) _48225_ ( .A(_source_stream_conv2d_16_source_29_pat_size_buf_0), .B(_source_stream_conv2d_16_source_29_pat_size_0), .S(_06746_), .Y(_25704_) );
  \$mux  #( .WIDTH(33) ) _48226_ ( .A(_25704_), .B(33'h000000000), .S(RST), .Y(_02136_) );
  \$mux  #( .WIDTH(33) ) _48227_ ( .A(_source_stream_conv2d_16_source_29_pat_count_3), .B(_28775_), .S(_06746_), .Y(_25705_) );
  \$mux  #( .WIDTH(33) ) _48228_ ( .A(_25705_), .B(_28782_), .S(_06749_), .Y(_25706_) );
  \$mux  #( .WIDTH(33) ) _48229_ ( .A(_25706_), .B(_28783_), .S(_06750_), .Y(_25707_) );
  \$mux  #( .WIDTH(33) ) _48230_ ( .A(_25707_), .B(33'h000000000), .S(RST), .Y(_02127_) );
  \$mux  #( .WIDTH(33) ) _48231_ ( .A(_source_stream_conv2d_16_source_29_pat_count_2), .B(_28774_), .S(_06746_), .Y(_25708_) );
  \$mux  #( .WIDTH(33) ) _48232_ ( .A(_25708_), .B(_28780_), .S(_06748_), .Y(_25709_) );
  \$mux  #( .WIDTH(33) ) _48233_ ( .A(_25709_), .B(_28781_), .S(_06749_), .Y(_25710_) );
  \$mux  #( .WIDTH(33) ) _48234_ ( .A(_25710_), .B(33'h000000000), .S(RST), .Y(_02126_) );
  \$mux  #( .WIDTH(33) ) _48235_ ( .A(_source_stream_conv2d_16_source_29_pat_count_1), .B(_28773_), .S(_06746_), .Y(_25711_) );
  \$mux  #( .WIDTH(33) ) _48236_ ( .A(_25711_), .B(_28778_), .S(_06747_), .Y(_25712_) );
  \$mux  #( .WIDTH(33) ) _48237_ ( .A(_25712_), .B(_28779_), .S(_06748_), .Y(_25713_) );
  \$mux  #( .WIDTH(33) ) _48238_ ( .A(_25713_), .B(33'h000000000), .S(RST), .Y(_02125_) );
  \$mux  #( .WIDTH(33) ) _48239_ ( .A(_source_stream_conv2d_16_source_29_pat_count_0), .B(_28772_), .S(_06746_), .Y(_25714_) );
  \$mux  #( .WIDTH(33) ) _48240_ ( .A(_28776_), .B(_25714_), .S(_05965_), .Y(_25715_) );
  \$mux  #( .WIDTH(33) ) _48241_ ( .A(_25715_), .B(_28777_), .S(_06747_), .Y(_25716_) );
  \$mux  #( .WIDTH(33) ) _48242_ ( .A(_25716_), .B(33'h000000000), .S(RST), .Y(_02124_) );
  \$mux  #( .WIDTH(32) ) _48243_ ( .A(_source_stream_conv2d_16_source_29_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25717_) );
  \$mux  #( .WIDTH(32) ) _48244_ ( .A(_25717_), .B(0), .S(RST), .Y(_02143_) );
  \$mux  #( .WIDTH(32) ) _48245_ ( .A(_source_stream_conv2d_16_source_29_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25718_) );
  \$mux  #( .WIDTH(32) ) _48246_ ( .A(_25718_), .B(0), .S(RST), .Y(_02142_) );
  \$mux  #( .WIDTH(32) ) _48247_ ( .A(_source_stream_conv2d_16_source_29_pat_stride_1), .B({ 26'h0000000, cparam_conv2d_16_filter_read_block }), .S(_set_flag_710), .Y(_25719_) );
  \$mux  #( .WIDTH(32) ) _48248_ ( .A(_25719_), .B(0), .S(RST), .Y(_02141_) );
  \$mux  #( .WIDTH(32) ) _48249_ ( .A(_source_stream_conv2d_16_source_29_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25720_) );
  \$mux  #( .WIDTH(32) ) _48250_ ( .A(_25720_), .B(0), .S(RST), .Y(_02140_) );
  \$mux  #( .WIDTH(33) ) _48251_ ( .A(_source_stream_conv2d_16_source_29_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25721_) );
  \$mux  #( .WIDTH(33) ) _48252_ ( .A(_25721_), .B(33'h000000000), .S(RST), .Y(_02135_) );
  \$mux  #( .WIDTH(33) ) _48253_ ( .A(_source_stream_conv2d_16_source_29_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25722_) );
  \$mux  #( .WIDTH(33) ) _48254_ ( .A(_25722_), .B(33'h000000000), .S(RST), .Y(_02134_) );
  \$mux  #( .WIDTH(33) ) _48255_ ( .A(_source_stream_conv2d_16_source_29_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25723_) );
  \$mux  #( .WIDTH(33) ) _48256_ ( .A(_25723_), .B(33'h000000000), .S(RST), .Y(_02133_) );
  \$mux  #( .WIDTH(33) ) _48257_ ( .A(_source_stream_conv2d_16_source_29_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25724_) );
  \$mux  #( .WIDTH(33) ) _48258_ ( .A(_25724_), .B(33'h000000000), .S(RST), .Y(_02132_) );
  \$mux  #( .WIDTH(32) ) _48259_ ( .A(_source_stream_conv2d_16_source_29_pat_cur_offset_3), .B(0), .S(_06746_), .Y(_25725_) );
  \$mux  #( .WIDTH(32) ) _48260_ ( .A(_25725_), .B(_24368_), .S(_06749_), .Y(_25726_) );
  \$mux  #( .WIDTH(32) ) _48261_ ( .A(_25726_), .B(0), .S(_06750_), .Y(_25727_) );
  \$mux  #( .WIDTH(32) ) _48262_ ( .A(_25727_), .B(0), .S(RST), .Y(_02131_) );
  \$mux  #( .WIDTH(32) ) _48263_ ( .A(_source_stream_conv2d_16_source_29_pat_cur_offset_2), .B(0), .S(_06746_), .Y(_25728_) );
  \$mux  #( .WIDTH(32) ) _48264_ ( .A(_25728_), .B(_24367_), .S(_06748_), .Y(_25729_) );
  \$mux  #( .WIDTH(32) ) _48265_ ( .A(_25729_), .B(0), .S(_06749_), .Y(_25730_) );
  \$mux  #( .WIDTH(32) ) _48266_ ( .A(_25730_), .B(0), .S(RST), .Y(_02130_) );
  \$mux  #( .WIDTH(32) ) _48267_ ( .A(_source_stream_conv2d_16_source_29_pat_cur_offset_1), .B(0), .S(_06746_), .Y(_25731_) );
  \$mux  #( .WIDTH(32) ) _48268_ ( .A(_25731_), .B(_24366_), .S(_06747_), .Y(_25732_) );
  \$mux  #( .WIDTH(32) ) _48269_ ( .A(_25732_), .B(0), .S(_06748_), .Y(_25733_) );
  \$mux  #( .WIDTH(32) ) _48270_ ( .A(_25733_), .B(0), .S(RST), .Y(_02129_) );
  \$mux  #( .WIDTH(32) ) _48271_ ( .A(_source_stream_conv2d_16_source_29_pat_cur_offset_0), .B(0), .S(_06746_), .Y(_25734_) );
  \$mux  #( .WIDTH(32) ) _48272_ ( .A(_24365_), .B(_25734_), .S(_05965_), .Y(_25735_) );
  \$mux  #( .WIDTH(32) ) _48273_ ( .A(_25735_), .B(0), .S(_06747_), .Y(_25736_) );
  \$mux  #( .WIDTH(32) ) _48274_ ( .A(_25736_), .B(0), .S(RST), .Y(_02128_) );
  \$mux  #( .WIDTH(4) ) _48275_ ( .A(__variable_wdata_502), .B(_stream_conv2d_16_source_28_source_ram_rdata), .S(_stream_conv2d_16_source_28_source_ram_rvalid), .Y(_25737_) );
  \$mux  #( .WIDTH(4) ) _48276_ ( .A(_25737_), .B(4'h0), .S(RST), .Y(_01430_) );
  \$mux  #( .WIDTH(1) ) _48277_ ( .A(_tmp_597), .B(1'h0), .S(RST), .Y(_01264_) );
  \$mux  #( .WIDTH(32) ) _48278_ ( .A(_source_stream_conv2d_16_source_28_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_28_pat_stride_3), .S(_06741_), .Y(_25738_) );
  \$mux  #( .WIDTH(32) ) _48279_ ( .A(_25738_), .B(0), .S(RST), .Y(_02123_) );
  \$mux  #( .WIDTH(32) ) _48280_ ( .A(_source_stream_conv2d_16_source_28_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_28_pat_stride_2), .S(_06741_), .Y(_25739_) );
  \$mux  #( .WIDTH(32) ) _48281_ ( .A(_25739_), .B(0), .S(RST), .Y(_02122_) );
  \$mux  #( .WIDTH(32) ) _48282_ ( .A(_source_stream_conv2d_16_source_28_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_28_pat_stride_1), .S(_06741_), .Y(_25740_) );
  \$mux  #( .WIDTH(32) ) _48283_ ( .A(_25740_), .B(0), .S(RST), .Y(_02121_) );
  \$mux  #( .WIDTH(32) ) _48284_ ( .A(_source_stream_conv2d_16_source_28_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_28_pat_stride_0), .S(_06741_), .Y(_25741_) );
  \$mux  #( .WIDTH(32) ) _48285_ ( .A(_25741_), .B(0), .S(RST), .Y(_02120_) );
  \$mux  #( .WIDTH(33) ) _48286_ ( .A(_source_stream_conv2d_16_source_28_pat_size_buf_3), .B(_source_stream_conv2d_16_source_28_pat_size_3), .S(_06741_), .Y(_25742_) );
  \$mux  #( .WIDTH(33) ) _48287_ ( .A(_25742_), .B(33'h000000000), .S(RST), .Y(_02115_) );
  \$mux  #( .WIDTH(33) ) _48288_ ( .A(_source_stream_conv2d_16_source_28_pat_size_buf_2), .B(_source_stream_conv2d_16_source_28_pat_size_2), .S(_06741_), .Y(_25743_) );
  \$mux  #( .WIDTH(33) ) _48289_ ( .A(_25743_), .B(33'h000000000), .S(RST), .Y(_02114_) );
  \$mux  #( .WIDTH(33) ) _48290_ ( .A(_source_stream_conv2d_16_source_28_pat_size_buf_1), .B(_source_stream_conv2d_16_source_28_pat_size_1), .S(_06741_), .Y(_25744_) );
  \$mux  #( .WIDTH(33) ) _48291_ ( .A(_25744_), .B(33'h000000000), .S(RST), .Y(_02113_) );
  \$mux  #( .WIDTH(33) ) _48292_ ( .A(_source_stream_conv2d_16_source_28_pat_size_buf_0), .B(_source_stream_conv2d_16_source_28_pat_size_0), .S(_06741_), .Y(_25745_) );
  \$mux  #( .WIDTH(33) ) _48293_ ( .A(_25745_), .B(33'h000000000), .S(RST), .Y(_02112_) );
  \$mux  #( .WIDTH(33) ) _48294_ ( .A(_source_stream_conv2d_16_source_28_pat_count_3), .B(_28763_), .S(_06741_), .Y(_25746_) );
  \$mux  #( .WIDTH(33) ) _48295_ ( .A(_25746_), .B(_28770_), .S(_06744_), .Y(_25747_) );
  \$mux  #( .WIDTH(33) ) _48296_ ( .A(_25747_), .B(_28771_), .S(_06745_), .Y(_25748_) );
  \$mux  #( .WIDTH(33) ) _48297_ ( .A(_25748_), .B(33'h000000000), .S(RST), .Y(_02103_) );
  \$mux  #( .WIDTH(33) ) _48298_ ( .A(_source_stream_conv2d_16_source_28_pat_count_2), .B(_28762_), .S(_06741_), .Y(_25749_) );
  \$mux  #( .WIDTH(33) ) _48299_ ( .A(_25749_), .B(_28768_), .S(_06743_), .Y(_25750_) );
  \$mux  #( .WIDTH(33) ) _48300_ ( .A(_25750_), .B(_28769_), .S(_06744_), .Y(_25751_) );
  \$mux  #( .WIDTH(33) ) _48301_ ( .A(_25751_), .B(33'h000000000), .S(RST), .Y(_02102_) );
  \$mux  #( .WIDTH(33) ) _48302_ ( .A(_source_stream_conv2d_16_source_28_pat_count_1), .B(_28761_), .S(_06741_), .Y(_25752_) );
  \$mux  #( .WIDTH(33) ) _48303_ ( .A(_25752_), .B(_28766_), .S(_06742_), .Y(_25753_) );
  \$mux  #( .WIDTH(33) ) _48304_ ( .A(_25753_), .B(_28767_), .S(_06743_), .Y(_25754_) );
  \$mux  #( .WIDTH(33) ) _48305_ ( .A(_25754_), .B(33'h000000000), .S(RST), .Y(_02101_) );
  \$mux  #( .WIDTH(33) ) _48306_ ( .A(_source_stream_conv2d_16_source_28_pat_count_0), .B(_28760_), .S(_06741_), .Y(_25755_) );
  \$mux  #( .WIDTH(33) ) _48307_ ( .A(_28764_), .B(_25755_), .S(_05966_), .Y(_25756_) );
  \$mux  #( .WIDTH(33) ) _48308_ ( .A(_25756_), .B(_28765_), .S(_06742_), .Y(_25757_) );
  \$mux  #( .WIDTH(33) ) _48309_ ( .A(_25757_), .B(33'h000000000), .S(RST), .Y(_02100_) );
  \$mux  #( .WIDTH(32) ) _48310_ ( .A(_source_stream_conv2d_16_source_28_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25758_) );
  \$mux  #( .WIDTH(32) ) _48311_ ( .A(_25758_), .B(0), .S(RST), .Y(_02119_) );
  \$mux  #( .WIDTH(32) ) _48312_ ( .A(_source_stream_conv2d_16_source_28_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25759_) );
  \$mux  #( .WIDTH(32) ) _48313_ ( .A(_25759_), .B(0), .S(RST), .Y(_02118_) );
  \$mux  #( .WIDTH(32) ) _48314_ ( .A(_source_stream_conv2d_16_source_28_pat_stride_1), .B({ 26'h0000000, cparam_conv2d_16_filter_read_block }), .S(_set_flag_710), .Y(_25760_) );
  \$mux  #( .WIDTH(32) ) _48315_ ( .A(_25760_), .B(0), .S(RST), .Y(_02117_) );
  \$mux  #( .WIDTH(32) ) _48316_ ( .A(_source_stream_conv2d_16_source_28_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25761_) );
  \$mux  #( .WIDTH(32) ) _48317_ ( .A(_25761_), .B(0), .S(RST), .Y(_02116_) );
  \$mux  #( .WIDTH(33) ) _48318_ ( .A(_source_stream_conv2d_16_source_28_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25762_) );
  \$mux  #( .WIDTH(33) ) _48319_ ( .A(_25762_), .B(33'h000000000), .S(RST), .Y(_02111_) );
  \$mux  #( .WIDTH(33) ) _48320_ ( .A(_source_stream_conv2d_16_source_28_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25763_) );
  \$mux  #( .WIDTH(33) ) _48321_ ( .A(_25763_), .B(33'h000000000), .S(RST), .Y(_02110_) );
  \$mux  #( .WIDTH(33) ) _48322_ ( .A(_source_stream_conv2d_16_source_28_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25764_) );
  \$mux  #( .WIDTH(33) ) _48323_ ( .A(_25764_), .B(33'h000000000), .S(RST), .Y(_02109_) );
  \$mux  #( .WIDTH(33) ) _48324_ ( .A(_source_stream_conv2d_16_source_28_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25765_) );
  \$mux  #( .WIDTH(33) ) _48325_ ( .A(_25765_), .B(33'h000000000), .S(RST), .Y(_02108_) );
  \$mux  #( .WIDTH(32) ) _48326_ ( .A(_source_stream_conv2d_16_source_28_pat_cur_offset_3), .B(0), .S(_06741_), .Y(_25766_) );
  \$mux  #( .WIDTH(32) ) _48327_ ( .A(_25766_), .B(_24364_), .S(_06744_), .Y(_25767_) );
  \$mux  #( .WIDTH(32) ) _48328_ ( .A(_25767_), .B(0), .S(_06745_), .Y(_25768_) );
  \$mux  #( .WIDTH(32) ) _48329_ ( .A(_25768_), .B(0), .S(RST), .Y(_02107_) );
  \$mux  #( .WIDTH(32) ) _48330_ ( .A(_source_stream_conv2d_16_source_28_pat_cur_offset_2), .B(0), .S(_06741_), .Y(_25769_) );
  \$mux  #( .WIDTH(32) ) _48331_ ( .A(_25769_), .B(_24363_), .S(_06743_), .Y(_25770_) );
  \$mux  #( .WIDTH(32) ) _48332_ ( .A(_25770_), .B(0), .S(_06744_), .Y(_25771_) );
  \$mux  #( .WIDTH(32) ) _48333_ ( .A(_25771_), .B(0), .S(RST), .Y(_02106_) );
  \$mux  #( .WIDTH(32) ) _48334_ ( .A(_source_stream_conv2d_16_source_28_pat_cur_offset_1), .B(0), .S(_06741_), .Y(_25772_) );
  \$mux  #( .WIDTH(32) ) _48335_ ( .A(_25772_), .B(_24362_), .S(_06742_), .Y(_25773_) );
  \$mux  #( .WIDTH(32) ) _48336_ ( .A(_25773_), .B(0), .S(_06743_), .Y(_25774_) );
  \$mux  #( .WIDTH(32) ) _48337_ ( .A(_25774_), .B(0), .S(RST), .Y(_02105_) );
  \$mux  #( .WIDTH(32) ) _48338_ ( .A(_source_stream_conv2d_16_source_28_pat_cur_offset_0), .B(0), .S(_06741_), .Y(_25775_) );
  \$mux  #( .WIDTH(32) ) _48339_ ( .A(_24361_), .B(_25775_), .S(_05966_), .Y(_25776_) );
  \$mux  #( .WIDTH(32) ) _48340_ ( .A(_25776_), .B(0), .S(_06742_), .Y(_25777_) );
  \$mux  #( .WIDTH(32) ) _48341_ ( .A(_25777_), .B(0), .S(RST), .Y(_02104_) );
  \$mux  #( .WIDTH(8) ) _48342_ ( .A(__variable_wdata_276), .B(_stream_conv2d_16_source_27_source_ram_rdata), .S(_stream_conv2d_16_source_27_source_ram_rvalid), .Y(_25778_) );
  \$mux  #( .WIDTH(8) ) _48343_ ( .A(_25778_), .B(8'h00), .S(RST), .Y(_01419_) );
  \$mux  #( .WIDTH(32) ) _48344_ ( .A(_source_stream_conv2d_16_source_27_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_27_pat_stride_3), .S(_06736_), .Y(_25779_) );
  \$mux  #( .WIDTH(32) ) _48345_ ( .A(_25779_), .B(0), .S(RST), .Y(_02099_) );
  \$mux  #( .WIDTH(32) ) _48346_ ( .A(_source_stream_conv2d_16_source_27_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_27_pat_stride_2), .S(_06736_), .Y(_25780_) );
  \$mux  #( .WIDTH(32) ) _48347_ ( .A(_25780_), .B(0), .S(RST), .Y(_02098_) );
  \$mux  #( .WIDTH(32) ) _48348_ ( .A(_source_stream_conv2d_16_source_27_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_27_pat_stride_1), .S(_06736_), .Y(_25781_) );
  \$mux  #( .WIDTH(32) ) _48349_ ( .A(_25781_), .B(0), .S(RST), .Y(_02097_) );
  \$mux  #( .WIDTH(32) ) _48350_ ( .A(_source_stream_conv2d_16_source_27_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_27_pat_stride_0), .S(_06736_), .Y(_25782_) );
  \$mux  #( .WIDTH(32) ) _48351_ ( .A(_25782_), .B(0), .S(RST), .Y(_02096_) );
  \$mux  #( .WIDTH(33) ) _48352_ ( .A(_source_stream_conv2d_16_source_27_pat_size_buf_3), .B(_source_stream_conv2d_16_source_27_pat_size_3), .S(_06736_), .Y(_25783_) );
  \$mux  #( .WIDTH(33) ) _48353_ ( .A(_25783_), .B(33'h000000000), .S(RST), .Y(_02091_) );
  \$mux  #( .WIDTH(33) ) _48354_ ( .A(_source_stream_conv2d_16_source_27_pat_size_buf_2), .B(_source_stream_conv2d_16_source_27_pat_size_2), .S(_06736_), .Y(_25784_) );
  \$mux  #( .WIDTH(33) ) _48355_ ( .A(_25784_), .B(33'h000000000), .S(RST), .Y(_02090_) );
  \$mux  #( .WIDTH(33) ) _48356_ ( .A(_source_stream_conv2d_16_source_27_pat_size_buf_1), .B(_source_stream_conv2d_16_source_27_pat_size_1), .S(_06736_), .Y(_25785_) );
  \$mux  #( .WIDTH(33) ) _48357_ ( .A(_25785_), .B(33'h000000000), .S(RST), .Y(_02089_) );
  \$mux  #( .WIDTH(33) ) _48358_ ( .A(_source_stream_conv2d_16_source_27_pat_size_buf_0), .B(_source_stream_conv2d_16_source_27_pat_size_0), .S(_06736_), .Y(_25786_) );
  \$mux  #( .WIDTH(33) ) _48359_ ( .A(_25786_), .B(33'h000000000), .S(RST), .Y(_02088_) );
  \$mux  #( .WIDTH(33) ) _48360_ ( .A(_source_stream_conv2d_16_source_27_pat_count_3), .B(_28751_), .S(_06736_), .Y(_25787_) );
  \$mux  #( .WIDTH(33) ) _48361_ ( .A(_25787_), .B(_28758_), .S(_06739_), .Y(_25788_) );
  \$mux  #( .WIDTH(33) ) _48362_ ( .A(_25788_), .B(_28759_), .S(_06740_), .Y(_25789_) );
  \$mux  #( .WIDTH(33) ) _48363_ ( .A(_25789_), .B(33'h000000000), .S(RST), .Y(_02079_) );
  \$mux  #( .WIDTH(33) ) _48364_ ( .A(_source_stream_conv2d_16_source_27_pat_count_2), .B(_28750_), .S(_06736_), .Y(_25790_) );
  \$mux  #( .WIDTH(33) ) _48365_ ( .A(_25790_), .B(_28756_), .S(_06738_), .Y(_25791_) );
  \$mux  #( .WIDTH(33) ) _48366_ ( .A(_25791_), .B(_28757_), .S(_06739_), .Y(_25792_) );
  \$mux  #( .WIDTH(33) ) _48367_ ( .A(_25792_), .B(33'h000000000), .S(RST), .Y(_02078_) );
  \$mux  #( .WIDTH(33) ) _48368_ ( .A(_source_stream_conv2d_16_source_27_pat_count_1), .B(_28749_), .S(_06736_), .Y(_25793_) );
  \$mux  #( .WIDTH(33) ) _48369_ ( .A(_25793_), .B(_28754_), .S(_06737_), .Y(_25794_) );
  \$mux  #( .WIDTH(33) ) _48370_ ( .A(_25794_), .B(_28755_), .S(_06738_), .Y(_25795_) );
  \$mux  #( .WIDTH(33) ) _48371_ ( .A(_25795_), .B(33'h000000000), .S(RST), .Y(_02077_) );
  \$mux  #( .WIDTH(33) ) _48372_ ( .A(_source_stream_conv2d_16_source_27_pat_count_0), .B(_28748_), .S(_06736_), .Y(_25796_) );
  \$mux  #( .WIDTH(33) ) _48373_ ( .A(_28752_), .B(_25796_), .S(_05968_), .Y(_25797_) );
  \$mux  #( .WIDTH(33) ) _48374_ ( .A(_25797_), .B(_28753_), .S(_06737_), .Y(_25798_) );
  \$mux  #( .WIDTH(33) ) _48375_ ( .A(_25798_), .B(33'h000000000), .S(RST), .Y(_02076_) );
  \$mux  #( .WIDTH(32) ) _48376_ ( .A(_source_stream_conv2d_16_source_27_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25799_) );
  \$mux  #( .WIDTH(32) ) _48377_ ( .A(_25799_), .B(0), .S(RST), .Y(_02095_) );
  \$mux  #( .WIDTH(32) ) _48378_ ( .A(_source_stream_conv2d_16_source_27_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25800_) );
  \$mux  #( .WIDTH(32) ) _48379_ ( .A(_25800_), .B(0), .S(RST), .Y(_02094_) );
  \$mux  #( .WIDTH(32) ) _48380_ ( .A(_source_stream_conv2d_16_source_27_pat_stride_1), .B(0), .S(_set_flag_710), .Y(_25801_) );
  \$mux  #( .WIDTH(32) ) _48381_ ( .A(_25801_), .B(0), .S(RST), .Y(_02093_) );
  \$mux  #( .WIDTH(32) ) _48382_ ( .A(_source_stream_conv2d_16_source_27_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25802_) );
  \$mux  #( .WIDTH(32) ) _48383_ ( .A(_25802_), .B(0), .S(RST), .Y(_02092_) );
  \$mux  #( .WIDTH(33) ) _48384_ ( .A(_source_stream_conv2d_16_source_27_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25803_) );
  \$mux  #( .WIDTH(33) ) _48385_ ( .A(_25803_), .B(33'h000000000), .S(RST), .Y(_02087_) );
  \$mux  #( .WIDTH(33) ) _48386_ ( .A(_source_stream_conv2d_16_source_27_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25804_) );
  \$mux  #( .WIDTH(33) ) _48387_ ( .A(_25804_), .B(33'h000000000), .S(RST), .Y(_02086_) );
  \$mux  #( .WIDTH(33) ) _48388_ ( .A(_source_stream_conv2d_16_source_27_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25805_) );
  \$mux  #( .WIDTH(33) ) _48389_ ( .A(_25805_), .B(33'h000000000), .S(RST), .Y(_02085_) );
  \$mux  #( .WIDTH(33) ) _48390_ ( .A(_source_stream_conv2d_16_source_27_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25806_) );
  \$mux  #( .WIDTH(33) ) _48391_ ( .A(_25806_), .B(33'h000000000), .S(RST), .Y(_02084_) );
  \$mux  #( .WIDTH(32) ) _48392_ ( .A(_source_stream_conv2d_16_source_27_pat_cur_offset_3), .B(0), .S(_06736_), .Y(_25807_) );
  \$mux  #( .WIDTH(32) ) _48393_ ( .A(_25807_), .B(_24360_), .S(_06739_), .Y(_25808_) );
  \$mux  #( .WIDTH(32) ) _48394_ ( .A(_25808_), .B(0), .S(_06740_), .Y(_25809_) );
  \$mux  #( .WIDTH(32) ) _48395_ ( .A(_25809_), .B(0), .S(RST), .Y(_02083_) );
  \$mux  #( .WIDTH(32) ) _48396_ ( .A(_source_stream_conv2d_16_source_27_pat_cur_offset_2), .B(0), .S(_06736_), .Y(_25810_) );
  \$mux  #( .WIDTH(32) ) _48397_ ( .A(_25810_), .B(_24359_), .S(_06738_), .Y(_25811_) );
  \$mux  #( .WIDTH(32) ) _48398_ ( .A(_25811_), .B(0), .S(_06739_), .Y(_25812_) );
  \$mux  #( .WIDTH(32) ) _48399_ ( .A(_25812_), .B(0), .S(RST), .Y(_02082_) );
  \$mux  #( .WIDTH(32) ) _48400_ ( .A(_source_stream_conv2d_16_source_27_pat_cur_offset_1), .B(0), .S(_06736_), .Y(_25813_) );
  \$mux  #( .WIDTH(32) ) _48401_ ( .A(_25813_), .B(_24358_), .S(_06737_), .Y(_25814_) );
  \$mux  #( .WIDTH(32) ) _48402_ ( .A(_25814_), .B(0), .S(_06738_), .Y(_25815_) );
  \$mux  #( .WIDTH(32) ) _48403_ ( .A(_25815_), .B(0), .S(RST), .Y(_02081_) );
  \$mux  #( .WIDTH(32) ) _48404_ ( .A(_source_stream_conv2d_16_source_27_pat_cur_offset_0), .B(0), .S(_06736_), .Y(_25816_) );
  \$mux  #( .WIDTH(32) ) _48405_ ( .A(_24357_), .B(_25816_), .S(_05968_), .Y(_25817_) );
  \$mux  #( .WIDTH(32) ) _48406_ ( .A(_25817_), .B(0), .S(_06737_), .Y(_25818_) );
  \$mux  #( .WIDTH(32) ) _48407_ ( .A(_25818_), .B(0), .S(RST), .Y(_02080_) );
  \$mux  #( .WIDTH(8) ) _48408_ ( .A(__variable_wdata_275), .B(_stream_conv2d_16_source_26_source_ram_rdata), .S(_stream_conv2d_16_source_26_source_ram_rvalid), .Y(_25819_) );
  \$mux  #( .WIDTH(8) ) _48409_ ( .A(_25819_), .B(8'h00), .S(RST), .Y(_01418_) );
  \$mux  #( .WIDTH(32) ) _48410_ ( .A(_source_stream_conv2d_16_source_26_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_26_pat_stride_3), .S(_06731_), .Y(_25820_) );
  \$mux  #( .WIDTH(32) ) _48411_ ( .A(_25820_), .B(0), .S(RST), .Y(_02075_) );
  \$mux  #( .WIDTH(32) ) _48412_ ( .A(_source_stream_conv2d_16_source_26_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_26_pat_stride_2), .S(_06731_), .Y(_25821_) );
  \$mux  #( .WIDTH(32) ) _48413_ ( .A(_25821_), .B(0), .S(RST), .Y(_02074_) );
  \$mux  #( .WIDTH(32) ) _48414_ ( .A(_source_stream_conv2d_16_source_26_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_26_pat_stride_1), .S(_06731_), .Y(_25822_) );
  \$mux  #( .WIDTH(32) ) _48415_ ( .A(_25822_), .B(0), .S(RST), .Y(_02073_) );
  \$mux  #( .WIDTH(32) ) _48416_ ( .A(_source_stream_conv2d_16_source_26_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_26_pat_stride_0), .S(_06731_), .Y(_25823_) );
  \$mux  #( .WIDTH(32) ) _48417_ ( .A(_25823_), .B(0), .S(RST), .Y(_02072_) );
  \$mux  #( .WIDTH(33) ) _48418_ ( .A(_source_stream_conv2d_16_source_26_pat_size_buf_3), .B(_source_stream_conv2d_16_source_26_pat_size_3), .S(_06731_), .Y(_25824_) );
  \$mux  #( .WIDTH(33) ) _48419_ ( .A(_25824_), .B(33'h000000000), .S(RST), .Y(_02067_) );
  \$mux  #( .WIDTH(33) ) _48420_ ( .A(_source_stream_conv2d_16_source_26_pat_size_buf_2), .B(_source_stream_conv2d_16_source_26_pat_size_2), .S(_06731_), .Y(_25825_) );
  \$mux  #( .WIDTH(33) ) _48421_ ( .A(_25825_), .B(33'h000000000), .S(RST), .Y(_02066_) );
  \$mux  #( .WIDTH(33) ) _48422_ ( .A(_source_stream_conv2d_16_source_26_pat_size_buf_1), .B(_source_stream_conv2d_16_source_26_pat_size_1), .S(_06731_), .Y(_25826_) );
  \$mux  #( .WIDTH(33) ) _48423_ ( .A(_25826_), .B(33'h000000000), .S(RST), .Y(_02065_) );
  \$mux  #( .WIDTH(33) ) _48424_ ( .A(_source_stream_conv2d_16_source_26_pat_size_buf_0), .B(_source_stream_conv2d_16_source_26_pat_size_0), .S(_06731_), .Y(_25827_) );
  \$mux  #( .WIDTH(33) ) _48425_ ( .A(_25827_), .B(33'h000000000), .S(RST), .Y(_02064_) );
  \$mux  #( .WIDTH(33) ) _48426_ ( .A(_source_stream_conv2d_16_source_26_pat_count_3), .B(_28739_), .S(_06731_), .Y(_25828_) );
  \$mux  #( .WIDTH(33) ) _48427_ ( .A(_25828_), .B(_28746_), .S(_06734_), .Y(_25829_) );
  \$mux  #( .WIDTH(33) ) _48428_ ( .A(_25829_), .B(_28747_), .S(_06735_), .Y(_25830_) );
  \$mux  #( .WIDTH(33) ) _48429_ ( .A(_25830_), .B(33'h000000000), .S(RST), .Y(_02055_) );
  \$mux  #( .WIDTH(33) ) _48430_ ( .A(_source_stream_conv2d_16_source_26_pat_count_2), .B(_28738_), .S(_06731_), .Y(_25831_) );
  \$mux  #( .WIDTH(33) ) _48431_ ( .A(_25831_), .B(_28744_), .S(_06733_), .Y(_25832_) );
  \$mux  #( .WIDTH(33) ) _48432_ ( .A(_25832_), .B(_28745_), .S(_06734_), .Y(_25833_) );
  \$mux  #( .WIDTH(33) ) _48433_ ( .A(_25833_), .B(33'h000000000), .S(RST), .Y(_02054_) );
  \$mux  #( .WIDTH(33) ) _48434_ ( .A(_source_stream_conv2d_16_source_26_pat_count_1), .B(_28737_), .S(_06731_), .Y(_25834_) );
  \$mux  #( .WIDTH(33) ) _48435_ ( .A(_25834_), .B(_28742_), .S(_06732_), .Y(_25835_) );
  \$mux  #( .WIDTH(33) ) _48436_ ( .A(_25835_), .B(_28743_), .S(_06733_), .Y(_25836_) );
  \$mux  #( .WIDTH(33) ) _48437_ ( .A(_25836_), .B(33'h000000000), .S(RST), .Y(_02053_) );
  \$mux  #( .WIDTH(33) ) _48438_ ( .A(_source_stream_conv2d_16_source_26_pat_count_0), .B(_28736_), .S(_06731_), .Y(_25837_) );
  \$mux  #( .WIDTH(33) ) _48439_ ( .A(_28740_), .B(_25837_), .S(_05971_), .Y(_25838_) );
  \$mux  #( .WIDTH(33) ) _48440_ ( .A(_25838_), .B(_28741_), .S(_06732_), .Y(_25839_) );
  \$mux  #( .WIDTH(33) ) _48441_ ( .A(_25839_), .B(33'h000000000), .S(RST), .Y(_02052_) );
  \$mux  #( .WIDTH(32) ) _48442_ ( .A(_source_stream_conv2d_16_source_26_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25840_) );
  \$mux  #( .WIDTH(32) ) _48443_ ( .A(_25840_), .B(0), .S(RST), .Y(_02071_) );
  \$mux  #( .WIDTH(32) ) _48444_ ( .A(_source_stream_conv2d_16_source_26_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25841_) );
  \$mux  #( .WIDTH(32) ) _48445_ ( .A(_25841_), .B(0), .S(RST), .Y(_02070_) );
  \$mux  #( .WIDTH(32) ) _48446_ ( .A(_source_stream_conv2d_16_source_26_pat_stride_1), .B(0), .S(_set_flag_710), .Y(_25842_) );
  \$mux  #( .WIDTH(32) ) _48447_ ( .A(_25842_), .B(0), .S(RST), .Y(_02069_) );
  \$mux  #( .WIDTH(32) ) _48448_ ( .A(_source_stream_conv2d_16_source_26_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25843_) );
  \$mux  #( .WIDTH(32) ) _48449_ ( .A(_25843_), .B(0), .S(RST), .Y(_02068_) );
  \$mux  #( .WIDTH(33) ) _48450_ ( .A(_source_stream_conv2d_16_source_26_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25844_) );
  \$mux  #( .WIDTH(33) ) _48451_ ( .A(_25844_), .B(33'h000000000), .S(RST), .Y(_02063_) );
  \$mux  #( .WIDTH(33) ) _48452_ ( .A(_source_stream_conv2d_16_source_26_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25845_) );
  \$mux  #( .WIDTH(33) ) _48453_ ( .A(_25845_), .B(33'h000000000), .S(RST), .Y(_02062_) );
  \$mux  #( .WIDTH(33) ) _48454_ ( .A(_source_stream_conv2d_16_source_26_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25846_) );
  \$mux  #( .WIDTH(33) ) _48455_ ( .A(_25846_), .B(33'h000000000), .S(RST), .Y(_02061_) );
  \$mux  #( .WIDTH(33) ) _48456_ ( .A(_source_stream_conv2d_16_source_26_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25847_) );
  \$mux  #( .WIDTH(33) ) _48457_ ( .A(_25847_), .B(33'h000000000), .S(RST), .Y(_02060_) );
  \$mux  #( .WIDTH(32) ) _48458_ ( .A(_source_stream_conv2d_16_source_26_pat_cur_offset_3), .B(0), .S(_06731_), .Y(_25848_) );
  \$mux  #( .WIDTH(32) ) _48459_ ( .A(_25848_), .B(_24355_), .S(_06734_), .Y(_25849_) );
  \$mux  #( .WIDTH(32) ) _48460_ ( .A(_25849_), .B(0), .S(_06735_), .Y(_25850_) );
  \$mux  #( .WIDTH(32) ) _48461_ ( .A(_25850_), .B(0), .S(RST), .Y(_02059_) );
  \$mux  #( .WIDTH(32) ) _48462_ ( .A(_source_stream_conv2d_16_source_26_pat_cur_offset_2), .B(0), .S(_06731_), .Y(_25851_) );
  \$mux  #( .WIDTH(32) ) _48463_ ( .A(_25851_), .B(_24354_), .S(_06733_), .Y(_25852_) );
  \$mux  #( .WIDTH(32) ) _48464_ ( .A(_25852_), .B(0), .S(_06734_), .Y(_25853_) );
  \$mux  #( .WIDTH(32) ) _48465_ ( .A(_25853_), .B(0), .S(RST), .Y(_02058_) );
  \$mux  #( .WIDTH(32) ) _48466_ ( .A(_source_stream_conv2d_16_source_26_pat_cur_offset_1), .B(0), .S(_06731_), .Y(_25854_) );
  \$mux  #( .WIDTH(32) ) _48467_ ( .A(_25854_), .B(_24353_), .S(_06732_), .Y(_25855_) );
  \$mux  #( .WIDTH(32) ) _48468_ ( .A(_25855_), .B(0), .S(_06733_), .Y(_25856_) );
  \$mux  #( .WIDTH(32) ) _48469_ ( .A(_25856_), .B(0), .S(RST), .Y(_02057_) );
  \$mux  #( .WIDTH(32) ) _48470_ ( .A(_source_stream_conv2d_16_source_26_pat_cur_offset_0), .B(0), .S(_06731_), .Y(_25857_) );
  \$mux  #( .WIDTH(32) ) _48471_ ( .A(_24352_), .B(_25857_), .S(_05971_), .Y(_25858_) );
  \$mux  #( .WIDTH(32) ) _48472_ ( .A(_25858_), .B(0), .S(_06732_), .Y(_25859_) );
  \$mux  #( .WIDTH(32) ) _48473_ ( .A(_25859_), .B(0), .S(RST), .Y(_02056_) );
  \$mux  #( .WIDTH(8) ) _48474_ ( .A(__variable_wdata_274), .B(_stream_conv2d_16_source_25_source_ram_rdata), .S(_stream_conv2d_16_source_25_source_ram_rvalid), .Y(_25860_) );
  \$mux  #( .WIDTH(8) ) _48475_ ( .A(_25860_), .B(8'h00), .S(RST), .Y(_01417_) );
  \$mux  #( .WIDTH(32) ) _48476_ ( .A(_source_stream_conv2d_16_source_25_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_25_pat_stride_3), .S(_06726_), .Y(_25861_) );
  \$mux  #( .WIDTH(32) ) _48477_ ( .A(_25861_), .B(0), .S(RST), .Y(_02051_) );
  \$mux  #( .WIDTH(32) ) _48478_ ( .A(_source_stream_conv2d_16_source_25_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_25_pat_stride_2), .S(_06726_), .Y(_25862_) );
  \$mux  #( .WIDTH(32) ) _48479_ ( .A(_25862_), .B(0), .S(RST), .Y(_02050_) );
  \$mux  #( .WIDTH(32) ) _48480_ ( .A(_source_stream_conv2d_16_source_25_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_25_pat_stride_1), .S(_06726_), .Y(_25863_) );
  \$mux  #( .WIDTH(32) ) _48481_ ( .A(_25863_), .B(0), .S(RST), .Y(_02049_) );
  \$mux  #( .WIDTH(32) ) _48482_ ( .A(_source_stream_conv2d_16_source_25_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_25_pat_stride_0), .S(_06726_), .Y(_25864_) );
  \$mux  #( .WIDTH(32) ) _48483_ ( .A(_25864_), .B(0), .S(RST), .Y(_02048_) );
  \$mux  #( .WIDTH(33) ) _48484_ ( .A(_source_stream_conv2d_16_source_25_pat_size_buf_3), .B(_source_stream_conv2d_16_source_25_pat_size_3), .S(_06726_), .Y(_25865_) );
  \$mux  #( .WIDTH(33) ) _48485_ ( .A(_25865_), .B(33'h000000000), .S(RST), .Y(_02043_) );
  \$mux  #( .WIDTH(33) ) _48486_ ( .A(_source_stream_conv2d_16_source_25_pat_size_buf_2), .B(_source_stream_conv2d_16_source_25_pat_size_2), .S(_06726_), .Y(_25866_) );
  \$mux  #( .WIDTH(33) ) _48487_ ( .A(_25866_), .B(33'h000000000), .S(RST), .Y(_02042_) );
  \$mux  #( .WIDTH(33) ) _48488_ ( .A(_source_stream_conv2d_16_source_25_pat_size_buf_1), .B(_source_stream_conv2d_16_source_25_pat_size_1), .S(_06726_), .Y(_25867_) );
  \$mux  #( .WIDTH(33) ) _48489_ ( .A(_25867_), .B(33'h000000000), .S(RST), .Y(_02041_) );
  \$mux  #( .WIDTH(33) ) _48490_ ( .A(_source_stream_conv2d_16_source_25_pat_size_buf_0), .B(_source_stream_conv2d_16_source_25_pat_size_0), .S(_06726_), .Y(_25868_) );
  \$mux  #( .WIDTH(33) ) _48491_ ( .A(_25868_), .B(33'h000000000), .S(RST), .Y(_02040_) );
  \$mux  #( .WIDTH(33) ) _48492_ ( .A(_source_stream_conv2d_16_source_25_pat_count_3), .B(_28727_), .S(_06726_), .Y(_25869_) );
  \$mux  #( .WIDTH(33) ) _48493_ ( .A(_25869_), .B(_28734_), .S(_06729_), .Y(_25870_) );
  \$mux  #( .WIDTH(33) ) _48494_ ( .A(_25870_), .B(_28735_), .S(_06730_), .Y(_25871_) );
  \$mux  #( .WIDTH(33) ) _48495_ ( .A(_25871_), .B(33'h000000000), .S(RST), .Y(_02031_) );
  \$mux  #( .WIDTH(33) ) _48496_ ( .A(_source_stream_conv2d_16_source_25_pat_count_2), .B(_28726_), .S(_06726_), .Y(_25872_) );
  \$mux  #( .WIDTH(33) ) _48497_ ( .A(_25872_), .B(_28732_), .S(_06728_), .Y(_25873_) );
  \$mux  #( .WIDTH(33) ) _48498_ ( .A(_25873_), .B(_28733_), .S(_06729_), .Y(_25874_) );
  \$mux  #( .WIDTH(33) ) _48499_ ( .A(_25874_), .B(33'h000000000), .S(RST), .Y(_02030_) );
  \$mux  #( .WIDTH(33) ) _48500_ ( .A(_source_stream_conv2d_16_source_25_pat_count_1), .B(_28725_), .S(_06726_), .Y(_25875_) );
  \$mux  #( .WIDTH(33) ) _48501_ ( .A(_25875_), .B(_28730_), .S(_06727_), .Y(_25876_) );
  \$mux  #( .WIDTH(33) ) _48502_ ( .A(_25876_), .B(_28731_), .S(_06728_), .Y(_25877_) );
  \$mux  #( .WIDTH(33) ) _48503_ ( .A(_25877_), .B(33'h000000000), .S(RST), .Y(_02029_) );
  \$mux  #( .WIDTH(33) ) _48504_ ( .A(_source_stream_conv2d_16_source_25_pat_count_0), .B(_28724_), .S(_06726_), .Y(_25878_) );
  \$mux  #( .WIDTH(33) ) _48505_ ( .A(_28728_), .B(_25878_), .S(_05974_), .Y(_25879_) );
  \$mux  #( .WIDTH(33) ) _48506_ ( .A(_25879_), .B(_28729_), .S(_06727_), .Y(_25880_) );
  \$mux  #( .WIDTH(33) ) _48507_ ( .A(_25880_), .B(33'h000000000), .S(RST), .Y(_02028_) );
  \$mux  #( .WIDTH(32) ) _48508_ ( .A(_source_stream_conv2d_16_source_25_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25881_) );
  \$mux  #( .WIDTH(32) ) _48509_ ( .A(_25881_), .B(0), .S(RST), .Y(_02047_) );
  \$mux  #( .WIDTH(32) ) _48510_ ( .A(_source_stream_conv2d_16_source_25_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25882_) );
  \$mux  #( .WIDTH(32) ) _48511_ ( .A(_25882_), .B(0), .S(RST), .Y(_02046_) );
  \$mux  #( .WIDTH(32) ) _48512_ ( .A(_source_stream_conv2d_16_source_25_pat_stride_1), .B(0), .S(_set_flag_710), .Y(_25883_) );
  \$mux  #( .WIDTH(32) ) _48513_ ( .A(_25883_), .B(0), .S(RST), .Y(_02045_) );
  \$mux  #( .WIDTH(32) ) _48514_ ( .A(_source_stream_conv2d_16_source_25_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25884_) );
  \$mux  #( .WIDTH(32) ) _48515_ ( .A(_25884_), .B(0), .S(RST), .Y(_02044_) );
  \$mux  #( .WIDTH(33) ) _48516_ ( .A(_source_stream_conv2d_16_source_25_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25885_) );
  \$mux  #( .WIDTH(33) ) _48517_ ( .A(_25885_), .B(33'h000000000), .S(RST), .Y(_02039_) );
  \$mux  #( .WIDTH(33) ) _48518_ ( .A(_source_stream_conv2d_16_source_25_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25886_) );
  \$mux  #( .WIDTH(33) ) _48519_ ( .A(_25886_), .B(33'h000000000), .S(RST), .Y(_02038_) );
  \$mux  #( .WIDTH(33) ) _48520_ ( .A(_source_stream_conv2d_16_source_25_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25887_) );
  \$mux  #( .WIDTH(33) ) _48521_ ( .A(_25887_), .B(33'h000000000), .S(RST), .Y(_02037_) );
  \$mux  #( .WIDTH(33) ) _48522_ ( .A(_source_stream_conv2d_16_source_25_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25888_) );
  \$mux  #( .WIDTH(33) ) _48523_ ( .A(_25888_), .B(33'h000000000), .S(RST), .Y(_02036_) );
  \$mux  #( .WIDTH(32) ) _48524_ ( .A(_source_stream_conv2d_16_source_25_pat_cur_offset_3), .B(0), .S(_06726_), .Y(_25889_) );
  \$mux  #( .WIDTH(32) ) _48525_ ( .A(_25889_), .B(_24350_), .S(_06729_), .Y(_25890_) );
  \$mux  #( .WIDTH(32) ) _48526_ ( .A(_25890_), .B(0), .S(_06730_), .Y(_25891_) );
  \$mux  #( .WIDTH(32) ) _48527_ ( .A(_25891_), .B(0), .S(RST), .Y(_02035_) );
  \$mux  #( .WIDTH(32) ) _48528_ ( .A(_source_stream_conv2d_16_source_25_pat_cur_offset_2), .B(0), .S(_06726_), .Y(_25892_) );
  \$mux  #( .WIDTH(32) ) _48529_ ( .A(_25892_), .B(_24349_), .S(_06728_), .Y(_25893_) );
  \$mux  #( .WIDTH(32) ) _48530_ ( .A(_25893_), .B(0), .S(_06729_), .Y(_25894_) );
  \$mux  #( .WIDTH(32) ) _48531_ ( .A(_25894_), .B(0), .S(RST), .Y(_02034_) );
  \$mux  #( .WIDTH(32) ) _48532_ ( .A(_source_stream_conv2d_16_source_25_pat_cur_offset_1), .B(0), .S(_06726_), .Y(_25895_) );
  \$mux  #( .WIDTH(32) ) _48533_ ( .A(_25895_), .B(_24348_), .S(_06727_), .Y(_25896_) );
  \$mux  #( .WIDTH(32) ) _48534_ ( .A(_25896_), .B(0), .S(_06728_), .Y(_25897_) );
  \$mux  #( .WIDTH(32) ) _48535_ ( .A(_25897_), .B(0), .S(RST), .Y(_02033_) );
  \$mux  #( .WIDTH(32) ) _48536_ ( .A(_source_stream_conv2d_16_source_25_pat_cur_offset_0), .B(0), .S(_06726_), .Y(_25898_) );
  \$mux  #( .WIDTH(32) ) _48537_ ( .A(_24347_), .B(_25898_), .S(_05974_), .Y(_25899_) );
  \$mux  #( .WIDTH(32) ) _48538_ ( .A(_25899_), .B(0), .S(_06727_), .Y(_25900_) );
  \$mux  #( .WIDTH(32) ) _48539_ ( .A(_25900_), .B(0), .S(RST), .Y(_02032_) );
  \$mux  #( .WIDTH(8) ) _48540_ ( .A(__variable_wdata_273), .B(_stream_conv2d_16_source_24_source_ram_rdata), .S(_stream_conv2d_16_source_24_source_ram_rvalid), .Y(_25901_) );
  \$mux  #( .WIDTH(8) ) _48541_ ( .A(_25901_), .B(8'h00), .S(RST), .Y(_01416_) );
  \$mux  #( .WIDTH(32) ) _48542_ ( .A(_source_stream_conv2d_16_source_24_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_24_pat_stride_3), .S(_06721_), .Y(_25902_) );
  \$mux  #( .WIDTH(32) ) _48543_ ( .A(_25902_), .B(0), .S(RST), .Y(_02027_) );
  \$mux  #( .WIDTH(32) ) _48544_ ( .A(_source_stream_conv2d_16_source_24_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_24_pat_stride_2), .S(_06721_), .Y(_25903_) );
  \$mux  #( .WIDTH(32) ) _48545_ ( .A(_25903_), .B(0), .S(RST), .Y(_02026_) );
  \$mux  #( .WIDTH(32) ) _48546_ ( .A(_source_stream_conv2d_16_source_24_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_24_pat_stride_1), .S(_06721_), .Y(_25904_) );
  \$mux  #( .WIDTH(32) ) _48547_ ( .A(_25904_), .B(0), .S(RST), .Y(_02025_) );
  \$mux  #( .WIDTH(32) ) _48548_ ( .A(_source_stream_conv2d_16_source_24_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_24_pat_stride_0), .S(_06721_), .Y(_25905_) );
  \$mux  #( .WIDTH(32) ) _48549_ ( .A(_25905_), .B(0), .S(RST), .Y(_02024_) );
  \$mux  #( .WIDTH(33) ) _48550_ ( .A(_source_stream_conv2d_16_source_24_pat_size_buf_3), .B(_source_stream_conv2d_16_source_24_pat_size_3), .S(_06721_), .Y(_25906_) );
  \$mux  #( .WIDTH(33) ) _48551_ ( .A(_25906_), .B(33'h000000000), .S(RST), .Y(_02019_) );
  \$mux  #( .WIDTH(33) ) _48552_ ( .A(_source_stream_conv2d_16_source_24_pat_size_buf_2), .B(_source_stream_conv2d_16_source_24_pat_size_2), .S(_06721_), .Y(_25907_) );
  \$mux  #( .WIDTH(33) ) _48553_ ( .A(_25907_), .B(33'h000000000), .S(RST), .Y(_02018_) );
  \$mux  #( .WIDTH(33) ) _48554_ ( .A(_source_stream_conv2d_16_source_24_pat_size_buf_1), .B(_source_stream_conv2d_16_source_24_pat_size_1), .S(_06721_), .Y(_25908_) );
  \$mux  #( .WIDTH(33) ) _48555_ ( .A(_25908_), .B(33'h000000000), .S(RST), .Y(_02017_) );
  \$mux  #( .WIDTH(33) ) _48556_ ( .A(_source_stream_conv2d_16_source_24_pat_size_buf_0), .B(_source_stream_conv2d_16_source_24_pat_size_0), .S(_06721_), .Y(_25909_) );
  \$mux  #( .WIDTH(33) ) _48557_ ( .A(_25909_), .B(33'h000000000), .S(RST), .Y(_02016_) );
  \$mux  #( .WIDTH(33) ) _48558_ ( .A(_source_stream_conv2d_16_source_24_pat_count_3), .B(_28715_), .S(_06721_), .Y(_25910_) );
  \$mux  #( .WIDTH(33) ) _48559_ ( .A(_25910_), .B(_28722_), .S(_06724_), .Y(_25911_) );
  \$mux  #( .WIDTH(33) ) _48560_ ( .A(_25911_), .B(_28723_), .S(_06725_), .Y(_25912_) );
  \$mux  #( .WIDTH(33) ) _48561_ ( .A(_25912_), .B(33'h000000000), .S(RST), .Y(_02007_) );
  \$mux  #( .WIDTH(33) ) _48562_ ( .A(_source_stream_conv2d_16_source_24_pat_count_2), .B(_28714_), .S(_06721_), .Y(_25913_) );
  \$mux  #( .WIDTH(33) ) _48563_ ( .A(_25913_), .B(_28720_), .S(_06723_), .Y(_25914_) );
  \$mux  #( .WIDTH(33) ) _48564_ ( .A(_25914_), .B(_28721_), .S(_06724_), .Y(_25915_) );
  \$mux  #( .WIDTH(33) ) _48565_ ( .A(_25915_), .B(33'h000000000), .S(RST), .Y(_02006_) );
  \$mux  #( .WIDTH(33) ) _48566_ ( .A(_source_stream_conv2d_16_source_24_pat_count_1), .B(_28713_), .S(_06721_), .Y(_25916_) );
  \$mux  #( .WIDTH(33) ) _48567_ ( .A(_25916_), .B(_28718_), .S(_06722_), .Y(_25917_) );
  \$mux  #( .WIDTH(33) ) _48568_ ( .A(_25917_), .B(_28719_), .S(_06723_), .Y(_25918_) );
  \$mux  #( .WIDTH(33) ) _48569_ ( .A(_25918_), .B(33'h000000000), .S(RST), .Y(_02005_) );
  \$mux  #( .WIDTH(33) ) _48570_ ( .A(_source_stream_conv2d_16_source_24_pat_count_0), .B(_28712_), .S(_06721_), .Y(_25919_) );
  \$mux  #( .WIDTH(33) ) _48571_ ( .A(_28716_), .B(_25919_), .S(_05972_), .Y(_25920_) );
  \$mux  #( .WIDTH(33) ) _48572_ ( .A(_25920_), .B(_28717_), .S(_06722_), .Y(_25921_) );
  \$mux  #( .WIDTH(33) ) _48573_ ( .A(_25921_), .B(33'h000000000), .S(RST), .Y(_02004_) );
  \$mux  #( .WIDTH(32) ) _48574_ ( .A(_source_stream_conv2d_16_source_24_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25922_) );
  \$mux  #( .WIDTH(32) ) _48575_ ( .A(_25922_), .B(0), .S(RST), .Y(_02023_) );
  \$mux  #( .WIDTH(32) ) _48576_ ( .A(_source_stream_conv2d_16_source_24_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25923_) );
  \$mux  #( .WIDTH(32) ) _48577_ ( .A(_25923_), .B(0), .S(RST), .Y(_02022_) );
  \$mux  #( .WIDTH(32) ) _48578_ ( .A(_source_stream_conv2d_16_source_24_pat_stride_1), .B(0), .S(_set_flag_710), .Y(_25924_) );
  \$mux  #( .WIDTH(32) ) _48579_ ( .A(_25924_), .B(0), .S(RST), .Y(_02021_) );
  \$mux  #( .WIDTH(32) ) _48580_ ( .A(_source_stream_conv2d_16_source_24_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25925_) );
  \$mux  #( .WIDTH(32) ) _48581_ ( .A(_25925_), .B(0), .S(RST), .Y(_02020_) );
  \$mux  #( .WIDTH(33) ) _48582_ ( .A(_source_stream_conv2d_16_source_24_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25926_) );
  \$mux  #( .WIDTH(33) ) _48583_ ( .A(_25926_), .B(33'h000000000), .S(RST), .Y(_02015_) );
  \$mux  #( .WIDTH(33) ) _48584_ ( .A(_source_stream_conv2d_16_source_24_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25927_) );
  \$mux  #( .WIDTH(33) ) _48585_ ( .A(_25927_), .B(33'h000000000), .S(RST), .Y(_02014_) );
  \$mux  #( .WIDTH(33) ) _48586_ ( .A(_source_stream_conv2d_16_source_24_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25928_) );
  \$mux  #( .WIDTH(33) ) _48587_ ( .A(_25928_), .B(33'h000000000), .S(RST), .Y(_02013_) );
  \$mux  #( .WIDTH(33) ) _48588_ ( .A(_source_stream_conv2d_16_source_24_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25929_) );
  \$mux  #( .WIDTH(33) ) _48589_ ( .A(_25929_), .B(33'h000000000), .S(RST), .Y(_02012_) );
  \$mux  #( .WIDTH(32) ) _48590_ ( .A(_source_stream_conv2d_16_source_24_pat_cur_offset_3), .B(0), .S(_06721_), .Y(_25930_) );
  \$mux  #( .WIDTH(32) ) _48591_ ( .A(_25930_), .B(_24345_), .S(_06724_), .Y(_25931_) );
  \$mux  #( .WIDTH(32) ) _48592_ ( .A(_25931_), .B(0), .S(_06725_), .Y(_25932_) );
  \$mux  #( .WIDTH(32) ) _48593_ ( .A(_25932_), .B(0), .S(RST), .Y(_02011_) );
  \$mux  #( .WIDTH(32) ) _48594_ ( .A(_source_stream_conv2d_16_source_24_pat_cur_offset_2), .B(0), .S(_06721_), .Y(_25933_) );
  \$mux  #( .WIDTH(32) ) _48595_ ( .A(_25933_), .B(_24344_), .S(_06723_), .Y(_25934_) );
  \$mux  #( .WIDTH(32) ) _48596_ ( .A(_25934_), .B(0), .S(_06724_), .Y(_25935_) );
  \$mux  #( .WIDTH(32) ) _48597_ ( .A(_25935_), .B(0), .S(RST), .Y(_02010_) );
  \$mux  #( .WIDTH(32) ) _48598_ ( .A(_source_stream_conv2d_16_source_24_pat_cur_offset_1), .B(0), .S(_06721_), .Y(_25936_) );
  \$mux  #( .WIDTH(32) ) _48599_ ( .A(_25936_), .B(_24343_), .S(_06722_), .Y(_25937_) );
  \$mux  #( .WIDTH(32) ) _48600_ ( .A(_25937_), .B(0), .S(_06723_), .Y(_25938_) );
  \$mux  #( .WIDTH(32) ) _48601_ ( .A(_25938_), .B(0), .S(RST), .Y(_02009_) );
  \$mux  #( .WIDTH(32) ) _48602_ ( .A(_source_stream_conv2d_16_source_24_pat_cur_offset_0), .B(0), .S(_06721_), .Y(_25939_) );
  \$mux  #( .WIDTH(32) ) _48603_ ( .A(_24342_), .B(_25939_), .S(_05972_), .Y(_25940_) );
  \$mux  #( .WIDTH(32) ) _48604_ ( .A(_25940_), .B(0), .S(_06722_), .Y(_25941_) );
  \$mux  #( .WIDTH(32) ) _48605_ ( .A(_25941_), .B(0), .S(RST), .Y(_02008_) );
  \$mux  #( .WIDTH(8) ) _48606_ ( .A(__variable_wdata_272), .B(_stream_conv2d_16_source_23_source_ram_rdata), .S(_stream_conv2d_16_source_23_source_ram_rvalid), .Y(_25942_) );
  \$mux  #( .WIDTH(8) ) _48607_ ( .A(_25942_), .B(8'h00), .S(RST), .Y(_01415_) );
  \$mux  #( .WIDTH(32) ) _48608_ ( .A(_source_stream_conv2d_16_source_23_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_23_pat_stride_3), .S(_06716_), .Y(_25943_) );
  \$mux  #( .WIDTH(32) ) _48609_ ( .A(_25943_), .B(0), .S(RST), .Y(_02003_) );
  \$mux  #( .WIDTH(32) ) _48610_ ( .A(_source_stream_conv2d_16_source_23_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_23_pat_stride_2), .S(_06716_), .Y(_25944_) );
  \$mux  #( .WIDTH(32) ) _48611_ ( .A(_25944_), .B(0), .S(RST), .Y(_02002_) );
  \$mux  #( .WIDTH(32) ) _48612_ ( .A(_source_stream_conv2d_16_source_23_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_23_pat_stride_1), .S(_06716_), .Y(_25945_) );
  \$mux  #( .WIDTH(32) ) _48613_ ( .A(_25945_), .B(0), .S(RST), .Y(_02001_) );
  \$mux  #( .WIDTH(32) ) _48614_ ( .A(_source_stream_conv2d_16_source_23_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_23_pat_stride_0), .S(_06716_), .Y(_25946_) );
  \$mux  #( .WIDTH(32) ) _48615_ ( .A(_25946_), .B(0), .S(RST), .Y(_02000_) );
  \$mux  #( .WIDTH(33) ) _48616_ ( .A(_source_stream_conv2d_16_source_23_pat_size_buf_3), .B(_source_stream_conv2d_16_source_23_pat_size_3), .S(_06716_), .Y(_25947_) );
  \$mux  #( .WIDTH(33) ) _48617_ ( .A(_25947_), .B(33'h000000000), .S(RST), .Y(_01995_) );
  \$mux  #( .WIDTH(33) ) _48618_ ( .A(_source_stream_conv2d_16_source_23_pat_size_buf_2), .B(_source_stream_conv2d_16_source_23_pat_size_2), .S(_06716_), .Y(_25948_) );
  \$mux  #( .WIDTH(33) ) _48619_ ( .A(_25948_), .B(33'h000000000), .S(RST), .Y(_01994_) );
  \$mux  #( .WIDTH(33) ) _48620_ ( .A(_source_stream_conv2d_16_source_23_pat_size_buf_1), .B(_source_stream_conv2d_16_source_23_pat_size_1), .S(_06716_), .Y(_25949_) );
  \$mux  #( .WIDTH(33) ) _48621_ ( .A(_25949_), .B(33'h000000000), .S(RST), .Y(_01993_) );
  \$mux  #( .WIDTH(33) ) _48622_ ( .A(_source_stream_conv2d_16_source_23_pat_size_buf_0), .B(_source_stream_conv2d_16_source_23_pat_size_0), .S(_06716_), .Y(_25950_) );
  \$mux  #( .WIDTH(33) ) _48623_ ( .A(_25950_), .B(33'h000000000), .S(RST), .Y(_01992_) );
  \$mux  #( .WIDTH(33) ) _48624_ ( .A(_source_stream_conv2d_16_source_23_pat_count_3), .B(_28703_), .S(_06716_), .Y(_25951_) );
  \$mux  #( .WIDTH(33) ) _48625_ ( .A(_25951_), .B(_28710_), .S(_06719_), .Y(_25952_) );
  \$mux  #( .WIDTH(33) ) _48626_ ( .A(_25952_), .B(_28711_), .S(_06720_), .Y(_25953_) );
  \$mux  #( .WIDTH(33) ) _48627_ ( .A(_25953_), .B(33'h000000000), .S(RST), .Y(_01983_) );
  \$mux  #( .WIDTH(33) ) _48628_ ( .A(_source_stream_conv2d_16_source_23_pat_count_2), .B(_28702_), .S(_06716_), .Y(_25954_) );
  \$mux  #( .WIDTH(33) ) _48629_ ( .A(_25954_), .B(_28708_), .S(_06718_), .Y(_25955_) );
  \$mux  #( .WIDTH(33) ) _48630_ ( .A(_25955_), .B(_28709_), .S(_06719_), .Y(_25956_) );
  \$mux  #( .WIDTH(33) ) _48631_ ( .A(_25956_), .B(33'h000000000), .S(RST), .Y(_01982_) );
  \$mux  #( .WIDTH(33) ) _48632_ ( .A(_source_stream_conv2d_16_source_23_pat_count_1), .B(_28701_), .S(_06716_), .Y(_25957_) );
  \$mux  #( .WIDTH(33) ) _48633_ ( .A(_25957_), .B(_28706_), .S(_06717_), .Y(_25958_) );
  \$mux  #( .WIDTH(33) ) _48634_ ( .A(_25958_), .B(_28707_), .S(_06718_), .Y(_25959_) );
  \$mux  #( .WIDTH(33) ) _48635_ ( .A(_25959_), .B(33'h000000000), .S(RST), .Y(_01981_) );
  \$mux  #( .WIDTH(33) ) _48636_ ( .A(_source_stream_conv2d_16_source_23_pat_count_0), .B(_28700_), .S(_06716_), .Y(_25960_) );
  \$mux  #( .WIDTH(33) ) _48637_ ( .A(_28704_), .B(_25960_), .S(_05977_), .Y(_25961_) );
  \$mux  #( .WIDTH(33) ) _48638_ ( .A(_25961_), .B(_28705_), .S(_06717_), .Y(_25962_) );
  \$mux  #( .WIDTH(33) ) _48639_ ( .A(_25962_), .B(33'h000000000), .S(RST), .Y(_01980_) );
  \$mux  #( .WIDTH(32) ) _48640_ ( .A(_source_stream_conv2d_16_source_23_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_25963_) );
  \$mux  #( .WIDTH(32) ) _48641_ ( .A(_25963_), .B(0), .S(RST), .Y(_01999_) );
  \$mux  #( .WIDTH(32) ) _48642_ ( .A(_source_stream_conv2d_16_source_23_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_25964_) );
  \$mux  #( .WIDTH(32) ) _48643_ ( .A(_25964_), .B(0), .S(RST), .Y(_01998_) );
  \$mux  #( .WIDTH(32) ) _48644_ ( .A(_source_stream_conv2d_16_source_23_pat_stride_1), .B(0), .S(_set_flag_710), .Y(_25965_) );
  \$mux  #( .WIDTH(32) ) _48645_ ( .A(_25965_), .B(0), .S(RST), .Y(_01997_) );
  \$mux  #( .WIDTH(32) ) _48646_ ( .A(_source_stream_conv2d_16_source_23_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_25966_) );
  \$mux  #( .WIDTH(32) ) _48647_ ( .A(_25966_), .B(0), .S(RST), .Y(_01996_) );
  \$mux  #( .WIDTH(33) ) _48648_ ( .A(_source_stream_conv2d_16_source_23_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_25967_) );
  \$mux  #( .WIDTH(33) ) _48649_ ( .A(_25967_), .B(33'h000000000), .S(RST), .Y(_01991_) );
  \$mux  #( .WIDTH(33) ) _48650_ ( .A(_source_stream_conv2d_16_source_23_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_25968_) );
  \$mux  #( .WIDTH(33) ) _48651_ ( .A(_25968_), .B(33'h000000000), .S(RST), .Y(_01990_) );
  \$mux  #( .WIDTH(33) ) _48652_ ( .A(_source_stream_conv2d_16_source_23_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_25969_) );
  \$mux  #( .WIDTH(33) ) _48653_ ( .A(_25969_), .B(33'h000000000), .S(RST), .Y(_01989_) );
  \$mux  #( .WIDTH(33) ) _48654_ ( .A(_source_stream_conv2d_16_source_23_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_25970_) );
  \$mux  #( .WIDTH(33) ) _48655_ ( .A(_25970_), .B(33'h000000000), .S(RST), .Y(_01988_) );
  \$mux  #( .WIDTH(32) ) _48656_ ( .A(_source_stream_conv2d_16_source_23_pat_cur_offset_3), .B(0), .S(_06716_), .Y(_25971_) );
  \$mux  #( .WIDTH(32) ) _48657_ ( .A(_25971_), .B(_24340_), .S(_06719_), .Y(_25972_) );
  \$mux  #( .WIDTH(32) ) _48658_ ( .A(_25972_), .B(0), .S(_06720_), .Y(_25973_) );
  \$mux  #( .WIDTH(32) ) _48659_ ( .A(_25973_), .B(0), .S(RST), .Y(_01987_) );
  \$mux  #( .WIDTH(32) ) _48660_ ( .A(_source_stream_conv2d_16_source_23_pat_cur_offset_2), .B(0), .S(_06716_), .Y(_25974_) );
  \$mux  #( .WIDTH(32) ) _48661_ ( .A(_25974_), .B(_24339_), .S(_06718_), .Y(_25975_) );
  \$mux  #( .WIDTH(32) ) _48662_ ( .A(_25975_), .B(0), .S(_06719_), .Y(_25976_) );
  \$mux  #( .WIDTH(32) ) _48663_ ( .A(_25976_), .B(0), .S(RST), .Y(_01986_) );
  \$mux  #( .WIDTH(32) ) _48664_ ( .A(_source_stream_conv2d_16_source_23_pat_cur_offset_1), .B(0), .S(_06716_), .Y(_25977_) );
  \$mux  #( .WIDTH(32) ) _48665_ ( .A(_25977_), .B(_24338_), .S(_06717_), .Y(_25978_) );
  \$mux  #( .WIDTH(32) ) _48666_ ( .A(_25978_), .B(0), .S(_06718_), .Y(_25979_) );
  \$mux  #( .WIDTH(32) ) _48667_ ( .A(_25979_), .B(0), .S(RST), .Y(_01985_) );
  \$mux  #( .WIDTH(32) ) _48668_ ( .A(_source_stream_conv2d_16_source_23_pat_cur_offset_0), .B(0), .S(_06716_), .Y(_25980_) );
  \$mux  #( .WIDTH(32) ) _48669_ ( .A(_24337_), .B(_25980_), .S(_05977_), .Y(_25981_) );
  \$mux  #( .WIDTH(32) ) _48670_ ( .A(_25981_), .B(0), .S(_06717_), .Y(_25982_) );
  \$mux  #( .WIDTH(32) ) _48671_ ( .A(_25982_), .B(0), .S(RST), .Y(_01984_) );
  \$mux  #( .WIDTH(8) ) _48672_ ( .A(__variable_wdata_271), .B(_stream_conv2d_16_source_22_source_ram_rdata), .S(_stream_conv2d_16_source_22_source_ram_rvalid), .Y(_25983_) );
  \$mux  #( .WIDTH(8) ) _48673_ ( .A(_25983_), .B(8'h00), .S(RST), .Y(_01414_) );
  \$mux  #( .WIDTH(32) ) _48674_ ( .A(_source_stream_conv2d_16_source_22_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_22_pat_stride_3), .S(_06711_), .Y(_25984_) );
  \$mux  #( .WIDTH(32) ) _48675_ ( .A(_25984_), .B(0), .S(RST), .Y(_01979_) );
  \$mux  #( .WIDTH(32) ) _48676_ ( .A(_source_stream_conv2d_16_source_22_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_22_pat_stride_2), .S(_06711_), .Y(_25985_) );
  \$mux  #( .WIDTH(32) ) _48677_ ( .A(_25985_), .B(0), .S(RST), .Y(_01978_) );
  \$mux  #( .WIDTH(32) ) _48678_ ( .A(_source_stream_conv2d_16_source_22_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_22_pat_stride_1), .S(_06711_), .Y(_25986_) );
  \$mux  #( .WIDTH(32) ) _48679_ ( .A(_25986_), .B(0), .S(RST), .Y(_01977_) );
  \$mux  #( .WIDTH(32) ) _48680_ ( .A(_source_stream_conv2d_16_source_22_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_22_pat_stride_0), .S(_06711_), .Y(_25987_) );
  \$mux  #( .WIDTH(32) ) _48681_ ( .A(_25987_), .B(0), .S(RST), .Y(_01976_) );
  \$mux  #( .WIDTH(33) ) _48682_ ( .A(_source_stream_conv2d_16_source_22_pat_size_buf_3), .B(_source_stream_conv2d_16_source_22_pat_size_3), .S(_06711_), .Y(_25988_) );
  \$mux  #( .WIDTH(33) ) _48683_ ( .A(_25988_), .B(33'h000000000), .S(RST), .Y(_01971_) );
  \$mux  #( .WIDTH(33) ) _48684_ ( .A(_source_stream_conv2d_16_source_22_pat_size_buf_2), .B(_source_stream_conv2d_16_source_22_pat_size_2), .S(_06711_), .Y(_25989_) );
  \$mux  #( .WIDTH(33) ) _48685_ ( .A(_25989_), .B(33'h000000000), .S(RST), .Y(_01970_) );
  \$mux  #( .WIDTH(33) ) _48686_ ( .A(_source_stream_conv2d_16_source_22_pat_size_buf_1), .B(_source_stream_conv2d_16_source_22_pat_size_1), .S(_06711_), .Y(_25990_) );
  \$mux  #( .WIDTH(33) ) _48687_ ( .A(_25990_), .B(33'h000000000), .S(RST), .Y(_01969_) );
  \$mux  #( .WIDTH(33) ) _48688_ ( .A(_source_stream_conv2d_16_source_22_pat_size_buf_0), .B(_source_stream_conv2d_16_source_22_pat_size_0), .S(_06711_), .Y(_25991_) );
  \$mux  #( .WIDTH(33) ) _48689_ ( .A(_25991_), .B(33'h000000000), .S(RST), .Y(_01968_) );
  \$mux  #( .WIDTH(33) ) _48690_ ( .A(_source_stream_conv2d_16_source_22_pat_count_3), .B(_28691_), .S(_06711_), .Y(_25992_) );
  \$mux  #( .WIDTH(33) ) _48691_ ( .A(_25992_), .B(_28698_), .S(_06714_), .Y(_25993_) );
  \$mux  #( .WIDTH(33) ) _48692_ ( .A(_25993_), .B(_28699_), .S(_06715_), .Y(_25994_) );
  \$mux  #( .WIDTH(33) ) _48693_ ( .A(_25994_), .B(33'h000000000), .S(RST), .Y(_01959_) );
  \$mux  #( .WIDTH(33) ) _48694_ ( .A(_source_stream_conv2d_16_source_22_pat_count_2), .B(_28690_), .S(_06711_), .Y(_25995_) );
  \$mux  #( .WIDTH(33) ) _48695_ ( .A(_25995_), .B(_28696_), .S(_06713_), .Y(_25996_) );
  \$mux  #( .WIDTH(33) ) _48696_ ( .A(_25996_), .B(_28697_), .S(_06714_), .Y(_25997_) );
  \$mux  #( .WIDTH(33) ) _48697_ ( .A(_25997_), .B(33'h000000000), .S(RST), .Y(_01958_) );
  \$mux  #( .WIDTH(33) ) _48698_ ( .A(_source_stream_conv2d_16_source_22_pat_count_1), .B(_28689_), .S(_06711_), .Y(_25998_) );
  \$mux  #( .WIDTH(33) ) _48699_ ( .A(_25998_), .B(_28694_), .S(_06712_), .Y(_25999_) );
  \$mux  #( .WIDTH(33) ) _48700_ ( .A(_25999_), .B(_28695_), .S(_06713_), .Y(_26000_) );
  \$mux  #( .WIDTH(33) ) _48701_ ( .A(_26000_), .B(33'h000000000), .S(RST), .Y(_01957_) );
  \$mux  #( .WIDTH(33) ) _48702_ ( .A(_source_stream_conv2d_16_source_22_pat_count_0), .B(_28688_), .S(_06711_), .Y(_26001_) );
  \$mux  #( .WIDTH(33) ) _48703_ ( .A(_28692_), .B(_26001_), .S(_05979_), .Y(_26002_) );
  \$mux  #( .WIDTH(33) ) _48704_ ( .A(_26002_), .B(_28693_), .S(_06712_), .Y(_26003_) );
  \$mux  #( .WIDTH(33) ) _48705_ ( .A(_26003_), .B(33'h000000000), .S(RST), .Y(_01956_) );
  \$mux  #( .WIDTH(32) ) _48706_ ( .A(_source_stream_conv2d_16_source_22_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_26004_) );
  \$mux  #( .WIDTH(32) ) _48707_ ( .A(_26004_), .B(0), .S(RST), .Y(_01975_) );
  \$mux  #( .WIDTH(32) ) _48708_ ( .A(_source_stream_conv2d_16_source_22_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_26005_) );
  \$mux  #( .WIDTH(32) ) _48709_ ( .A(_26005_), .B(0), .S(RST), .Y(_01974_) );
  \$mux  #( .WIDTH(32) ) _48710_ ( .A(_source_stream_conv2d_16_source_22_pat_stride_1), .B(0), .S(_set_flag_710), .Y(_26006_) );
  \$mux  #( .WIDTH(32) ) _48711_ ( .A(_26006_), .B(0), .S(RST), .Y(_01973_) );
  \$mux  #( .WIDTH(32) ) _48712_ ( .A(_source_stream_conv2d_16_source_22_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_26007_) );
  \$mux  #( .WIDTH(32) ) _48713_ ( .A(_26007_), .B(0), .S(RST), .Y(_01972_) );
  \$mux  #( .WIDTH(33) ) _48714_ ( .A(_source_stream_conv2d_16_source_22_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_26008_) );
  \$mux  #( .WIDTH(33) ) _48715_ ( .A(_26008_), .B(33'h000000000), .S(RST), .Y(_01967_) );
  \$mux  #( .WIDTH(33) ) _48716_ ( .A(_source_stream_conv2d_16_source_22_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_26009_) );
  \$mux  #( .WIDTH(33) ) _48717_ ( .A(_26009_), .B(33'h000000000), .S(RST), .Y(_01966_) );
  \$mux  #( .WIDTH(33) ) _48718_ ( .A(_source_stream_conv2d_16_source_22_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_26010_) );
  \$mux  #( .WIDTH(33) ) _48719_ ( .A(_26010_), .B(33'h000000000), .S(RST), .Y(_01965_) );
  \$mux  #( .WIDTH(33) ) _48720_ ( .A(_source_stream_conv2d_16_source_22_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_26011_) );
  \$mux  #( .WIDTH(33) ) _48721_ ( .A(_26011_), .B(33'h000000000), .S(RST), .Y(_01964_) );
  \$mux  #( .WIDTH(32) ) _48722_ ( .A(_source_stream_conv2d_16_source_22_pat_cur_offset_3), .B(0), .S(_06711_), .Y(_26012_) );
  \$mux  #( .WIDTH(32) ) _48723_ ( .A(_26012_), .B(_24335_), .S(_06714_), .Y(_26013_) );
  \$mux  #( .WIDTH(32) ) _48724_ ( .A(_26013_), .B(0), .S(_06715_), .Y(_26014_) );
  \$mux  #( .WIDTH(32) ) _48725_ ( .A(_26014_), .B(0), .S(RST), .Y(_01963_) );
  \$mux  #( .WIDTH(32) ) _48726_ ( .A(_source_stream_conv2d_16_source_22_pat_cur_offset_2), .B(0), .S(_06711_), .Y(_26015_) );
  \$mux  #( .WIDTH(32) ) _48727_ ( .A(_26015_), .B(_24334_), .S(_06713_), .Y(_26016_) );
  \$mux  #( .WIDTH(32) ) _48728_ ( .A(_26016_), .B(0), .S(_06714_), .Y(_26017_) );
  \$mux  #( .WIDTH(32) ) _48729_ ( .A(_26017_), .B(0), .S(RST), .Y(_01962_) );
  \$mux  #( .WIDTH(32) ) _48730_ ( .A(_source_stream_conv2d_16_source_22_pat_cur_offset_1), .B(0), .S(_06711_), .Y(_26018_) );
  \$mux  #( .WIDTH(32) ) _48731_ ( .A(_26018_), .B(_24333_), .S(_06712_), .Y(_26019_) );
  \$mux  #( .WIDTH(32) ) _48732_ ( .A(_26019_), .B(0), .S(_06713_), .Y(_26020_) );
  \$mux  #( .WIDTH(32) ) _48733_ ( .A(_26020_), .B(0), .S(RST), .Y(_01961_) );
  \$mux  #( .WIDTH(32) ) _48734_ ( .A(_source_stream_conv2d_16_source_22_pat_cur_offset_0), .B(0), .S(_06711_), .Y(_26021_) );
  \$mux  #( .WIDTH(32) ) _48735_ ( .A(_24332_), .B(_26021_), .S(_05979_), .Y(_26022_) );
  \$mux  #( .WIDTH(32) ) _48736_ ( .A(_26022_), .B(0), .S(_06712_), .Y(_26023_) );
  \$mux  #( .WIDTH(32) ) _48737_ ( .A(_26023_), .B(0), .S(RST), .Y(_01960_) );
  \$mux  #( .WIDTH(8) ) _48738_ ( .A(__variable_wdata_270), .B(_stream_conv2d_16_source_21_source_ram_rdata), .S(_stream_conv2d_16_source_21_source_ram_rvalid), .Y(_26024_) );
  \$mux  #( .WIDTH(8) ) _48739_ ( .A(_26024_), .B(8'h00), .S(RST), .Y(_01413_) );
  \$mux  #( .WIDTH(32) ) _48740_ ( .A(_source_stream_conv2d_16_source_21_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_21_pat_stride_3), .S(_06706_), .Y(_26025_) );
  \$mux  #( .WIDTH(32) ) _48741_ ( .A(_26025_), .B(0), .S(RST), .Y(_01955_) );
  \$mux  #( .WIDTH(32) ) _48742_ ( .A(_source_stream_conv2d_16_source_21_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_21_pat_stride_2), .S(_06706_), .Y(_26026_) );
  \$mux  #( .WIDTH(32) ) _48743_ ( .A(_26026_), .B(0), .S(RST), .Y(_01954_) );
  \$mux  #( .WIDTH(32) ) _48744_ ( .A(_source_stream_conv2d_16_source_21_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_21_pat_stride_1), .S(_06706_), .Y(_26027_) );
  \$mux  #( .WIDTH(32) ) _48745_ ( .A(_26027_), .B(0), .S(RST), .Y(_01953_) );
  \$mux  #( .WIDTH(32) ) _48746_ ( .A(_source_stream_conv2d_16_source_21_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_21_pat_stride_0), .S(_06706_), .Y(_26028_) );
  \$mux  #( .WIDTH(32) ) _48747_ ( .A(_26028_), .B(0), .S(RST), .Y(_01952_) );
  \$mux  #( .WIDTH(33) ) _48748_ ( .A(_source_stream_conv2d_16_source_21_pat_size_buf_3), .B(_source_stream_conv2d_16_source_21_pat_size_3), .S(_06706_), .Y(_26029_) );
  \$mux  #( .WIDTH(33) ) _48749_ ( .A(_26029_), .B(33'h000000000), .S(RST), .Y(_01947_) );
  \$mux  #( .WIDTH(33) ) _48750_ ( .A(_source_stream_conv2d_16_source_21_pat_size_buf_2), .B(_source_stream_conv2d_16_source_21_pat_size_2), .S(_06706_), .Y(_26030_) );
  \$mux  #( .WIDTH(33) ) _48751_ ( .A(_26030_), .B(33'h000000000), .S(RST), .Y(_01946_) );
  \$mux  #( .WIDTH(33) ) _48752_ ( .A(_source_stream_conv2d_16_source_21_pat_size_buf_1), .B(_source_stream_conv2d_16_source_21_pat_size_1), .S(_06706_), .Y(_26031_) );
  \$mux  #( .WIDTH(33) ) _48753_ ( .A(_26031_), .B(33'h000000000), .S(RST), .Y(_01945_) );
  \$mux  #( .WIDTH(33) ) _48754_ ( .A(_source_stream_conv2d_16_source_21_pat_size_buf_0), .B(_source_stream_conv2d_16_source_21_pat_size_0), .S(_06706_), .Y(_26032_) );
  \$mux  #( .WIDTH(33) ) _48755_ ( .A(_26032_), .B(33'h000000000), .S(RST), .Y(_01944_) );
  \$mux  #( .WIDTH(33) ) _48756_ ( .A(_source_stream_conv2d_16_source_21_pat_count_3), .B(_28679_), .S(_06706_), .Y(_26033_) );
  \$mux  #( .WIDTH(33) ) _48757_ ( .A(_26033_), .B(_28686_), .S(_06709_), .Y(_26034_) );
  \$mux  #( .WIDTH(33) ) _48758_ ( .A(_26034_), .B(_28687_), .S(_06710_), .Y(_26035_) );
  \$mux  #( .WIDTH(33) ) _48759_ ( .A(_26035_), .B(33'h000000000), .S(RST), .Y(_01935_) );
  \$mux  #( .WIDTH(33) ) _48760_ ( .A(_source_stream_conv2d_16_source_21_pat_count_2), .B(_28678_), .S(_06706_), .Y(_26036_) );
  \$mux  #( .WIDTH(33) ) _48761_ ( .A(_26036_), .B(_28684_), .S(_06708_), .Y(_26037_) );
  \$mux  #( .WIDTH(33) ) _48762_ ( .A(_26037_), .B(_28685_), .S(_06709_), .Y(_26038_) );
  \$mux  #( .WIDTH(33) ) _48763_ ( .A(_26038_), .B(33'h000000000), .S(RST), .Y(_01934_) );
  \$mux  #( .WIDTH(33) ) _48764_ ( .A(_source_stream_conv2d_16_source_21_pat_count_1), .B(_28677_), .S(_06706_), .Y(_26039_) );
  \$mux  #( .WIDTH(33) ) _48765_ ( .A(_26039_), .B(_28682_), .S(_06707_), .Y(_26040_) );
  \$mux  #( .WIDTH(33) ) _48766_ ( .A(_26040_), .B(_28683_), .S(_06708_), .Y(_26041_) );
  \$mux  #( .WIDTH(33) ) _48767_ ( .A(_26041_), .B(33'h000000000), .S(RST), .Y(_01933_) );
  \$mux  #( .WIDTH(33) ) _48768_ ( .A(_source_stream_conv2d_16_source_21_pat_count_0), .B(_28676_), .S(_06706_), .Y(_26042_) );
  \$mux  #( .WIDTH(33) ) _48769_ ( .A(_28680_), .B(_26042_), .S(_05981_), .Y(_26043_) );
  \$mux  #( .WIDTH(33) ) _48770_ ( .A(_26043_), .B(_28681_), .S(_06707_), .Y(_26044_) );
  \$mux  #( .WIDTH(33) ) _48771_ ( .A(_26044_), .B(33'h000000000), .S(RST), .Y(_01932_) );
  \$mux  #( .WIDTH(32) ) _48772_ ( .A(_source_stream_conv2d_16_source_21_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_26045_) );
  \$mux  #( .WIDTH(32) ) _48773_ ( .A(_26045_), .B(0), .S(RST), .Y(_01951_) );
  \$mux  #( .WIDTH(32) ) _48774_ ( .A(_source_stream_conv2d_16_source_21_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_26046_) );
  \$mux  #( .WIDTH(32) ) _48775_ ( .A(_26046_), .B(0), .S(RST), .Y(_01950_) );
  \$mux  #( .WIDTH(32) ) _48776_ ( .A(_source_stream_conv2d_16_source_21_pat_stride_1), .B(0), .S(_set_flag_710), .Y(_26047_) );
  \$mux  #( .WIDTH(32) ) _48777_ ( .A(_26047_), .B(0), .S(RST), .Y(_01949_) );
  \$mux  #( .WIDTH(32) ) _48778_ ( .A(_source_stream_conv2d_16_source_21_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_26048_) );
  \$mux  #( .WIDTH(32) ) _48779_ ( .A(_26048_), .B(0), .S(RST), .Y(_01948_) );
  \$mux  #( .WIDTH(33) ) _48780_ ( .A(_source_stream_conv2d_16_source_21_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_26049_) );
  \$mux  #( .WIDTH(33) ) _48781_ ( .A(_26049_), .B(33'h000000000), .S(RST), .Y(_01943_) );
  \$mux  #( .WIDTH(33) ) _48782_ ( .A(_source_stream_conv2d_16_source_21_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_26050_) );
  \$mux  #( .WIDTH(33) ) _48783_ ( .A(_26050_), .B(33'h000000000), .S(RST), .Y(_01942_) );
  \$mux  #( .WIDTH(33) ) _48784_ ( .A(_source_stream_conv2d_16_source_21_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_26051_) );
  \$mux  #( .WIDTH(33) ) _48785_ ( .A(_26051_), .B(33'h000000000), .S(RST), .Y(_01941_) );
  \$mux  #( .WIDTH(33) ) _48786_ ( .A(_source_stream_conv2d_16_source_21_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_26052_) );
  \$mux  #( .WIDTH(33) ) _48787_ ( .A(_26052_), .B(33'h000000000), .S(RST), .Y(_01940_) );
  \$mux  #( .WIDTH(32) ) _48788_ ( .A(_source_stream_conv2d_16_source_21_pat_cur_offset_3), .B(0), .S(_06706_), .Y(_26053_) );
  \$mux  #( .WIDTH(32) ) _48789_ ( .A(_26053_), .B(_24330_), .S(_06709_), .Y(_26054_) );
  \$mux  #( .WIDTH(32) ) _48790_ ( .A(_26054_), .B(0), .S(_06710_), .Y(_26055_) );
  \$mux  #( .WIDTH(32) ) _48791_ ( .A(_26055_), .B(0), .S(RST), .Y(_01939_) );
  \$mux  #( .WIDTH(32) ) _48792_ ( .A(_source_stream_conv2d_16_source_21_pat_cur_offset_2), .B(0), .S(_06706_), .Y(_26056_) );
  \$mux  #( .WIDTH(32) ) _48793_ ( .A(_26056_), .B(_24329_), .S(_06708_), .Y(_26057_) );
  \$mux  #( .WIDTH(32) ) _48794_ ( .A(_26057_), .B(0), .S(_06709_), .Y(_26058_) );
  \$mux  #( .WIDTH(32) ) _48795_ ( .A(_26058_), .B(0), .S(RST), .Y(_01938_) );
  \$mux  #( .WIDTH(32) ) _48796_ ( .A(_source_stream_conv2d_16_source_21_pat_cur_offset_1), .B(0), .S(_06706_), .Y(_26059_) );
  \$mux  #( .WIDTH(32) ) _48797_ ( .A(_26059_), .B(_24328_), .S(_06707_), .Y(_26060_) );
  \$mux  #( .WIDTH(32) ) _48798_ ( .A(_26060_), .B(0), .S(_06708_), .Y(_26061_) );
  \$mux  #( .WIDTH(32) ) _48799_ ( .A(_26061_), .B(0), .S(RST), .Y(_01937_) );
  \$mux  #( .WIDTH(32) ) _48800_ ( .A(_source_stream_conv2d_16_source_21_pat_cur_offset_0), .B(0), .S(_06706_), .Y(_26062_) );
  \$mux  #( .WIDTH(32) ) _48801_ ( .A(_24327_), .B(_26062_), .S(_05981_), .Y(_26063_) );
  \$mux  #( .WIDTH(32) ) _48802_ ( .A(_26063_), .B(0), .S(_06707_), .Y(_26064_) );
  \$mux  #( .WIDTH(32) ) _48803_ ( .A(_26064_), .B(0), .S(RST), .Y(_01936_) );
  \$mux  #( .WIDTH(8) ) _48804_ ( .A(__variable_wdata_269), .B(_stream_conv2d_16_source_20_source_ram_rdata), .S(_stream_conv2d_16_source_20_source_ram_rvalid), .Y(_26065_) );
  \$mux  #( .WIDTH(8) ) _48805_ ( .A(_26065_), .B(8'h00), .S(RST), .Y(_01411_) );
  \$mux  #( .WIDTH(32) ) _48806_ ( .A(_source_stream_conv2d_16_source_20_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_20_pat_stride_3), .S(_06701_), .Y(_26066_) );
  \$mux  #( .WIDTH(32) ) _48807_ ( .A(_26066_), .B(0), .S(RST), .Y(_01931_) );
  \$mux  #( .WIDTH(32) ) _48808_ ( .A(_source_stream_conv2d_16_source_20_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_20_pat_stride_2), .S(_06701_), .Y(_26067_) );
  \$mux  #( .WIDTH(32) ) _48809_ ( .A(_26067_), .B(0), .S(RST), .Y(_01930_) );
  \$mux  #( .WIDTH(32) ) _48810_ ( .A(_source_stream_conv2d_16_source_20_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_20_pat_stride_1), .S(_06701_), .Y(_26068_) );
  \$mux  #( .WIDTH(32) ) _48811_ ( .A(_26068_), .B(0), .S(RST), .Y(_01929_) );
  \$mux  #( .WIDTH(32) ) _48812_ ( .A(_source_stream_conv2d_16_source_20_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_20_pat_stride_0), .S(_06701_), .Y(_26069_) );
  \$mux  #( .WIDTH(32) ) _48813_ ( .A(_26069_), .B(0), .S(RST), .Y(_01928_) );
  \$mux  #( .WIDTH(33) ) _48814_ ( .A(_source_stream_conv2d_16_source_20_pat_size_buf_3), .B(_source_stream_conv2d_16_source_20_pat_size_3), .S(_06701_), .Y(_26070_) );
  \$mux  #( .WIDTH(33) ) _48815_ ( .A(_26070_), .B(33'h000000000), .S(RST), .Y(_01923_) );
  \$mux  #( .WIDTH(33) ) _48816_ ( .A(_source_stream_conv2d_16_source_20_pat_size_buf_2), .B(_source_stream_conv2d_16_source_20_pat_size_2), .S(_06701_), .Y(_26071_) );
  \$mux  #( .WIDTH(33) ) _48817_ ( .A(_26071_), .B(33'h000000000), .S(RST), .Y(_01922_) );
  \$mux  #( .WIDTH(33) ) _48818_ ( .A(_source_stream_conv2d_16_source_20_pat_size_buf_1), .B(_source_stream_conv2d_16_source_20_pat_size_1), .S(_06701_), .Y(_26072_) );
  \$mux  #( .WIDTH(33) ) _48819_ ( .A(_26072_), .B(33'h000000000), .S(RST), .Y(_01921_) );
  \$mux  #( .WIDTH(33) ) _48820_ ( .A(_source_stream_conv2d_16_source_20_pat_size_buf_0), .B(_source_stream_conv2d_16_source_20_pat_size_0), .S(_06701_), .Y(_26073_) );
  \$mux  #( .WIDTH(33) ) _48821_ ( .A(_26073_), .B(33'h000000000), .S(RST), .Y(_01920_) );
  \$mux  #( .WIDTH(33) ) _48822_ ( .A(_source_stream_conv2d_16_source_20_pat_count_3), .B(_28667_), .S(_06701_), .Y(_26074_) );
  \$mux  #( .WIDTH(33) ) _48823_ ( .A(_26074_), .B(_28674_), .S(_06704_), .Y(_26075_) );
  \$mux  #( .WIDTH(33) ) _48824_ ( .A(_26075_), .B(_28675_), .S(_06705_), .Y(_26076_) );
  \$mux  #( .WIDTH(33) ) _48825_ ( .A(_26076_), .B(33'h000000000), .S(RST), .Y(_01911_) );
  \$mux  #( .WIDTH(33) ) _48826_ ( .A(_source_stream_conv2d_16_source_20_pat_count_2), .B(_28666_), .S(_06701_), .Y(_26077_) );
  \$mux  #( .WIDTH(33) ) _48827_ ( .A(_26077_), .B(_28672_), .S(_06703_), .Y(_26078_) );
  \$mux  #( .WIDTH(33) ) _48828_ ( .A(_26078_), .B(_28673_), .S(_06704_), .Y(_26079_) );
  \$mux  #( .WIDTH(33) ) _48829_ ( .A(_26079_), .B(33'h000000000), .S(RST), .Y(_01910_) );
  \$mux  #( .WIDTH(33) ) _48830_ ( .A(_source_stream_conv2d_16_source_20_pat_count_1), .B(_28665_), .S(_06701_), .Y(_26080_) );
  \$mux  #( .WIDTH(33) ) _48831_ ( .A(_26080_), .B(_28670_), .S(_06702_), .Y(_26081_) );
  \$mux  #( .WIDTH(33) ) _48832_ ( .A(_26081_), .B(_28671_), .S(_06703_), .Y(_26082_) );
  \$mux  #( .WIDTH(33) ) _48833_ ( .A(_26082_), .B(33'h000000000), .S(RST), .Y(_01909_) );
  \$mux  #( .WIDTH(33) ) _48834_ ( .A(_source_stream_conv2d_16_source_20_pat_count_0), .B(_28664_), .S(_06701_), .Y(_26083_) );
  \$mux  #( .WIDTH(33) ) _48835_ ( .A(_28668_), .B(_26083_), .S(_05982_), .Y(_26084_) );
  \$mux  #( .WIDTH(33) ) _48836_ ( .A(_26084_), .B(_28669_), .S(_06702_), .Y(_26085_) );
  \$mux  #( .WIDTH(33) ) _48837_ ( .A(_26085_), .B(33'h000000000), .S(RST), .Y(_01908_) );
  \$mux  #( .WIDTH(32) ) _48838_ ( .A(_source_stream_conv2d_16_source_20_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_26086_) );
  \$mux  #( .WIDTH(32) ) _48839_ ( .A(_26086_), .B(0), .S(RST), .Y(_01927_) );
  \$mux  #( .WIDTH(32) ) _48840_ ( .A(_source_stream_conv2d_16_source_20_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_26087_) );
  \$mux  #( .WIDTH(32) ) _48841_ ( .A(_26087_), .B(0), .S(RST), .Y(_01926_) );
  \$mux  #( .WIDTH(32) ) _48842_ ( .A(_source_stream_conv2d_16_source_20_pat_stride_1), .B(0), .S(_set_flag_710), .Y(_26088_) );
  \$mux  #( .WIDTH(32) ) _48843_ ( .A(_26088_), .B(0), .S(RST), .Y(_01925_) );
  \$mux  #( .WIDTH(32) ) _48844_ ( .A(_source_stream_conv2d_16_source_20_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_26089_) );
  \$mux  #( .WIDTH(32) ) _48845_ ( .A(_26089_), .B(0), .S(RST), .Y(_01924_) );
  \$mux  #( .WIDTH(33) ) _48846_ ( .A(_source_stream_conv2d_16_source_20_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_26090_) );
  \$mux  #( .WIDTH(33) ) _48847_ ( .A(_26090_), .B(33'h000000000), .S(RST), .Y(_01919_) );
  \$mux  #( .WIDTH(33) ) _48848_ ( .A(_source_stream_conv2d_16_source_20_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_26091_) );
  \$mux  #( .WIDTH(33) ) _48849_ ( .A(_26091_), .B(33'h000000000), .S(RST), .Y(_01918_) );
  \$mux  #( .WIDTH(33) ) _48850_ ( .A(_source_stream_conv2d_16_source_20_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_26092_) );
  \$mux  #( .WIDTH(33) ) _48851_ ( .A(_26092_), .B(33'h000000000), .S(RST), .Y(_01917_) );
  \$mux  #( .WIDTH(33) ) _48852_ ( .A(_source_stream_conv2d_16_source_20_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_26093_) );
  \$mux  #( .WIDTH(33) ) _48853_ ( .A(_26093_), .B(33'h000000000), .S(RST), .Y(_01916_) );
  \$mux  #( .WIDTH(32) ) _48854_ ( .A(_source_stream_conv2d_16_source_20_pat_cur_offset_3), .B(0), .S(_06701_), .Y(_26094_) );
  \$mux  #( .WIDTH(32) ) _48855_ ( .A(_26094_), .B(_24325_), .S(_06704_), .Y(_26095_) );
  \$mux  #( .WIDTH(32) ) _48856_ ( .A(_26095_), .B(0), .S(_06705_), .Y(_26096_) );
  \$mux  #( .WIDTH(32) ) _48857_ ( .A(_26096_), .B(0), .S(RST), .Y(_01915_) );
  \$mux  #( .WIDTH(32) ) _48858_ ( .A(_source_stream_conv2d_16_source_20_pat_cur_offset_2), .B(0), .S(_06701_), .Y(_26097_) );
  \$mux  #( .WIDTH(32) ) _48859_ ( .A(_26097_), .B(_24324_), .S(_06703_), .Y(_26098_) );
  \$mux  #( .WIDTH(32) ) _48860_ ( .A(_26098_), .B(0), .S(_06704_), .Y(_26099_) );
  \$mux  #( .WIDTH(32) ) _48861_ ( .A(_26099_), .B(0), .S(RST), .Y(_01914_) );
  \$mux  #( .WIDTH(32) ) _48862_ ( .A(_source_stream_conv2d_16_source_20_pat_cur_offset_1), .B(0), .S(_06701_), .Y(_26100_) );
  \$mux  #( .WIDTH(32) ) _48863_ ( .A(_26100_), .B(_24323_), .S(_06702_), .Y(_26101_) );
  \$mux  #( .WIDTH(32) ) _48864_ ( .A(_26101_), .B(0), .S(_06703_), .Y(_26102_) );
  \$mux  #( .WIDTH(32) ) _48865_ ( .A(_26102_), .B(0), .S(RST), .Y(_01913_) );
  \$mux  #( .WIDTH(32) ) _48866_ ( .A(_source_stream_conv2d_16_source_20_pat_cur_offset_0), .B(0), .S(_06701_), .Y(_26103_) );
  \$mux  #( .WIDTH(32) ) _48867_ ( .A(_24322_), .B(_26103_), .S(_05982_), .Y(_26104_) );
  \$mux  #( .WIDTH(32) ) _48868_ ( .A(_26104_), .B(0), .S(_06702_), .Y(_26105_) );
  \$mux  #( .WIDTH(32) ) _48869_ ( .A(_26105_), .B(0), .S(RST), .Y(_01912_) );
  \$mux  #( .WIDTH(8) ) _48870_ ( .A(__variable_wdata_268), .B(_stream_conv2d_16_source_19_source_ram_rdata), .S(_stream_conv2d_16_source_19_source_ram_rvalid), .Y(_26106_) );
  \$mux  #( .WIDTH(8) ) _48871_ ( .A(_26106_), .B(8'h00), .S(RST), .Y(_01410_) );
  \$mux  #( .WIDTH(32) ) _48872_ ( .A(_source_stream_conv2d_16_source_19_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_19_pat_stride_3), .S(_06696_), .Y(_26107_) );
  \$mux  #( .WIDTH(32) ) _48873_ ( .A(_26107_), .B(0), .S(RST), .Y(_01907_) );
  \$mux  #( .WIDTH(32) ) _48874_ ( .A(_source_stream_conv2d_16_source_19_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_19_pat_stride_2), .S(_06696_), .Y(_26108_) );
  \$mux  #( .WIDTH(32) ) _48875_ ( .A(_26108_), .B(0), .S(RST), .Y(_01906_) );
  \$mux  #( .WIDTH(32) ) _48876_ ( .A(_source_stream_conv2d_16_source_19_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_19_pat_stride_1), .S(_06696_), .Y(_26109_) );
  \$mux  #( .WIDTH(32) ) _48877_ ( .A(_26109_), .B(0), .S(RST), .Y(_01905_) );
  \$mux  #( .WIDTH(32) ) _48878_ ( .A(_source_stream_conv2d_16_source_19_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_19_pat_stride_0), .S(_06696_), .Y(_26110_) );
  \$mux  #( .WIDTH(32) ) _48879_ ( .A(_26110_), .B(0), .S(RST), .Y(_01904_) );
  \$mux  #( .WIDTH(33) ) _48880_ ( .A(_source_stream_conv2d_16_source_19_pat_size_buf_3), .B(_source_stream_conv2d_16_source_19_pat_size_3), .S(_06696_), .Y(_26111_) );
  \$mux  #( .WIDTH(33) ) _48881_ ( .A(_26111_), .B(33'h000000000), .S(RST), .Y(_01899_) );
  \$mux  #( .WIDTH(33) ) _48882_ ( .A(_source_stream_conv2d_16_source_19_pat_size_buf_2), .B(_source_stream_conv2d_16_source_19_pat_size_2), .S(_06696_), .Y(_26112_) );
  \$mux  #( .WIDTH(33) ) _48883_ ( .A(_26112_), .B(33'h000000000), .S(RST), .Y(_01898_) );
  \$mux  #( .WIDTH(33) ) _48884_ ( .A(_source_stream_conv2d_16_source_19_pat_size_buf_1), .B(_source_stream_conv2d_16_source_19_pat_size_1), .S(_06696_), .Y(_26113_) );
  \$mux  #( .WIDTH(33) ) _48885_ ( .A(_26113_), .B(33'h000000000), .S(RST), .Y(_01897_) );
  \$mux  #( .WIDTH(33) ) _48886_ ( .A(_source_stream_conv2d_16_source_19_pat_size_buf_0), .B(_source_stream_conv2d_16_source_19_pat_size_0), .S(_06696_), .Y(_26114_) );
  \$mux  #( .WIDTH(33) ) _48887_ ( .A(_26114_), .B(33'h000000000), .S(RST), .Y(_01896_) );
  \$mux  #( .WIDTH(33) ) _48888_ ( .A(_source_stream_conv2d_16_source_19_pat_count_3), .B(_28655_), .S(_06696_), .Y(_26115_) );
  \$mux  #( .WIDTH(33) ) _48889_ ( .A(_26115_), .B(_28662_), .S(_06699_), .Y(_26116_) );
  \$mux  #( .WIDTH(33) ) _48890_ ( .A(_26116_), .B(_28663_), .S(_06700_), .Y(_26117_) );
  \$mux  #( .WIDTH(33) ) _48891_ ( .A(_26117_), .B(33'h000000000), .S(RST), .Y(_01887_) );
  \$mux  #( .WIDTH(33) ) _48892_ ( .A(_source_stream_conv2d_16_source_19_pat_count_2), .B(_28654_), .S(_06696_), .Y(_26118_) );
  \$mux  #( .WIDTH(33) ) _48893_ ( .A(_26118_), .B(_28660_), .S(_06698_), .Y(_26119_) );
  \$mux  #( .WIDTH(33) ) _48894_ ( .A(_26119_), .B(_28661_), .S(_06699_), .Y(_26120_) );
  \$mux  #( .WIDTH(33) ) _48895_ ( .A(_26120_), .B(33'h000000000), .S(RST), .Y(_01886_) );
  \$mux  #( .WIDTH(33) ) _48896_ ( .A(_source_stream_conv2d_16_source_19_pat_count_1), .B(_28653_), .S(_06696_), .Y(_26121_) );
  \$mux  #( .WIDTH(33) ) _48897_ ( .A(_26121_), .B(_28658_), .S(_06697_), .Y(_26122_) );
  \$mux  #( .WIDTH(33) ) _48898_ ( .A(_26122_), .B(_28659_), .S(_06698_), .Y(_26123_) );
  \$mux  #( .WIDTH(33) ) _48899_ ( .A(_26123_), .B(33'h000000000), .S(RST), .Y(_01885_) );
  \$mux  #( .WIDTH(33) ) _48900_ ( .A(_source_stream_conv2d_16_source_19_pat_count_0), .B(_28652_), .S(_06696_), .Y(_26124_) );
  \$mux  #( .WIDTH(33) ) _48901_ ( .A(_28656_), .B(_26124_), .S(_05983_), .Y(_26125_) );
  \$mux  #( .WIDTH(33) ) _48902_ ( .A(_26125_), .B(_28657_), .S(_06697_), .Y(_26126_) );
  \$mux  #( .WIDTH(33) ) _48903_ ( .A(_26126_), .B(33'h000000000), .S(RST), .Y(_01884_) );
  \$mux  #( .WIDTH(32) ) _48904_ ( .A(_source_stream_conv2d_16_source_19_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_26127_) );
  \$mux  #( .WIDTH(32) ) _48905_ ( .A(_26127_), .B(0), .S(RST), .Y(_01903_) );
  \$mux  #( .WIDTH(32) ) _48906_ ( .A(_source_stream_conv2d_16_source_19_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_26128_) );
  \$mux  #( .WIDTH(32) ) _48907_ ( .A(_26128_), .B(0), .S(RST), .Y(_01902_) );
  \$mux  #( .WIDTH(32) ) _48908_ ( .A(_source_stream_conv2d_16_source_19_pat_stride_1), .B(0), .S(_set_flag_710), .Y(_26129_) );
  \$mux  #( .WIDTH(32) ) _48909_ ( .A(_26129_), .B(0), .S(RST), .Y(_01901_) );
  \$mux  #( .WIDTH(32) ) _48910_ ( .A(_source_stream_conv2d_16_source_19_pat_stride_0), .B(1), .S(_set_flag_710), .Y(_26130_) );
  \$mux  #( .WIDTH(32) ) _48911_ ( .A(_26130_), .B(0), .S(RST), .Y(_01900_) );
  \$mux  #( .WIDTH(33) ) _48912_ ( .A(_source_stream_conv2d_16_source_19_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_26131_) );
  \$mux  #( .WIDTH(33) ) _48913_ ( .A(_26131_), .B(33'h000000000), .S(RST), .Y(_01895_) );
  \$mux  #( .WIDTH(33) ) _48914_ ( .A(_source_stream_conv2d_16_source_19_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_26132_) );
  \$mux  #( .WIDTH(33) ) _48915_ ( .A(_26132_), .B(33'h000000000), .S(RST), .Y(_01894_) );
  \$mux  #( .WIDTH(33) ) _48916_ ( .A(_source_stream_conv2d_16_source_19_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_26133_) );
  \$mux  #( .WIDTH(33) ) _48917_ ( .A(_26133_), .B(33'h000000000), .S(RST), .Y(_01893_) );
  \$mux  #( .WIDTH(33) ) _48918_ ( .A(_source_stream_conv2d_16_source_19_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_26134_) );
  \$mux  #( .WIDTH(33) ) _48919_ ( .A(_26134_), .B(33'h000000000), .S(RST), .Y(_01892_) );
  \$mux  #( .WIDTH(32) ) _48920_ ( .A(_source_stream_conv2d_16_source_19_pat_cur_offset_3), .B(0), .S(_06696_), .Y(_26135_) );
  \$mux  #( .WIDTH(32) ) _48921_ ( .A(_26135_), .B(_24320_), .S(_06699_), .Y(_26136_) );
  \$mux  #( .WIDTH(32) ) _48922_ ( .A(_26136_), .B(0), .S(_06700_), .Y(_26137_) );
  \$mux  #( .WIDTH(32) ) _48923_ ( .A(_26137_), .B(0), .S(RST), .Y(_01891_) );
  \$mux  #( .WIDTH(32) ) _48924_ ( .A(_source_stream_conv2d_16_source_19_pat_cur_offset_2), .B(0), .S(_06696_), .Y(_26138_) );
  \$mux  #( .WIDTH(32) ) _48925_ ( .A(_26138_), .B(_24319_), .S(_06698_), .Y(_26139_) );
  \$mux  #( .WIDTH(32) ) _48926_ ( .A(_26139_), .B(0), .S(_06699_), .Y(_26140_) );
  \$mux  #( .WIDTH(32) ) _48927_ ( .A(_26140_), .B(0), .S(RST), .Y(_01890_) );
  \$mux  #( .WIDTH(32) ) _48928_ ( .A(_source_stream_conv2d_16_source_19_pat_cur_offset_1), .B(0), .S(_06696_), .Y(_26141_) );
  \$mux  #( .WIDTH(32) ) _48929_ ( .A(_26141_), .B(_24318_), .S(_06697_), .Y(_26142_) );
  \$mux  #( .WIDTH(32) ) _48930_ ( .A(_26142_), .B(0), .S(_06698_), .Y(_26143_) );
  \$mux  #( .WIDTH(32) ) _48931_ ( .A(_26143_), .B(0), .S(RST), .Y(_01889_) );
  \$mux  #( .WIDTH(32) ) _48932_ ( .A(_source_stream_conv2d_16_source_19_pat_cur_offset_0), .B(0), .S(_06696_), .Y(_26144_) );
  \$mux  #( .WIDTH(32) ) _48933_ ( .A(_24317_), .B(_26144_), .S(_05983_), .Y(_26145_) );
  \$mux  #( .WIDTH(32) ) _48934_ ( .A(_26145_), .B(0), .S(_06697_), .Y(_26146_) );
  \$mux  #( .WIDTH(32) ) _48935_ ( .A(_26146_), .B(0), .S(RST), .Y(_01888_) );
  \$mux  #( .WIDTH(4) ) _48936_ ( .A(__variable_wdata_266), .B(_stream_conv2d_16_constant_17_next_constant_data), .S(_stream_conv2d_16_start), .Y(_26147_) );
  \$mux  #( .WIDTH(4) ) _48937_ ( .A(_26147_), .B(4'h0), .S(RST), .Y(_01409_) );
  \$mux  #( .WIDTH(1) ) _48938_ ( .A(__variable_wdata_265), .B(_stream_conv2d_16_constant_16_next_constant_data), .S(_stream_conv2d_16_start), .Y(_26148_) );
  \$mux  #( .WIDTH(1) ) _48939_ ( .A(_26148_), .B(1'h0), .S(RST), .Y(_01408_) );
  \$mux  #( .WIDTH(1) ) _48940_ ( .A(__variable_wdata_264), .B(_stream_conv2d_16_constant_15_next_constant_data), .S(_stream_conv2d_16_start), .Y(_26149_) );
  \$mux  #( .WIDTH(1) ) _48941_ ( .A(_26149_), .B(1'h0), .S(RST), .Y(_01407_) );
  \$mux  #( .WIDTH(8) ) _48942_ ( .A(__variable_wdata_258), .B(_stream_conv2d_16_source_14_source_empty_data), .S(_stream_conv2d_16_start), .Y(_26150_) );
  \$mux  #( .WIDTH(8) ) _48943_ ( .A(_26150_), .B(8'h00), .S(RST), .Y(_01405_) );
  \$mux  #( .WIDTH(8) ) _48944_ ( .A(__variable_wdata_251), .B(_stream_conv2d_16_source_12_source_empty_data), .S(_stream_conv2d_16_start), .Y(_26151_) );
  \$mux  #( .WIDTH(8) ) _48945_ ( .A(_26151_), .B(8'h00), .S(RST), .Y(_01404_) );
  \$mux  #( .WIDTH(8) ) _48946_ ( .A(__variable_wdata_244), .B(_stream_conv2d_16_source_10_source_empty_data), .S(_stream_conv2d_16_start), .Y(_26152_) );
  \$mux  #( .WIDTH(8) ) _48947_ ( .A(_26152_), .B(8'h00), .S(RST), .Y(_01402_) );
  \$mux  #( .WIDTH(8) ) _48948_ ( .A(__variable_wdata_237), .B(_stream_conv2d_16_source_8_source_ram_rdata), .S(_stream_conv2d_16_source_8_source_ram_rvalid), .Y(_26153_) );
  \$mux  #( .WIDTH(8) ) _48949_ ( .A(_26153_), .B(8'h00), .S(RST), .Y(_01401_) );
  \$mux  #( .WIDTH(32) ) _48950_ ( .A(_source_stream_conv2d_16_source_8_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_8_pat_stride_3), .S(_06691_), .Y(_26154_) );
  \$mux  #( .WIDTH(32) ) _48951_ ( .A(_26154_), .B(0), .S(RST), .Y(_02363_) );
  \$mux  #( .WIDTH(32) ) _48952_ ( .A(_source_stream_conv2d_16_source_8_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_8_pat_stride_2), .S(_06691_), .Y(_26155_) );
  \$mux  #( .WIDTH(32) ) _48953_ ( .A(_26155_), .B(0), .S(RST), .Y(_02362_) );
  \$mux  #( .WIDTH(32) ) _48954_ ( .A(_source_stream_conv2d_16_source_8_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_8_pat_stride_1), .S(_06691_), .Y(_26156_) );
  \$mux  #( .WIDTH(32) ) _48955_ ( .A(_26156_), .B(0), .S(RST), .Y(_02361_) );
  \$mux  #( .WIDTH(32) ) _48956_ ( .A(_source_stream_conv2d_16_source_8_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_8_pat_stride_0), .S(_06691_), .Y(_26157_) );
  \$mux  #( .WIDTH(32) ) _48957_ ( .A(_26157_), .B(0), .S(RST), .Y(_02360_) );
  \$mux  #( .WIDTH(33) ) _48958_ ( .A(_source_stream_conv2d_16_source_8_pat_size_buf_3), .B(_source_stream_conv2d_16_source_8_pat_size_3), .S(_06691_), .Y(_26158_) );
  \$mux  #( .WIDTH(33) ) _48959_ ( .A(_26158_), .B(33'h000000000), .S(RST), .Y(_02355_) );
  \$mux  #( .WIDTH(33) ) _48960_ ( .A(_source_stream_conv2d_16_source_8_pat_size_buf_2), .B(_source_stream_conv2d_16_source_8_pat_size_2), .S(_06691_), .Y(_26159_) );
  \$mux  #( .WIDTH(33) ) _48961_ ( .A(_26159_), .B(33'h000000000), .S(RST), .Y(_02354_) );
  \$mux  #( .WIDTH(33) ) _48962_ ( .A(_source_stream_conv2d_16_source_8_pat_size_buf_1), .B(_source_stream_conv2d_16_source_8_pat_size_1), .S(_06691_), .Y(_26160_) );
  \$mux  #( .WIDTH(33) ) _48963_ ( .A(_26160_), .B(33'h000000000), .S(RST), .Y(_02353_) );
  \$mux  #( .WIDTH(33) ) _48964_ ( .A(_source_stream_conv2d_16_source_8_pat_size_buf_0), .B(_source_stream_conv2d_16_source_8_pat_size_0), .S(_06691_), .Y(_26161_) );
  \$mux  #( .WIDTH(33) ) _48965_ ( .A(_26161_), .B(33'h000000000), .S(RST), .Y(_02352_) );
  \$mux  #( .WIDTH(33) ) _48966_ ( .A(_source_stream_conv2d_16_source_8_pat_count_3), .B(_28643_), .S(_06691_), .Y(_26162_) );
  \$mux  #( .WIDTH(33) ) _48967_ ( .A(_26162_), .B(_28650_), .S(_06694_), .Y(_26163_) );
  \$mux  #( .WIDTH(33) ) _48968_ ( .A(_26163_), .B(_28651_), .S(_06695_), .Y(_26164_) );
  \$mux  #( .WIDTH(33) ) _48969_ ( .A(_26164_), .B(33'h000000000), .S(RST), .Y(_02343_) );
  \$mux  #( .WIDTH(33) ) _48970_ ( .A(_source_stream_conv2d_16_source_8_pat_count_2), .B(_28642_), .S(_06691_), .Y(_26165_) );
  \$mux  #( .WIDTH(33) ) _48971_ ( .A(_26165_), .B(_28648_), .S(_06693_), .Y(_26166_) );
  \$mux  #( .WIDTH(33) ) _48972_ ( .A(_26166_), .B(_28649_), .S(_06694_), .Y(_26167_) );
  \$mux  #( .WIDTH(33) ) _48973_ ( .A(_26167_), .B(33'h000000000), .S(RST), .Y(_02342_) );
  \$mux  #( .WIDTH(33) ) _48974_ ( .A(_source_stream_conv2d_16_source_8_pat_count_1), .B(_28641_), .S(_06691_), .Y(_26168_) );
  \$mux  #( .WIDTH(33) ) _48975_ ( .A(_26168_), .B(_28646_), .S(_06692_), .Y(_26169_) );
  \$mux  #( .WIDTH(33) ) _48976_ ( .A(_26169_), .B(_28647_), .S(_06693_), .Y(_26170_) );
  \$mux  #( .WIDTH(33) ) _48977_ ( .A(_26170_), .B(33'h000000000), .S(RST), .Y(_02341_) );
  \$mux  #( .WIDTH(33) ) _48978_ ( .A(_source_stream_conv2d_16_source_8_pat_count_0), .B(_28640_), .S(_06691_), .Y(_26171_) );
  \$mux  #( .WIDTH(33) ) _48979_ ( .A(_28644_), .B(_26171_), .S(_05986_), .Y(_26172_) );
  \$mux  #( .WIDTH(33) ) _48980_ ( .A(_26172_), .B(_28645_), .S(_06692_), .Y(_26173_) );
  \$mux  #( .WIDTH(33) ) _48981_ ( .A(_26173_), .B(33'h000000000), .S(RST), .Y(_02340_) );
  \$mux  #( .WIDTH(32) ) _48982_ ( .A(_source_stream_conv2d_16_source_8_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_26174_) );
  \$mux  #( .WIDTH(32) ) _48983_ ( .A(_26174_), .B(0), .S(RST), .Y(_02359_) );
  \$mux  #( .WIDTH(32) ) _48984_ ( .A(_source_stream_conv2d_16_source_8_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_26175_) );
  \$mux  #( .WIDTH(32) ) _48985_ ( .A(_26175_), .B(0), .S(RST), .Y(_02358_) );
  \$mux  #( .WIDTH(32) ) _48986_ ( .A(_source_stream_conv2d_16_source_8_pat_stride_1), .B(0), .S(_set_flag_710), .Y(_26176_) );
  \$mux  #( .WIDTH(32) ) _48987_ ( .A(_26176_), .B(0), .S(RST), .Y(_02357_) );
  \$mux  #( .WIDTH(32) ) _48988_ ( .A(_source_stream_conv2d_16_source_8_pat_stride_0), .B(0), .S(_set_flag_710), .Y(_26177_) );
  \$mux  #( .WIDTH(32) ) _48989_ ( .A(_26177_), .B(0), .S(RST), .Y(_02356_) );
  \$mux  #( .WIDTH(33) ) _48990_ ( .A(_source_stream_conv2d_16_source_8_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_26178_) );
  \$mux  #( .WIDTH(33) ) _48991_ ( .A(_26178_), .B(33'h000000000), .S(RST), .Y(_02351_) );
  \$mux  #( .WIDTH(33) ) _48992_ ( .A(_source_stream_conv2d_16_source_8_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_26179_) );
  \$mux  #( .WIDTH(33) ) _48993_ ( .A(_26179_), .B(33'h000000000), .S(RST), .Y(_02350_) );
  \$mux  #( .WIDTH(33) ) _48994_ ( .A(_source_stream_conv2d_16_source_8_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_26180_) );
  \$mux  #( .WIDTH(33) ) _48995_ ( .A(_26180_), .B(33'h000000000), .S(RST), .Y(_02349_) );
  \$mux  #( .WIDTH(33) ) _48996_ ( .A(_source_stream_conv2d_16_source_8_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_26181_) );
  \$mux  #( .WIDTH(33) ) _48997_ ( .A(_26181_), .B(33'h000000000), .S(RST), .Y(_02348_) );
  \$mux  #( .WIDTH(32) ) _48998_ ( .A(_source_stream_conv2d_16_source_8_pat_cur_offset_3), .B(0), .S(_06691_), .Y(_26182_) );
  \$mux  #( .WIDTH(32) ) _48999_ ( .A(_26182_), .B(_24315_), .S(_06694_), .Y(_26183_) );
  \$mux  #( .WIDTH(32) ) _49000_ ( .A(_26183_), .B(0), .S(_06695_), .Y(_26184_) );
  \$mux  #( .WIDTH(32) ) _49001_ ( .A(_26184_), .B(0), .S(RST), .Y(_02347_) );
  \$mux  #( .WIDTH(32) ) _49002_ ( .A(_source_stream_conv2d_16_source_8_pat_cur_offset_2), .B(0), .S(_06691_), .Y(_26185_) );
  \$mux  #( .WIDTH(32) ) _49003_ ( .A(_26185_), .B(_24314_), .S(_06693_), .Y(_26186_) );
  \$mux  #( .WIDTH(32) ) _49004_ ( .A(_26186_), .B(0), .S(_06694_), .Y(_26187_) );
  \$mux  #( .WIDTH(32) ) _49005_ ( .A(_26187_), .B(0), .S(RST), .Y(_02346_) );
  \$mux  #( .WIDTH(32) ) _49006_ ( .A(_source_stream_conv2d_16_source_8_pat_cur_offset_1), .B(0), .S(_06691_), .Y(_26188_) );
  \$mux  #( .WIDTH(32) ) _49007_ ( .A(_26188_), .B(_24313_), .S(_06692_), .Y(_26189_) );
  \$mux  #( .WIDTH(32) ) _49008_ ( .A(_26189_), .B(0), .S(_06693_), .Y(_26190_) );
  \$mux  #( .WIDTH(32) ) _49009_ ( .A(_26190_), .B(0), .S(RST), .Y(_02345_) );
  \$mux  #( .WIDTH(32) ) _49010_ ( .A(_source_stream_conv2d_16_source_8_pat_cur_offset_0), .B(0), .S(_06691_), .Y(_26191_) );
  \$mux  #( .WIDTH(32) ) _49011_ ( .A(_24312_), .B(_26191_), .S(_05986_), .Y(_26192_) );
  \$mux  #( .WIDTH(32) ) _49012_ ( .A(_26192_), .B(0), .S(_06692_), .Y(_26193_) );
  \$mux  #( .WIDTH(32) ) _49013_ ( .A(_26193_), .B(0), .S(RST), .Y(_02344_) );
  \$mux  #( .WIDTH(8) ) _49014_ ( .A(__variable_wdata_230), .B(_stream_conv2d_16_source_6_source_ram_rdata), .S(_stream_conv2d_16_source_6_source_ram_rvalid), .Y(_26194_) );
  \$mux  #( .WIDTH(8) ) _49015_ ( .A(_26194_), .B(8'h00), .S(RST), .Y(_01400_) );
  \$mux  #( .WIDTH(32) ) _49016_ ( .A(_source_stream_conv2d_16_source_6_pat_stride_buf_3), .B(_source_stream_conv2d_16_source_6_pat_stride_3), .S(_06686_), .Y(_26195_) );
  \$mux  #( .WIDTH(32) ) _49017_ ( .A(_26195_), .B(0), .S(RST), .Y(_02339_) );
  \$mux  #( .WIDTH(32) ) _49018_ ( .A(_source_stream_conv2d_16_source_6_pat_stride_buf_2), .B(_source_stream_conv2d_16_source_6_pat_stride_2), .S(_06686_), .Y(_26196_) );
  \$mux  #( .WIDTH(32) ) _49019_ ( .A(_26196_), .B(0), .S(RST), .Y(_02338_) );
  \$mux  #( .WIDTH(32) ) _49020_ ( .A(_source_stream_conv2d_16_source_6_pat_stride_buf_1), .B(_source_stream_conv2d_16_source_6_pat_stride_1), .S(_06686_), .Y(_26197_) );
  \$mux  #( .WIDTH(32) ) _49021_ ( .A(_26197_), .B(0), .S(RST), .Y(_02337_) );
  \$mux  #( .WIDTH(32) ) _49022_ ( .A(_source_stream_conv2d_16_source_6_pat_stride_buf_0), .B(_source_stream_conv2d_16_source_6_pat_stride_0), .S(_06686_), .Y(_26198_) );
  \$mux  #( .WIDTH(32) ) _49023_ ( .A(_26198_), .B(0), .S(RST), .Y(_02336_) );
  \$mux  #( .WIDTH(33) ) _49024_ ( .A(_source_stream_conv2d_16_source_6_pat_size_buf_3), .B(_source_stream_conv2d_16_source_6_pat_size_3), .S(_06686_), .Y(_26199_) );
  \$mux  #( .WIDTH(33) ) _49025_ ( .A(_26199_), .B(33'h000000000), .S(RST), .Y(_02331_) );
  \$mux  #( .WIDTH(33) ) _49026_ ( .A(_source_stream_conv2d_16_source_6_pat_size_buf_2), .B(_source_stream_conv2d_16_source_6_pat_size_2), .S(_06686_), .Y(_26200_) );
  \$mux  #( .WIDTH(33) ) _49027_ ( .A(_26200_), .B(33'h000000000), .S(RST), .Y(_02330_) );
  \$mux  #( .WIDTH(33) ) _49028_ ( .A(_source_stream_conv2d_16_source_6_pat_size_buf_1), .B(_source_stream_conv2d_16_source_6_pat_size_1), .S(_06686_), .Y(_26201_) );
  \$mux  #( .WIDTH(33) ) _49029_ ( .A(_26201_), .B(33'h000000000), .S(RST), .Y(_02329_) );
  \$mux  #( .WIDTH(33) ) _49030_ ( .A(_source_stream_conv2d_16_source_6_pat_size_buf_0), .B(_source_stream_conv2d_16_source_6_pat_size_0), .S(_06686_), .Y(_26202_) );
  \$mux  #( .WIDTH(33) ) _49031_ ( .A(_26202_), .B(33'h000000000), .S(RST), .Y(_02328_) );
  \$mux  #( .WIDTH(33) ) _49032_ ( .A(_source_stream_conv2d_16_source_6_pat_count_3), .B(_28631_), .S(_06686_), .Y(_26203_) );
  \$mux  #( .WIDTH(33) ) _49033_ ( .A(_26203_), .B(_28638_), .S(_06689_), .Y(_26204_) );
  \$mux  #( .WIDTH(33) ) _49034_ ( .A(_26204_), .B(_28639_), .S(_06690_), .Y(_26205_) );
  \$mux  #( .WIDTH(33) ) _49035_ ( .A(_26205_), .B(33'h000000000), .S(RST), .Y(_02319_) );
  \$mux  #( .WIDTH(33) ) _49036_ ( .A(_source_stream_conv2d_16_source_6_pat_count_2), .B(_28630_), .S(_06686_), .Y(_26206_) );
  \$mux  #( .WIDTH(33) ) _49037_ ( .A(_26206_), .B(_28636_), .S(_06688_), .Y(_26207_) );
  \$mux  #( .WIDTH(33) ) _49038_ ( .A(_26207_), .B(_28637_), .S(_06689_), .Y(_26208_) );
  \$mux  #( .WIDTH(33) ) _49039_ ( .A(_26208_), .B(33'h000000000), .S(RST), .Y(_02318_) );
  \$mux  #( .WIDTH(33) ) _49040_ ( .A(_source_stream_conv2d_16_source_6_pat_count_1), .B(_28629_), .S(_06686_), .Y(_26209_) );
  \$mux  #( .WIDTH(33) ) _49041_ ( .A(_26209_), .B(_28634_), .S(_06687_), .Y(_26210_) );
  \$mux  #( .WIDTH(33) ) _49042_ ( .A(_26210_), .B(_28635_), .S(_06688_), .Y(_26211_) );
  \$mux  #( .WIDTH(33) ) _49043_ ( .A(_26211_), .B(33'h000000000), .S(RST), .Y(_02317_) );
  \$mux  #( .WIDTH(33) ) _49044_ ( .A(_source_stream_conv2d_16_source_6_pat_count_0), .B(_28628_), .S(_06686_), .Y(_26212_) );
  \$mux  #( .WIDTH(33) ) _49045_ ( .A(_28632_), .B(_26212_), .S(_05987_), .Y(_26213_) );
  \$mux  #( .WIDTH(33) ) _49046_ ( .A(_26213_), .B(_28633_), .S(_06687_), .Y(_26214_) );
  \$mux  #( .WIDTH(33) ) _49047_ ( .A(_26214_), .B(33'h000000000), .S(RST), .Y(_02316_) );
  \$mux  #( .WIDTH(32) ) _49048_ ( .A(_source_stream_conv2d_16_source_6_pat_stride_3), .B(0), .S(_set_flag_710), .Y(_26215_) );
  \$mux  #( .WIDTH(32) ) _49049_ ( .A(_26215_), .B(0), .S(RST), .Y(_02335_) );
  \$mux  #( .WIDTH(32) ) _49050_ ( .A(_source_stream_conv2d_16_source_6_pat_stride_2), .B(0), .S(_set_flag_710), .Y(_26216_) );
  \$mux  #( .WIDTH(32) ) _49051_ ( .A(_26216_), .B(0), .S(RST), .Y(_02334_) );
  \$mux  #( .WIDTH(32) ) _49052_ ( .A(_source_stream_conv2d_16_source_6_pat_stride_1), .B(_29232_), .S(_set_flag_710), .Y(_26217_) );
  \$mux  #( .WIDTH(32) ) _49053_ ( .A(_26217_), .B(0), .S(RST), .Y(_02333_) );
  \$mux  #( .WIDTH(32) ) _49054_ ( .A(_source_stream_conv2d_16_source_6_pat_stride_0), .B(0), .S(_set_flag_710), .Y(_26218_) );
  \$mux  #( .WIDTH(32) ) _49055_ ( .A(_26218_), .B(0), .S(RST), .Y(_02332_) );
  \$mux  #( .WIDTH(33) ) _49056_ ( .A(_source_stream_conv2d_16_source_6_pat_size_3), .B(33'h000000001), .S(_set_flag_710), .Y(_26219_) );
  \$mux  #( .WIDTH(33) ) _49057_ ( .A(_26219_), .B(33'h000000000), .S(RST), .Y(_02327_) );
  \$mux  #( .WIDTH(33) ) _49058_ ( .A(_source_stream_conv2d_16_source_6_pat_size_2), .B(33'h000000001), .S(_set_flag_710), .Y(_26220_) );
  \$mux  #( .WIDTH(33) ) _49059_ ( .A(_26220_), .B(33'h000000000), .S(RST), .Y(_02326_) );
  \$mux  #( .WIDTH(33) ) _49060_ ( .A(_source_stream_conv2d_16_source_6_pat_size_1), .B({ 1'h0, conv2d_16_next_stream_num_ops }), .S(_set_flag_710), .Y(_26221_) );
  \$mux  #( .WIDTH(33) ) _49061_ ( .A(_26221_), .B(33'h000000000), .S(RST), .Y(_02325_) );
  \$mux  #( .WIDTH(33) ) _49062_ ( .A(_source_stream_conv2d_16_source_6_pat_size_0), .B({ 27'h0000000, cparam_conv2d_16_stream_reduce_size }), .S(_set_flag_710), .Y(_26222_) );
  \$mux  #( .WIDTH(33) ) _49063_ ( .A(_26222_), .B(33'h000000000), .S(RST), .Y(_02324_) );
  \$mux  #( .WIDTH(32) ) _49064_ ( .A(_source_stream_conv2d_16_source_6_pat_cur_offset_3), .B(0), .S(_06686_), .Y(_26223_) );
  \$mux  #( .WIDTH(32) ) _49065_ ( .A(_26223_), .B(_24311_), .S(_06689_), .Y(_26224_) );
  \$mux  #( .WIDTH(32) ) _49066_ ( .A(_26224_), .B(0), .S(_06690_), .Y(_26225_) );
  \$mux  #( .WIDTH(32) ) _49067_ ( .A(_26225_), .B(0), .S(RST), .Y(_02323_) );
  \$mux  #( .WIDTH(32) ) _49068_ ( .A(_source_stream_conv2d_16_source_6_pat_cur_offset_2), .B(0), .S(_06686_), .Y(_26226_) );
  \$mux  #( .WIDTH(32) ) _49069_ ( .A(_26226_), .B(_24310_), .S(_06688_), .Y(_26227_) );
  \$mux  #( .WIDTH(32) ) _49070_ ( .A(_26227_), .B(0), .S(_06689_), .Y(_26228_) );
  \$mux  #( .WIDTH(32) ) _49071_ ( .A(_26228_), .B(0), .S(RST), .Y(_02322_) );
  \$mux  #( .WIDTH(32) ) _49072_ ( .A(_source_stream_conv2d_16_source_6_pat_cur_offset_1), .B(0), .S(_06686_), .Y(_26229_) );
  \$mux  #( .WIDTH(32) ) _49073_ ( .A(_26229_), .B(_24309_), .S(_06687_), .Y(_26230_) );
  \$mux  #( .WIDTH(32) ) _49074_ ( .A(_26230_), .B(0), .S(_06688_), .Y(_26231_) );
  \$mux  #( .WIDTH(32) ) _49075_ ( .A(_26231_), .B(0), .S(RST), .Y(_02321_) );
  \$mux  #( .WIDTH(32) ) _49076_ ( .A(_source_stream_conv2d_16_source_6_pat_cur_offset_0), .B(0), .S(_06686_), .Y(_26232_) );
  \$mux  #( .WIDTH(32) ) _49077_ ( .A(_24308_), .B(_26232_), .S(_05987_), .Y(_26233_) );
  \$mux  #( .WIDTH(32) ) _49078_ ( .A(_26233_), .B(0), .S(_06687_), .Y(_26234_) );
  \$mux  #( .WIDTH(32) ) _49079_ ( .A(_26234_), .B(0), .S(RST), .Y(_02320_) );
  \$mux  #( .WIDTH(9) ) _49080_ ( .A(__variable_wdata_217), .B(_stream_conv2d_16_constant_3_next_constant_data), .S(_stream_conv2d_16_start), .Y(_26235_) );
  \$mux  #( .WIDTH(9) ) _49081_ ( .A(_26235_), .B(9'h000), .S(RST), .Y(_01398_) );
  \$mux  #( .WIDTH(2) ) _49082_ ( .A(__variable_wdata_216), .B(_stream_conv2d_16_constant_2_next_constant_data), .S(_stream_conv2d_16_start), .Y(_26236_) );
  \$mux  #( .WIDTH(2) ) _49083_ ( .A(_26236_), .B(2'h0), .S(RST), .Y(_01397_) );
  \$mux  #( .WIDTH(2) ) _49084_ ( .A(__variable_wdata_215), .B(_stream_conv2d_16_constant_1_next_constant_data), .S(_stream_conv2d_16_start), .Y(_26237_) );
  \$mux  #( .WIDTH(2) ) _49085_ ( .A(_26237_), .B(2'h0), .S(RST), .Y(_01396_) );
  \$mux  #( .WIDTH(6) ) _49086_ ( .A(__variable_wdata_214), .B(_stream_conv2d_16_constant_0_next_constant_data), .S(_stream_conv2d_16_start), .Y(_26238_) );
  \$mux  #( .WIDTH(6) ) _49087_ ( .A(_26238_), .B(6'h00), .S(RST), .Y(_01395_) );
  \$mux  #( .WIDTH(1) ) _49088_ ( .A(1'h1), .B(1'h0), .S(_05989_), .Y(_25408_) );
  \$mux  #( .WIDTH(1) ) _49089_ ( .A(_25408_), .B(1'h0), .S(RST), .Y(_01873_) );
  \$mux  #( .WIDTH(1) ) _49090_ ( .A(__delay_data_1613), .B(1'h0), .S(RST), .Y(_00291_) );
  \$mux  #( .WIDTH(8) ) _49091_ ( .A(_29230_), .B(8'h00), .S(RST), .Y(_01547_) );
  \$mux  #( .WIDTH(1) ) _49092_ ( .A(__delay_data_1612), .B(1'h0), .S(RST), .Y(_00290_) );
  \$mux  #( .WIDTH(8) ) _49093_ ( .A(__substreamoutput_data_886), .B(8'h00), .S(RST), .Y(_00278_) );
  \$mux  #( .WIDTH(1) ) _49094_ ( .A(_06174_), .B(1'h0), .S(RST), .Y(_01701_) );
  \$mux  #( .WIDTH(1) ) _49095_ ( .A(__delay_data_1611), .B(1'h0), .S(RST), .Y(_00289_) );
  \$mux  #( .WIDTH(8) ) _49096_ ( .A(_cond_data_53), .B(8'h00), .S(RST), .Y(_01101_) );
  \$mux  #( .WIDTH(1) ) _49097_ ( .A(__delay_data_1610), .B(1'h0), .S(RST), .Y(_00288_) );
  \$mux  #( .WIDTH(1) ) _49098_ ( .A(__delay_data_1609), .B(1'h0), .S(RST), .Y(_00287_) );
  \$mux  #( .WIDTH(1) ) _49099_ ( .A(__delay_data_1608), .B(1'h0), .S(RST), .Y(_00286_) );
  \$mux  #( .WIDTH(1) ) _49100_ ( .A(__delay_data_1607), .B(1'h0), .S(RST), .Y(_00285_) );
  \$mux  #( .WIDTH(1) ) _49101_ ( .A(__delay_data_1606), .B(1'h0), .S(RST), .Y(_00284_) );
  \$mux  #( .WIDTH(1) ) _49102_ ( .A(__delay_data_1605), .B(1'h0), .S(RST), .Y(_00283_) );
  \$mux  #( .WIDTH(1) ) _49103_ ( .A(__delay_data_1604), .B(1'h0), .S(RST), .Y(_00282_) );
  \$mux  #( .WIDTH(1) ) _49104_ ( .A(__delay_data_1603), .B(1'h0), .S(RST), .Y(_00281_) );
  \$mux  #( .WIDTH(1) ) _49105_ ( .A(__delay_data_1602), .B(1'h0), .S(RST), .Y(_00280_) );
  \$mux  #( .WIDTH(1) ) _49106_ ( .A(__substreamoutput_data_882), .B(1'h0), .S(RST), .Y(_00279_) );
  \$mux  #( .WIDTH(8) ) _49107_ ( .A(__delay_data_1395), .B(8'h00), .S(RST), .Y(_00277_) );
  \$mux  #( .WIDTH(8) ) _49108_ ( .A(__delay_data_1367), .B(8'h00), .S(RST), .Y(_00249_) );
  \$mux  #( .WIDTH(32) ) _49109_ ( .A(_24307_), .B(0), .S(RST), .Y(_01813_) );
  \$mux  #( .WIDTH(8) ) _49110_ ( .A(__delay_data_1394), .B(8'h00), .S(RST), .Y(_00276_) );
  \$mux  #( .WIDTH(8) ) _49111_ ( .A(__delay_data_1366), .B(8'h00), .S(RST), .Y(_00248_) );
  \$mux  #( .WIDTH(8) ) _49112_ ( .A(__delay_data_1337), .B(8'h00), .S(RST), .Y(_00219_) );
  \$mux  #( .WIDTH(1) ) _49113_ ( .A(__delay_data_758), .B(1'h0), .S(RST), .Y(_01100_) );
  \$mux  #( .WIDTH(32) ) _49114_ ( .A(_sra_data_21), .B(0), .S(RST), .Y(_01099_) );
  \$mux  #( .WIDTH(8) ) _49115_ ( .A(__delay_data_1393), .B(8'h00), .S(RST), .Y(_00275_) );
  \$mux  #( .WIDTH(8) ) _49116_ ( .A(__delay_data_1365), .B(8'h00), .S(RST), .Y(_00247_) );
  \$mux  #( .WIDTH(8) ) _49117_ ( .A(__delay_data_1336), .B(8'h00), .S(RST), .Y(_00218_) );
  \$mux  #( .WIDTH(8) ) _49118_ ( .A(__delay_data_1392), .B(8'h00), .S(RST), .Y(_00274_) );
  \$mux  #( .WIDTH(8) ) _49119_ ( .A(__delay_data_1364), .B(8'h00), .S(RST), .Y(_00246_) );
  \$mux  #( .WIDTH(8) ) _49120_ ( .A(__delay_data_1335), .B(8'h00), .S(RST), .Y(_00217_) );
  \$mux  #( .WIDTH(8) ) _49121_ ( .A(__delay_data_1391), .B(8'h00), .S(RST), .Y(_00273_) );
  \$mux  #( .WIDTH(8) ) _49122_ ( .A(__delay_data_1363), .B(8'h00), .S(RST), .Y(_00245_) );
  \$mux  #( .WIDTH(8) ) _49123_ ( .A(__delay_data_1334), .B(8'h00), .S(RST), .Y(_00216_) );
  \$mux  #( .WIDTH(8) ) _49124_ ( .A(__delay_data_1390), .B(8'h00), .S(RST), .Y(_00272_) );
  \$mux  #( .WIDTH(8) ) _49125_ ( .A(__delay_data_1362), .B(8'h00), .S(RST), .Y(_00244_) );
  \$mux  #( .WIDTH(8) ) _49126_ ( .A(__delay_data_1333), .B(8'h00), .S(RST), .Y(_00215_) );
  \$mux  #( .WIDTH(8) ) _49127_ ( .A(__delay_data_1389), .B(8'h00), .S(RST), .Y(_00271_) );
  \$mux  #( .WIDTH(8) ) _49128_ ( .A(__delay_data_1361), .B(8'h00), .S(RST), .Y(_00243_) );
  \$mux  #( .WIDTH(8) ) _49129_ ( .A(__delay_data_1332), .B(8'h00), .S(RST), .Y(_00214_) );
  \$mux  #( .WIDTH(8) ) _49130_ ( .A(__delay_data_1388), .B(8'h00), .S(RST), .Y(_00270_) );
  \$mux  #( .WIDTH(8) ) _49131_ ( .A(__delay_data_1360), .B(8'h00), .S(RST), .Y(_00242_) );
  \$mux  #( .WIDTH(8) ) _49132_ ( .A(__delay_data_1331), .B(8'h00), .S(RST), .Y(_00213_) );
  \$mux  #( .WIDTH(8) ) _49133_ ( .A(__delay_data_1387), .B(8'h00), .S(RST), .Y(_00269_) );
  \$mux  #( .WIDTH(8) ) _49134_ ( .A(__delay_data_1359), .B(8'h00), .S(RST), .Y(_00241_) );
  \$mux  #( .WIDTH(8) ) _49135_ ( .A(__delay_data_1330), .B(8'h00), .S(RST), .Y(_00212_) );
  \$mux  #( .WIDTH(6) ) _49136_ ( .A(__delay_data_1309), .B(6'h00), .S(RST), .Y(_00191_) );
  \$mux  #( .WIDTH(8) ) _49137_ ( .A(__delay_data_1287), .B(8'h00), .S(RST), .Y(_00169_) );
  \$mux  #( .WIDTH(32) ) _49138_ ( .A(__plusn_data_37), .B(0), .S(RST), .Y(_01098_) );
  \$mux  #( .WIDTH(8) ) _49139_ ( .A(__delay_data_1386), .B(8'h00), .S(RST), .Y(_00268_) );
  \$mux  #( .WIDTH(8) ) _49140_ ( .A(__delay_data_1358), .B(8'h00), .S(RST), .Y(_00240_) );
  \$mux  #( .WIDTH(8) ) _49141_ ( .A(__delay_data_1329), .B(8'h00), .S(RST), .Y(_00211_) );
  \$mux  #( .WIDTH(6) ) _49142_ ( .A(__delay_data_1308), .B(6'h00), .S(RST), .Y(_00190_) );
  \$mux  #( .WIDTH(8) ) _49143_ ( .A(__delay_data_1286), .B(8'h00), .S(RST), .Y(_00168_) );
  \$mux  #( .WIDTH(8) ) _49144_ ( .A(__delay_data_1385), .B(8'h00), .S(RST), .Y(_00267_) );
  \$mux  #( .WIDTH(8) ) _49145_ ( .A(__delay_data_1357), .B(8'h00), .S(RST), .Y(_00239_) );
  \$mux  #( .WIDTH(8) ) _49146_ ( .A(__delay_data_1328), .B(8'h00), .S(RST), .Y(_00210_) );
  \$mux  #( .WIDTH(6) ) _49147_ ( .A(__delay_data_1307), .B(6'h00), .S(RST), .Y(_00189_) );
  \$mux  #( .WIDTH(8) ) _49148_ ( .A(__delay_data_1285), .B(8'h00), .S(RST), .Y(_00167_) );
  \$mux  #( .WIDTH(8) ) _49149_ ( .A(__delay_data_1384), .B(8'h00), .S(RST), .Y(_00266_) );
  \$mux  #( .WIDTH(8) ) _49150_ ( .A(__delay_data_1356), .B(8'h00), .S(RST), .Y(_00238_) );
  \$mux  #( .WIDTH(8) ) _49151_ ( .A(__delay_data_1327), .B(8'h00), .S(RST), .Y(_00209_) );
  \$mux  #( .WIDTH(6) ) _49152_ ( .A(__delay_data_1306), .B(6'h00), .S(RST), .Y(_00188_) );
  \$mux  #( .WIDTH(8) ) _49153_ ( .A(__delay_data_1284), .B(8'h00), .S(RST), .Y(_00166_) );
  \$mux  #( .WIDTH(8) ) _49154_ ( .A(__delay_data_1383), .B(8'h00), .S(RST), .Y(_00265_) );
  \$mux  #( .WIDTH(8) ) _49155_ ( .A(__delay_data_1355), .B(8'h00), .S(RST), .Y(_00237_) );
  \$mux  #( .WIDTH(8) ) _49156_ ( .A(__delay_data_1326), .B(8'h00), .S(RST), .Y(_00208_) );
  \$mux  #( .WIDTH(6) ) _49157_ ( .A(__delay_data_1305), .B(6'h00), .S(RST), .Y(_00187_) );
  \$mux  #( .WIDTH(8) ) _49158_ ( .A(__delay_data_1283), .B(8'h00), .S(RST), .Y(_00165_) );
  \$mux  #( .WIDTH(12) ) _49159_ ( .A(_sra_data_206), .B(12'h000), .S(RST), .Y(_01097_) );
  \$mux  #( .WIDTH(12) ) _49160_ ( .A(_sra_data_189), .B(12'h000), .S(RST), .Y(_01096_) );
  \$mux  #( .WIDTH(12) ) _49161_ ( .A(_sra_data_172), .B(12'h000), .S(RST), .Y(_01095_) );
  \$mux  #( .WIDTH(12) ) _49162_ ( .A(_sra_data_155), .B(12'h000), .S(RST), .Y(_01094_) );
  \$mux  #( .WIDTH(12) ) _49163_ ( .A(_sra_data_138), .B(12'h000), .S(RST), .Y(_01093_) );
  \$mux  #( .WIDTH(12) ) _49164_ ( .A(_sra_data_121), .B(12'h000), .S(RST), .Y(_01092_) );
  \$mux  #( .WIDTH(12) ) _49165_ ( .A(_sra_data_104), .B(12'h000), .S(RST), .Y(_01091_) );
  \$mux  #( .WIDTH(12) ) _49166_ ( .A(_sra_data_87), .B(12'h000), .S(RST), .Y(_01090_) );
  \$mux  #( .WIDTH(12) ) _49167_ ( .A(_sra_data_70), .B(12'h000), .S(RST), .Y(_01089_) );
  \$mux  #( .WIDTH(8) ) _49168_ ( .A(__delay_data_1382), .B(8'h00), .S(RST), .Y(_00264_) );
  \$mux  #( .WIDTH(8) ) _49169_ ( .A(__delay_data_1354), .B(8'h00), .S(RST), .Y(_00236_) );
  \$mux  #( .WIDTH(8) ) _49170_ ( .A(__delay_data_1325), .B(8'h00), .S(RST), .Y(_00207_) );
  \$mux  #( .WIDTH(6) ) _49171_ ( .A(__delay_data_1304), .B(6'h00), .S(RST), .Y(_00186_) );
  \$mux  #( .WIDTH(8) ) _49172_ ( .A(__delay_data_1282), .B(8'h00), .S(RST), .Y(_00164_) );
  \$mux  #( .WIDTH(8) ) _49173_ ( .A(__delay_data_1381), .B(8'h00), .S(RST), .Y(_00263_) );
  \$mux  #( .WIDTH(8) ) _49174_ ( .A(__delay_data_1353), .B(8'h00), .S(RST), .Y(_00235_) );
  \$mux  #( .WIDTH(8) ) _49175_ ( .A(__delay_data_1324), .B(8'h00), .S(RST), .Y(_00206_) );
  \$mux  #( .WIDTH(6) ) _49176_ ( .A(__delay_data_1303), .B(6'h00), .S(RST), .Y(_00185_) );
  \$mux  #( .WIDTH(8) ) _49177_ ( .A(__delay_data_1281), .B(8'h00), .S(RST), .Y(_00163_) );
  \$mux  #( .WIDTH(8) ) _49178_ ( .A(__delay_data_1380), .B(8'h00), .S(RST), .Y(_00262_) );
  \$mux  #( .WIDTH(8) ) _49179_ ( .A(__delay_data_1352), .B(8'h00), .S(RST), .Y(_00234_) );
  \$mux  #( .WIDTH(8) ) _49180_ ( .A(__delay_data_1323), .B(8'h00), .S(RST), .Y(_00205_) );
  \$mux  #( .WIDTH(6) ) _49181_ ( .A(__delay_data_1302), .B(6'h00), .S(RST), .Y(_00184_) );
  \$mux  #( .WIDTH(8) ) _49182_ ( .A(__delay_data_1280), .B(8'h00), .S(RST), .Y(_00162_) );
  \$mux  #( .WIDTH(8) ) _49183_ ( .A(__delay_data_1379), .B(8'h00), .S(RST), .Y(_00261_) );
  \$mux  #( .WIDTH(8) ) _49184_ ( .A(__delay_data_1351), .B(8'h00), .S(RST), .Y(_00233_) );
  \$mux  #( .WIDTH(8) ) _49185_ ( .A(__delay_data_1322), .B(8'h00), .S(RST), .Y(_00204_) );
  \$mux  #( .WIDTH(6) ) _49186_ ( .A(__delay_data_1301), .B(6'h00), .S(RST), .Y(_00183_) );
  \$mux  #( .WIDTH(8) ) _49187_ ( .A(__delay_data_1279), .B(8'h00), .S(RST), .Y(_00161_) );
  \$mux  #( .WIDTH(8) ) _49188_ ( .A(__delay_data_1378), .B(8'h00), .S(RST), .Y(_00260_) );
  \$mux  #( .WIDTH(8) ) _49189_ ( .A(__delay_data_1350), .B(8'h00), .S(RST), .Y(_00232_) );
  \$mux  #( .WIDTH(8) ) _49190_ ( .A(__delay_data_1321), .B(8'h00), .S(RST), .Y(_00203_) );
  \$mux  #( .WIDTH(6) ) _49191_ ( .A(__delay_data_1300), .B(6'h00), .S(RST), .Y(_00182_) );
  \$mux  #( .WIDTH(8) ) _49192_ ( .A(__delay_data_1278), .B(8'h00), .S(RST), .Y(_00160_) );
  \$mux  #( .WIDTH(8) ) _49193_ ( .A(__delay_data_1377), .B(8'h00), .S(RST), .Y(_00259_) );
  \$mux  #( .WIDTH(8) ) _49194_ ( .A(__delay_data_1349), .B(8'h00), .S(RST), .Y(_00231_) );
  \$mux  #( .WIDTH(8) ) _49195_ ( .A(__delay_data_1320), .B(8'h00), .S(RST), .Y(_00202_) );
  \$mux  #( .WIDTH(6) ) _49196_ ( .A(__delay_data_1299), .B(6'h00), .S(RST), .Y(_00181_) );
  \$mux  #( .WIDTH(8) ) _49197_ ( .A(__delay_data_1277), .B(8'h00), .S(RST), .Y(_00159_) );
  \$mux  #( .WIDTH(8) ) _49198_ ( .A(__delay_data_1376), .B(8'h00), .S(RST), .Y(_00258_) );
  \$mux  #( .WIDTH(8) ) _49199_ ( .A(__delay_data_1348), .B(8'h00), .S(RST), .Y(_00230_) );
  \$mux  #( .WIDTH(8) ) _49200_ ( .A(__delay_data_1319), .B(8'h00), .S(RST), .Y(_00201_) );
  \$mux  #( .WIDTH(6) ) _49201_ ( .A(__delay_data_1298), .B(6'h00), .S(RST), .Y(_00180_) );
  \$mux  #( .WIDTH(8) ) _49202_ ( .A(__delay_data_1276), .B(8'h00), .S(RST), .Y(_00158_) );
  \$mux  #( .WIDTH(8) ) _49203_ ( .A(__delay_data_1375), .B(8'h00), .S(RST), .Y(_00257_) );
  \$mux  #( .WIDTH(8) ) _49204_ ( .A(__delay_data_1347), .B(8'h00), .S(RST), .Y(_00229_) );
  \$mux  #( .WIDTH(8) ) _49205_ ( .A(__delay_data_1318), .B(8'h00), .S(RST), .Y(_00200_) );
  \$mux  #( .WIDTH(6) ) _49206_ ( .A(__delay_data_1297), .B(6'h00), .S(RST), .Y(_00179_) );
  \$mux  #( .WIDTH(8) ) _49207_ ( .A(__delay_data_1275), .B(8'h00), .S(RST), .Y(_00157_) );
  \$mux  #( .WIDTH(8) ) _49208_ ( .A(__delay_data_1374), .B(8'h00), .S(RST), .Y(_00256_) );
  \$mux  #( .WIDTH(8) ) _49209_ ( .A(__delay_data_1346), .B(8'h00), .S(RST), .Y(_00228_) );
  \$mux  #( .WIDTH(8) ) _49210_ ( .A(__delay_data_1317), .B(8'h00), .S(RST), .Y(_00199_) );
  \$mux  #( .WIDTH(6) ) _49211_ ( .A(__delay_data_1296), .B(6'h00), .S(RST), .Y(_00178_) );
  \$mux  #( .WIDTH(8) ) _49212_ ( .A(__delay_data_1274), .B(8'h00), .S(RST), .Y(_00156_) );
  \$mux  #( .WIDTH(8) ) _49213_ ( .A(__delay_data_1373), .B(8'h00), .S(RST), .Y(_00255_) );
  \$mux  #( .WIDTH(8) ) _49214_ ( .A(__delay_data_1345), .B(8'h00), .S(RST), .Y(_00227_) );
  \$mux  #( .WIDTH(8) ) _49215_ ( .A(__delay_data_1316), .B(8'h00), .S(RST), .Y(_00198_) );
  \$mux  #( .WIDTH(6) ) _49216_ ( .A(__delay_data_1295), .B(6'h00), .S(RST), .Y(_00177_) );
  \$mux  #( .WIDTH(8) ) _49217_ ( .A(__delay_data_1273), .B(8'h00), .S(RST), .Y(_00155_) );
  \$mux  #( .WIDTH(4) ) _49218_ ( .A(__delay_data_1260), .B(4'h0), .S(RST), .Y(_00148_) );
  \$mux  #( .WIDTH(4) ) _49219_ ( .A(__delay_data_1226), .B(4'h0), .S(RST), .Y(_00132_) );
  \$mux  #( .WIDTH(4) ) _49220_ ( .A(__delay_data_1192), .B(4'h0), .S(RST), .Y(_00116_) );
  \$mux  #( .WIDTH(4) ) _49221_ ( .A(__delay_data_1158), .B(4'h0), .S(RST), .Y(_00100_) );
  \$mux  #( .WIDTH(4) ) _49222_ ( .A(__delay_data_1123), .B(4'h0), .S(RST), .Y(_00083_) );
  \$mux  #( .WIDTH(4) ) _49223_ ( .A(__delay_data_1088), .B(4'h0), .S(RST), .Y(_00066_) );
  \$mux  #( .WIDTH(4) ) _49224_ ( .A(__delay_data_1053), .B(4'h0), .S(RST), .Y(_00049_) );
  \$mux  #( .WIDTH(4) ) _49225_ ( .A(__delay_data_1005), .B(4'h0), .S(RST), .Y(_00007_) );
  \$mux  #( .WIDTH(8) ) _49226_ ( .A(__delay_data_1266), .B(8'h00), .S(RST), .Y(_00013_) );
  \$mux  #( .WIDTH(4) ) _49227_ ( .A(__delay_data_954), .B(4'h0), .S(RST), .Y(_00663_) );
  \$mux  #( .WIDTH(8) ) _49228_ ( .A(_29229_), .B(8'h00), .S(RST), .Y(_01545_) );
  \$mux  #( .WIDTH(8) ) _49229_ ( .A(_29228_), .B(8'h00), .S(RST), .Y(_01544_) );
  \$mux  #( .WIDTH(8) ) _49230_ ( .A(_29227_), .B(8'h00), .S(RST), .Y(_01543_) );
  \$mux  #( .WIDTH(8) ) _49231_ ( .A(_29226_), .B(8'h00), .S(RST), .Y(_01542_) );
  \$mux  #( .WIDTH(8) ) _49232_ ( .A(_29225_), .B(8'h00), .S(RST), .Y(_01541_) );
  \$mux  #( .WIDTH(8) ) _49233_ ( .A(_29224_), .B(8'h00), .S(RST), .Y(_01540_) );
  \$mux  #( .WIDTH(8) ) _49234_ ( .A(_29223_), .B(8'h00), .S(RST), .Y(_01539_) );
  \$mux  #( .WIDTH(8) ) _49235_ ( .A(_29222_), .B(8'h00), .S(RST), .Y(_01538_) );
  \$mux  #( .WIDTH(8) ) _49236_ ( .A(_29221_), .B(8'h00), .S(RST), .Y(_01537_) );
  \$mux  #( .WIDTH(8) ) _49237_ ( .A(__delay_data_1372), .B(8'h00), .S(RST), .Y(_00254_) );
  \$mux  #( .WIDTH(8) ) _49238_ ( .A(__delay_data_1344), .B(8'h00), .S(RST), .Y(_00226_) );
  \$mux  #( .WIDTH(8) ) _49239_ ( .A(__delay_data_1315), .B(8'h00), .S(RST), .Y(_00197_) );
  \$mux  #( .WIDTH(6) ) _49240_ ( .A(__delay_data_1294), .B(6'h00), .S(RST), .Y(_00176_) );
  \$mux  #( .WIDTH(8) ) _49241_ ( .A(__delay_data_1272), .B(8'h00), .S(RST), .Y(_00154_) );
  \$mux  #( .WIDTH(4) ) _49242_ ( .A(__delay_data_1259), .B(4'h0), .S(RST), .Y(_00147_) );
  \$mux  #( .WIDTH(1) ) _49243_ ( .A(__delay_data_1252), .B(1'h0), .S(RST), .Y(_00140_) );
  \$mux  #( .WIDTH(4) ) _49244_ ( .A(__delay_data_1225), .B(4'h0), .S(RST), .Y(_00131_) );
  \$mux  #( .WIDTH(1) ) _49245_ ( .A(__delay_data_1218), .B(1'h0), .S(RST), .Y(_00124_) );
  \$mux  #( .WIDTH(4) ) _49246_ ( .A(__delay_data_1191), .B(4'h0), .S(RST), .Y(_00115_) );
  \$mux  #( .WIDTH(1) ) _49247_ ( .A(__delay_data_1184), .B(1'h0), .S(RST), .Y(_00108_) );
  \$mux  #( .WIDTH(4) ) _49248_ ( .A(__delay_data_1157), .B(4'h0), .S(RST), .Y(_00099_) );
  \$mux  #( .WIDTH(1) ) _49249_ ( .A(__delay_data_1150), .B(1'h0), .S(RST), .Y(_00092_) );
  \$mux  #( .WIDTH(4) ) _49250_ ( .A(__delay_data_1122), .B(4'h0), .S(RST), .Y(_00082_) );
  \$mux  #( .WIDTH(1) ) _49251_ ( .A(__delay_data_1115), .B(1'h0), .S(RST), .Y(_00075_) );
  \$mux  #( .WIDTH(4) ) _49252_ ( .A(__delay_data_1087), .B(4'h0), .S(RST), .Y(_00065_) );
  \$mux  #( .WIDTH(1) ) _49253_ ( .A(__delay_data_1080), .B(1'h0), .S(RST), .Y(_00058_) );
  \$mux  #( .WIDTH(4) ) _49254_ ( .A(__delay_data_1052), .B(4'h0), .S(RST), .Y(_00048_) );
  \$mux  #( .WIDTH(1) ) _49255_ ( .A(__delay_data_1045), .B(1'h0), .S(RST), .Y(_00041_) );
  \$mux  #( .WIDTH(4) ) _49256_ ( .A(__delay_data_1004), .B(4'h0), .S(RST), .Y(_00006_) );
  \$mux  #( .WIDTH(1) ) _49257_ ( .A(__delay_data_997), .B(1'h0), .S(RST), .Y(_00679_) );
  \$mux  #( .WIDTH(8) ) _49258_ ( .A(__delay_data_1265), .B(8'h00), .S(RST), .Y(_00012_) );
  \$mux  #( .WIDTH(4) ) _49259_ ( .A(__delay_data_953), .B(4'h0), .S(RST), .Y(_00662_) );
  \$mux  #( .WIDTH(1) ) _49260_ ( .A(__delay_data_945), .B(1'h0), .S(RST), .Y(_00654_) );
  \$mux  #( .WIDTH(8) ) _49261_ ( .A(_29220_), .B(8'h00), .S(RST), .Y(_01533_) );
  \$mux  #( .WIDTH(8) ) _49262_ ( .A(_29219_), .B(8'h00), .S(RST), .Y(_01530_) );
  \$mux  #( .WIDTH(8) ) _49263_ ( .A(_29218_), .B(8'h00), .S(RST), .Y(_01527_) );
  \$mux  #( .WIDTH(8) ) _49264_ ( .A(_29217_), .B(8'h00), .S(RST), .Y(_01524_) );
  \$mux  #( .WIDTH(8) ) _49265_ ( .A(_29216_), .B(8'h00), .S(RST), .Y(_01521_) );
  \$mux  #( .WIDTH(8) ) _49266_ ( .A(_29215_), .B(8'h00), .S(RST), .Y(_01518_) );
  \$mux  #( .WIDTH(8) ) _49267_ ( .A(_29214_), .B(8'h00), .S(RST), .Y(_01515_) );
  \$mux  #( .WIDTH(8) ) _49268_ ( .A(_29213_), .B(8'h00), .S(RST), .Y(_01512_) );
  \$mux  #( .WIDTH(8) ) _49269_ ( .A(_29212_), .B(8'h00), .S(RST), .Y(_01509_) );
  \$mux  #( .WIDTH(8) ) _49270_ ( .A(__delay_data_1371), .B(8'h00), .S(RST), .Y(_00253_) );
  \$mux  #( .WIDTH(8) ) _49271_ ( .A(__delay_data_1343), .B(8'h00), .S(RST), .Y(_00225_) );
  \$mux  #( .WIDTH(8) ) _49272_ ( .A(__delay_data_1314), .B(8'h00), .S(RST), .Y(_00196_) );
  \$mux  #( .WIDTH(6) ) _49273_ ( .A(__delay_data_1293), .B(6'h00), .S(RST), .Y(_00175_) );
  \$mux  #( .WIDTH(8) ) _49274_ ( .A(__delay_data_1271), .B(8'h00), .S(RST), .Y(_00153_) );
  \$mux  #( .WIDTH(4) ) _49275_ ( .A(__delay_data_1258), .B(4'h0), .S(RST), .Y(_00146_) );
  \$mux  #( .WIDTH(1) ) _49276_ ( .A(__delay_data_1251), .B(1'h0), .S(RST), .Y(_00139_) );
  \$mux  #( .WIDTH(8) ) _49277_ ( .A(__delay_data_1138), .B(8'h00), .S(RST), .Y(_00133_) );
  \$mux  #( .WIDTH(4) ) _49278_ ( .A(__delay_data_1224), .B(4'h0), .S(RST), .Y(_00130_) );
  \$mux  #( .WIDTH(1) ) _49279_ ( .A(__delay_data_1217), .B(1'h0), .S(RST), .Y(_00123_) );
  \$mux  #( .WIDTH(8) ) _49280_ ( .A(__delay_data_1103), .B(8'h00), .S(RST), .Y(_00117_) );
  \$mux  #( .WIDTH(4) ) _49281_ ( .A(__delay_data_1190), .B(4'h0), .S(RST), .Y(_00114_) );
  \$mux  #( .WIDTH(1) ) _49282_ ( .A(__delay_data_1183), .B(1'h0), .S(RST), .Y(_00107_) );
  \$mux  #( .WIDTH(8) ) _49283_ ( .A(__delay_data_1068), .B(8'h00), .S(RST), .Y(_00101_) );
  \$mux  #( .WIDTH(4) ) _49284_ ( .A(__delay_data_1156), .B(4'h0), .S(RST), .Y(_00098_) );
  \$mux  #( .WIDTH(1) ) _49285_ ( .A(__delay_data_1149), .B(1'h0), .S(RST), .Y(_00091_) );
  \$mux  #( .WIDTH(8) ) _49286_ ( .A(__delay_data_1032), .B(8'h00), .S(RST), .Y(_00085_) );
  \$mux  #( .WIDTH(4) ) _49287_ ( .A(__delay_data_1121), .B(4'h0), .S(RST), .Y(_00081_) );
  \$mux  #( .WIDTH(1) ) _49288_ ( .A(__delay_data_1114), .B(1'h0), .S(RST), .Y(_00074_) );
  \$mux  #( .WIDTH(8) ) _49289_ ( .A(__delay_data_984), .B(8'h00), .S(RST), .Y(_00068_) );
  \$mux  #( .WIDTH(4) ) _49290_ ( .A(__delay_data_1086), .B(4'h0), .S(RST), .Y(_00064_) );
  \$mux  #( .WIDTH(1) ) _49291_ ( .A(__delay_data_1079), .B(1'h0), .S(RST), .Y(_00057_) );
  \$mux  #( .WIDTH(8) ) _49292_ ( .A(__delay_data_932), .B(8'h00), .S(RST), .Y(_00051_) );
  \$mux  #( .WIDTH(4) ) _49293_ ( .A(__delay_data_1051), .B(4'h0), .S(RST), .Y(_00047_) );
  \$mux  #( .WIDTH(1) ) _49294_ ( .A(__delay_data_1044), .B(1'h0), .S(RST), .Y(_00040_) );
  \$mux  #( .WIDTH(8) ) _49295_ ( .A(__delay_data_1038), .B(8'h00), .S(RST), .Y(_00034_) );
  \$mux  #( .WIDTH(4) ) _49296_ ( .A(__delay_data_1003), .B(4'h0), .S(RST), .Y(_00005_) );
  \$mux  #( .WIDTH(1) ) _49297_ ( .A(__delay_data_996), .B(1'h0), .S(RST), .Y(_00678_) );
  \$mux  #( .WIDTH(8) ) _49298_ ( .A(__delay_data_990), .B(8'h00), .S(RST), .Y(_00672_) );
  \$mux  #( .WIDTH(8) ) _49299_ ( .A(__delay_data_1264), .B(8'h00), .S(RST), .Y(_00011_) );
  \$mux  #( .WIDTH(4) ) _49300_ ( .A(__delay_data_952), .B(4'h0), .S(RST), .Y(_00661_) );
  \$mux  #( .WIDTH(1) ) _49301_ ( .A(__delay_data_944), .B(1'h0), .S(RST), .Y(_00653_) );
  \$mux  #( .WIDTH(8) ) _49302_ ( .A(__delay_data_938), .B(8'h00), .S(RST), .Y(_00647_) );
  \$mux  #( .WIDTH(1) ) _49303_ ( .A(__delay_data_1244), .B(1'h0), .S(RST), .Y(_00032_) );
  \$mux  #( .WIDTH(8) ) _49304_ ( .A(_29211_), .B(8'h00), .S(RST), .Y(_01532_) );
  \$mux  #( .WIDTH(8) ) _49305_ ( .A(_29210_), .B(8'h00), .S(RST), .Y(_01529_) );
  \$mux  #( .WIDTH(8) ) _49306_ ( .A(_29209_), .B(8'h00), .S(RST), .Y(_01526_) );
  \$mux  #( .WIDTH(8) ) _49307_ ( .A(_29208_), .B(8'h00), .S(RST), .Y(_01523_) );
  \$mux  #( .WIDTH(8) ) _49308_ ( .A(_29207_), .B(8'h00), .S(RST), .Y(_01520_) );
  \$mux  #( .WIDTH(8) ) _49309_ ( .A(_29206_), .B(8'h00), .S(RST), .Y(_01517_) );
  \$mux  #( .WIDTH(8) ) _49310_ ( .A(_29205_), .B(8'h00), .S(RST), .Y(_01514_) );
  \$mux  #( .WIDTH(8) ) _49311_ ( .A(_29204_), .B(8'h00), .S(RST), .Y(_01511_) );
  \$mux  #( .WIDTH(8) ) _49312_ ( .A(_29203_), .B(8'h00), .S(RST), .Y(_01508_) );
  \$mux  #( .WIDTH(8) ) _49313_ ( .A(__delay_data_1370), .B(8'h00), .S(RST), .Y(_00252_) );
  \$mux  #( .WIDTH(8) ) _49314_ ( .A(__delay_data_1342), .B(8'h00), .S(RST), .Y(_00224_) );
  \$mux  #( .WIDTH(8) ) _49315_ ( .A(__delay_data_1313), .B(8'h00), .S(RST), .Y(_00195_) );
  \$mux  #( .WIDTH(6) ) _49316_ ( .A(__delay_data_1292), .B(6'h00), .S(RST), .Y(_00174_) );
  \$mux  #( .WIDTH(8) ) _49317_ ( .A(__delay_data_1270), .B(8'h00), .S(RST), .Y(_00152_) );
  \$mux  #( .WIDTH(4) ) _49318_ ( .A(__delay_data_1257), .B(4'h0), .S(RST), .Y(_00145_) );
  \$mux  #( .WIDTH(1) ) _49319_ ( .A(__delay_data_1250), .B(1'h0), .S(RST), .Y(_00138_) );
  \$mux  #( .WIDTH(4) ) _49320_ ( .A(__delay_data_1223), .B(4'h0), .S(RST), .Y(_00129_) );
  \$mux  #( .WIDTH(1) ) _49321_ ( .A(__delay_data_1216), .B(1'h0), .S(RST), .Y(_00122_) );
  \$mux  #( .WIDTH(4) ) _49322_ ( .A(__delay_data_1189), .B(4'h0), .S(RST), .Y(_00113_) );
  \$mux  #( .WIDTH(1) ) _49323_ ( .A(__delay_data_1182), .B(1'h0), .S(RST), .Y(_00106_) );
  \$mux  #( .WIDTH(4) ) _49324_ ( .A(__delay_data_1155), .B(4'h0), .S(RST), .Y(_00097_) );
  \$mux  #( .WIDTH(1) ) _49325_ ( .A(__delay_data_1148), .B(1'h0), .S(RST), .Y(_00090_) );
  \$mux  #( .WIDTH(8) ) _49326_ ( .A(_cond_data_366), .B(8'h00), .S(RST), .Y(_00084_) );
  \$mux  #( .WIDTH(4) ) _49327_ ( .A(__delay_data_1120), .B(4'h0), .S(RST), .Y(_00080_) );
  \$mux  #( .WIDTH(1) ) _49328_ ( .A(__delay_data_1113), .B(1'h0), .S(RST), .Y(_00073_) );
  \$mux  #( .WIDTH(8) ) _49329_ ( .A(_cond_data_356), .B(8'h00), .S(RST), .Y(_00067_) );
  \$mux  #( .WIDTH(4) ) _49330_ ( .A(__delay_data_1085), .B(4'h0), .S(RST), .Y(_00063_) );
  \$mux  #( .WIDTH(1) ) _49331_ ( .A(__delay_data_1078), .B(1'h0), .S(RST), .Y(_00056_) );
  \$mux  #( .WIDTH(8) ) _49332_ ( .A(_cond_data_346), .B(8'h00), .S(RST), .Y(_00050_) );
  \$mux  #( .WIDTH(4) ) _49333_ ( .A(__delay_data_1050), .B(4'h0), .S(RST), .Y(_00046_) );
  \$mux  #( .WIDTH(1) ) _49334_ ( .A(__delay_data_1043), .B(1'h0), .S(RST), .Y(_00039_) );
  \$mux  #( .WIDTH(8) ) _49335_ ( .A(_cond_data_306), .B(8'h00), .S(RST), .Y(_00033_) );
  \$mux  #( .WIDTH(8) ) _49336_ ( .A(_cond_data_336), .B(8'h00), .S(RST), .Y(_00027_) );
  \$mux  #( .WIDTH(4) ) _49337_ ( .A(__delay_data_1002), .B(4'h0), .S(RST), .Y(_00004_) );
  \$mux  #( .WIDTH(1) ) _49338_ ( .A(__delay_data_995), .B(1'h0), .S(RST), .Y(_00677_) );
  \$mux  #( .WIDTH(8) ) _49339_ ( .A(_cond_data_296), .B(8'h00), .S(RST), .Y(_00671_) );
  \$mux  #( .WIDTH(8) ) _49340_ ( .A(_cond_data_326), .B(8'h00), .S(RST), .Y(_00670_) );
  \$mux  #( .WIDTH(8) ) _49341_ ( .A(__delay_data_1263), .B(8'h00), .S(RST), .Y(_00010_) );
  \$mux  #( .WIDTH(4) ) _49342_ ( .A(__delay_data_951), .B(4'h0), .S(RST), .Y(_00660_) );
  \$mux  #( .WIDTH(1) ) _49343_ ( .A(__delay_data_943), .B(1'h0), .S(RST), .Y(_00652_) );
  \$mux  #( .WIDTH(8) ) _49344_ ( .A(_cond_data_286), .B(8'h00), .S(RST), .Y(_00646_) );
  \$mux  #( .WIDTH(1) ) _49345_ ( .A(__delay_data_1243), .B(1'h0), .S(RST), .Y(_00031_) );
  \$mux  #( .WIDTH(8) ) _49346_ ( .A(_cond_data_316), .B(8'h00), .S(RST), .Y(_00645_) );
  \$mux  #( .WIDTH(1) ) _49347_ ( .A(__delay_data_1239), .B(1'h0), .S(RST), .Y(_00026_) );
  \$mux  #( .WIDTH(8) ) _49348_ ( .A(_29202_), .B(8'h00), .S(RST), .Y(_01531_) );
  \$mux  #( .WIDTH(8) ) _49349_ ( .A(_29201_), .B(8'h00), .S(RST), .Y(_01528_) );
  \$mux  #( .WIDTH(8) ) _49350_ ( .A(_29200_), .B(8'h00), .S(RST), .Y(_01525_) );
  \$mux  #( .WIDTH(8) ) _49351_ ( .A(_29199_), .B(8'h00), .S(RST), .Y(_01522_) );
  \$mux  #( .WIDTH(8) ) _49352_ ( .A(_29198_), .B(8'h00), .S(RST), .Y(_01519_) );
  \$mux  #( .WIDTH(8) ) _49353_ ( .A(_29197_), .B(8'h00), .S(RST), .Y(_01516_) );
  \$mux  #( .WIDTH(8) ) _49354_ ( .A(_29196_), .B(8'h00), .S(RST), .Y(_01513_) );
  \$mux  #( .WIDTH(8) ) _49355_ ( .A(_29195_), .B(8'h00), .S(RST), .Y(_01510_) );
  \$mux  #( .WIDTH(8) ) _49356_ ( .A(_29194_), .B(8'h00), .S(RST), .Y(_01507_) );
  \$mux  #( .WIDTH(8) ) _49357_ ( .A(__delay_data_1369), .B(8'h00), .S(RST), .Y(_00251_) );
  \$mux  #( .WIDTH(8) ) _49358_ ( .A(__delay_data_1341), .B(8'h00), .S(RST), .Y(_00223_) );
  \$mux  #( .WIDTH(8) ) _49359_ ( .A(__delay_data_1312), .B(8'h00), .S(RST), .Y(_00194_) );
  \$mux  #( .WIDTH(6) ) _49360_ ( .A(__delay_data_1291), .B(6'h00), .S(RST), .Y(_00173_) );
  \$mux  #( .WIDTH(8) ) _49361_ ( .A(__delay_data_1269), .B(8'h00), .S(RST), .Y(_00151_) );
  \$mux  #( .WIDTH(4) ) _49362_ ( .A(__delay_data_1256), .B(4'h0), .S(RST), .Y(_00144_) );
  \$mux  #( .WIDTH(1) ) _49363_ ( .A(__delay_data_1249), .B(1'h0), .S(RST), .Y(_00137_) );
  \$mux  #( .WIDTH(4) ) _49364_ ( .A(__delay_data_1222), .B(4'h0), .S(RST), .Y(_00128_) );
  \$mux  #( .WIDTH(1) ) _49365_ ( .A(__delay_data_1215), .B(1'h0), .S(RST), .Y(_00121_) );
  \$mux  #( .WIDTH(4) ) _49366_ ( .A(__delay_data_1188), .B(4'h0), .S(RST), .Y(_00112_) );
  \$mux  #( .WIDTH(1) ) _49367_ ( .A(__delay_data_1181), .B(1'h0), .S(RST), .Y(_00105_) );
  \$mux  #( .WIDTH(4) ) _49368_ ( .A(__delay_data_1154), .B(4'h0), .S(RST), .Y(_00096_) );
  \$mux  #( .WIDTH(1) ) _49369_ ( .A(__delay_data_1147), .B(1'h0), .S(RST), .Y(_00089_) );
  \$mux  #( .WIDTH(4) ) _49370_ ( .A(__delay_data_1119), .B(4'h0), .S(RST), .Y(_00079_) );
  \$mux  #( .WIDTH(1) ) _49371_ ( .A(__delay_data_1112), .B(1'h0), .S(RST), .Y(_00072_) );
  \$mux  #( .WIDTH(4) ) _49372_ ( .A(__delay_data_1084), .B(4'h0), .S(RST), .Y(_00062_) );
  \$mux  #( .WIDTH(1) ) _49373_ ( .A(__delay_data_1077), .B(1'h0), .S(RST), .Y(_00055_) );
  \$mux  #( .WIDTH(4) ) _49374_ ( .A(__delay_data_1049), .B(4'h0), .S(RST), .Y(_00045_) );
  \$mux  #( .WIDTH(1) ) _49375_ ( .A(__delay_data_1042), .B(1'h0), .S(RST), .Y(_00038_) );
  \$mux  #( .WIDTH(4) ) _49376_ ( .A(__delay_data_1001), .B(4'h0), .S(RST), .Y(_00003_) );
  \$mux  #( .WIDTH(1) ) _49377_ ( .A(__delay_data_994), .B(1'h0), .S(RST), .Y(_00676_) );
  \$mux  #( .WIDTH(8) ) _49378_ ( .A(__delay_data_1262), .B(8'h00), .S(RST), .Y(_00009_) );
  \$mux  #( .WIDTH(4) ) _49379_ ( .A(__delay_data_950), .B(4'h0), .S(RST), .Y(_00659_) );
  \$mux  #( .WIDTH(1) ) _49380_ ( .A(__delay_data_942), .B(1'h0), .S(RST), .Y(_00651_) );
  \$mux  #( .WIDTH(1) ) _49381_ ( .A(__delay_data_1242), .B(1'h0), .S(RST), .Y(_00030_) );
  \$mux  #( .WIDTH(1) ) _49382_ ( .A(__delay_data_1238), .B(1'h0), .S(RST), .Y(_00025_) );
  \$mux  #( .WIDTH(1) ) _49383_ ( .A(__delay_data_1235), .B(1'h0), .S(RST), .Y(_00022_) );
  \$mux  #( .WIDTH(8) ) _49384_ ( .A(_29193_), .B(8'h00), .S(RST), .Y(_01506_) );
  \$mux  #( .WIDTH(8) ) _49385_ ( .A(_29192_), .B(8'h00), .S(RST), .Y(_01503_) );
  \$mux  #( .WIDTH(8) ) _49386_ ( .A(_29191_), .B(8'h00), .S(RST), .Y(_01500_) );
  \$mux  #( .WIDTH(8) ) _49387_ ( .A(_29190_), .B(8'h00), .S(RST), .Y(_01497_) );
  \$mux  #( .WIDTH(8) ) _49388_ ( .A(_29189_), .B(8'h00), .S(RST), .Y(_01494_) );
  \$mux  #( .WIDTH(8) ) _49389_ ( .A(_29188_), .B(8'h00), .S(RST), .Y(_01491_) );
  \$mux  #( .WIDTH(8) ) _49390_ ( .A(_29187_), .B(8'h00), .S(RST), .Y(_01488_) );
  \$mux  #( .WIDTH(8) ) _49391_ ( .A(_29186_), .B(8'h00), .S(RST), .Y(_01485_) );
  \$mux  #( .WIDTH(8) ) _49392_ ( .A(_29185_), .B(8'h00), .S(RST), .Y(_01482_) );
  \$mux  #( .WIDTH(8) ) _49393_ ( .A(_plus_data_770), .B(8'h00), .S(RST), .Y(_00250_) );
  \$mux  #( .WIDTH(8) ) _49394_ ( .A(__delay_data_1340), .B(8'h00), .S(RST), .Y(_00222_) );
  \$mux  #( .WIDTH(8) ) _49395_ ( .A(__delay_data_1311), .B(8'h00), .S(RST), .Y(_00193_) );
  \$mux  #( .WIDTH(6) ) _49396_ ( .A(__delay_data_1290), .B(6'h00), .S(RST), .Y(_00172_) );
  \$mux  #( .WIDTH(8) ) _49397_ ( .A(_plus_data_759), .B(8'h00), .S(RST), .Y(_00150_) );
  \$mux  #( .WIDTH(4) ) _49398_ ( .A(__delay_data_1255), .B(4'h0), .S(RST), .Y(_00143_) );
  \$mux  #( .WIDTH(1) ) _49399_ ( .A(__delay_data_1248), .B(1'h0), .S(RST), .Y(_00136_) );
  \$mux  #( .WIDTH(4) ) _49400_ ( .A(__delay_data_1221), .B(4'h0), .S(RST), .Y(_00127_) );
  \$mux  #( .WIDTH(1) ) _49401_ ( .A(__delay_data_1214), .B(1'h0), .S(RST), .Y(_00120_) );
  \$mux  #( .WIDTH(4) ) _49402_ ( .A(__delay_data_1187), .B(4'h0), .S(RST), .Y(_00111_) );
  \$mux  #( .WIDTH(1) ) _49403_ ( .A(__delay_data_1180), .B(1'h0), .S(RST), .Y(_00104_) );
  \$mux  #( .WIDTH(4) ) _49404_ ( .A(__delay_data_1153), .B(4'h0), .S(RST), .Y(_00095_) );
  \$mux  #( .WIDTH(1) ) _49405_ ( .A(__delay_data_1146), .B(1'h0), .S(RST), .Y(_00088_) );
  \$mux  #( .WIDTH(4) ) _49406_ ( .A(__delay_data_1118), .B(4'h0), .S(RST), .Y(_00078_) );
  \$mux  #( .WIDTH(1) ) _49407_ ( .A(__delay_data_1111), .B(1'h0), .S(RST), .Y(_00071_) );
  \$mux  #( .WIDTH(4) ) _49408_ ( .A(__delay_data_1083), .B(4'h0), .S(RST), .Y(_00061_) );
  \$mux  #( .WIDTH(1) ) _49409_ ( .A(__delay_data_1076), .B(1'h0), .S(RST), .Y(_00054_) );
  \$mux  #( .WIDTH(4) ) _49410_ ( .A(__delay_data_1048), .B(4'h0), .S(RST), .Y(_00044_) );
  \$mux  #( .WIDTH(1) ) _49411_ ( .A(__delay_data_1041), .B(1'h0), .S(RST), .Y(_00037_) );
  \$mux  #( .WIDTH(8) ) _49412_ ( .A(__delay_data_973), .B(8'h00), .S(RST), .Y(_00019_) );
  \$mux  #( .WIDTH(8) ) _49413_ ( .A(__delay_data_968), .B(8'h00), .S(RST), .Y(_00018_) );
  \$mux  #( .WIDTH(8) ) _49414_ ( .A(__delay_data_963), .B(8'h00), .S(RST), .Y(_00017_) );
  \$mux  #( .WIDTH(4) ) _49415_ ( .A(__delay_data_1000), .B(4'h0), .S(RST), .Y(_00002_) );
  \$mux  #( .WIDTH(1) ) _49416_ ( .A(__delay_data_993), .B(1'h0), .S(RST), .Y(_00675_) );
  \$mux  #( .WIDTH(8) ) _49417_ ( .A(__delay_data_919), .B(8'h00), .S(RST), .Y(_00669_) );
  \$mux  #( .WIDTH(8) ) _49418_ ( .A(__delay_data_910), .B(8'h00), .S(RST), .Y(_00667_) );
  \$mux  #( .WIDTH(8) ) _49419_ ( .A(__delay_data_901), .B(8'h00), .S(RST), .Y(_00665_) );
  \$mux  #( .WIDTH(8) ) _49420_ ( .A(_plus_data_743), .B(8'h00), .S(RST), .Y(_00008_) );
  \$mux  #( .WIDTH(4) ) _49421_ ( .A(__delay_data_949), .B(4'h0), .S(RST), .Y(_00658_) );
  \$mux  #( .WIDTH(1) ) _49422_ ( .A(__delay_data_941), .B(1'h0), .S(RST), .Y(_00650_) );
  \$mux  #( .WIDTH(1) ) _49423_ ( .A(__delay_data_1241), .B(1'h0), .S(RST), .Y(_00029_) );
  \$mux  #( .WIDTH(1) ) _49424_ ( .A(__delay_data_1237), .B(1'h0), .S(RST), .Y(_00024_) );
  \$mux  #( .WIDTH(1) ) _49425_ ( .A(__delay_data_1234), .B(1'h0), .S(RST), .Y(_00021_) );
  \$mux  #( .WIDTH(8) ) _49426_ ( .A(__delay_data_923), .B(8'h00), .S(RST), .Y(_00644_) );
  \$mux  #( .WIDTH(8) ) _49427_ ( .A(__delay_data_914), .B(8'h00), .S(RST), .Y(_00638_) );
  \$mux  #( .WIDTH(8) ) _49428_ ( .A(__delay_data_905), .B(8'h00), .S(RST), .Y(_00632_) );
  \$mux  #( .WIDTH(1) ) _49429_ ( .A(__delay_data_1022), .B(1'h0), .S(RST), .Y(_00016_) );
  \$mux  #( .WIDTH(8) ) _49430_ ( .A(_29184_), .B(8'h00), .S(RST), .Y(_01505_) );
  \$mux  #( .WIDTH(8) ) _49431_ ( .A(_29183_), .B(8'h00), .S(RST), .Y(_01502_) );
  \$mux  #( .WIDTH(8) ) _49432_ ( .A(_29182_), .B(8'h00), .S(RST), .Y(_01499_) );
  \$mux  #( .WIDTH(8) ) _49433_ ( .A(_29181_), .B(8'h00), .S(RST), .Y(_01496_) );
  \$mux  #( .WIDTH(8) ) _49434_ ( .A(_29180_), .B(8'h00), .S(RST), .Y(_01493_) );
  \$mux  #( .WIDTH(8) ) _49435_ ( .A(_29179_), .B(8'h00), .S(RST), .Y(_01490_) );
  \$mux  #( .WIDTH(8) ) _49436_ ( .A(_29178_), .B(8'h00), .S(RST), .Y(_01487_) );
  \$mux  #( .WIDTH(8) ) _49437_ ( .A(_29177_), .B(8'h00), .S(RST), .Y(_01484_) );
  \$mux  #( .WIDTH(8) ) _49438_ ( .A(_29176_), .B(8'h00), .S(RST), .Y(_01481_) );
  \$mux  #( .WIDTH(8) ) _49439_ ( .A(_cond_data_242), .B(8'h00), .S(RST), .Y(_00221_) );
  \$mux  #( .WIDTH(8) ) _49440_ ( .A(_cond_data_235), .B(8'h00), .S(RST), .Y(_00192_) );
  \$mux  #( .WIDTH(6) ) _49441_ ( .A(__delay_data_1289), .B(6'h00), .S(RST), .Y(_00171_) );
  \$mux  #( .WIDTH(4) ) _49442_ ( .A(__delay_data_1254), .B(4'h0), .S(RST), .Y(_00142_) );
  \$mux  #( .WIDTH(1) ) _49443_ ( .A(__delay_data_1247), .B(1'h0), .S(RST), .Y(_00135_) );
  \$mux  #( .WIDTH(4) ) _49444_ ( .A(__delay_data_1220), .B(4'h0), .S(RST), .Y(_00126_) );
  \$mux  #( .WIDTH(1) ) _49445_ ( .A(__delay_data_1213), .B(1'h0), .S(RST), .Y(_00119_) );
  \$mux  #( .WIDTH(4) ) _49446_ ( .A(__delay_data_1186), .B(4'h0), .S(RST), .Y(_00110_) );
  \$mux  #( .WIDTH(1) ) _49447_ ( .A(__delay_data_1179), .B(1'h0), .S(RST), .Y(_00103_) );
  \$mux  #( .WIDTH(4) ) _49448_ ( .A(__delay_data_1152), .B(4'h0), .S(RST), .Y(_00094_) );
  \$mux  #( .WIDTH(1) ) _49449_ ( .A(__delay_data_1145), .B(1'h0), .S(RST), .Y(_00087_) );
  \$mux  #( .WIDTH(4) ) _49450_ ( .A(__delay_data_1117), .B(4'h0), .S(RST), .Y(_00077_) );
  \$mux  #( .WIDTH(1) ) _49451_ ( .A(__delay_data_1110), .B(1'h0), .S(RST), .Y(_00070_) );
  \$mux  #( .WIDTH(4) ) _49452_ ( .A(__delay_data_1082), .B(4'h0), .S(RST), .Y(_00060_) );
  \$mux  #( .WIDTH(1) ) _49453_ ( .A(__delay_data_1075), .B(1'h0), .S(RST), .Y(_00053_) );
  \$mux  #( .WIDTH(4) ) _49454_ ( .A(__delay_data_1047), .B(4'h0), .S(RST), .Y(_00043_) );
  \$mux  #( .WIDTH(1) ) _49455_ ( .A(__delay_data_1040), .B(1'h0), .S(RST), .Y(_00036_) );
  \$mux  #( .WIDTH(4) ) _49456_ ( .A(__delay_data_999), .B(4'h0), .S(RST), .Y(_00001_) );
  \$mux  #( .WIDTH(1) ) _49457_ ( .A(__delay_data_992), .B(1'h0), .S(RST), .Y(_00674_) );
  \$mux  #( .WIDTH(8) ) _49458_ ( .A(__delay_data_916), .B(8'h00), .S(RST), .Y(_00668_) );
  \$mux  #( .WIDTH(8) ) _49459_ ( .A(__delay_data_907), .B(8'h00), .S(RST), .Y(_00666_) );
  \$mux  #( .WIDTH(8) ) _49460_ ( .A(__delay_data_898), .B(8'h00), .S(RST), .Y(_00664_) );
  \$mux  #( .WIDTH(4) ) _49461_ ( .A(__delay_data_948), .B(4'h0), .S(RST), .Y(_00657_) );
  \$mux  #( .WIDTH(1) ) _49462_ ( .A(__delay_data_940), .B(1'h0), .S(RST), .Y(_00649_) );
  \$mux  #( .WIDTH(1) ) _49463_ ( .A(_eq_data_454), .B(1'h0), .S(RST), .Y(_00028_) );
  \$mux  #( .WIDTH(1) ) _49464_ ( .A(_eq_data_451), .B(1'h0), .S(RST), .Y(_00023_) );
  \$mux  #( .WIDTH(1) ) _49465_ ( .A(_eq_data_447), .B(1'h0), .S(RST), .Y(_00020_) );
  \$mux  #( .WIDTH(8) ) _49466_ ( .A(__delay_data_922), .B(8'h00), .S(RST), .Y(_00643_) );
  \$mux  #( .WIDTH(8) ) _49467_ ( .A(__delay_data_918), .B(8'h00), .S(RST), .Y(_00641_) );
  \$mux  #( .WIDTH(8) ) _49468_ ( .A(__delay_data_913), .B(8'h00), .S(RST), .Y(_00637_) );
  \$mux  #( .WIDTH(8) ) _49469_ ( .A(__delay_data_909), .B(8'h00), .S(RST), .Y(_00635_) );
  \$mux  #( .WIDTH(8) ) _49470_ ( .A(__delay_data_904), .B(8'h00), .S(RST), .Y(_00631_) );
  \$mux  #( .WIDTH(1) ) _49471_ ( .A(_eq_data_364), .B(1'h0), .S(RST), .Y(_00015_) );
  \$mux  #( .WIDTH(8) ) _49472_ ( .A(__delay_data_900), .B(8'h00), .S(RST), .Y(_00629_) );
  \$mux  #( .WIDTH(1) ) _49473_ ( .A(_eq_data_361), .B(1'h0), .S(RST), .Y(_00014_) );
  \$mux  #( .WIDTH(8) ) _49474_ ( .A(_24306_), .B(8'h00), .S(RST), .Y(_01814_) );
  \$mux  #( .WIDTH(8) ) _49475_ ( .A(_24305_), .B(8'h00), .S(RST), .Y(_01812_) );
  \$mux  #( .WIDTH(8) ) _49476_ ( .A(_24304_), .B(8'h00), .S(RST), .Y(_01811_) );
  \$mux  #( .WIDTH(8) ) _49477_ ( .A(_29175_), .B(8'h00), .S(RST), .Y(_01504_) );
  \$mux  #( .WIDTH(8) ) _49478_ ( .A(_29174_), .B(8'h00), .S(RST), .Y(_01501_) );
  \$mux  #( .WIDTH(8) ) _49479_ ( .A(_29173_), .B(8'h00), .S(RST), .Y(_01498_) );
  \$mux  #( .WIDTH(8) ) _49480_ ( .A(_29172_), .B(8'h00), .S(RST), .Y(_01495_) );
  \$mux  #( .WIDTH(8) ) _49481_ ( .A(_29171_), .B(8'h00), .S(RST), .Y(_01492_) );
  \$mux  #( .WIDTH(8) ) _49482_ ( .A(_29170_), .B(8'h00), .S(RST), .Y(_01489_) );
  \$mux  #( .WIDTH(8) ) _49483_ ( .A(_29169_), .B(8'h00), .S(RST), .Y(_01486_) );
  \$mux  #( .WIDTH(8) ) _49484_ ( .A(_29168_), .B(8'h00), .S(RST), .Y(_01483_) );
  \$mux  #( .WIDTH(8) ) _49485_ ( .A(_29167_), .B(8'h00), .S(RST), .Y(_01480_) );
  \$mux  #( .WIDTH(4) ) _49486_ ( .A(__variable_wdata_266), .B(4'h0), .S(RST), .Y(_00220_) );
  \$mux  #( .WIDTH(6) ) _49487_ ( .A(__variable_wdata_214), .B(6'h00), .S(RST), .Y(_00170_) );
  \$mux  #( .WIDTH(1) ) _49488_ ( .A(__variable_wdata_265), .B(1'h0), .S(RST), .Y(_00149_) );
  \$mux  #( .WIDTH(4) ) _49489_ ( .A(__variable_wdata_510), .B(4'h0), .S(RST), .Y(_00141_) );
  \$mux  #( .WIDTH(1) ) _49490_ ( .A(__variable_wdata_217[8]), .B(1'h0), .S(RST), .Y(_00134_) );
  \$mux  #( .WIDTH(4) ) _49491_ ( .A(__variable_wdata_509), .B(4'h0), .S(RST), .Y(_00125_) );
  \$mux  #( .WIDTH(1) ) _49492_ ( .A(__variable_wdata_217[7]), .B(1'h0), .S(RST), .Y(_00118_) );
  \$mux  #( .WIDTH(4) ) _49493_ ( .A(__variable_wdata_508), .B(4'h0), .S(RST), .Y(_00109_) );
  \$mux  #( .WIDTH(1) ) _49494_ ( .A(__variable_wdata_217[6]), .B(1'h0), .S(RST), .Y(_00102_) );
  \$mux  #( .WIDTH(4) ) _49495_ ( .A(__variable_wdata_507), .B(4'h0), .S(RST), .Y(_00093_) );
  \$mux  #( .WIDTH(1) ) _49496_ ( .A(__variable_wdata_217[5]), .B(1'h0), .S(RST), .Y(_00086_) );
  \$mux  #( .WIDTH(4) ) _49497_ ( .A(__variable_wdata_506), .B(4'h0), .S(RST), .Y(_00076_) );
  \$mux  #( .WIDTH(1) ) _49498_ ( .A(__variable_wdata_217[4]), .B(1'h0), .S(RST), .Y(_00069_) );
  \$mux  #( .WIDTH(4) ) _49499_ ( .A(__variable_wdata_505), .B(4'h0), .S(RST), .Y(_00059_) );
  \$mux  #( .WIDTH(1) ) _49500_ ( .A(__variable_wdata_217[3]), .B(1'h0), .S(RST), .Y(_00052_) );
  \$mux  #( .WIDTH(4) ) _49501_ ( .A(__variable_wdata_504), .B(4'h0), .S(RST), .Y(_00042_) );
  \$mux  #( .WIDTH(1) ) _49502_ ( .A(__variable_wdata_217[2]), .B(1'h0), .S(RST), .Y(_00035_) );
  \$mux  #( .WIDTH(4) ) _49503_ ( .A(__variable_wdata_503), .B(4'h0), .S(RST), .Y(_00680_) );
  \$mux  #( .WIDTH(1) ) _49504_ ( .A(__variable_wdata_217[1]), .B(1'h0), .S(RST), .Y(_00673_) );
  \$mux  #( .WIDTH(4) ) _49505_ ( .A(__variable_wdata_502), .B(4'h0), .S(RST), .Y(_00656_) );
  \$mux  #( .WIDTH(1) ) _49506_ ( .A(__variable_wdata_264), .B(1'h0), .S(RST), .Y(_00655_) );
  \$mux  #( .WIDTH(1) ) _49507_ ( .A(__variable_wdata_217[0]), .B(1'h0), .S(RST), .Y(_00648_) );
  \$mux  #( .WIDTH(8) ) _49508_ ( .A(__variable_wdata_274), .B(8'h00), .S(RST), .Y(_00642_) );
  \$mux  #( .WIDTH(8) ) _49509_ ( .A(__variable_wdata_275), .B(8'h00), .S(RST), .Y(_00640_) );
  \$mux  #( .WIDTH(8) ) _49510_ ( .A(__variable_wdata_276), .B(8'h00), .S(RST), .Y(_00639_) );
  \$mux  #( .WIDTH(8) ) _49511_ ( .A(__variable_wdata_271), .B(8'h00), .S(RST), .Y(_00636_) );
  \$mux  #( .WIDTH(8) ) _49512_ ( .A(__variable_wdata_272), .B(8'h00), .S(RST), .Y(_00634_) );
  \$mux  #( .WIDTH(8) ) _49513_ ( .A(__variable_wdata_273), .B(8'h00), .S(RST), .Y(_00633_) );
  \$mux  #( .WIDTH(8) ) _49514_ ( .A(__variable_wdata_268), .B(8'h00), .S(RST), .Y(_00630_) );
  \$mux  #( .WIDTH(8) ) _49515_ ( .A(__variable_wdata_269), .B(8'h00), .S(RST), .Y(_00628_) );
  \$mux  #( .WIDTH(8) ) _49516_ ( .A(__variable_wdata_270), .B(8'h00), .S(RST), .Y(_00627_) );
  \$mux  #( .WIDTH(1) ) _49517_ ( .A(_06141_), .B(1'h0), .S(RST), .Y(_01685_) );
  \$mux  #( .WIDTH(1) ) _49518_ ( .A(_06140_), .B(1'h0), .S(RST), .Y(_01684_) );
  \$mux  #( .WIDTH(1) ) _49519_ ( .A(_06139_), .B(1'h0), .S(RST), .Y(_01683_) );
  \$mux  #( .WIDTH(1) ) _49520_ ( .A(_06138_), .B(1'h0), .S(RST), .Y(_01682_) );
  \$mux  #( .WIDTH(1) ) _49521_ ( .A(_06137_), .B(1'h0), .S(RST), .Y(_01681_) );
  \$mux  #( .WIDTH(1) ) _49522_ ( .A(_06136_), .B(1'h0), .S(RST), .Y(_01680_) );
  \$mux  #( .WIDTH(8) ) _49523_ ( .A(__variable_wdata_258), .B(8'h00), .S(RST), .Y(_01479_) );
  \$mux  #( .WIDTH(8) ) _49524_ ( .A(__variable_wdata_251), .B(8'h00), .S(RST), .Y(_01478_) );
  \$mux  #( .WIDTH(8) ) _49525_ ( .A(__variable_wdata_244), .B(8'h00), .S(RST), .Y(_01477_) );
  \$mux  #( .WIDTH(8) ) _49526_ ( .A(__variable_wdata_237), .B(8'h00), .S(RST), .Y(_01476_) );
  \$mux  #( .WIDTH(8) ) _49527_ ( .A(__variable_wdata_230), .B(8'h00), .S(RST), .Y(_01475_) );
  \$mux  #( .WIDTH(8) ) _49528_ ( .A(_stream_conv2d_16_sink_37_sink_wdata), .B(_cond_data_890), .S(_06787_), .Y(_26239_) );
  \$mux  #( .WIDTH(8) ) _49529_ ( .A(_26239_), .B(8'h00), .S(RST), .Y(_02513_) );
  \$mux  #( .WIDTH(1) ) _49530_ ( .A(1'h0), .B(1'h1), .S(_06787_), .Y(_26240_) );
  \$mux  #( .WIDTH(1) ) _49531_ ( .A(_26240_), .B(1'h0), .S(RST), .Y(_02514_) );
  \$mux  #( .WIDTH(32) ) _49532_ ( .A(_stream_conv2d_16_sink_37_sink_waddr), .B(_28868_), .S(_06786_), .Y(_26241_) );
  \$mux  #( .WIDTH(32) ) _49533_ ( .A(_26241_), .B(_24398_), .S(_06787_), .Y(_26242_) );
  \$mux  #( .WIDTH(32) ) _49534_ ( .A(_26242_), .B(0), .S(RST), .Y(_02512_) );
  \$mux  #( .WIDTH(8) ) _49535_ ( .A(_stream_conv2d_16_sink_37_sink_ram_sel), .B(8'h15), .S(__set_flag_710_45), .Y(_26243_) );
  \$mux  #( .WIDTH(8) ) _49536_ ( .A(_26243_), .B(8'h00), .S(RST), .Y(_02508_) );
  \$mux  #( .WIDTH(32) ) _49537_ ( .A(_stream_conv2d_16_sink_37_sink_stride_buf), .B(_stream_conv2d_16_sink_37_sink_stride), .S(_06786_), .Y(_26244_) );
  \$mux  #( .WIDTH(32) ) _49538_ ( .A(_26244_), .B(0), .S(RST), .Y(_02511_) );
  \$mux  #( .WIDTH(33) ) _49539_ ( .A(_stream_conv2d_16_sink_37_sink_count), .B(_stream_conv2d_16_sink_37_sink_size), .S(_06786_), .Y(_26245_) );
  \$mux  #( .WIDTH(33) ) _49540_ ( .A(_26245_), .B(_28869_), .S(_06787_), .Y(_26246_) );
  \$mux  #( .WIDTH(33) ) _49541_ ( .A(_26246_), .B(33'h000000000), .S(RST), .Y(_02504_) );
  \$mux  #( .WIDTH(32) ) _49542_ ( .A(_stream_conv2d_16_sink_37_sink_stride), .B(1), .S(__set_flag_710_45), .Y(_26247_) );
  \$mux  #( .WIDTH(32) ) _49543_ ( .A(_26247_), .B(0), .S(RST), .Y(_02510_) );
  \$mux  #( .WIDTH(33) ) _49544_ ( .A(_stream_conv2d_16_sink_37_sink_size), .B(__stream_conv2d_16_sink_37_sink_size_1_45), .S(__set_flag_710_45), .Y(_26248_) );
  \$mux  #( .WIDTH(33) ) _49545_ ( .A(_26248_), .B(33'h000000000), .S(RST), .Y(_02509_) );
  \$mux  #( .WIDTH(32) ) _49546_ ( .A(_stream_conv2d_16_sink_37_sink_offset), .B(__stream_conv2d_16_sink_37_sink_offset_0_45), .S(__set_flag_710_45), .Y(_26249_) );
  \$mux  #( .WIDTH(32) ) _49547_ ( .A(_26249_), .B(0), .S(RST), .Y(_02507_) );
  \$mux  #( .WIDTH(3) ) _49548_ ( .A(_stream_conv2d_16_sink_37_sink_mode), .B(3'h1), .S(__set_flag_710_45), .Y(_26250_) );
  \$mux  #( .WIDTH(3) ) _49549_ ( .A(_26250_), .B(3'h0), .S(RST), .Y(_02506_) );
  \$mux  #( .WIDTH(1) ) _49550_ ( .A(1'h0), .B(1'h1), .S(_ram_w4_l8192_id8_0_cond_1_1), .Y(_26251_) );
  \$mux  #( .WIDTH(1) ) _49551_ ( .A(_26251_), .B(1'h0), .S(RST), .Y(_02681_) );
  \$mux  #( .WIDTH(1) ) _49552_ ( .A(1'h1), .B(_stream_conv2d_16_source_36_source_ram_renable), .S(_05949_), .Y(_26252_) );
  \$mux  #( .WIDTH(1) ) _49553_ ( .A(1'h0), .B(_26252_), .S(_05950_), .Y(_26253_) );
  \$mux  #( .WIDTH(1) ) _49554_ ( .A(_26253_), .B(1'h0), .S(RST), .Y(_02680_) );
  \$mux  #( .WIDTH(32) ) _49555_ ( .A(_stream_conv2d_16_source_36_source_pat_all_offset), .B(_stream_conv2d_16_source_36_source_ram_raddr), .S(_05949_), .Y(_26254_) );
  \$mux  #( .WIDTH(32) ) _49556_ ( .A(_26254_), .B(0), .S(RST), .Y(_02679_) );
  \$mux  #( .WIDTH(8) ) _49557_ ( .A(_stream_conv2d_16_source_36_source_ram_sel), .B(8'h14), .S(_set_flag_710), .Y(_26255_) );
  \$mux  #( .WIDTH(8) ) _49558_ ( .A(_26255_), .B(8'h00), .S(RST), .Y(_02682_) );
  \$mux  #( .WIDTH(32) ) _49559_ ( .A(_stream_conv2d_16_source_36_source_offset_buf), .B(_stream_conv2d_16_source_36_source_offset), .S(_06781_), .Y(_26256_) );
  \$mux  #( .WIDTH(32) ) _49560_ ( .A(_26256_), .B(0), .S(RST), .Y(_02677_) );
  \$mux  #( .WIDTH(32) ) _49561_ ( .A(_stream_conv2d_16_source_36_source_offset), .B(conv2d_16_filter_page_comp_offset_buf), .S(_set_flag_710), .Y(_26257_) );
  \$mux  #( .WIDTH(32) ) _49562_ ( .A(_26257_), .B(0), .S(RST), .Y(_02676_) );
  \$mux  #( .WIDTH(3) ) _49563_ ( .A(_stream_conv2d_16_source_36_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26258_) );
  \$mux  #( .WIDTH(3) ) _49564_ ( .A(_26258_), .B(3'h0), .S(RST), .Y(_02675_) );
  \$mux  #( .WIDTH(1) ) _49565_ ( .A(_stream_conv2d_16_source_36_idle), .B(1'h0), .S(_06781_), .Y(_26259_) );
  \$mux  #( .WIDTH(1) ) _49566_ ( .A(1'h1), .B(_26259_), .S(_05950_), .Y(_26260_) );
  \$mux  #( .WIDTH(1) ) _49567_ ( .A(_26260_), .B(1'h1), .S(RST), .Y(_02674_) );
  \$mux  #( .WIDTH(1) ) _49568_ ( .A(1'h0), .B(1'h1), .S(_ram_w4_l8192_id7_7_cond_1_1), .Y(_26261_) );
  \$mux  #( .WIDTH(1) ) _49569_ ( .A(_26261_), .B(1'h0), .S(RST), .Y(_02672_) );
  \$mux  #( .WIDTH(1) ) _49570_ ( .A(1'h1), .B(_stream_conv2d_16_source_35_source_ram_renable), .S(_05952_), .Y(_26262_) );
  \$mux  #( .WIDTH(1) ) _49571_ ( .A(1'h0), .B(_26262_), .S(_05951_), .Y(_26263_) );
  \$mux  #( .WIDTH(1) ) _49572_ ( .A(_26263_), .B(1'h0), .S(RST), .Y(_02671_) );
  \$mux  #( .WIDTH(32) ) _49573_ ( .A(_stream_conv2d_16_source_35_source_pat_all_offset), .B(_stream_conv2d_16_source_35_source_ram_raddr), .S(_05952_), .Y(_26264_) );
  \$mux  #( .WIDTH(32) ) _49574_ ( .A(_26264_), .B(0), .S(RST), .Y(_02670_) );
  \$mux  #( .WIDTH(8) ) _49575_ ( .A(_stream_conv2d_16_source_35_source_ram_sel), .B(8'h13), .S(_set_flag_710), .Y(_26265_) );
  \$mux  #( .WIDTH(8) ) _49576_ ( .A(_26265_), .B(8'h00), .S(RST), .Y(_02673_) );
  \$mux  #( .WIDTH(32) ) _49577_ ( .A(_stream_conv2d_16_source_35_source_offset_buf), .B(_stream_conv2d_16_source_35_source_offset), .S(_06776_), .Y(_26266_) );
  \$mux  #( .WIDTH(32) ) _49578_ ( .A(_26266_), .B(0), .S(RST), .Y(_02668_) );
  \$mux  #( .WIDTH(32) ) _49579_ ( .A(_stream_conv2d_16_source_35_source_offset), .B(conv2d_16_filter_page_comp_offset_buf), .S(_set_flag_710), .Y(_26267_) );
  \$mux  #( .WIDTH(32) ) _49580_ ( .A(_26267_), .B(0), .S(RST), .Y(_02667_) );
  \$mux  #( .WIDTH(3) ) _49581_ ( .A(_stream_conv2d_16_source_35_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26268_) );
  \$mux  #( .WIDTH(3) ) _49582_ ( .A(_26268_), .B(3'h0), .S(RST), .Y(_02666_) );
  \$mux  #( .WIDTH(1) ) _49583_ ( .A(_stream_conv2d_16_source_35_idle), .B(1'h0), .S(_06776_), .Y(_26269_) );
  \$mux  #( .WIDTH(1) ) _49584_ ( .A(1'h1), .B(_26269_), .S(_05951_), .Y(_26270_) );
  \$mux  #( .WIDTH(1) ) _49585_ ( .A(_26270_), .B(1'h1), .S(RST), .Y(_02665_) );
  \$mux  #( .WIDTH(1) ) _49586_ ( .A(1'h0), .B(1'h1), .S(_ram_w4_l8192_id6_2_cond_1_1), .Y(_26271_) );
  \$mux  #( .WIDTH(1) ) _49587_ ( .A(_26271_), .B(1'h0), .S(RST), .Y(_02663_) );
  \$mux  #( .WIDTH(1) ) _49588_ ( .A(1'h1), .B(_stream_conv2d_16_source_34_source_ram_renable), .S(_05954_), .Y(_26272_) );
  \$mux  #( .WIDTH(1) ) _49589_ ( .A(1'h0), .B(_26272_), .S(_05953_), .Y(_26273_) );
  \$mux  #( .WIDTH(1) ) _49590_ ( .A(_26273_), .B(1'h0), .S(RST), .Y(_02662_) );
  \$mux  #( .WIDTH(32) ) _49591_ ( .A(_stream_conv2d_16_source_34_source_pat_all_offset), .B(_stream_conv2d_16_source_34_source_ram_raddr), .S(_05954_), .Y(_26274_) );
  \$mux  #( .WIDTH(32) ) _49592_ ( .A(_26274_), .B(0), .S(RST), .Y(_02661_) );
  \$mux  #( .WIDTH(8) ) _49593_ ( .A(_stream_conv2d_16_source_34_source_ram_sel), .B(8'h12), .S(_set_flag_710), .Y(_26275_) );
  \$mux  #( .WIDTH(8) ) _49594_ ( .A(_26275_), .B(8'h00), .S(RST), .Y(_02664_) );
  \$mux  #( .WIDTH(32) ) _49595_ ( .A(_stream_conv2d_16_source_34_source_offset_buf), .B(_stream_conv2d_16_source_34_source_offset), .S(_06771_), .Y(_26276_) );
  \$mux  #( .WIDTH(32) ) _49596_ ( .A(_26276_), .B(0), .S(RST), .Y(_02659_) );
  \$mux  #( .WIDTH(32) ) _49597_ ( .A(_stream_conv2d_16_source_34_source_offset), .B(conv2d_16_filter_page_comp_offset_buf), .S(_set_flag_710), .Y(_26277_) );
  \$mux  #( .WIDTH(32) ) _49598_ ( .A(_26277_), .B(0), .S(RST), .Y(_02658_) );
  \$mux  #( .WIDTH(3) ) _49599_ ( .A(_stream_conv2d_16_source_34_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26278_) );
  \$mux  #( .WIDTH(3) ) _49600_ ( .A(_26278_), .B(3'h0), .S(RST), .Y(_02657_) );
  \$mux  #( .WIDTH(1) ) _49601_ ( .A(_stream_conv2d_16_source_34_idle), .B(1'h0), .S(_06771_), .Y(_26279_) );
  \$mux  #( .WIDTH(1) ) _49602_ ( .A(1'h1), .B(_26279_), .S(_05953_), .Y(_26280_) );
  \$mux  #( .WIDTH(1) ) _49603_ ( .A(_26280_), .B(1'h1), .S(RST), .Y(_02656_) );
  \$mux  #( .WIDTH(1) ) _49604_ ( .A(1'h0), .B(1'h1), .S(_ram_w4_l8192_id5_7_cond_2_1), .Y(_26281_) );
  \$mux  #( .WIDTH(1) ) _49605_ ( .A(_26281_), .B(1'h0), .S(RST), .Y(_02654_) );
  \$mux  #( .WIDTH(1) ) _49606_ ( .A(1'h1), .B(_stream_conv2d_16_source_33_source_ram_renable), .S(_05956_), .Y(_26282_) );
  \$mux  #( .WIDTH(1) ) _49607_ ( .A(1'h0), .B(_26282_), .S(_05955_), .Y(_26283_) );
  \$mux  #( .WIDTH(1) ) _49608_ ( .A(_26283_), .B(1'h0), .S(RST), .Y(_02653_) );
  \$mux  #( .WIDTH(32) ) _49609_ ( .A(_stream_conv2d_16_source_33_source_pat_all_offset), .B(_stream_conv2d_16_source_33_source_ram_raddr), .S(_05956_), .Y(_26284_) );
  \$mux  #( .WIDTH(32) ) _49610_ ( .A(_26284_), .B(0), .S(RST), .Y(_02652_) );
  \$mux  #( .WIDTH(8) ) _49611_ ( .A(_stream_conv2d_16_source_33_source_ram_sel), .B(8'h11), .S(_set_flag_710), .Y(_26285_) );
  \$mux  #( .WIDTH(8) ) _49612_ ( .A(_26285_), .B(8'h00), .S(RST), .Y(_02655_) );
  \$mux  #( .WIDTH(32) ) _49613_ ( .A(_stream_conv2d_16_source_33_source_offset_buf), .B(_stream_conv2d_16_source_33_source_offset), .S(_06766_), .Y(_26286_) );
  \$mux  #( .WIDTH(32) ) _49614_ ( .A(_26286_), .B(0), .S(RST), .Y(_02650_) );
  \$mux  #( .WIDTH(32) ) _49615_ ( .A(_stream_conv2d_16_source_33_source_offset), .B(conv2d_16_filter_page_comp_offset_buf), .S(_set_flag_710), .Y(_26287_) );
  \$mux  #( .WIDTH(32) ) _49616_ ( .A(_26287_), .B(0), .S(RST), .Y(_02649_) );
  \$mux  #( .WIDTH(3) ) _49617_ ( .A(_stream_conv2d_16_source_33_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26288_) );
  \$mux  #( .WIDTH(3) ) _49618_ ( .A(_26288_), .B(3'h0), .S(RST), .Y(_02648_) );
  \$mux  #( .WIDTH(1) ) _49619_ ( .A(_stream_conv2d_16_source_33_idle), .B(1'h0), .S(_06766_), .Y(_26289_) );
  \$mux  #( .WIDTH(1) ) _49620_ ( .A(1'h1), .B(_26289_), .S(_05955_), .Y(_26290_) );
  \$mux  #( .WIDTH(1) ) _49621_ ( .A(_26290_), .B(1'h1), .S(RST), .Y(_02647_) );
  \$mux  #( .WIDTH(1) ) _49622_ ( .A(1'h0), .B(1'h1), .S(_ram_w4_l8192_id4_7_cond_1_1), .Y(_26291_) );
  \$mux  #( .WIDTH(1) ) _49623_ ( .A(_26291_), .B(1'h0), .S(RST), .Y(_02645_) );
  \$mux  #( .WIDTH(1) ) _49624_ ( .A(1'h1), .B(_stream_conv2d_16_source_32_source_ram_renable), .S(_05959_), .Y(_26292_) );
  \$mux  #( .WIDTH(1) ) _49625_ ( .A(1'h0), .B(_26292_), .S(_05957_), .Y(_26293_) );
  \$mux  #( .WIDTH(1) ) _49626_ ( .A(_26293_), .B(1'h0), .S(RST), .Y(_02644_) );
  \$mux  #( .WIDTH(32) ) _49627_ ( .A(_stream_conv2d_16_source_32_source_pat_all_offset), .B(_stream_conv2d_16_source_32_source_ram_raddr), .S(_05959_), .Y(_26294_) );
  \$mux  #( .WIDTH(32) ) _49628_ ( .A(_26294_), .B(0), .S(RST), .Y(_02643_) );
  \$mux  #( .WIDTH(8) ) _49629_ ( .A(_stream_conv2d_16_source_32_source_ram_sel), .B(8'h10), .S(_set_flag_710), .Y(_26295_) );
  \$mux  #( .WIDTH(8) ) _49630_ ( .A(_26295_), .B(8'h00), .S(RST), .Y(_02646_) );
  \$mux  #( .WIDTH(32) ) _49631_ ( .A(_stream_conv2d_16_source_32_source_offset_buf), .B(_stream_conv2d_16_source_32_source_offset), .S(_06761_), .Y(_26296_) );
  \$mux  #( .WIDTH(32) ) _49632_ ( .A(_26296_), .B(0), .S(RST), .Y(_02641_) );
  \$mux  #( .WIDTH(32) ) _49633_ ( .A(_stream_conv2d_16_source_32_source_offset), .B(conv2d_16_filter_page_comp_offset_buf), .S(_set_flag_710), .Y(_26297_) );
  \$mux  #( .WIDTH(32) ) _49634_ ( .A(_26297_), .B(0), .S(RST), .Y(_02640_) );
  \$mux  #( .WIDTH(3) ) _49635_ ( .A(_stream_conv2d_16_source_32_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26298_) );
  \$mux  #( .WIDTH(3) ) _49636_ ( .A(_26298_), .B(3'h0), .S(RST), .Y(_02639_) );
  \$mux  #( .WIDTH(1) ) _49637_ ( .A(_stream_conv2d_16_source_32_idle), .B(1'h0), .S(_06761_), .Y(_26299_) );
  \$mux  #( .WIDTH(1) ) _49638_ ( .A(1'h1), .B(_26299_), .S(_05957_), .Y(_26300_) );
  \$mux  #( .WIDTH(1) ) _49639_ ( .A(_26300_), .B(1'h1), .S(RST), .Y(_02638_) );
  \$mux  #( .WIDTH(1) ) _49640_ ( .A(1'h0), .B(1'h1), .S(_ram_w4_l8192_id3_7_cond_1_1), .Y(_26301_) );
  \$mux  #( .WIDTH(1) ) _49641_ ( .A(_26301_), .B(1'h0), .S(RST), .Y(_02636_) );
  \$mux  #( .WIDTH(1) ) _49642_ ( .A(1'h1), .B(_stream_conv2d_16_source_31_source_ram_renable), .S(_05962_), .Y(_26302_) );
  \$mux  #( .WIDTH(1) ) _49643_ ( .A(1'h0), .B(_26302_), .S(_05958_), .Y(_26303_) );
  \$mux  #( .WIDTH(1) ) _49644_ ( .A(_26303_), .B(1'h0), .S(RST), .Y(_02635_) );
  \$mux  #( .WIDTH(32) ) _49645_ ( .A(_stream_conv2d_16_source_31_source_pat_all_offset), .B(_stream_conv2d_16_source_31_source_ram_raddr), .S(_05962_), .Y(_26304_) );
  \$mux  #( .WIDTH(32) ) _49646_ ( .A(_26304_), .B(0), .S(RST), .Y(_02634_) );
  \$mux  #( .WIDTH(8) ) _49647_ ( .A(_stream_conv2d_16_source_31_source_ram_sel), .B(8'h0f), .S(_set_flag_710), .Y(_26305_) );
  \$mux  #( .WIDTH(8) ) _49648_ ( .A(_26305_), .B(8'h00), .S(RST), .Y(_02637_) );
  \$mux  #( .WIDTH(32) ) _49649_ ( .A(_stream_conv2d_16_source_31_source_offset_buf), .B(_stream_conv2d_16_source_31_source_offset), .S(_06756_), .Y(_26306_) );
  \$mux  #( .WIDTH(32) ) _49650_ ( .A(_26306_), .B(0), .S(RST), .Y(_02632_) );
  \$mux  #( .WIDTH(32) ) _49651_ ( .A(_stream_conv2d_16_source_31_source_offset), .B(conv2d_16_filter_page_comp_offset_buf), .S(_set_flag_710), .Y(_26307_) );
  \$mux  #( .WIDTH(32) ) _49652_ ( .A(_26307_), .B(0), .S(RST), .Y(_02631_) );
  \$mux  #( .WIDTH(3) ) _49653_ ( .A(_stream_conv2d_16_source_31_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26308_) );
  \$mux  #( .WIDTH(3) ) _49654_ ( .A(_26308_), .B(3'h0), .S(RST), .Y(_02630_) );
  \$mux  #( .WIDTH(1) ) _49655_ ( .A(_stream_conv2d_16_source_31_idle), .B(1'h0), .S(_06756_), .Y(_26309_) );
  \$mux  #( .WIDTH(1) ) _49656_ ( .A(1'h1), .B(_26309_), .S(_05958_), .Y(_26310_) );
  \$mux  #( .WIDTH(1) ) _49657_ ( .A(_26310_), .B(1'h1), .S(RST), .Y(_02629_) );
  \$mux  #( .WIDTH(1) ) _49658_ ( .A(1'h0), .B(1'h1), .S(_ram_w4_l8192_id2_7_cond_1_1), .Y(_26311_) );
  \$mux  #( .WIDTH(1) ) _49659_ ( .A(_26311_), .B(1'h0), .S(RST), .Y(_02627_) );
  \$mux  #( .WIDTH(1) ) _49660_ ( .A(1'h1), .B(_stream_conv2d_16_source_30_source_ram_renable), .S(_05960_), .Y(_26312_) );
  \$mux  #( .WIDTH(1) ) _49661_ ( .A(1'h0), .B(_26312_), .S(_05961_), .Y(_26313_) );
  \$mux  #( .WIDTH(1) ) _49662_ ( .A(_26313_), .B(1'h0), .S(RST), .Y(_02626_) );
  \$mux  #( .WIDTH(32) ) _49663_ ( .A(_stream_conv2d_16_source_30_source_pat_all_offset), .B(_stream_conv2d_16_source_30_source_ram_raddr), .S(_05960_), .Y(_26314_) );
  \$mux  #( .WIDTH(32) ) _49664_ ( .A(_26314_), .B(0), .S(RST), .Y(_02625_) );
  \$mux  #( .WIDTH(8) ) _49665_ ( .A(_stream_conv2d_16_source_30_source_ram_sel), .B(8'h0e), .S(_set_flag_710), .Y(_26315_) );
  \$mux  #( .WIDTH(8) ) _49666_ ( .A(_26315_), .B(8'h00), .S(RST), .Y(_02628_) );
  \$mux  #( .WIDTH(32) ) _49667_ ( .A(_stream_conv2d_16_source_30_source_offset_buf), .B(_stream_conv2d_16_source_30_source_offset), .S(_06751_), .Y(_26316_) );
  \$mux  #( .WIDTH(32) ) _49668_ ( .A(_26316_), .B(0), .S(RST), .Y(_02623_) );
  \$mux  #( .WIDTH(32) ) _49669_ ( .A(_stream_conv2d_16_source_30_source_offset), .B(conv2d_16_filter_page_comp_offset_buf), .S(_set_flag_710), .Y(_26317_) );
  \$mux  #( .WIDTH(32) ) _49670_ ( .A(_26317_), .B(0), .S(RST), .Y(_02622_) );
  \$mux  #( .WIDTH(3) ) _49671_ ( .A(_stream_conv2d_16_source_30_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26318_) );
  \$mux  #( .WIDTH(3) ) _49672_ ( .A(_26318_), .B(3'h0), .S(RST), .Y(_02621_) );
  \$mux  #( .WIDTH(1) ) _49673_ ( .A(_stream_conv2d_16_source_30_idle), .B(1'h0), .S(_06751_), .Y(_26319_) );
  \$mux  #( .WIDTH(1) ) _49674_ ( .A(1'h1), .B(_26319_), .S(_05961_), .Y(_26320_) );
  \$mux  #( .WIDTH(1) ) _49675_ ( .A(_26320_), .B(1'h1), .S(RST), .Y(_02620_) );
  \$mux  #( .WIDTH(1) ) _49676_ ( .A(1'h0), .B(1'h1), .S(_ram_w4_l8192_id1_7_cond_1_1), .Y(_26321_) );
  \$mux  #( .WIDTH(1) ) _49677_ ( .A(_26321_), .B(1'h0), .S(RST), .Y(_02618_) );
  \$mux  #( .WIDTH(1) ) _49678_ ( .A(1'h1), .B(_stream_conv2d_16_source_29_source_ram_renable), .S(_05965_), .Y(_26322_) );
  \$mux  #( .WIDTH(1) ) _49679_ ( .A(1'h0), .B(_26322_), .S(_05963_), .Y(_26323_) );
  \$mux  #( .WIDTH(1) ) _49680_ ( .A(_26323_), .B(1'h0), .S(RST), .Y(_02617_) );
  \$mux  #( .WIDTH(32) ) _49681_ ( .A(_stream_conv2d_16_source_29_source_pat_all_offset), .B(_stream_conv2d_16_source_29_source_ram_raddr), .S(_05965_), .Y(_26324_) );
  \$mux  #( .WIDTH(32) ) _49682_ ( .A(_26324_), .B(0), .S(RST), .Y(_02616_) );
  \$mux  #( .WIDTH(8) ) _49683_ ( .A(_stream_conv2d_16_source_29_source_ram_sel), .B(8'h0d), .S(_set_flag_710), .Y(_26325_) );
  \$mux  #( .WIDTH(8) ) _49684_ ( .A(_26325_), .B(8'h00), .S(RST), .Y(_02619_) );
  \$mux  #( .WIDTH(32) ) _49685_ ( .A(_stream_conv2d_16_source_29_source_offset_buf), .B(_stream_conv2d_16_source_29_source_offset), .S(_06746_), .Y(_26326_) );
  \$mux  #( .WIDTH(32) ) _49686_ ( .A(_26326_), .B(0), .S(RST), .Y(_02614_) );
  \$mux  #( .WIDTH(32) ) _49687_ ( .A(_stream_conv2d_16_source_29_source_offset), .B(conv2d_16_filter_page_comp_offset_buf), .S(_set_flag_710), .Y(_26327_) );
  \$mux  #( .WIDTH(32) ) _49688_ ( .A(_26327_), .B(0), .S(RST), .Y(_02613_) );
  \$mux  #( .WIDTH(3) ) _49689_ ( .A(_stream_conv2d_16_source_29_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26328_) );
  \$mux  #( .WIDTH(3) ) _49690_ ( .A(_26328_), .B(3'h0), .S(RST), .Y(_02612_) );
  \$mux  #( .WIDTH(1) ) _49691_ ( .A(_stream_conv2d_16_source_29_idle), .B(1'h0), .S(_06746_), .Y(_26329_) );
  \$mux  #( .WIDTH(1) ) _49692_ ( .A(1'h1), .B(_26329_), .S(_05963_), .Y(_26330_) );
  \$mux  #( .WIDTH(1) ) _49693_ ( .A(_26330_), .B(1'h1), .S(RST), .Y(_02611_) );
  \$mux  #( .WIDTH(1) ) _49694_ ( .A(1'h0), .B(1'h1), .S(_ram_w4_l8192_id0_7_cond_2_1), .Y(_26331_) );
  \$mux  #( .WIDTH(1) ) _49695_ ( .A(_26331_), .B(1'h0), .S(RST), .Y(_02609_) );
  \$mux  #( .WIDTH(1) ) _49696_ ( .A(1'h1), .B(_stream_conv2d_16_source_28_source_ram_renable), .S(_05966_), .Y(_26332_) );
  \$mux  #( .WIDTH(1) ) _49697_ ( .A(1'h0), .B(_26332_), .S(_05964_), .Y(_26333_) );
  \$mux  #( .WIDTH(1) ) _49698_ ( .A(_26333_), .B(1'h0), .S(RST), .Y(_02608_) );
  \$mux  #( .WIDTH(32) ) _49699_ ( .A(_stream_conv2d_16_source_28_source_pat_all_offset), .B(_stream_conv2d_16_source_28_source_ram_raddr), .S(_05966_), .Y(_26334_) );
  \$mux  #( .WIDTH(32) ) _49700_ ( .A(_26334_), .B(0), .S(RST), .Y(_02607_) );
  \$mux  #( .WIDTH(8) ) _49701_ ( .A(_stream_conv2d_16_source_28_source_ram_sel), .B(8'h0c), .S(_set_flag_710), .Y(_26335_) );
  \$mux  #( .WIDTH(8) ) _49702_ ( .A(_26335_), .B(8'h00), .S(RST), .Y(_02610_) );
  \$mux  #( .WIDTH(32) ) _49703_ ( .A(_stream_conv2d_16_source_28_source_offset_buf), .B(_stream_conv2d_16_source_28_source_offset), .S(_06741_), .Y(_26336_) );
  \$mux  #( .WIDTH(32) ) _49704_ ( .A(_26336_), .B(0), .S(RST), .Y(_02605_) );
  \$mux  #( .WIDTH(32) ) _49705_ ( .A(_stream_conv2d_16_source_28_source_offset), .B(conv2d_16_filter_page_comp_offset_buf), .S(_set_flag_710), .Y(_26337_) );
  \$mux  #( .WIDTH(32) ) _49706_ ( .A(_26337_), .B(0), .S(RST), .Y(_02604_) );
  \$mux  #( .WIDTH(3) ) _49707_ ( .A(_stream_conv2d_16_source_28_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26338_) );
  \$mux  #( .WIDTH(3) ) _49708_ ( .A(_26338_), .B(3'h0), .S(RST), .Y(_02603_) );
  \$mux  #( .WIDTH(1) ) _49709_ ( .A(_stream_conv2d_16_source_28_idle), .B(1'h0), .S(_06741_), .Y(_26339_) );
  \$mux  #( .WIDTH(1) ) _49710_ ( .A(1'h1), .B(_26339_), .S(_05964_), .Y(_26340_) );
  \$mux  #( .WIDTH(1) ) _49711_ ( .A(_26340_), .B(1'h1), .S(RST), .Y(_02602_) );
  \$mux  #( .WIDTH(1) ) _49712_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id10_0_cond_2_1), .Y(_26341_) );
  \$mux  #( .WIDTH(1) ) _49713_ ( .A(_26341_), .B(1'h0), .S(RST), .Y(_02600_) );
  \$mux  #( .WIDTH(1) ) _49714_ ( .A(1'h1), .B(_stream_conv2d_16_source_27_source_ram_renable), .S(_05968_), .Y(_26342_) );
  \$mux  #( .WIDTH(1) ) _49715_ ( .A(1'h0), .B(_26342_), .S(_05967_), .Y(_26343_) );
  \$mux  #( .WIDTH(1) ) _49716_ ( .A(_26343_), .B(1'h0), .S(RST), .Y(_02599_) );
  \$mux  #( .WIDTH(32) ) _49717_ ( .A(_stream_conv2d_16_source_27_source_pat_all_offset), .B(_stream_conv2d_16_source_27_source_ram_raddr), .S(_05968_), .Y(_26344_) );
  \$mux  #( .WIDTH(32) ) _49718_ ( .A(_26344_), .B(0), .S(RST), .Y(_02598_) );
  \$mux  #( .WIDTH(8) ) _49719_ ( .A(_stream_conv2d_16_source_27_source_ram_sel), .B(8'h0b), .S(_set_flag_710), .Y(_26345_) );
  \$mux  #( .WIDTH(8) ) _49720_ ( .A(_26345_), .B(8'h00), .S(RST), .Y(_02601_) );
  \$mux  #( .WIDTH(32) ) _49721_ ( .A(_stream_conv2d_16_source_27_source_offset_buf), .B(_stream_conv2d_16_source_27_source_offset), .S(_06736_), .Y(_26346_) );
  \$mux  #( .WIDTH(32) ) _49722_ ( .A(_26346_), .B(0), .S(RST), .Y(_02596_) );
  \$mux  #( .WIDTH(32) ) _49723_ ( .A(_stream_conv2d_16_source_27_source_offset), .B(_24356_), .S(_set_flag_710), .Y(_26347_) );
  \$mux  #( .WIDTH(32) ) _49724_ ( .A(_26347_), .B(0), .S(RST), .Y(_02595_) );
  \$mux  #( .WIDTH(3) ) _49725_ ( .A(_stream_conv2d_16_source_27_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26348_) );
  \$mux  #( .WIDTH(3) ) _49726_ ( .A(_26348_), .B(3'h0), .S(RST), .Y(_02594_) );
  \$mux  #( .WIDTH(1) ) _49727_ ( .A(_stream_conv2d_16_source_27_idle), .B(1'h0), .S(_06736_), .Y(_26349_) );
  \$mux  #( .WIDTH(1) ) _49728_ ( .A(1'h1), .B(_26349_), .S(_05967_), .Y(_26350_) );
  \$mux  #( .WIDTH(1) ) _49729_ ( .A(_26350_), .B(1'h1), .S(RST), .Y(_02593_) );
  \$mux  #( .WIDTH(1) ) _49730_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id9_0_cond_2_1), .Y(_26351_) );
  \$mux  #( .WIDTH(1) ) _49731_ ( .A(_26351_), .B(1'h0), .S(RST), .Y(_02591_) );
  \$mux  #( .WIDTH(1) ) _49732_ ( .A(1'h1), .B(_stream_conv2d_16_source_26_source_ram_renable), .S(_05971_), .Y(_26352_) );
  \$mux  #( .WIDTH(1) ) _49733_ ( .A(1'h0), .B(_26352_), .S(_05969_), .Y(_26353_) );
  \$mux  #( .WIDTH(1) ) _49734_ ( .A(_26353_), .B(1'h0), .S(RST), .Y(_02590_) );
  \$mux  #( .WIDTH(32) ) _49735_ ( .A(_stream_conv2d_16_source_26_source_pat_all_offset), .B(_stream_conv2d_16_source_26_source_ram_raddr), .S(_05971_), .Y(_26354_) );
  \$mux  #( .WIDTH(32) ) _49736_ ( .A(_26354_), .B(0), .S(RST), .Y(_02589_) );
  \$mux  #( .WIDTH(8) ) _49737_ ( .A(_stream_conv2d_16_source_26_source_ram_sel), .B(8'h0a), .S(_set_flag_710), .Y(_26355_) );
  \$mux  #( .WIDTH(8) ) _49738_ ( .A(_26355_), .B(8'h00), .S(RST), .Y(_02592_) );
  \$mux  #( .WIDTH(32) ) _49739_ ( .A(_stream_conv2d_16_source_26_source_offset_buf), .B(_stream_conv2d_16_source_26_source_offset), .S(_06731_), .Y(_26356_) );
  \$mux  #( .WIDTH(32) ) _49740_ ( .A(_26356_), .B(0), .S(RST), .Y(_02587_) );
  \$mux  #( .WIDTH(32) ) _49741_ ( .A(_stream_conv2d_16_source_26_source_offset), .B(_24351_), .S(_set_flag_710), .Y(_26357_) );
  \$mux  #( .WIDTH(32) ) _49742_ ( .A(_26357_), .B(0), .S(RST), .Y(_02586_) );
  \$mux  #( .WIDTH(3) ) _49743_ ( .A(_stream_conv2d_16_source_26_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26358_) );
  \$mux  #( .WIDTH(3) ) _49744_ ( .A(_26358_), .B(3'h0), .S(RST), .Y(_02585_) );
  \$mux  #( .WIDTH(1) ) _49745_ ( .A(_stream_conv2d_16_source_26_idle), .B(1'h0), .S(_06731_), .Y(_26359_) );
  \$mux  #( .WIDTH(1) ) _49746_ ( .A(1'h1), .B(_26359_), .S(_05969_), .Y(_26360_) );
  \$mux  #( .WIDTH(1) ) _49747_ ( .A(_26360_), .B(1'h1), .S(RST), .Y(_02584_) );
  \$mux  #( .WIDTH(1) ) _49748_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id8_0_cond_3_1), .Y(_26361_) );
  \$mux  #( .WIDTH(1) ) _49749_ ( .A(_26361_), .B(1'h0), .S(RST), .Y(_02582_) );
  \$mux  #( .WIDTH(1) ) _49750_ ( .A(1'h1), .B(_stream_conv2d_16_source_25_source_ram_renable), .S(_05974_), .Y(_26362_) );
  \$mux  #( .WIDTH(1) ) _49751_ ( .A(1'h0), .B(_26362_), .S(_05970_), .Y(_26363_) );
  \$mux  #( .WIDTH(1) ) _49752_ ( .A(_26363_), .B(1'h0), .S(RST), .Y(_02581_) );
  \$mux  #( .WIDTH(32) ) _49753_ ( .A(_stream_conv2d_16_source_25_source_pat_all_offset), .B(_stream_conv2d_16_source_25_source_ram_raddr), .S(_05974_), .Y(_26364_) );
  \$mux  #( .WIDTH(32) ) _49754_ ( .A(_26364_), .B(0), .S(RST), .Y(_02580_) );
  \$mux  #( .WIDTH(8) ) _49755_ ( .A(_stream_conv2d_16_source_25_source_ram_sel), .B(8'h09), .S(_set_flag_710), .Y(_26365_) );
  \$mux  #( .WIDTH(8) ) _49756_ ( .A(_26365_), .B(8'h00), .S(RST), .Y(_02583_) );
  \$mux  #( .WIDTH(32) ) _49757_ ( .A(_stream_conv2d_16_source_25_source_offset_buf), .B(_stream_conv2d_16_source_25_source_offset), .S(_06726_), .Y(_26366_) );
  \$mux  #( .WIDTH(32) ) _49758_ ( .A(_26366_), .B(0), .S(RST), .Y(_02578_) );
  \$mux  #( .WIDTH(32) ) _49759_ ( .A(_stream_conv2d_16_source_25_source_offset), .B(_24346_), .S(_set_flag_710), .Y(_26367_) );
  \$mux  #( .WIDTH(32) ) _49760_ ( .A(_26367_), .B(0), .S(RST), .Y(_02577_) );
  \$mux  #( .WIDTH(3) ) _49761_ ( .A(_stream_conv2d_16_source_25_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26368_) );
  \$mux  #( .WIDTH(3) ) _49762_ ( .A(_26368_), .B(3'h0), .S(RST), .Y(_02576_) );
  \$mux  #( .WIDTH(1) ) _49763_ ( .A(_stream_conv2d_16_source_25_idle), .B(1'h0), .S(_06726_), .Y(_26369_) );
  \$mux  #( .WIDTH(1) ) _49764_ ( .A(1'h1), .B(_26369_), .S(_05970_), .Y(_26370_) );
  \$mux  #( .WIDTH(1) ) _49765_ ( .A(_26370_), .B(1'h1), .S(RST), .Y(_02575_) );
  \$mux  #( .WIDTH(1) ) _49766_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id7_0_cond_2_1), .Y(_26371_) );
  \$mux  #( .WIDTH(1) ) _49767_ ( .A(_26371_), .B(1'h0), .S(RST), .Y(_02573_) );
  \$mux  #( .WIDTH(1) ) _49768_ ( .A(1'h1), .B(_stream_conv2d_16_source_24_source_ram_renable), .S(_05972_), .Y(_26372_) );
  \$mux  #( .WIDTH(1) ) _49769_ ( .A(1'h0), .B(_26372_), .S(_05973_), .Y(_26373_) );
  \$mux  #( .WIDTH(1) ) _49770_ ( .A(_26373_), .B(1'h0), .S(RST), .Y(_02572_) );
  \$mux  #( .WIDTH(32) ) _49771_ ( .A(_stream_conv2d_16_source_24_source_pat_all_offset), .B(_stream_conv2d_16_source_24_source_ram_raddr), .S(_05972_), .Y(_26374_) );
  \$mux  #( .WIDTH(32) ) _49772_ ( .A(_26374_), .B(0), .S(RST), .Y(_02571_) );
  \$mux  #( .WIDTH(8) ) _49773_ ( .A(_stream_conv2d_16_source_24_source_ram_sel), .B(8'h08), .S(_set_flag_710), .Y(_26375_) );
  \$mux  #( .WIDTH(8) ) _49774_ ( .A(_26375_), .B(8'h00), .S(RST), .Y(_02574_) );
  \$mux  #( .WIDTH(32) ) _49775_ ( .A(_stream_conv2d_16_source_24_source_offset_buf), .B(_stream_conv2d_16_source_24_source_offset), .S(_06721_), .Y(_26376_) );
  \$mux  #( .WIDTH(32) ) _49776_ ( .A(_26376_), .B(0), .S(RST), .Y(_02569_) );
  \$mux  #( .WIDTH(32) ) _49777_ ( .A(_stream_conv2d_16_source_24_source_offset), .B(_24341_), .S(_set_flag_710), .Y(_26377_) );
  \$mux  #( .WIDTH(32) ) _49778_ ( .A(_26377_), .B(0), .S(RST), .Y(_02568_) );
  \$mux  #( .WIDTH(3) ) _49779_ ( .A(_stream_conv2d_16_source_24_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26378_) );
  \$mux  #( .WIDTH(3) ) _49780_ ( .A(_26378_), .B(3'h0), .S(RST), .Y(_02567_) );
  \$mux  #( .WIDTH(1) ) _49781_ ( .A(_stream_conv2d_16_source_24_idle), .B(1'h0), .S(_06721_), .Y(_26379_) );
  \$mux  #( .WIDTH(1) ) _49782_ ( .A(1'h1), .B(_26379_), .S(_05973_), .Y(_26380_) );
  \$mux  #( .WIDTH(1) ) _49783_ ( .A(_26380_), .B(1'h1), .S(RST), .Y(_02566_) );
  \$mux  #( .WIDTH(1) ) _49784_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id6_0_cond_2_1), .Y(_26381_) );
  \$mux  #( .WIDTH(1) ) _49785_ ( .A(_26381_), .B(1'h0), .S(RST), .Y(_02564_) );
  \$mux  #( .WIDTH(1) ) _49786_ ( .A(1'h1), .B(_stream_conv2d_16_source_23_source_ram_renable), .S(_05977_), .Y(_26382_) );
  \$mux  #( .WIDTH(1) ) _49787_ ( .A(1'h0), .B(_26382_), .S(_05975_), .Y(_26383_) );
  \$mux  #( .WIDTH(1) ) _49788_ ( .A(_26383_), .B(1'h0), .S(RST), .Y(_02563_) );
  \$mux  #( .WIDTH(32) ) _49789_ ( .A(_stream_conv2d_16_source_23_source_pat_all_offset), .B(_stream_conv2d_16_source_23_source_ram_raddr), .S(_05977_), .Y(_26384_) );
  \$mux  #( .WIDTH(32) ) _49790_ ( .A(_26384_), .B(0), .S(RST), .Y(_02562_) );
  \$mux  #( .WIDTH(8) ) _49791_ ( .A(_stream_conv2d_16_source_23_source_ram_sel), .B(8'h07), .S(_set_flag_710), .Y(_26385_) );
  \$mux  #( .WIDTH(8) ) _49792_ ( .A(_26385_), .B(8'h00), .S(RST), .Y(_02565_) );
  \$mux  #( .WIDTH(32) ) _49793_ ( .A(_stream_conv2d_16_source_23_source_offset_buf), .B(_stream_conv2d_16_source_23_source_offset), .S(_06716_), .Y(_26386_) );
  \$mux  #( .WIDTH(32) ) _49794_ ( .A(_26386_), .B(0), .S(RST), .Y(_02560_) );
  \$mux  #( .WIDTH(32) ) _49795_ ( .A(_stream_conv2d_16_source_23_source_offset), .B(_24336_), .S(_set_flag_710), .Y(_26387_) );
  \$mux  #( .WIDTH(32) ) _49796_ ( .A(_26387_), .B(0), .S(RST), .Y(_02559_) );
  \$mux  #( .WIDTH(3) ) _49797_ ( .A(_stream_conv2d_16_source_23_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26388_) );
  \$mux  #( .WIDTH(3) ) _49798_ ( .A(_26388_), .B(3'h0), .S(RST), .Y(_02558_) );
  \$mux  #( .WIDTH(1) ) _49799_ ( .A(_stream_conv2d_16_source_23_idle), .B(1'h0), .S(_06716_), .Y(_26389_) );
  \$mux  #( .WIDTH(1) ) _49800_ ( .A(1'h1), .B(_26389_), .S(_05975_), .Y(_26390_) );
  \$mux  #( .WIDTH(1) ) _49801_ ( .A(_26390_), .B(1'h1), .S(RST), .Y(_02557_) );
  \$mux  #( .WIDTH(1) ) _49802_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id5_0_cond_3_1), .Y(_26391_) );
  \$mux  #( .WIDTH(1) ) _49803_ ( .A(_26391_), .B(1'h0), .S(RST), .Y(_02555_) );
  \$mux  #( .WIDTH(1) ) _49804_ ( .A(1'h1), .B(_stream_conv2d_16_source_22_source_ram_renable), .S(_05979_), .Y(_26392_) );
  \$mux  #( .WIDTH(1) ) _49805_ ( .A(1'h0), .B(_26392_), .S(_05976_), .Y(_26393_) );
  \$mux  #( .WIDTH(1) ) _49806_ ( .A(_26393_), .B(1'h0), .S(RST), .Y(_02554_) );
  \$mux  #( .WIDTH(32) ) _49807_ ( .A(_stream_conv2d_16_source_22_source_pat_all_offset), .B(_stream_conv2d_16_source_22_source_ram_raddr), .S(_05979_), .Y(_26394_) );
  \$mux  #( .WIDTH(32) ) _49808_ ( .A(_26394_), .B(0), .S(RST), .Y(_02553_) );
  \$mux  #( .WIDTH(8) ) _49809_ ( .A(_stream_conv2d_16_source_22_source_ram_sel), .B(8'h06), .S(_set_flag_710), .Y(_26395_) );
  \$mux  #( .WIDTH(8) ) _49810_ ( .A(_26395_), .B(8'h00), .S(RST), .Y(_02556_) );
  \$mux  #( .WIDTH(32) ) _49811_ ( .A(_stream_conv2d_16_source_22_source_offset_buf), .B(_stream_conv2d_16_source_22_source_offset), .S(_06711_), .Y(_26396_) );
  \$mux  #( .WIDTH(32) ) _49812_ ( .A(_26396_), .B(0), .S(RST), .Y(_02551_) );
  \$mux  #( .WIDTH(32) ) _49813_ ( .A(_stream_conv2d_16_source_22_source_offset), .B(_24331_), .S(_set_flag_710), .Y(_26397_) );
  \$mux  #( .WIDTH(32) ) _49814_ ( .A(_26397_), .B(0), .S(RST), .Y(_02550_) );
  \$mux  #( .WIDTH(3) ) _49815_ ( .A(_stream_conv2d_16_source_22_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26398_) );
  \$mux  #( .WIDTH(3) ) _49816_ ( .A(_26398_), .B(3'h0), .S(RST), .Y(_02549_) );
  \$mux  #( .WIDTH(1) ) _49817_ ( .A(_stream_conv2d_16_source_22_idle), .B(1'h0), .S(_06711_), .Y(_26399_) );
  \$mux  #( .WIDTH(1) ) _49818_ ( .A(1'h1), .B(_26399_), .S(_05976_), .Y(_26400_) );
  \$mux  #( .WIDTH(1) ) _49819_ ( .A(_26400_), .B(1'h1), .S(RST), .Y(_02548_) );
  \$mux  #( .WIDTH(1) ) _49820_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id4_0_cond_2_1), .Y(_26401_) );
  \$mux  #( .WIDTH(1) ) _49821_ ( .A(_26401_), .B(1'h0), .S(RST), .Y(_02546_) );
  \$mux  #( .WIDTH(1) ) _49822_ ( .A(1'h1), .B(_stream_conv2d_16_source_21_source_ram_renable), .S(_05981_), .Y(_26402_) );
  \$mux  #( .WIDTH(1) ) _49823_ ( .A(1'h0), .B(_26402_), .S(_05978_), .Y(_26403_) );
  \$mux  #( .WIDTH(1) ) _49824_ ( .A(_26403_), .B(1'h0), .S(RST), .Y(_02545_) );
  \$mux  #( .WIDTH(32) ) _49825_ ( .A(_stream_conv2d_16_source_21_source_pat_all_offset), .B(_stream_conv2d_16_source_21_source_ram_raddr), .S(_05981_), .Y(_26404_) );
  \$mux  #( .WIDTH(32) ) _49826_ ( .A(_26404_), .B(0), .S(RST), .Y(_02544_) );
  \$mux  #( .WIDTH(8) ) _49827_ ( .A(_stream_conv2d_16_source_21_source_ram_sel), .B(8'h05), .S(_set_flag_710), .Y(_26405_) );
  \$mux  #( .WIDTH(8) ) _49828_ ( .A(_26405_), .B(8'h00), .S(RST), .Y(_02547_) );
  \$mux  #( .WIDTH(32) ) _49829_ ( .A(_stream_conv2d_16_source_21_source_offset_buf), .B(_stream_conv2d_16_source_21_source_offset), .S(_06706_), .Y(_26406_) );
  \$mux  #( .WIDTH(32) ) _49830_ ( .A(_26406_), .B(0), .S(RST), .Y(_02542_) );
  \$mux  #( .WIDTH(32) ) _49831_ ( .A(_stream_conv2d_16_source_21_source_offset), .B(_24326_), .S(_set_flag_710), .Y(_26407_) );
  \$mux  #( .WIDTH(32) ) _49832_ ( .A(_26407_), .B(0), .S(RST), .Y(_02541_) );
  \$mux  #( .WIDTH(3) ) _49833_ ( .A(_stream_conv2d_16_source_21_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26408_) );
  \$mux  #( .WIDTH(3) ) _49834_ ( .A(_26408_), .B(3'h0), .S(RST), .Y(_02540_) );
  \$mux  #( .WIDTH(1) ) _49835_ ( .A(_stream_conv2d_16_source_21_idle), .B(1'h0), .S(_06706_), .Y(_26409_) );
  \$mux  #( .WIDTH(1) ) _49836_ ( .A(1'h1), .B(_26409_), .S(_05978_), .Y(_26410_) );
  \$mux  #( .WIDTH(1) ) _49837_ ( .A(_26410_), .B(1'h1), .S(RST), .Y(_02539_) );
  \$mux  #( .WIDTH(1) ) _49838_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id3_0_cond_2_1), .Y(_26411_) );
  \$mux  #( .WIDTH(1) ) _49839_ ( .A(_26411_), .B(1'h0), .S(RST), .Y(_02537_) );
  \$mux  #( .WIDTH(1) ) _49840_ ( .A(1'h1), .B(_stream_conv2d_16_source_20_source_ram_renable), .S(_05982_), .Y(_26412_) );
  \$mux  #( .WIDTH(1) ) _49841_ ( .A(1'h0), .B(_26412_), .S(_05980_), .Y(_26413_) );
  \$mux  #( .WIDTH(1) ) _49842_ ( .A(_26413_), .B(1'h0), .S(RST), .Y(_02536_) );
  \$mux  #( .WIDTH(32) ) _49843_ ( .A(_stream_conv2d_16_source_20_source_pat_all_offset), .B(_stream_conv2d_16_source_20_source_ram_raddr), .S(_05982_), .Y(_26414_) );
  \$mux  #( .WIDTH(32) ) _49844_ ( .A(_26414_), .B(0), .S(RST), .Y(_02535_) );
  \$mux  #( .WIDTH(8) ) _49845_ ( .A(_stream_conv2d_16_source_20_source_ram_sel), .B(8'h04), .S(_set_flag_710), .Y(_26415_) );
  \$mux  #( .WIDTH(8) ) _49846_ ( .A(_26415_), .B(8'h00), .S(RST), .Y(_02538_) );
  \$mux  #( .WIDTH(32) ) _49847_ ( .A(_stream_conv2d_16_source_20_source_offset_buf), .B(_stream_conv2d_16_source_20_source_offset), .S(_06701_), .Y(_26416_) );
  \$mux  #( .WIDTH(32) ) _49848_ ( .A(_26416_), .B(0), .S(RST), .Y(_02533_) );
  \$mux  #( .WIDTH(32) ) _49849_ ( .A(_stream_conv2d_16_source_20_source_offset), .B(_24321_), .S(_set_flag_710), .Y(_26417_) );
  \$mux  #( .WIDTH(32) ) _49850_ ( .A(_26417_), .B(0), .S(RST), .Y(_02532_) );
  \$mux  #( .WIDTH(3) ) _49851_ ( .A(_stream_conv2d_16_source_20_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26418_) );
  \$mux  #( .WIDTH(3) ) _49852_ ( .A(_26418_), .B(3'h0), .S(RST), .Y(_02531_) );
  \$mux  #( .WIDTH(1) ) _49853_ ( .A(_stream_conv2d_16_source_20_idle), .B(1'h0), .S(_06701_), .Y(_26419_) );
  \$mux  #( .WIDTH(1) ) _49854_ ( .A(1'h1), .B(_26419_), .S(_05980_), .Y(_26420_) );
  \$mux  #( .WIDTH(1) ) _49855_ ( .A(_26420_), .B(1'h1), .S(RST), .Y(_02530_) );
  \$mux  #( .WIDTH(1) ) _49856_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id2_0_cond_3_1), .Y(_26421_) );
  \$mux  #( .WIDTH(1) ) _49857_ ( .A(_26421_), .B(1'h0), .S(RST), .Y(_02528_) );
  \$mux  #( .WIDTH(1) ) _49858_ ( .A(1'h1), .B(_stream_conv2d_16_source_19_source_ram_renable), .S(_05983_), .Y(_26422_) );
  \$mux  #( .WIDTH(1) ) _49859_ ( .A(1'h0), .B(_26422_), .S(_05984_), .Y(_26423_) );
  \$mux  #( .WIDTH(1) ) _49860_ ( .A(_26423_), .B(1'h0), .S(RST), .Y(_02527_) );
  \$mux  #( .WIDTH(32) ) _49861_ ( .A(_stream_conv2d_16_source_19_source_pat_all_offset), .B(_stream_conv2d_16_source_19_source_ram_raddr), .S(_05983_), .Y(_26424_) );
  \$mux  #( .WIDTH(32) ) _49862_ ( .A(_26424_), .B(0), .S(RST), .Y(_02526_) );
  \$mux  #( .WIDTH(8) ) _49863_ ( .A(_stream_conv2d_16_source_19_source_ram_sel), .B(8'h03), .S(_set_flag_710), .Y(_26425_) );
  \$mux  #( .WIDTH(8) ) _49864_ ( .A(_26425_), .B(8'h00), .S(RST), .Y(_02529_) );
  \$mux  #( .WIDTH(32) ) _49865_ ( .A(_stream_conv2d_16_source_19_source_offset_buf), .B(_stream_conv2d_16_source_19_source_offset), .S(_06696_), .Y(_26426_) );
  \$mux  #( .WIDTH(32) ) _49866_ ( .A(_26426_), .B(0), .S(RST), .Y(_02524_) );
  \$mux  #( .WIDTH(32) ) _49867_ ( .A(_stream_conv2d_16_source_19_source_offset), .B(_24316_), .S(_set_flag_710), .Y(_26427_) );
  \$mux  #( .WIDTH(32) ) _49868_ ( .A(_26427_), .B(0), .S(RST), .Y(_02523_) );
  \$mux  #( .WIDTH(3) ) _49869_ ( .A(_stream_conv2d_16_source_19_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26428_) );
  \$mux  #( .WIDTH(3) ) _49870_ ( .A(_26428_), .B(3'h0), .S(RST), .Y(_02522_) );
  \$mux  #( .WIDTH(1) ) _49871_ ( .A(_stream_conv2d_16_source_19_idle), .B(1'h0), .S(_06696_), .Y(_26429_) );
  \$mux  #( .WIDTH(1) ) _49872_ ( .A(1'h1), .B(_26429_), .S(_05984_), .Y(_26430_) );
  \$mux  #( .WIDTH(1) ) _49873_ ( .A(_26430_), .B(1'h1), .S(RST), .Y(_02521_) );
  \$mux  #( .WIDTH(4) ) _49874_ ( .A(_stream_conv2d_16_constant_17_next_constant_data), .B(cparam_conv2d_16_cshamt_out_value), .S(_set_flag_710), .Y(_26431_) );
  \$mux  #( .WIDTH(4) ) _49875_ ( .A(_26431_), .B(4'h0), .S(RST), .Y(_02498_) );
  \$mux  #( .WIDTH(1) ) _49876_ ( .A(_stream_conv2d_16_constant_16_next_constant_data), .B(1'h0), .S(_set_flag_710), .Y(_26432_) );
  \$mux  #( .WIDTH(1) ) _49877_ ( .A(_26432_), .B(1'h0), .S(RST), .Y(_02497_) );
  \$mux  #( .WIDTH(1) ) _49878_ ( .A(_stream_conv2d_16_constant_15_next_constant_data), .B(1'h0), .S(_set_flag_710), .Y(_26433_) );
  \$mux  #( .WIDTH(1) ) _49879_ ( .A(_26433_), .B(1'h0), .S(RST), .Y(_02496_) );
  \$mux  #( .WIDTH(8) ) _49880_ ( .A(_stream_conv2d_16_source_14_source_empty_data), .B(8'h00), .S(_set_flag_710), .Y(_26434_) );
  \$mux  #( .WIDTH(8) ) _49881_ ( .A(_26434_), .B(8'h00), .S(RST), .Y(_02520_) );
  \$mux  #( .WIDTH(1) ) _49882_ ( .A(_stream_conv2d_16_source_14_idle), .B(1'h1), .S(_stream_conv2d_16_start), .Y(_26435_) );
  \$mux  #( .WIDTH(1) ) _49883_ ( .A(_26435_), .B(1'h1), .S(RST), .Y(_02519_) );
  \$mux  #( .WIDTH(8) ) _49884_ ( .A(_stream_conv2d_16_source_12_source_empty_data), .B(8'h00), .S(_set_flag_710), .Y(_26436_) );
  \$mux  #( .WIDTH(8) ) _49885_ ( .A(_26436_), .B(8'h00), .S(RST), .Y(_02518_) );
  \$mux  #( .WIDTH(1) ) _49886_ ( .A(_stream_conv2d_16_source_12_idle), .B(1'h1), .S(_stream_conv2d_16_start), .Y(_26437_) );
  \$mux  #( .WIDTH(1) ) _49887_ ( .A(_26437_), .B(1'h1), .S(RST), .Y(_02517_) );
  \$mux  #( .WIDTH(8) ) _49888_ ( .A(_stream_conv2d_16_source_10_source_empty_data), .B(8'h00), .S(_set_flag_710), .Y(_26438_) );
  \$mux  #( .WIDTH(8) ) _49889_ ( .A(_26438_), .B(8'h00), .S(RST), .Y(_02516_) );
  \$mux  #( .WIDTH(1) ) _49890_ ( .A(_stream_conv2d_16_source_10_idle), .B(1'h1), .S(_stream_conv2d_16_start), .Y(_26439_) );
  \$mux  #( .WIDTH(1) ) _49891_ ( .A(_26439_), .B(1'h1), .S(RST), .Y(_02515_) );
  \$mux  #( .WIDTH(1) ) _49892_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id0_3_cond_2_1), .Y(_26440_) );
  \$mux  #( .WIDTH(1) ) _49893_ ( .A(_26440_), .B(1'h0), .S(RST), .Y(_02699_) );
  \$mux  #( .WIDTH(1) ) _49894_ ( .A(1'h1), .B(_stream_conv2d_16_source_8_source_ram_renable), .S(_05986_), .Y(_26441_) );
  \$mux  #( .WIDTH(1) ) _49895_ ( .A(1'h0), .B(_26441_), .S(_05985_), .Y(_26442_) );
  \$mux  #( .WIDTH(1) ) _49896_ ( .A(_26442_), .B(1'h0), .S(RST), .Y(_02698_) );
  \$mux  #( .WIDTH(32) ) _49897_ ( .A(_stream_conv2d_16_source_8_source_pat_all_offset), .B(_stream_conv2d_16_source_8_source_ram_raddr), .S(_05986_), .Y(_26443_) );
  \$mux  #( .WIDTH(32) ) _49898_ ( .A(_26443_), .B(0), .S(RST), .Y(_02697_) );
  \$mux  #( .WIDTH(8) ) _49899_ ( .A(_stream_conv2d_16_source_8_source_ram_sel), .B(8'h02), .S(_set_flag_710), .Y(_26444_) );
  \$mux  #( .WIDTH(8) ) _49900_ ( .A(_26444_), .B(8'h00), .S(RST), .Y(_02700_) );
  \$mux  #( .WIDTH(32) ) _49901_ ( .A(_stream_conv2d_16_source_8_source_offset_buf), .B(_stream_conv2d_16_source_8_source_offset), .S(_06691_), .Y(_26445_) );
  \$mux  #( .WIDTH(32) ) _49902_ ( .A(_26445_), .B(0), .S(RST), .Y(_02695_) );
  \$mux  #( .WIDTH(32) ) _49903_ ( .A(_stream_conv2d_16_source_8_source_offset), .B(0), .S(_set_flag_710), .Y(_26446_) );
  \$mux  #( .WIDTH(32) ) _49904_ ( .A(_26446_), .B(0), .S(RST), .Y(_02694_) );
  \$mux  #( .WIDTH(3) ) _49905_ ( .A(_stream_conv2d_16_source_8_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26447_) );
  \$mux  #( .WIDTH(3) ) _49906_ ( .A(_26447_), .B(3'h0), .S(RST), .Y(_02693_) );
  \$mux  #( .WIDTH(1) ) _49907_ ( .A(_stream_conv2d_16_source_8_idle), .B(1'h0), .S(_06691_), .Y(_26448_) );
  \$mux  #( .WIDTH(1) ) _49908_ ( .A(1'h1), .B(_26448_), .S(_05985_), .Y(_26449_) );
  \$mux  #( .WIDTH(1) ) _49909_ ( .A(_26449_), .B(1'h1), .S(RST), .Y(_02692_) );
  \$mux  #( .WIDTH(1) ) _49910_ ( .A(1'h0), .B(1'h1), .S(_ram_w8_l2048_id1_0_cond_2_1), .Y(_26450_) );
  \$mux  #( .WIDTH(1) ) _49911_ ( .A(_26450_), .B(1'h0), .S(RST), .Y(_02690_) );
  \$mux  #( .WIDTH(1) ) _49912_ ( .A(1'h1), .B(_stream_conv2d_16_source_6_source_ram_renable), .S(_05987_), .Y(_26451_) );
  \$mux  #( .WIDTH(1) ) _49913_ ( .A(1'h0), .B(_26451_), .S(_05988_), .Y(_26452_) );
  \$mux  #( .WIDTH(1) ) _49914_ ( .A(_26452_), .B(1'h0), .S(RST), .Y(_02689_) );
  \$mux  #( .WIDTH(32) ) _49915_ ( .A(_stream_conv2d_16_source_6_source_pat_all_offset), .B(_stream_conv2d_16_source_6_source_ram_raddr), .S(_05987_), .Y(_26453_) );
  \$mux  #( .WIDTH(32) ) _49916_ ( .A(_26453_), .B(0), .S(RST), .Y(_02688_) );
  \$mux  #( .WIDTH(8) ) _49917_ ( .A(_stream_conv2d_16_source_6_source_ram_sel), .B(8'h01), .S(_set_flag_710), .Y(_26454_) );
  \$mux  #( .WIDTH(8) ) _49918_ ( .A(_26454_), .B(8'h00), .S(RST), .Y(_02691_) );
  \$mux  #( .WIDTH(32) ) _49919_ ( .A(_stream_conv2d_16_source_6_source_offset_buf), .B(_stream_conv2d_16_source_6_source_offset), .S(_06686_), .Y(_26455_) );
  \$mux  #( .WIDTH(32) ) _49920_ ( .A(_26455_), .B(0), .S(RST), .Y(_02686_) );
  \$mux  #( .WIDTH(32) ) _49921_ ( .A(_stream_conv2d_16_source_6_source_offset), .B(_29231_), .S(_set_flag_710), .Y(_26456_) );
  \$mux  #( .WIDTH(32) ) _49922_ ( .A(_26456_), .B(0), .S(RST), .Y(_02685_) );
  \$mux  #( .WIDTH(3) ) _49923_ ( .A(_stream_conv2d_16_source_6_source_mode), .B(3'h2), .S(_set_flag_710), .Y(_26457_) );
  \$mux  #( .WIDTH(3) ) _49924_ ( .A(_26457_), .B(3'h0), .S(RST), .Y(_02684_) );
  \$mux  #( .WIDTH(1) ) _49925_ ( .A(_stream_conv2d_16_source_6_idle), .B(1'h0), .S(_06686_), .Y(_26458_) );
  \$mux  #( .WIDTH(1) ) _49926_ ( .A(1'h1), .B(_26458_), .S(_05988_), .Y(_26459_) );
  \$mux  #( .WIDTH(1) ) _49927_ ( .A(_26459_), .B(1'h1), .S(RST), .Y(_02683_) );
  \$mux  #( .WIDTH(9) ) _49928_ ( .A(_stream_conv2d_16_constant_3_next_constant_data), .B(conv2d_16_stream_pad_masks), .S(_set_flag_710), .Y(_26460_) );
  \$mux  #( .WIDTH(9) ) _49929_ ( .A(_26460_), .B(9'h000), .S(RST), .Y(_02501_) );
  \$mux  #( .WIDTH(2) ) _49930_ ( .A(_stream_conv2d_16_constant_2_next_constant_data), .B(conv2d_16_row_select_buf), .S(_set_flag_710), .Y(_26461_) );
  \$mux  #( .WIDTH(2) ) _49931_ ( .A(_26461_), .B(2'h0), .S(RST), .Y(_02500_) );
  \$mux  #( .WIDTH(2) ) _49932_ ( .A(_stream_conv2d_16_constant_1_next_constant_data), .B(conv2d_16_col_select), .S(_set_flag_710), .Y(_26462_) );
  \$mux  #( .WIDTH(2) ) _49933_ ( .A(_26462_), .B(2'h0), .S(RST), .Y(_02499_) );
  \$mux  #( .WIDTH(6) ) _49934_ ( .A(_stream_conv2d_16_constant_0_next_constant_data), .B(cparam_conv2d_16_stream_reduce_size), .S(_set_flag_710), .Y(_26463_) );
  \$mux  #( .WIDTH(6) ) _49935_ ( .A(_26463_), .B(6'h00), .S(RST), .Y(_02495_) );
  \$mux  #( .WIDTH(1) ) _49936_ ( .A(_substream__reduce_max_13_size_data_cond_792_43), .B(1'h1), .S(__tmp_1046_7), .Y(_26464_) );
  \$mux  #( .WIDTH(1) ) _49937_ ( .A(_26464_), .B(1'h0), .S(__tmp_1060_4), .Y(_26465_) );
  \$mux  #( .WIDTH(1) ) _49938_ ( .A(_26465_), .B(1'h0), .S(RST), .Y(_02798_) );
  \$mux  #( .WIDTH(1) ) _49939_ ( .A(_substream__reduce_max_13_x_data_cond_792_42), .B(1'h1), .S(__tmp_1046_7), .Y(_26466_) );
  \$mux  #( .WIDTH(1) ) _49940_ ( .A(_26466_), .B(1'h0), .S(__tmp_1060_4), .Y(_26467_) );
  \$mux  #( .WIDTH(1) ) _49941_ ( .A(_26467_), .B(1'h0), .S(RST), .Y(_02799_) );
  \$mux  #( .WIDTH(1) ) _49942_ ( .A(__reduce_max_13_reduce_reset), .B(1'h0), .S(__tmp_1042_9), .Y(_26468_) );
  \$mux  #( .WIDTH(1) ) _49943_ ( .A(_26468_), .B(1'h1), .S(__tmp_1060_5), .Y(_26469_) );
  \$mux  #( .WIDTH(1) ) _49944_ ( .A(_26469_), .B(1'h1), .S(RST), .Y(_00705_) );
  \$mux  #( .WIDTH(1) ) _49945_ ( .A(__tmp_1060_4), .B(1'h0), .S(RST), .Y(_01125_) );
  \$mux  #( .WIDTH(1) ) _49946_ ( .A(__tmp_1060_3), .B(1'h0), .S(RST), .Y(_01124_) );
  \$mux  #( .WIDTH(1) ) _49947_ ( .A(__tmp_1060_2), .B(1'h0), .S(RST), .Y(_01123_) );
  \$mux  #( .WIDTH(1) ) _49948_ ( .A(__tmp_1060_1), .B(1'h0), .S(RST), .Y(_01122_) );
  \$mux  #( .WIDTH(1) ) _49949_ ( .A(_tmp_1056), .B(1'h0), .S(RST), .Y(_01121_) );
  \$mux  #( .WIDTH(8) ) _49950_ ( .A(__variable_wdata_208), .B({ 5'h00, __delay_data_1416 }), .S(_substream__reduce_max_13_size_data_cond_792_43), .Y(_26470_) );
  \$mux  #( .WIDTH(8) ) _49951_ ( .A(_26470_), .B(8'h00), .S(RST), .Y(_01394_) );
  \$mux  #( .WIDTH(8) ) _49952_ ( .A(__variable_wdata_207), .B(_cond_data_791[7:0]), .S(_substream__reduce_max_13_x_data_cond_792_42), .Y(_26471_) );
  \$mux  #( .WIDTH(8) ) _49953_ ( .A(_26471_), .B(8'h00), .S(RST), .Y(_01393_) );
  \$mux  #( .WIDTH(9) ) _49954_ ( .A(_29166_[8:0]), .B(9'h000), .S(__reduce_max_13_reduce_reset), .Y(_26472_) );
  \$mux  #( .WIDTH(9) ) _49955_ ( .A(_26472_), .B(9'h000), .S(RST), .Y(_01821_) );
  \$mux  #( .WIDTH(1) ) _49956_ ( .A(_06151_), .B(1'h0), .S(RST), .Y(_01823_) );
  \$mux  #( .WIDTH(9) ) _49957_ ( .A(_29164_[8:0]), .B(9'h000), .S(__reduce_max_13_reduce_reset), .Y(_26473_) );
  \$mux  #( .WIDTH(9) ) _49958_ ( .A(_26473_), .B(9'h000), .S(RST), .Y(_01839_) );
  \$mux  #( .WIDTH(8) ) _49959_ ( .A(_29163_), .B(_29165_[7:0]), .S(__reduce_max_13_reduce_reset), .Y(_26474_) );
  \$mux  #( .WIDTH(8) ) _49960_ ( .A(_29165_[7:0]), .B(_26474_), .S(_05721_), .Y(_26475_) );
  \$mux  #( .WIDTH(8) ) _49961_ ( .A(_26475_), .B(8'h80), .S(RST), .Y(_01840_) );
  \$mux  #( .WIDTH(1) ) _49962_ ( .A(_substream_mul_12_rshift_data_cond_728_26), .B(1'h1), .S(__tmp_799_12), .Y(_26476_) );
  \$mux  #( .WIDTH(1) ) _49963_ ( .A(_26476_), .B(1'h0), .S(__tmp_947_9), .Y(_26477_) );
  \$mux  #( .WIDTH(1) ) _49964_ ( .A(_26477_), .B(1'h0), .S(RST), .Y(_02822_) );
  \$mux  #( .WIDTH(1) ) _49965_ ( .A(_substream_mul_12_y_data_cond_728_25), .B(1'h1), .S(__tmp_799_12), .Y(_26478_) );
  \$mux  #( .WIDTH(1) ) _49966_ ( .A(_26478_), .B(1'h0), .S(__tmp_947_9), .Y(_26479_) );
  \$mux  #( .WIDTH(1) ) _49967_ ( .A(_26479_), .B(1'h0), .S(RST), .Y(_02824_) );
  \$mux  #( .WIDTH(1) ) _49968_ ( .A(_substream_mul_12_x_data_cond_728_24), .B(1'h1), .S(__tmp_799_12), .Y(_26480_) );
  \$mux  #( .WIDTH(1) ) _49969_ ( .A(_26480_), .B(1'h0), .S(__tmp_947_9), .Y(_26481_) );
  \$mux  #( .WIDTH(1) ) _49970_ ( .A(_26481_), .B(1'h0), .S(RST), .Y(_02823_) );
  \$mux  #( .WIDTH(4) ) _49971_ ( .A(__variable_wdata_192), .B(__delay_data_1267[3:0]), .S(_substream_mul_12_rshift_data_cond_728_26), .Y(_26482_) );
  \$mux  #( .WIDTH(4) ) _49972_ ( .A(_26482_), .B(4'h0), .S(RST), .Y(_01391_) );
  \$mux  #( .WIDTH(4) ) _49973_ ( .A(__variable_wdata_191), .B(__delay_data_1261), .S(_substream_mul_12_y_data_cond_728_25), .Y(_26483_) );
  \$mux  #( .WIDTH(4) ) _49974_ ( .A(_26483_), .B(4'h0), .S(RST), .Y(_01390_) );
  \$mux  #( .WIDTH(8) ) _49975_ ( .A(__variable_wdata_190), .B(_cond_data_591), .S(_substream_mul_12_x_data_cond_728_24), .Y(_26484_) );
  \$mux  #( .WIDTH(8) ) _49976_ ( .A(_26484_), .B(8'h00), .S(RST), .Y(_01389_) );
  \$mux  #( .WIDTH(12) ) _49977_ ( .A(_28531_), .B(12'h000), .S(RST), .Y(_02490_) );
  \$mux  #( .WIDTH(4) ) _49978_ ( .A(__delay_data_741), .B(4'h0), .S(RST), .Y(_00609_) );
  \$mux  #( .WIDTH(4) ) _49979_ ( .A(__delay_data_740), .B(4'h0), .S(RST), .Y(_00608_) );
  \$mux  #( .WIDTH(4) ) _49980_ ( .A(__delay_data_739), .B(4'h0), .S(RST), .Y(_00607_) );
  \$mux  #( .WIDTH(4) ) _49981_ ( .A(__delay_data_738), .B(4'h0), .S(RST), .Y(_00606_) );
  \$mux  #( .WIDTH(12) ) _49982_ ( .A(\__muladd_madd_205.madd._pipe_madd1 ), .B(12'h000), .S(RST), .Y(_00698_) );
  \$mux  #( .WIDTH(4) ) _49983_ ( .A(__delay_data_737), .B(4'h0), .S(RST), .Y(_00605_) );
  \$mux  #( .WIDTH(4) ) _49984_ ( .A(__delay_data_734), .B(4'h0), .S(RST), .Y(_00602_) );
  \$mux  #( .WIDTH(8) ) _49985_ ( .A(__delay_data_731), .B(8'h00), .S(RST), .Y(_00599_) );
  \$mux  #( .WIDTH(12) ) _49986_ ( .A(_29162_[11:0]), .B(12'h000), .S(RST), .Y(_01474_) );
  \$mux  #( .WIDTH(4) ) _49987_ ( .A(__delay_data_736), .B(4'h0), .S(RST), .Y(_00604_) );
  \$mux  #( .WIDTH(4) ) _49988_ ( .A(__delay_data_733), .B(4'h0), .S(RST), .Y(_00601_) );
  \$mux  #( .WIDTH(8) ) _49989_ ( .A(__delay_data_730), .B(8'h00), .S(RST), .Y(_00598_) );
  \$mux  #( .WIDTH(1) ) _49990_ ( .A(_greaterthan_data_193), .B(1'h0), .S(RST), .Y(_00596_) );
  \$mux  #( .WIDTH(18) ) _49991_ ( .A(_28518_), .B(18'h00000), .S(RST), .Y(_01879_) );
  \$mux  #( .WIDTH(4) ) _49992_ ( .A(__variable_wdata_192), .B(4'h0), .S(RST), .Y(_00603_) );
  \$mux  #( .WIDTH(4) ) _49993_ ( .A(__variable_wdata_191), .B(4'h0), .S(RST), .Y(_00600_) );
  \$mux  #( .WIDTH(8) ) _49994_ ( .A(__variable_wdata_190), .B(8'h00), .S(RST), .Y(_00597_) );
  \$mux  #( .WIDTH(4) ) _49995_ ( .A(_28627_), .B(4'h0), .S(RST), .Y(_01805_) );
  \$mux  #( .WIDTH(1) ) _49996_ ( .A(_06173_), .B(1'h0), .S(RST), .Y(_01696_) );
  \$mux  #( .WIDTH(1) ) _49997_ ( .A(_substream_mul_11_rshift_data_cond_711_23), .B(1'h1), .S(__tmp_799_12), .Y(_26485_) );
  \$mux  #( .WIDTH(1) ) _49998_ ( .A(_26485_), .B(1'h0), .S(__tmp_947_9), .Y(_26486_) );
  \$mux  #( .WIDTH(1) ) _49999_ ( .A(_26486_), .B(1'h0), .S(RST), .Y(_02819_) );
  \$mux  #( .WIDTH(1) ) _50000_ ( .A(_substream_mul_11_y_data_cond_711_22), .B(1'h1), .S(__tmp_799_12), .Y(_26487_) );
  \$mux  #( .WIDTH(1) ) _50001_ ( .A(_26487_), .B(1'h0), .S(__tmp_947_9), .Y(_26488_) );
  \$mux  #( .WIDTH(1) ) _50002_ ( .A(_26488_), .B(1'h0), .S(RST), .Y(_02821_) );
  \$mux  #( .WIDTH(1) ) _50003_ ( .A(_substream_mul_11_x_data_cond_711_21), .B(1'h1), .S(__tmp_799_12), .Y(_26489_) );
  \$mux  #( .WIDTH(1) ) _50004_ ( .A(_26489_), .B(1'h0), .S(__tmp_947_9), .Y(_26490_) );
  \$mux  #( .WIDTH(1) ) _50005_ ( .A(_26490_), .B(1'h0), .S(RST), .Y(_02820_) );
  \$mux  #( .WIDTH(4) ) _50006_ ( .A(__variable_wdata_175), .B(__delay_data_1267[3:0]), .S(_substream_mul_11_rshift_data_cond_711_23), .Y(_26491_) );
  \$mux  #( .WIDTH(4) ) _50007_ ( .A(_26491_), .B(4'h0), .S(RST), .Y(_01388_) );
  \$mux  #( .WIDTH(4) ) _50008_ ( .A(__variable_wdata_174), .B(__delay_data_1227), .S(_substream_mul_11_y_data_cond_711_22), .Y(_26492_) );
  \$mux  #( .WIDTH(4) ) _50009_ ( .A(_26492_), .B(4'h0), .S(RST), .Y(_01387_) );
  \$mux  #( .WIDTH(8) ) _50010_ ( .A(__variable_wdata_173), .B(_cond_data_589), .S(_substream_mul_11_x_data_cond_711_21), .Y(_26493_) );
  \$mux  #( .WIDTH(8) ) _50011_ ( .A(_26493_), .B(8'h00), .S(RST), .Y(_01386_) );
  \$mux  #( .WIDTH(12) ) _50012_ ( .A(_28530_), .B(12'h000), .S(RST), .Y(_02489_) );
  \$mux  #( .WIDTH(4) ) _50013_ ( .A(__delay_data_724), .B(4'h0), .S(RST), .Y(_00595_) );
  \$mux  #( .WIDTH(4) ) _50014_ ( .A(__delay_data_723), .B(4'h0), .S(RST), .Y(_00594_) );
  \$mux  #( .WIDTH(4) ) _50015_ ( .A(__delay_data_722), .B(4'h0), .S(RST), .Y(_00593_) );
  \$mux  #( .WIDTH(4) ) _50016_ ( .A(__delay_data_721), .B(4'h0), .S(RST), .Y(_00592_) );
  \$mux  #( .WIDTH(12) ) _50017_ ( .A(\__muladd_madd_188.madd._pipe_madd1 ), .B(12'h000), .S(RST), .Y(_00697_) );
  \$mux  #( .WIDTH(4) ) _50018_ ( .A(__delay_data_720), .B(4'h0), .S(RST), .Y(_00591_) );
  \$mux  #( .WIDTH(4) ) _50019_ ( .A(__delay_data_717), .B(4'h0), .S(RST), .Y(_00588_) );
  \$mux  #( .WIDTH(8) ) _50020_ ( .A(__delay_data_714), .B(8'h00), .S(RST), .Y(_00585_) );
  \$mux  #( .WIDTH(12) ) _50021_ ( .A(_29161_[11:0]), .B(12'h000), .S(RST), .Y(_01473_) );
  \$mux  #( .WIDTH(4) ) _50022_ ( .A(__delay_data_719), .B(4'h0), .S(RST), .Y(_00590_) );
  \$mux  #( .WIDTH(4) ) _50023_ ( .A(__delay_data_716), .B(4'h0), .S(RST), .Y(_00587_) );
  \$mux  #( .WIDTH(8) ) _50024_ ( .A(__delay_data_713), .B(8'h00), .S(RST), .Y(_00584_) );
  \$mux  #( .WIDTH(1) ) _50025_ ( .A(_greaterthan_data_176), .B(1'h0), .S(RST), .Y(_00582_) );
  \$mux  #( .WIDTH(18) ) _50026_ ( .A(_28517_), .B(18'h00000), .S(RST), .Y(_01878_) );
  \$mux  #( .WIDTH(4) ) _50027_ ( .A(__variable_wdata_175), .B(4'h0), .S(RST), .Y(_00589_) );
  \$mux  #( .WIDTH(4) ) _50028_ ( .A(__variable_wdata_174), .B(4'h0), .S(RST), .Y(_00586_) );
  \$mux  #( .WIDTH(8) ) _50029_ ( .A(__variable_wdata_173), .B(8'h00), .S(RST), .Y(_00583_) );
  \$mux  #( .WIDTH(4) ) _50030_ ( .A(_28626_), .B(4'h0), .S(RST), .Y(_01804_) );
  \$mux  #( .WIDTH(1) ) _50031_ ( .A(_06172_), .B(1'h0), .S(RST), .Y(_01695_) );
  \$mux  #( .WIDTH(1) ) _50032_ ( .A(_substream_mul_10_rshift_data_cond_694_20), .B(1'h1), .S(__tmp_799_12), .Y(_26494_) );
  \$mux  #( .WIDTH(1) ) _50033_ ( .A(_26494_), .B(1'h0), .S(__tmp_947_9), .Y(_26495_) );
  \$mux  #( .WIDTH(1) ) _50034_ ( .A(_26495_), .B(1'h0), .S(RST), .Y(_02816_) );
  \$mux  #( .WIDTH(1) ) _50035_ ( .A(_substream_mul_10_y_data_cond_694_19), .B(1'h1), .S(__tmp_799_12), .Y(_26496_) );
  \$mux  #( .WIDTH(1) ) _50036_ ( .A(_26496_), .B(1'h0), .S(__tmp_947_9), .Y(_26497_) );
  \$mux  #( .WIDTH(1) ) _50037_ ( .A(_26497_), .B(1'h0), .S(RST), .Y(_02818_) );
  \$mux  #( .WIDTH(1) ) _50038_ ( .A(_substream_mul_10_x_data_cond_694_18), .B(1'h1), .S(__tmp_799_12), .Y(_26498_) );
  \$mux  #( .WIDTH(1) ) _50039_ ( .A(_26498_), .B(1'h0), .S(__tmp_947_9), .Y(_26499_) );
  \$mux  #( .WIDTH(1) ) _50040_ ( .A(_26499_), .B(1'h0), .S(RST), .Y(_02817_) );
  \$mux  #( .WIDTH(4) ) _50041_ ( .A(__variable_wdata_158), .B(__delay_data_1267[3:0]), .S(_substream_mul_10_rshift_data_cond_694_20), .Y(_26500_) );
  \$mux  #( .WIDTH(4) ) _50042_ ( .A(_26500_), .B(4'h0), .S(RST), .Y(_01385_) );
  \$mux  #( .WIDTH(4) ) _50043_ ( .A(__variable_wdata_157), .B(__delay_data_1193), .S(_substream_mul_10_y_data_cond_694_19), .Y(_26501_) );
  \$mux  #( .WIDTH(4) ) _50044_ ( .A(_26501_), .B(4'h0), .S(RST), .Y(_01384_) );
  \$mux  #( .WIDTH(8) ) _50045_ ( .A(__variable_wdata_156), .B(_cond_data_587), .S(_substream_mul_10_x_data_cond_694_18), .Y(_26502_) );
  \$mux  #( .WIDTH(8) ) _50046_ ( .A(_26502_), .B(8'h00), .S(RST), .Y(_01383_) );
  \$mux  #( .WIDTH(12) ) _50047_ ( .A(_28529_), .B(12'h000), .S(RST), .Y(_02488_) );
  \$mux  #( .WIDTH(4) ) _50048_ ( .A(__delay_data_707), .B(4'h0), .S(RST), .Y(_00581_) );
  \$mux  #( .WIDTH(4) ) _50049_ ( .A(__delay_data_706), .B(4'h0), .S(RST), .Y(_00580_) );
  \$mux  #( .WIDTH(4) ) _50050_ ( .A(__delay_data_705), .B(4'h0), .S(RST), .Y(_00579_) );
  \$mux  #( .WIDTH(4) ) _50051_ ( .A(__delay_data_704), .B(4'h0), .S(RST), .Y(_00578_) );
  \$mux  #( .WIDTH(12) ) _50052_ ( .A(\__muladd_madd_171.madd._pipe_madd1 ), .B(12'h000), .S(RST), .Y(_00696_) );
  \$mux  #( .WIDTH(4) ) _50053_ ( .A(__delay_data_703), .B(4'h0), .S(RST), .Y(_00577_) );
  \$mux  #( .WIDTH(4) ) _50054_ ( .A(__delay_data_700), .B(4'h0), .S(RST), .Y(_00574_) );
  \$mux  #( .WIDTH(8) ) _50055_ ( .A(__delay_data_697), .B(8'h00), .S(RST), .Y(_00571_) );
  \$mux  #( .WIDTH(12) ) _50056_ ( .A(_29160_[11:0]), .B(12'h000), .S(RST), .Y(_01472_) );
  \$mux  #( .WIDTH(4) ) _50057_ ( .A(__delay_data_702), .B(4'h0), .S(RST), .Y(_00576_) );
  \$mux  #( .WIDTH(4) ) _50058_ ( .A(__delay_data_699), .B(4'h0), .S(RST), .Y(_00573_) );
  \$mux  #( .WIDTH(8) ) _50059_ ( .A(__delay_data_696), .B(8'h00), .S(RST), .Y(_00570_) );
  \$mux  #( .WIDTH(1) ) _50060_ ( .A(_greaterthan_data_159), .B(1'h0), .S(RST), .Y(_00568_) );
  \$mux  #( .WIDTH(18) ) _50061_ ( .A(_28516_), .B(18'h00000), .S(RST), .Y(_01877_) );
  \$mux  #( .WIDTH(4) ) _50062_ ( .A(__variable_wdata_158), .B(4'h0), .S(RST), .Y(_00575_) );
  \$mux  #( .WIDTH(4) ) _50063_ ( .A(__variable_wdata_157), .B(4'h0), .S(RST), .Y(_00572_) );
  \$mux  #( .WIDTH(8) ) _50064_ ( .A(__variable_wdata_156), .B(8'h00), .S(RST), .Y(_00569_) );
  \$mux  #( .WIDTH(4) ) _50065_ ( .A(_28625_), .B(4'h0), .S(RST), .Y(_01803_) );
  \$mux  #( .WIDTH(1) ) _50066_ ( .A(_06171_), .B(1'h0), .S(RST), .Y(_01694_) );
  \$mux  #( .WIDTH(1) ) _50067_ ( .A(_substream_mul_9_rshift_data_cond_677_17), .B(1'h1), .S(__tmp_799_12), .Y(_26503_) );
  \$mux  #( .WIDTH(1) ) _50068_ ( .A(_26503_), .B(1'h0), .S(__tmp_947_9), .Y(_26504_) );
  \$mux  #( .WIDTH(1) ) _50069_ ( .A(_26504_), .B(1'h0), .S(RST), .Y(_02843_) );
  \$mux  #( .WIDTH(1) ) _50070_ ( .A(_substream_mul_9_y_data_cond_677_16), .B(1'h1), .S(__tmp_799_12), .Y(_26505_) );
  \$mux  #( .WIDTH(1) ) _50071_ ( .A(_26505_), .B(1'h0), .S(__tmp_947_9), .Y(_26506_) );
  \$mux  #( .WIDTH(1) ) _50072_ ( .A(_26506_), .B(1'h0), .S(RST), .Y(_02845_) );
  \$mux  #( .WIDTH(1) ) _50073_ ( .A(_substream_mul_9_x_data_cond_677_15), .B(1'h1), .S(__tmp_799_12), .Y(_26507_) );
  \$mux  #( .WIDTH(1) ) _50074_ ( .A(_26507_), .B(1'h0), .S(__tmp_947_9), .Y(_26508_) );
  \$mux  #( .WIDTH(1) ) _50075_ ( .A(_26508_), .B(1'h0), .S(RST), .Y(_02844_) );
  \$mux  #( .WIDTH(1) ) _50076_ ( .A(__tmp_959_11), .B(1'h0), .S(RST), .Y(_01334_) );
  \$mux  #( .WIDTH(1) ) _50077_ ( .A(__tmp_959_10), .B(1'h0), .S(RST), .Y(_01333_) );
  \$mux  #( .WIDTH(1) ) _50078_ ( .A(__tmp_947_9), .B(1'h0), .S(RST), .Y(_01332_) );
  \$mux  #( .WIDTH(1) ) _50079_ ( .A(__tmp_947_8), .B(1'h0), .S(RST), .Y(_01331_) );
  \$mux  #( .WIDTH(1) ) _50080_ ( .A(__tmp_947_7), .B(1'h0), .S(RST), .Y(_01330_) );
  \$mux  #( .WIDTH(1) ) _50081_ ( .A(__tmp_947_5), .B(1'h0), .S(RST), .Y(_01328_) );
  \$mux  #( .WIDTH(4) ) _50082_ ( .A(__variable_wdata_141), .B(__delay_data_1267[3:0]), .S(_substream_mul_9_rshift_data_cond_677_17), .Y(_26509_) );
  \$mux  #( .WIDTH(4) ) _50083_ ( .A(_26509_), .B(4'h0), .S(RST), .Y(_01382_) );
  \$mux  #( .WIDTH(4) ) _50084_ ( .A(__variable_wdata_140), .B(__delay_data_1159), .S(_substream_mul_9_y_data_cond_677_16), .Y(_26510_) );
  \$mux  #( .WIDTH(4) ) _50085_ ( .A(_26510_), .B(4'h0), .S(RST), .Y(_01381_) );
  \$mux  #( .WIDTH(8) ) _50086_ ( .A(__variable_wdata_139), .B(_cond_data_585), .S(_substream_mul_9_x_data_cond_677_15), .Y(_26511_) );
  \$mux  #( .WIDTH(8) ) _50087_ ( .A(_26511_), .B(8'h00), .S(RST), .Y(_01380_) );
  \$mux  #( .WIDTH(12) ) _50088_ ( .A(_28528_), .B(12'h000), .S(RST), .Y(_02487_) );
  \$mux  #( .WIDTH(4) ) _50089_ ( .A(__delay_data_690), .B(4'h0), .S(RST), .Y(_00567_) );
  \$mux  #( .WIDTH(4) ) _50090_ ( .A(__delay_data_689), .B(4'h0), .S(RST), .Y(_00566_) );
  \$mux  #( .WIDTH(4) ) _50091_ ( .A(__delay_data_688), .B(4'h0), .S(RST), .Y(_00565_) );
  \$mux  #( .WIDTH(4) ) _50092_ ( .A(__delay_data_687), .B(4'h0), .S(RST), .Y(_00564_) );
  \$mux  #( .WIDTH(12) ) _50093_ ( .A(\__muladd_madd_154.madd._pipe_madd1 ), .B(12'h000), .S(RST), .Y(_00695_) );
  \$mux  #( .WIDTH(4) ) _50094_ ( .A(__delay_data_686), .B(4'h0), .S(RST), .Y(_00563_) );
  \$mux  #( .WIDTH(4) ) _50095_ ( .A(__delay_data_683), .B(4'h0), .S(RST), .Y(_00560_) );
  \$mux  #( .WIDTH(8) ) _50096_ ( .A(__delay_data_680), .B(8'h00), .S(RST), .Y(_00557_) );
  \$mux  #( .WIDTH(12) ) _50097_ ( .A(_29159_[11:0]), .B(12'h000), .S(RST), .Y(_01471_) );
  \$mux  #( .WIDTH(4) ) _50098_ ( .A(__delay_data_685), .B(4'h0), .S(RST), .Y(_00562_) );
  \$mux  #( .WIDTH(4) ) _50099_ ( .A(__delay_data_682), .B(4'h0), .S(RST), .Y(_00559_) );
  \$mux  #( .WIDTH(8) ) _50100_ ( .A(__delay_data_679), .B(8'h00), .S(RST), .Y(_00556_) );
  \$mux  #( .WIDTH(1) ) _50101_ ( .A(_greaterthan_data_142), .B(1'h0), .S(RST), .Y(_00554_) );
  \$mux  #( .WIDTH(18) ) _50102_ ( .A(_28515_), .B(18'h00000), .S(RST), .Y(_01876_) );
  \$mux  #( .WIDTH(4) ) _50103_ ( .A(__variable_wdata_141), .B(4'h0), .S(RST), .Y(_00561_) );
  \$mux  #( .WIDTH(4) ) _50104_ ( .A(__variable_wdata_140), .B(4'h0), .S(RST), .Y(_00558_) );
  \$mux  #( .WIDTH(8) ) _50105_ ( .A(__variable_wdata_139), .B(8'h00), .S(RST), .Y(_00555_) );
  \$mux  #( .WIDTH(4) ) _50106_ ( .A(_28624_), .B(4'h0), .S(RST), .Y(_01802_) );
  \$mux  #( .WIDTH(1) ) _50107_ ( .A(_06170_), .B(1'h0), .S(RST), .Y(_01693_) );
  \$mux  #( .WIDTH(1) ) _50108_ ( .A(_substream_mul_8_rshift_data_cond_660_14), .B(1'h1), .S(__tmp_799_12), .Y(_26512_) );
  \$mux  #( .WIDTH(1) ) _50109_ ( .A(_26512_), .B(1'h0), .S(__tmp_947_9), .Y(_26513_) );
  \$mux  #( .WIDTH(1) ) _50110_ ( .A(_26513_), .B(1'h0), .S(RST), .Y(_02840_) );
  \$mux  #( .WIDTH(1) ) _50111_ ( .A(_substream_mul_8_y_data_cond_660_13), .B(1'h1), .S(__tmp_799_12), .Y(_26514_) );
  \$mux  #( .WIDTH(1) ) _50112_ ( .A(_26514_), .B(1'h0), .S(__tmp_947_9), .Y(_26515_) );
  \$mux  #( .WIDTH(1) ) _50113_ ( .A(_26515_), .B(1'h0), .S(RST), .Y(_02842_) );
  \$mux  #( .WIDTH(1) ) _50114_ ( .A(_substream_mul_8_x_data_cond_660_12), .B(1'h1), .S(__tmp_799_12), .Y(_26516_) );
  \$mux  #( .WIDTH(1) ) _50115_ ( .A(_26516_), .B(1'h0), .S(__tmp_947_9), .Y(_26517_) );
  \$mux  #( .WIDTH(1) ) _50116_ ( .A(_26517_), .B(1'h0), .S(RST), .Y(_02841_) );
  \$mux  #( .WIDTH(4) ) _50117_ ( .A(__variable_wdata_124), .B(__delay_data_1267[3:0]), .S(_substream_mul_8_rshift_data_cond_660_14), .Y(_26518_) );
  \$mux  #( .WIDTH(4) ) _50118_ ( .A(_26518_), .B(4'h0), .S(RST), .Y(_01379_) );
  \$mux  #( .WIDTH(4) ) _50119_ ( .A(__variable_wdata_123), .B(__delay_data_1124), .S(_substream_mul_8_y_data_cond_660_13), .Y(_26519_) );
  \$mux  #( .WIDTH(4) ) _50120_ ( .A(_26519_), .B(4'h0), .S(RST), .Y(_01378_) );
  \$mux  #( .WIDTH(8) ) _50121_ ( .A(__variable_wdata_122), .B(_cond_data_583), .S(_substream_mul_8_x_data_cond_660_12), .Y(_26520_) );
  \$mux  #( .WIDTH(8) ) _50122_ ( .A(_26520_), .B(8'h00), .S(RST), .Y(_01377_) );
  \$mux  #( .WIDTH(12) ) _50123_ ( .A(_28527_), .B(12'h000), .S(RST), .Y(_02486_) );
  \$mux  #( .WIDTH(4) ) _50124_ ( .A(__delay_data_673), .B(4'h0), .S(RST), .Y(_00553_) );
  \$mux  #( .WIDTH(4) ) _50125_ ( .A(__delay_data_672), .B(4'h0), .S(RST), .Y(_00552_) );
  \$mux  #( .WIDTH(4) ) _50126_ ( .A(__delay_data_671), .B(4'h0), .S(RST), .Y(_00551_) );
  \$mux  #( .WIDTH(4) ) _50127_ ( .A(__delay_data_670), .B(4'h0), .S(RST), .Y(_00550_) );
  \$mux  #( .WIDTH(12) ) _50128_ ( .A(\__muladd_madd_137.madd._pipe_madd1 ), .B(12'h000), .S(RST), .Y(_00694_) );
  \$mux  #( .WIDTH(4) ) _50129_ ( .A(__delay_data_669), .B(4'h0), .S(RST), .Y(_00549_) );
  \$mux  #( .WIDTH(4) ) _50130_ ( .A(__delay_data_666), .B(4'h0), .S(RST), .Y(_00546_) );
  \$mux  #( .WIDTH(8) ) _50131_ ( .A(__delay_data_663), .B(8'h00), .S(RST), .Y(_00543_) );
  \$mux  #( .WIDTH(12) ) _50132_ ( .A(_29158_[11:0]), .B(12'h000), .S(RST), .Y(_01469_) );
  \$mux  #( .WIDTH(4) ) _50133_ ( .A(__delay_data_668), .B(4'h0), .S(RST), .Y(_00548_) );
  \$mux  #( .WIDTH(4) ) _50134_ ( .A(__delay_data_665), .B(4'h0), .S(RST), .Y(_00545_) );
  \$mux  #( .WIDTH(8) ) _50135_ ( .A(__delay_data_662), .B(8'h00), .S(RST), .Y(_00542_) );
  \$mux  #( .WIDTH(1) ) _50136_ ( .A(_greaterthan_data_125), .B(1'h0), .S(RST), .Y(_00540_) );
  \$mux  #( .WIDTH(18) ) _50137_ ( .A(_28514_), .B(18'h00000), .S(RST), .Y(_01875_) );
  \$mux  #( .WIDTH(4) ) _50138_ ( .A(__variable_wdata_124), .B(4'h0), .S(RST), .Y(_00547_) );
  \$mux  #( .WIDTH(4) ) _50139_ ( .A(__variable_wdata_123), .B(4'h0), .S(RST), .Y(_00544_) );
  \$mux  #( .WIDTH(8) ) _50140_ ( .A(__variable_wdata_122), .B(8'h00), .S(RST), .Y(_00541_) );
  \$mux  #( .WIDTH(4) ) _50141_ ( .A(_28623_), .B(4'h0), .S(RST), .Y(_01801_) );
  \$mux  #( .WIDTH(1) ) _50142_ ( .A(_06169_), .B(1'h0), .S(RST), .Y(_01692_) );
  \$mux  #( .WIDTH(1) ) _50143_ ( .A(_substream_mul_7_rshift_data_cond_643_11), .B(1'h1), .S(__tmp_799_12), .Y(_26521_) );
  \$mux  #( .WIDTH(1) ) _50144_ ( .A(_26521_), .B(1'h0), .S(__tmp_947_9), .Y(_26522_) );
  \$mux  #( .WIDTH(1) ) _50145_ ( .A(_26522_), .B(1'h0), .S(RST), .Y(_02837_) );
  \$mux  #( .WIDTH(1) ) _50146_ ( .A(_substream_mul_7_y_data_cond_643_10), .B(1'h1), .S(__tmp_799_12), .Y(_26523_) );
  \$mux  #( .WIDTH(1) ) _50147_ ( .A(_26523_), .B(1'h0), .S(__tmp_947_9), .Y(_26524_) );
  \$mux  #( .WIDTH(1) ) _50148_ ( .A(_26524_), .B(1'h0), .S(RST), .Y(_02839_) );
  \$mux  #( .WIDTH(1) ) _50149_ ( .A(_substream_mul_7_x_data_cond_643_9), .B(1'h1), .S(__tmp_799_12), .Y(_26525_) );
  \$mux  #( .WIDTH(1) ) _50150_ ( .A(_26525_), .B(1'h0), .S(__tmp_947_9), .Y(_26526_) );
  \$mux  #( .WIDTH(1) ) _50151_ ( .A(_26526_), .B(1'h0), .S(RST), .Y(_02838_) );
  \$mux  #( .WIDTH(4) ) _50152_ ( .A(__variable_wdata_107), .B(__delay_data_1267[3:0]), .S(_substream_mul_7_rshift_data_cond_643_11), .Y(_26527_) );
  \$mux  #( .WIDTH(4) ) _50153_ ( .A(_26527_), .B(4'h0), .S(RST), .Y(_01376_) );
  \$mux  #( .WIDTH(4) ) _50154_ ( .A(__variable_wdata_106), .B(__delay_data_1089), .S(_substream_mul_7_y_data_cond_643_10), .Y(_26528_) );
  \$mux  #( .WIDTH(4) ) _50155_ ( .A(_26528_), .B(4'h0), .S(RST), .Y(_01375_) );
  \$mux  #( .WIDTH(8) ) _50156_ ( .A(__variable_wdata_105), .B(_cond_data_581), .S(_substream_mul_7_x_data_cond_643_9), .Y(_26529_) );
  \$mux  #( .WIDTH(8) ) _50157_ ( .A(_26529_), .B(8'h00), .S(RST), .Y(_01374_) );
  \$mux  #( .WIDTH(12) ) _50158_ ( .A(_28526_), .B(12'h000), .S(RST), .Y(_02485_) );
  \$mux  #( .WIDTH(4) ) _50159_ ( .A(__delay_data_656), .B(4'h0), .S(RST), .Y(_00539_) );
  \$mux  #( .WIDTH(4) ) _50160_ ( .A(__delay_data_655), .B(4'h0), .S(RST), .Y(_00538_) );
  \$mux  #( .WIDTH(4) ) _50161_ ( .A(__delay_data_654), .B(4'h0), .S(RST), .Y(_00537_) );
  \$mux  #( .WIDTH(4) ) _50162_ ( .A(__delay_data_653), .B(4'h0), .S(RST), .Y(_00536_) );
  \$mux  #( .WIDTH(12) ) _50163_ ( .A(\__muladd_madd_120.madd._pipe_madd1 ), .B(12'h000), .S(RST), .Y(_00693_) );
  \$mux  #( .WIDTH(4) ) _50164_ ( .A(__delay_data_652), .B(4'h0), .S(RST), .Y(_00535_) );
  \$mux  #( .WIDTH(4) ) _50165_ ( .A(__delay_data_649), .B(4'h0), .S(RST), .Y(_00532_) );
  \$mux  #( .WIDTH(8) ) _50166_ ( .A(__delay_data_646), .B(8'h00), .S(RST), .Y(_00529_) );
  \$mux  #( .WIDTH(12) ) _50167_ ( .A(_29157_[11:0]), .B(12'h000), .S(RST), .Y(_01468_) );
  \$mux  #( .WIDTH(4) ) _50168_ ( .A(__delay_data_651), .B(4'h0), .S(RST), .Y(_00534_) );
  \$mux  #( .WIDTH(4) ) _50169_ ( .A(__delay_data_648), .B(4'h0), .S(RST), .Y(_00531_) );
  \$mux  #( .WIDTH(8) ) _50170_ ( .A(__delay_data_645), .B(8'h00), .S(RST), .Y(_00528_) );
  \$mux  #( .WIDTH(1) ) _50171_ ( .A(_greaterthan_data_108), .B(1'h0), .S(RST), .Y(_00526_) );
  \$mux  #( .WIDTH(18) ) _50172_ ( .A(_28513_), .B(18'h00000), .S(RST), .Y(_01874_) );
  \$mux  #( .WIDTH(4) ) _50173_ ( .A(__variable_wdata_107), .B(4'h0), .S(RST), .Y(_00533_) );
  \$mux  #( .WIDTH(4) ) _50174_ ( .A(__variable_wdata_106), .B(4'h0), .S(RST), .Y(_00530_) );
  \$mux  #( .WIDTH(8) ) _50175_ ( .A(__variable_wdata_105), .B(8'h00), .S(RST), .Y(_00527_) );
  \$mux  #( .WIDTH(4) ) _50176_ ( .A(_28622_), .B(4'h0), .S(RST), .Y(_01800_) );
  \$mux  #( .WIDTH(1) ) _50177_ ( .A(_06168_), .B(1'h0), .S(RST), .Y(_01691_) );
  \$mux  #( .WIDTH(1) ) _50178_ ( .A(_substream_mul_6_rshift_data_cond_626_8), .B(1'h1), .S(__tmp_799_12), .Y(_26530_) );
  \$mux  #( .WIDTH(1) ) _50179_ ( .A(_26530_), .B(1'h0), .S(__tmp_947_9), .Y(_26531_) );
  \$mux  #( .WIDTH(1) ) _50180_ ( .A(_26531_), .B(1'h0), .S(RST), .Y(_02834_) );
  \$mux  #( .WIDTH(1) ) _50181_ ( .A(_substream_mul_6_y_data_cond_626_7), .B(1'h1), .S(__tmp_799_12), .Y(_26532_) );
  \$mux  #( .WIDTH(1) ) _50182_ ( .A(_26532_), .B(1'h0), .S(__tmp_947_9), .Y(_26533_) );
  \$mux  #( .WIDTH(1) ) _50183_ ( .A(_26533_), .B(1'h0), .S(RST), .Y(_02836_) );
  \$mux  #( .WIDTH(1) ) _50184_ ( .A(_substream_mul_6_x_data_cond_626_6), .B(1'h1), .S(__tmp_799_12), .Y(_26534_) );
  \$mux  #( .WIDTH(1) ) _50185_ ( .A(_26534_), .B(1'h0), .S(__tmp_947_9), .Y(_26535_) );
  \$mux  #( .WIDTH(1) ) _50186_ ( .A(_26535_), .B(1'h0), .S(RST), .Y(_02835_) );
  \$mux  #( .WIDTH(4) ) _50187_ ( .A(__variable_wdata_90), .B(__delay_data_1267[3:0]), .S(_substream_mul_6_rshift_data_cond_626_8), .Y(_26536_) );
  \$mux  #( .WIDTH(4) ) _50188_ ( .A(_26536_), .B(4'h0), .S(RST), .Y(_01465_) );
  \$mux  #( .WIDTH(4) ) _50189_ ( .A(__variable_wdata_89), .B(__delay_data_1054), .S(_substream_mul_6_y_data_cond_626_7), .Y(_26537_) );
  \$mux  #( .WIDTH(4) ) _50190_ ( .A(_26537_), .B(4'h0), .S(RST), .Y(_01464_) );
  \$mux  #( .WIDTH(8) ) _50191_ ( .A(__variable_wdata_88), .B(_cond_data_579), .S(_substream_mul_6_x_data_cond_626_6), .Y(_26538_) );
  \$mux  #( .WIDTH(8) ) _50192_ ( .A(_26538_), .B(8'h00), .S(RST), .Y(_01463_) );
  \$mux  #( .WIDTH(12) ) _50193_ ( .A(_28525_), .B(12'h000), .S(RST), .Y(_02484_) );
  \$mux  #( .WIDTH(4) ) _50194_ ( .A(__delay_data_639), .B(4'h0), .S(RST), .Y(_00525_) );
  \$mux  #( .WIDTH(4) ) _50195_ ( .A(__delay_data_638), .B(4'h0), .S(RST), .Y(_00524_) );
  \$mux  #( .WIDTH(4) ) _50196_ ( .A(__delay_data_637), .B(4'h0), .S(RST), .Y(_00523_) );
  \$mux  #( .WIDTH(4) ) _50197_ ( .A(__delay_data_636), .B(4'h0), .S(RST), .Y(_00522_) );
  \$mux  #( .WIDTH(12) ) _50198_ ( .A(\__muladd_madd_103.madd._pipe_madd1 ), .B(12'h000), .S(RST), .Y(_00692_) );
  \$mux  #( .WIDTH(4) ) _50199_ ( .A(__delay_data_635), .B(4'h0), .S(RST), .Y(_00521_) );
  \$mux  #( .WIDTH(4) ) _50200_ ( .A(__delay_data_632), .B(4'h0), .S(RST), .Y(_00518_) );
  \$mux  #( .WIDTH(8) ) _50201_ ( .A(__delay_data_629), .B(8'h00), .S(RST), .Y(_00515_) );
  \$mux  #( .WIDTH(12) ) _50202_ ( .A(_29156_[11:0]), .B(12'h000), .S(RST), .Y(_01467_) );
  \$mux  #( .WIDTH(4) ) _50203_ ( .A(__delay_data_634), .B(4'h0), .S(RST), .Y(_00520_) );
  \$mux  #( .WIDTH(4) ) _50204_ ( .A(__delay_data_631), .B(4'h0), .S(RST), .Y(_00517_) );
  \$mux  #( .WIDTH(8) ) _50205_ ( .A(__delay_data_628), .B(8'h00), .S(RST), .Y(_00514_) );
  \$mux  #( .WIDTH(1) ) _50206_ ( .A(_greaterthan_data_91), .B(1'h0), .S(RST), .Y(_00512_) );
  \$mux  #( .WIDTH(18) ) _50207_ ( .A(_28512_), .B(18'h00000), .S(RST), .Y(_01883_) );
  \$mux  #( .WIDTH(4) ) _50208_ ( .A(__variable_wdata_90), .B(4'h0), .S(RST), .Y(_00519_) );
  \$mux  #( .WIDTH(4) ) _50209_ ( .A(__variable_wdata_89), .B(4'h0), .S(RST), .Y(_00516_) );
  \$mux  #( .WIDTH(8) ) _50210_ ( .A(__variable_wdata_88), .B(8'h00), .S(RST), .Y(_00513_) );
  \$mux  #( .WIDTH(4) ) _50211_ ( .A(_28621_), .B(4'h0), .S(RST), .Y(_01809_) );
  \$mux  #( .WIDTH(1) ) _50212_ ( .A(_06167_), .B(1'h0), .S(RST), .Y(_01702_) );
  \$mux  #( .WIDTH(1) ) _50213_ ( .A(_substream_mul_5_rshift_data_cond_609_5), .B(1'h1), .S(__tmp_799_12), .Y(_26539_) );
  \$mux  #( .WIDTH(1) ) _50214_ ( .A(_26539_), .B(1'h0), .S(__tmp_947_9), .Y(_26540_) );
  \$mux  #( .WIDTH(1) ) _50215_ ( .A(_26540_), .B(1'h0), .S(RST), .Y(_02831_) );
  \$mux  #( .WIDTH(1) ) _50216_ ( .A(_substream_mul_5_y_data_cond_609_4), .B(1'h1), .S(__tmp_799_12), .Y(_26541_) );
  \$mux  #( .WIDTH(1) ) _50217_ ( .A(_26541_), .B(1'h0), .S(__tmp_947_9), .Y(_26542_) );
  \$mux  #( .WIDTH(1) ) _50218_ ( .A(_26542_), .B(1'h0), .S(RST), .Y(_02833_) );
  \$mux  #( .WIDTH(1) ) _50219_ ( .A(_substream_mul_5_x_data_cond_609_3), .B(1'h1), .S(__tmp_799_12), .Y(_26543_) );
  \$mux  #( .WIDTH(1) ) _50220_ ( .A(_26543_), .B(1'h0), .S(__tmp_947_9), .Y(_26544_) );
  \$mux  #( .WIDTH(1) ) _50221_ ( .A(_26544_), .B(1'h0), .S(RST), .Y(_02832_) );
  \$mux  #( .WIDTH(4) ) _50222_ ( .A(__variable_wdata_73), .B(__delay_data_1267[3:0]), .S(_substream_mul_5_rshift_data_cond_609_5), .Y(_26545_) );
  \$mux  #( .WIDTH(4) ) _50223_ ( .A(_26545_), .B(4'h0), .S(RST), .Y(_01444_) );
  \$mux  #( .WIDTH(4) ) _50224_ ( .A(__variable_wdata_72), .B(__delay_data_1006), .S(_substream_mul_5_y_data_cond_609_4), .Y(_26546_) );
  \$mux  #( .WIDTH(4) ) _50225_ ( .A(_26546_), .B(4'h0), .S(RST), .Y(_01443_) );
  \$mux  #( .WIDTH(8) ) _50226_ ( .A(__variable_wdata_71), .B(_cond_data_577), .S(_substream_mul_5_x_data_cond_609_3), .Y(_26547_) );
  \$mux  #( .WIDTH(8) ) _50227_ ( .A(_26547_), .B(8'h00), .S(RST), .Y(_01442_) );
  \$mux  #( .WIDTH(12) ) _50228_ ( .A(_28524_), .B(12'h000), .S(RST), .Y(_02494_) );
  \$mux  #( .WIDTH(4) ) _50229_ ( .A(__delay_data_622), .B(4'h0), .S(RST), .Y(_00511_) );
  \$mux  #( .WIDTH(4) ) _50230_ ( .A(__delay_data_621), .B(4'h0), .S(RST), .Y(_00510_) );
  \$mux  #( .WIDTH(4) ) _50231_ ( .A(__delay_data_620), .B(4'h0), .S(RST), .Y(_00509_) );
  \$mux  #( .WIDTH(4) ) _50232_ ( .A(__delay_data_619), .B(4'h0), .S(RST), .Y(_00508_) );
  \$mux  #( .WIDTH(12) ) _50233_ ( .A(\__muladd_madd_86.madd._pipe_madd1 ), .B(12'h000), .S(RST), .Y(_00700_) );
  \$mux  #( .WIDTH(4) ) _50234_ ( .A(__delay_data_618), .B(4'h0), .S(RST), .Y(_00507_) );
  \$mux  #( .WIDTH(4) ) _50235_ ( .A(__delay_data_615), .B(4'h0), .S(RST), .Y(_00504_) );
  \$mux  #( .WIDTH(8) ) _50236_ ( .A(__delay_data_612), .B(8'h00), .S(RST), .Y(_00501_) );
  \$mux  #( .WIDTH(12) ) _50237_ ( .A(_29155_[11:0]), .B(12'h000), .S(RST), .Y(_01554_) );
  \$mux  #( .WIDTH(4) ) _50238_ ( .A(__delay_data_617), .B(4'h0), .S(RST), .Y(_00506_) );
  \$mux  #( .WIDTH(4) ) _50239_ ( .A(__delay_data_614), .B(4'h0), .S(RST), .Y(_00503_) );
  \$mux  #( .WIDTH(8) ) _50240_ ( .A(__delay_data_611), .B(8'h00), .S(RST), .Y(_00500_) );
  \$mux  #( .WIDTH(1) ) _50241_ ( .A(_greaterthan_data_74), .B(1'h0), .S(RST), .Y(_00498_) );
  \$mux  #( .WIDTH(18) ) _50242_ ( .A(_28511_), .B(18'h00000), .S(RST), .Y(_01881_) );
  \$mux  #( .WIDTH(4) ) _50243_ ( .A(__variable_wdata_73), .B(4'h0), .S(RST), .Y(_00505_) );
  \$mux  #( .WIDTH(4) ) _50244_ ( .A(__variable_wdata_72), .B(4'h0), .S(RST), .Y(_00502_) );
  \$mux  #( .WIDTH(8) ) _50245_ ( .A(__variable_wdata_71), .B(8'h00), .S(RST), .Y(_00499_) );
  \$mux  #( .WIDTH(4) ) _50246_ ( .A(_28620_), .B(4'h0), .S(RST), .Y(_01808_) );
  \$mux  #( .WIDTH(1) ) _50247_ ( .A(_06166_), .B(1'h0), .S(RST), .Y(_01700_) );
  \$mux  #( .WIDTH(1) ) _50248_ ( .A(_substream_mul_4_rshift_data_cond_874_46), .B(1'h1), .S(__tmp_1249_8), .Y(_26548_) );
  \$mux  #( .WIDTH(1) ) _50249_ ( .A(_26548_), .B(1'h0), .S(__tmp_1299_5), .Y(_26549_) );
  \$mux  #( .WIDTH(1) ) _50250_ ( .A(_26549_), .B(1'h0), .S(RST), .Y(_02826_) );
  \$mux  #( .WIDTH(1) ) _50251_ ( .A(_substream_mul_4_y_data_cond_874_45), .B(1'h1), .S(__tmp_1249_8), .Y(_26550_) );
  \$mux  #( .WIDTH(1) ) _50252_ ( .A(_26550_), .B(1'h0), .S(__tmp_1299_5), .Y(_26551_) );
  \$mux  #( .WIDTH(1) ) _50253_ ( .A(_26551_), .B(1'h0), .S(RST), .Y(_02830_) );
  \$mux  #( .WIDTH(1) ) _50254_ ( .A(_substream_mul_4_x_data_cond_874_44), .B(1'h1), .S(__tmp_1249_8), .Y(_26552_) );
  \$mux  #( .WIDTH(1) ) _50255_ ( .A(_26552_), .B(1'h0), .S(__tmp_1299_5), .Y(_26553_) );
  \$mux  #( .WIDTH(1) ) _50256_ ( .A(_26553_), .B(1'h0), .S(RST), .Y(_02828_) );
  \$mux  #( .WIDTH(1) ) _50257_ ( .A(_substream_mul_4_rshift_data_cond_592_2), .B(1'h1), .S(__tmp_799_12), .Y(_26554_) );
  \$mux  #( .WIDTH(1) ) _50258_ ( .A(_26554_), .B(1'h0), .S(__tmp_947_9), .Y(_26555_) );
  \$mux  #( .WIDTH(1) ) _50259_ ( .A(_26555_), .B(1'h0), .S(RST), .Y(_02825_) );
  \$mux  #( .WIDTH(1) ) _50260_ ( .A(_substream_mul_4_y_data_cond_592_1), .B(1'h1), .S(__tmp_799_12), .Y(_26556_) );
  \$mux  #( .WIDTH(1) ) _50261_ ( .A(_26556_), .B(1'h0), .S(__tmp_947_9), .Y(_26557_) );
  \$mux  #( .WIDTH(1) ) _50262_ ( .A(_26557_), .B(1'h0), .S(RST), .Y(_02829_) );
  \$mux  #( .WIDTH(1) ) _50263_ ( .A(_substream_mul_4_x_data_cond_592_0), .B(1'h1), .S(__tmp_799_12), .Y(_26558_) );
  \$mux  #( .WIDTH(1) ) _50264_ ( .A(_26558_), .B(1'h0), .S(__tmp_947_9), .Y(_26559_) );
  \$mux  #( .WIDTH(1) ) _50265_ ( .A(_26559_), .B(1'h0), .S(RST), .Y(_02827_) );
  \$mux  #( .WIDTH(1) ) _50266_ ( .A(__tmp_1299_11), .B(1'h0), .S(RST), .Y(_01186_) );
  \$mux  #( .WIDTH(1) ) _50267_ ( .A(__tmp_1299_10), .B(1'h0), .S(RST), .Y(_01185_) );
  \$mux  #( .WIDTH(1) ) _50268_ ( .A(__tmp_1299_9), .B(1'h0), .S(RST), .Y(_01184_) );
  \$mux  #( .WIDTH(1) ) _50269_ ( .A(__tmp_1299_8), .B(1'h0), .S(RST), .Y(_01190_) );
  \$mux  #( .WIDTH(1) ) _50270_ ( .A(__tmp_1299_7), .B(1'h0), .S(RST), .Y(_01189_) );
  \$mux  #( .WIDTH(1) ) _50271_ ( .A(__tmp_1299_6), .B(1'h0), .S(RST), .Y(_01188_) );
  \$mux  #( .WIDTH(1) ) _50272_ ( .A(__tmp_1299_5), .B(1'h0), .S(RST), .Y(_01187_) );
  \$mux  #( .WIDTH(1) ) _50273_ ( .A(__tmp_1299_4), .B(1'h0), .S(RST), .Y(_01183_) );
  \$mux  #( .WIDTH(1) ) _50274_ ( .A(__tmp_1299_3), .B(1'h0), .S(RST), .Y(_01182_) );
  \$mux  #( .WIDTH(1) ) _50275_ ( .A(__tmp_947_6), .B(1'h0), .S(RST), .Y(_01329_) );
  \$mux  #( .WIDTH(1) ) _50276_ ( .A(__tmp_947_4), .B(1'h0), .S(RST), .Y(_01327_) );
  \$mux  #( .WIDTH(1) ) _50277_ ( .A(__tmp_947_3), .B(1'h0), .S(RST), .Y(_01326_) );
  \$mux  #( .WIDTH(4) ) _50278_ ( .A(__variable_wdata_56), .B(__delay_data_1267[3:0]), .S(_substream_mul_4_rshift_data_cond_592_2), .Y(_26560_) );
  \$mux  #( .WIDTH(4) ) _50279_ ( .A(_26560_), .B(__delay_data_1428[3:0]), .S(_substream_mul_4_rshift_data_cond_874_46), .Y(_26561_) );
  \$mux  #( .WIDTH(4) ) _50280_ ( .A(_26561_), .B(4'h0), .S(RST), .Y(_01441_) );
  \$mux  #( .WIDTH(4) ) _50281_ ( .A(__variable_wdata_55), .B(__delay_data_955), .S(_substream_mul_4_y_data_cond_592_1), .Y(_26562_) );
  \$mux  #( .WIDTH(4) ) _50282_ ( .A(_26562_), .B(__delay_data_1426), .S(_substream_mul_4_y_data_cond_874_45), .Y(_26563_) );
  \$mux  #( .WIDTH(4) ) _50283_ ( .A(_26563_), .B(4'h0), .S(RST), .Y(_01440_) );
  \$mux  #( .WIDTH(8) ) _50284_ ( .A(__variable_wdata_54), .B(_cond_data_575), .S(_substream_mul_4_x_data_cond_592_0), .Y(_26564_) );
  \$mux  #( .WIDTH(8) ) _50285_ ( .A(_26564_), .B(_cond_data_873), .S(_substream_mul_4_x_data_cond_874_44), .Y(_26565_) );
  \$mux  #( .WIDTH(8) ) _50286_ ( .A(_26565_), .B(8'h00), .S(RST), .Y(_01439_) );
  \$mux  #( .WIDTH(12) ) _50287_ ( .A(_28523_), .B(12'h000), .S(RST), .Y(_02493_) );
  \$mux  #( .WIDTH(4) ) _50288_ ( .A(__delay_data_605), .B(4'h0), .S(RST), .Y(_00497_) );
  \$mux  #( .WIDTH(4) ) _50289_ ( .A(__delay_data_604), .B(4'h0), .S(RST), .Y(_00496_) );
  \$mux  #( .WIDTH(4) ) _50290_ ( .A(__delay_data_603), .B(4'h0), .S(RST), .Y(_00495_) );
  \$mux  #( .WIDTH(4) ) _50291_ ( .A(__delay_data_602), .B(4'h0), .S(RST), .Y(_00494_) );
  \$mux  #( .WIDTH(12) ) _50292_ ( .A(\__muladd_madd_69.madd._pipe_madd1 ), .B(12'h000), .S(RST), .Y(_00699_) );
  \$mux  #( .WIDTH(4) ) _50293_ ( .A(__delay_data_601), .B(4'h0), .S(RST), .Y(_00493_) );
  \$mux  #( .WIDTH(4) ) _50294_ ( .A(__delay_data_598), .B(4'h0), .S(RST), .Y(_00490_) );
  \$mux  #( .WIDTH(8) ) _50295_ ( .A(__delay_data_595), .B(8'h00), .S(RST), .Y(_00487_) );
  \$mux  #( .WIDTH(12) ) _50296_ ( .A(_29154_[11:0]), .B(12'h000), .S(RST), .Y(_01546_) );
  \$mux  #( .WIDTH(4) ) _50297_ ( .A(__delay_data_600), .B(4'h0), .S(RST), .Y(_00492_) );
  \$mux  #( .WIDTH(4) ) _50298_ ( .A(__delay_data_597), .B(4'h0), .S(RST), .Y(_00489_) );
  \$mux  #( .WIDTH(8) ) _50299_ ( .A(__delay_data_594), .B(8'h00), .S(RST), .Y(_00486_) );
  \$mux  #( .WIDTH(1) ) _50300_ ( .A(_greaterthan_data_57), .B(1'h0), .S(RST), .Y(_00484_) );
  \$mux  #( .WIDTH(18) ) _50301_ ( .A(_28510_), .B(18'h00000), .S(RST), .Y(_01880_) );
  \$mux  #( .WIDTH(4) ) _50302_ ( .A(__variable_wdata_56), .B(4'h0), .S(RST), .Y(_00491_) );
  \$mux  #( .WIDTH(4) ) _50303_ ( .A(__variable_wdata_55), .B(4'h0), .S(RST), .Y(_00488_) );
  \$mux  #( .WIDTH(8) ) _50304_ ( .A(__variable_wdata_54), .B(8'h00), .S(RST), .Y(_00485_) );
  \$mux  #( .WIDTH(4) ) _50305_ ( .A(_28619_), .B(4'h0), .S(RST), .Y(_01806_) );
  \$mux  #( .WIDTH(1) ) _50306_ ( .A(_06165_), .B(1'h0), .S(RST), .Y(_01699_) );
  \$mux  #( .WIDTH(1) ) _50307_ ( .A(_substream_mul_rshift_clip_3_rshift_data_cond_884_53), .B(1'h1), .S(__tmp_1249_28), .Y(_26566_) );
  \$mux  #( .WIDTH(1) ) _50308_ ( .A(_26566_), .B(1'h0), .S(__tmp_1291_25), .Y(_26567_) );
  \$mux  #( .WIDTH(1) ) _50309_ ( .A(_26567_), .B(1'h0), .S(RST), .Y(_02847_) );
  \$mux  #( .WIDTH(1) ) _50310_ ( .A(_substream_mul_rshift_clip_3_y_data_cond_884_52), .B(1'h1), .S(__tmp_1249_28), .Y(_26568_) );
  \$mux  #( .WIDTH(1) ) _50311_ ( .A(_26568_), .B(1'h0), .S(__tmp_1291_25), .Y(_26569_) );
  \$mux  #( .WIDTH(1) ) _50312_ ( .A(_26569_), .B(1'h0), .S(RST), .Y(_02851_) );
  \$mux  #( .WIDTH(1) ) _50313_ ( .A(_substream_mul_rshift_clip_3_x_data_cond_884_51), .B(1'h1), .S(__tmp_1249_28), .Y(_26570_) );
  \$mux  #( .WIDTH(1) ) _50314_ ( .A(_26570_), .B(1'h0), .S(__tmp_1291_25), .Y(_26571_) );
  \$mux  #( .WIDTH(1) ) _50315_ ( .A(_26571_), .B(1'h0), .S(RST), .Y(_02849_) );
  \$mux  #( .WIDTH(1) ) _50316_ ( .A(_substream_mul_rshift_clip_3_rshift_data_cond_763_41), .B(1'h1), .S(__tmp_799_34), .Y(_26572_) );
  \$mux  #( .WIDTH(1) ) _50317_ ( .A(_26572_), .B(1'h0), .S(__tmp_969_31), .Y(_26573_) );
  \$mux  #( .WIDTH(1) ) _50318_ ( .A(_26573_), .B(1'h0), .S(RST), .Y(_02846_) );
  \$mux  #( .WIDTH(1) ) _50319_ ( .A(_substream_mul_rshift_clip_3_y_data_cond_763_40), .B(1'h1), .S(__tmp_799_34), .Y(_26574_) );
  \$mux  #( .WIDTH(1) ) _50320_ ( .A(_26574_), .B(1'h0), .S(__tmp_969_31), .Y(_26575_) );
  \$mux  #( .WIDTH(1) ) _50321_ ( .A(_26575_), .B(1'h0), .S(RST), .Y(_02850_) );
  \$mux  #( .WIDTH(1) ) _50322_ ( .A(_substream_mul_rshift_clip_3_x_data_cond_763_39), .B(1'h1), .S(__tmp_799_34), .Y(_26576_) );
  \$mux  #( .WIDTH(1) ) _50323_ ( .A(_26576_), .B(1'h0), .S(__tmp_969_31), .Y(_26577_) );
  \$mux  #( .WIDTH(1) ) _50324_ ( .A(_26577_), .B(1'h0), .S(RST), .Y(_02848_) );
  \$mux  #( .WIDTH(6) ) _50325_ ( .A(__variable_wdata_40), .B(__delay_data_1396[5:0]), .S(_substream_mul_rshift_clip_3_rshift_data_cond_763_41), .Y(_26578_) );
  \$mux  #( .WIDTH(6) ) _50326_ ( .A(_26578_), .B(__delay_data_1527[5:0]), .S(_substream_mul_rshift_clip_3_rshift_data_cond_884_53), .Y(_26579_) );
  \$mux  #( .WIDTH(6) ) _50327_ ( .A(_26579_), .B(6'h00), .S(RST), .Y(_01429_) );
  \$mux  #( .WIDTH(8) ) _50328_ ( .A(__variable_wdata_39), .B(__delay_data_1368), .S(_substream_mul_rshift_clip_3_y_data_cond_763_40), .Y(_26580_) );
  \$mux  #( .WIDTH(8) ) _50329_ ( .A(_26580_), .B(__delay_data_1505), .S(_substream_mul_rshift_clip_3_y_data_cond_884_52), .Y(_26581_) );
  \$mux  #( .WIDTH(8) ) _50330_ ( .A(_26581_), .B(8'h00), .S(RST), .Y(_01428_) );
  \$mux  #( .WIDTH(32) ) _50331_ ( .A(__variable_wdata_38), .B(_plus_data_762), .S(_substream_mul_rshift_clip_3_x_data_cond_763_39), .Y(_26582_) );
  \$mux  #( .WIDTH(32) ) _50332_ ( .A(_26582_), .B(_plus_data_883), .S(_substream_mul_rshift_clip_3_x_data_cond_884_51), .Y(_26583_) );
  \$mux  #( .WIDTH(32) ) _50333_ ( .A(_26583_), .B(0), .S(RST), .Y(_01427_) );
  \$mux  #( .WIDTH(8) ) _50334_ ( .A(_29153_[7:0]), .B(8'h00), .S(RST), .Y(_01536_) );
  \$mux  #( .WIDTH(1) ) _50335_ ( .A(_greatereq_data_51), .B(1'h0), .S(RST), .Y(_00626_) );
  \$mux  #( .WIDTH(40) ) _50336_ ( .A(_29152_), .B(40'h0000000000), .S(RST), .Y(_01535_) );
  \$mux  #( .WIDTH(40) ) _50337_ ( .A(_29151_), .B(40'h0000000000), .S(RST), .Y(_01534_) );
  \$mux  #( .WIDTH(40) ) _50338_ ( .A(_sra_data_42), .B(40'h0000000000), .S(RST), .Y(_00625_) );
  \$mux  #( .WIDTH(1) ) _50339_ ( .A(_06149_), .B(1'h0), .S(RST), .Y(_01690_) );
  \$mux  #( .WIDTH(1) ) _50340_ ( .A(_06883_), .B(1'h0), .S(RST), .Y(_01703_) );
  \$mux  #( .WIDTH(1) ) _50341_ ( .A(_06164_), .B(1'h0), .S(RST), .Y(_01698_) );
  \$mux  #( .WIDTH(40) ) _50342_ ( .A(_28522_), .B(40'h0000000000), .S(RST), .Y(_02492_) );
  \$mux  #( .WIDTH(6) ) _50343_ ( .A(__delay_data_766), .B(6'h00), .S(RST), .Y(_00624_) );
  \$mux  #( .WIDTH(6) ) _50344_ ( .A(__delay_data_765), .B(6'h00), .S(RST), .Y(_00623_) );
  \$mux  #( .WIDTH(6) ) _50345_ ( .A(__delay_data_764), .B(6'h00), .S(RST), .Y(_00622_) );
  \$mux  #( .WIDTH(6) ) _50346_ ( .A(__variable_wdata_40), .B(6'h00), .S(RST), .Y(_00621_) );
  \$mux  #( .WIDTH(40) ) _50347_ ( .A(\_times_mul_41.mult._pipe_mul1 ), .B(40'h0000000000), .S(RST), .Y(_02852_) );
  \$mux  #( .WIDTH(1) ) _50348_ ( .A(_substream_add_tree_2_var8_data_cond_745_35), .B(1'h1), .S(__tmp_799_22), .Y(_26584_) );
  \$mux  #( .WIDTH(1) ) _50349_ ( .A(_26584_), .B(1'h0), .S(__tmp_969_19), .Y(_26585_) );
  \$mux  #( .WIDTH(1) ) _50350_ ( .A(_26585_), .B(1'h0), .S(RST), .Y(_02815_) );
  \$mux  #( .WIDTH(1) ) _50351_ ( .A(_substream_add_tree_2_var7_data_cond_745_34), .B(1'h1), .S(__tmp_799_22), .Y(_26586_) );
  \$mux  #( .WIDTH(1) ) _50352_ ( .A(_26586_), .B(1'h0), .S(__tmp_969_19), .Y(_26587_) );
  \$mux  #( .WIDTH(1) ) _50353_ ( .A(_26587_), .B(1'h0), .S(RST), .Y(_02814_) );
  \$mux  #( .WIDTH(1) ) _50354_ ( .A(_substream_add_tree_2_var6_data_cond_745_33), .B(1'h1), .S(__tmp_799_22), .Y(_26588_) );
  \$mux  #( .WIDTH(1) ) _50355_ ( .A(_26588_), .B(1'h0), .S(__tmp_969_19), .Y(_26589_) );
  \$mux  #( .WIDTH(1) ) _50356_ ( .A(_26589_), .B(1'h0), .S(RST), .Y(_02813_) );
  \$mux  #( .WIDTH(1) ) _50357_ ( .A(_substream_add_tree_2_var5_data_cond_745_32), .B(1'h1), .S(__tmp_799_22), .Y(_26590_) );
  \$mux  #( .WIDTH(1) ) _50358_ ( .A(_26590_), .B(1'h0), .S(__tmp_969_19), .Y(_26591_) );
  \$mux  #( .WIDTH(1) ) _50359_ ( .A(_26591_), .B(1'h0), .S(RST), .Y(_02812_) );
  \$mux  #( .WIDTH(1) ) _50360_ ( .A(_substream_add_tree_2_var4_data_cond_745_31), .B(1'h1), .S(__tmp_799_22), .Y(_26592_) );
  \$mux  #( .WIDTH(1) ) _50361_ ( .A(_26592_), .B(1'h0), .S(__tmp_969_19), .Y(_26593_) );
  \$mux  #( .WIDTH(1) ) _50362_ ( .A(_26593_), .B(1'h0), .S(RST), .Y(_02811_) );
  \$mux  #( .WIDTH(1) ) _50363_ ( .A(_substream_add_tree_2_var3_data_cond_745_30), .B(1'h1), .S(__tmp_799_22), .Y(_26594_) );
  \$mux  #( .WIDTH(1) ) _50364_ ( .A(_26594_), .B(1'h0), .S(__tmp_969_19), .Y(_26595_) );
  \$mux  #( .WIDTH(1) ) _50365_ ( .A(_26595_), .B(1'h0), .S(RST), .Y(_02810_) );
  \$mux  #( .WIDTH(1) ) _50366_ ( .A(_substream_add_tree_2_var2_data_cond_745_29), .B(1'h1), .S(__tmp_799_22), .Y(_26596_) );
  \$mux  #( .WIDTH(1) ) _50367_ ( .A(_26596_), .B(1'h0), .S(__tmp_969_19), .Y(_26597_) );
  \$mux  #( .WIDTH(1) ) _50368_ ( .A(_26597_), .B(1'h0), .S(RST), .Y(_02809_) );
  \$mux  #( .WIDTH(1) ) _50369_ ( .A(_substream_add_tree_2_var1_data_cond_745_28), .B(1'h1), .S(__tmp_799_22), .Y(_26598_) );
  \$mux  #( .WIDTH(1) ) _50370_ ( .A(_26598_), .B(1'h0), .S(__tmp_969_19), .Y(_26599_) );
  \$mux  #( .WIDTH(1) ) _50371_ ( .A(_26599_), .B(1'h0), .S(RST), .Y(_02808_) );
  \$mux  #( .WIDTH(1) ) _50372_ ( .A(_substream_add_tree_2_var0_data_cond_745_27), .B(1'h1), .S(__tmp_799_22), .Y(_26600_) );
  \$mux  #( .WIDTH(1) ) _50373_ ( .A(_26600_), .B(1'h0), .S(__tmp_969_19), .Y(_26601_) );
  \$mux  #( .WIDTH(1) ) _50374_ ( .A(_26601_), .B(1'h0), .S(RST), .Y(_02807_) );
  \$mux  #( .WIDTH(32) ) _50375_ ( .A(__variable_wdata_32), .B({ __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744[11], __substreamoutput_data_744 }), .S(_substream_add_tree_2_var8_data_cond_745_35), .Y(_26602_) );
  \$mux  #( .WIDTH(32) ) _50376_ ( .A(_26602_), .B(0), .S(RST), .Y(_01426_) );
  \$mux  #( .WIDTH(32) ) _50377_ ( .A(__variable_wdata_31), .B({ __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727[11], __substreamoutput_data_727 }), .S(_substream_add_tree_2_var7_data_cond_745_34), .Y(_26603_) );
  \$mux  #( .WIDTH(32) ) _50378_ ( .A(_26603_), .B(0), .S(RST), .Y(_01425_) );
  \$mux  #( .WIDTH(32) ) _50379_ ( .A(__variable_wdata_30), .B({ __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710[11], __substreamoutput_data_710 }), .S(_substream_add_tree_2_var6_data_cond_745_33), .Y(_26604_) );
  \$mux  #( .WIDTH(32) ) _50380_ ( .A(_26604_), .B(0), .S(RST), .Y(_01424_) );
  \$mux  #( .WIDTH(32) ) _50381_ ( .A(__variable_wdata_29), .B({ __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693[11], __substreamoutput_data_693 }), .S(_substream_add_tree_2_var5_data_cond_745_32), .Y(_26605_) );
  \$mux  #( .WIDTH(32) ) _50382_ ( .A(_26605_), .B(0), .S(RST), .Y(_01422_) );
  \$mux  #( .WIDTH(32) ) _50383_ ( .A(__variable_wdata_28), .B({ __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676[11], __substreamoutput_data_676 }), .S(_substream_add_tree_2_var4_data_cond_745_31), .Y(_26606_) );
  \$mux  #( .WIDTH(32) ) _50384_ ( .A(_26606_), .B(0), .S(RST), .Y(_01421_) );
  \$mux  #( .WIDTH(32) ) _50385_ ( .A(__variable_wdata_27), .B({ __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659[11], __substreamoutput_data_659 }), .S(_substream_add_tree_2_var3_data_cond_745_30), .Y(_26607_) );
  \$mux  #( .WIDTH(32) ) _50386_ ( .A(_26607_), .B(0), .S(RST), .Y(_01420_) );
  \$mux  #( .WIDTH(32) ) _50387_ ( .A(__variable_wdata_26), .B({ __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642[11], __substreamoutput_data_642 }), .S(_substream_add_tree_2_var2_data_cond_745_29), .Y(_26608_) );
  \$mux  #( .WIDTH(32) ) _50388_ ( .A(_26608_), .B(0), .S(RST), .Y(_01412_) );
  \$mux  #( .WIDTH(32) ) _50389_ ( .A(__variable_wdata_25), .B({ __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625[11], __substreamoutput_data_625 }), .S(_substream_add_tree_2_var1_data_cond_745_28), .Y(_26609_) );
  \$mux  #( .WIDTH(32) ) _50390_ ( .A(_26609_), .B(0), .S(RST), .Y(_01406_) );
  \$mux  #( .WIDTH(32) ) _50391_ ( .A(__variable_wdata_24), .B({ __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876 }), .S(_substream_add_tree_2_var0_data_cond_745_27), .Y(_26610_) );
  \$mux  #( .WIDTH(32) ) _50392_ ( .A(_26610_), .B(0), .S(RST), .Y(_01403_) );
  \$mux  #( .WIDTH(32) ) _50393_ ( .A(_24301_), .B(0), .S(RST), .Y(_00704_) );
  \$mux  #( .WIDTH(32) ) _50394_ ( .A(_24299_), .B(0), .S(RST), .Y(_00703_) );
  \$mux  #( .WIDTH(32) ) _50395_ ( .A(_24297_), .B(0), .S(RST), .Y(_00702_) );
  \$mux  #( .WIDTH(32) ) _50396_ ( .A(_24295_), .B(0), .S(RST), .Y(_00701_) );
  \$mux  #( .WIDTH(1) ) _50397_ ( .A(_substream_add_tree_1_var0_data_cond_877_47), .B(1'h1), .S(__tmp_1249_18), .Y(_26611_) );
  \$mux  #( .WIDTH(1) ) _50398_ ( .A(_26611_), .B(1'h0), .S(__tmp_1299_15), .Y(_26612_) );
  \$mux  #( .WIDTH(1) ) _50399_ ( .A(_26612_), .B(1'h0), .S(RST), .Y(_02806_) );
  \$mux  #( .WIDTH(32) ) _50400_ ( .A(__variable_wdata_22), .B({ __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876[11], __substreamoutput_data_876 }), .S(_substream_add_tree_1_var0_data_cond_877_47), .Y(_26613_) );
  \$mux  #( .WIDTH(32) ) _50401_ ( .A(_26613_), .B(0), .S(RST), .Y(_01399_) );
  \$mux  #( .WIDTH(1) ) _50402_ ( .A(_substream_acc_0_size_data_cond_879_50), .B(1'h1), .S(__tmp_1249_20), .Y(_26614_) );
  \$mux  #( .WIDTH(1) ) _50403_ ( .A(_26614_), .B(1'h0), .S(__tmp_1299_17), .Y(_26615_) );
  \$mux  #( .WIDTH(1) ) _50404_ ( .A(_26615_), .B(1'h0), .S(RST), .Y(_02803_) );
  \$mux  #( .WIDTH(1) ) _50405_ ( .A(_substream_acc_0_rshift_data_cond_879_49), .B(1'h1), .S(__tmp_1249_20), .Y(_26616_) );
  \$mux  #( .WIDTH(1) ) _50406_ ( .A(_26616_), .B(1'h0), .S(__tmp_1299_17), .Y(_26617_) );
  \$mux  #( .WIDTH(1) ) _50407_ ( .A(_26617_), .B(1'h0), .S(RST), .Y(_02801_) );
  \$mux  #( .WIDTH(1) ) _50408_ ( .A(_substream_acc_0_x_data_cond_879_48), .B(1'h1), .S(__tmp_1249_20), .Y(_26618_) );
  \$mux  #( .WIDTH(1) ) _50409_ ( .A(_26618_), .B(1'h0), .S(__tmp_1299_17), .Y(_26619_) );
  \$mux  #( .WIDTH(1) ) _50410_ ( .A(_26619_), .B(1'h0), .S(RST), .Y(_02805_) );
  \$mux  #( .WIDTH(1) ) _50411_ ( .A(_substream_acc_0_size_data_cond_747_38), .B(1'h1), .S(__tmp_799_26), .Y(_26620_) );
  \$mux  #( .WIDTH(1) ) _50412_ ( .A(_26620_), .B(1'h0), .S(__tmp_969_23), .Y(_26621_) );
  \$mux  #( .WIDTH(1) ) _50413_ ( .A(_26621_), .B(1'h0), .S(RST), .Y(_02802_) );
  \$mux  #( .WIDTH(1) ) _50414_ ( .A(_substream_acc_0_rshift_data_cond_747_37), .B(1'h1), .S(__tmp_799_26), .Y(_26622_) );
  \$mux  #( .WIDTH(1) ) _50415_ ( .A(_26622_), .B(1'h0), .S(__tmp_969_23), .Y(_26623_) );
  \$mux  #( .WIDTH(1) ) _50416_ ( .A(_26623_), .B(1'h0), .S(RST), .Y(_02800_) );
  \$mux  #( .WIDTH(1) ) _50417_ ( .A(_substream_acc_0_x_data_cond_747_36), .B(1'h1), .S(__tmp_799_26), .Y(_26624_) );
  \$mux  #( .WIDTH(1) ) _50418_ ( .A(_26624_), .B(1'h0), .S(__tmp_969_23), .Y(_26625_) );
  \$mux  #( .WIDTH(1) ) _50419_ ( .A(_26625_), .B(1'h0), .S(RST), .Y(_02804_) );
  \$mux  #( .WIDTH(1) ) _50420_ ( .A(_acc_0_reduce_reset), .B(1'h0), .S(__tmp_799_28), .Y(_26626_) );
  \$mux  #( .WIDTH(1) ) _50421_ ( .A(_26626_), .B(1'h1), .S(__tmp_969_24), .Y(_26627_) );
  \$mux  #( .WIDTH(1) ) _50422_ ( .A(_26627_), .B(1'h0), .S(__tmp_1249_22), .Y(_26628_) );
  \$mux  #( .WIDTH(1) ) _50423_ ( .A(_26628_), .B(1'h1), .S(__tmp_1299_18), .Y(_26629_) );
  \$mux  #( .WIDTH(1) ) _50424_ ( .A(_26629_), .B(1'h1), .S(RST), .Y(_01466_) );
  \$mux  #( .WIDTH(1) ) _50425_ ( .A(__tmp_1299_2), .B(1'h0), .S(RST), .Y(_01181_) );
  \$mux  #( .WIDTH(1) ) _50426_ ( .A(__tmp_1299_1), .B(1'h0), .S(RST), .Y(_01180_) );
  \$mux  #( .WIDTH(1) ) _50427_ ( .A(_tmp_1281), .B(1'h0), .S(RST), .Y(_01179_) );
  \$mux  #( .WIDTH(1) ) _50428_ ( .A(__tmp_947_2), .B(1'h0), .S(RST), .Y(_01325_) );
  \$mux  #( .WIDTH(1) ) _50429_ ( .A(__tmp_947_1), .B(1'h0), .S(RST), .Y(_01324_) );
  \$mux  #( .WIDTH(1) ) _50430_ ( .A(_tmp_943), .B(1'h0), .S(RST), .Y(_01323_) );
  \$mux  #( .WIDTH(32) ) _50431_ ( .A(__variable_wdata_2), .B({ 26'h0000000, __delay_data_1310 }), .S(_substream_acc_0_size_data_cond_747_38), .Y(_26630_) );
  \$mux  #( .WIDTH(32) ) _50432_ ( .A(_26630_), .B({ 21'h000000, __delay_data_1459 }), .S(_substream_acc_0_size_data_cond_879_50), .Y(_26631_) );
  \$mux  #( .WIDTH(32) ) _50433_ ( .A(_26631_), .B(0), .S(RST), .Y(_01423_) );
  \$mux  #( .WIDTH(6) ) _50434_ ( .A(__variable_wdata_1), .B(__delay_data_1288[5:0]), .S(_substream_acc_0_rshift_data_cond_747_37), .Y(_26632_) );
  \$mux  #( .WIDTH(6) ) _50435_ ( .A(_26632_), .B(__delay_data_1443[5:0]), .S(_substream_acc_0_rshift_data_cond_879_49), .Y(_26633_) );
  \$mux  #( .WIDTH(6) ) _50436_ ( .A(_26633_), .B(6'h00), .S(RST), .Y(_01392_) );
  \$mux  #( .WIDTH(32) ) _50437_ ( .A(__variable_wdata_0), .B(__substreamoutput_data_746), .S(_substream_acc_0_x_data_cond_747_36), .Y(_26634_) );
  \$mux  #( .WIDTH(32) ) _50438_ ( .A(_26634_), .B(__substreamoutput_data_878), .S(_substream_acc_0_x_data_cond_879_48), .Y(_26635_) );
  \$mux  #( .WIDTH(32) ) _50439_ ( .A(_26635_), .B(0), .S(RST), .Y(_01373_) );
  \$mux  #( .WIDTH(1) ) _50440_ ( .A(__delay_data_757), .B(1'h0), .S(RST), .Y(_00620_) );
  \$mux  #( .WIDTH(32) ) _50441_ ( .A(_28521_), .B(0), .S(RST), .Y(_02491_) );
  \$mux  #( .WIDTH(1) ) _50442_ ( .A(__delay_data_756), .B(1'h0), .S(RST), .Y(_00619_) );
  \$mux  #( .WIDTH(6) ) _50443_ ( .A(__delay_data_753), .B(6'h00), .S(RST), .Y(_00616_) );
  \$mux  #( .WIDTH(32) ) _50444_ ( .A(_24293_), .B(0), .S(RST), .Y(_01810_) );
  \$mux  #( .WIDTH(1) ) _50445_ ( .A(__delay_data_755), .B(1'h0), .S(RST), .Y(_00618_) );
  \$mux  #( .WIDTH(6) ) _50446_ ( .A(__delay_data_752), .B(6'h00), .S(RST), .Y(_00615_) );
  \$mux  #( .WIDTH(32) ) _50447_ ( .A(__delay_data_749), .B(0), .S(RST), .Y(_00612_) );
  \$mux  #( .WIDTH(32) ) _50448_ ( .A(_29150_[31:0]), .B(0), .S(RST), .Y(_01470_) );
  \$mux  #( .WIDTH(1) ) _50449_ ( .A(_pulse_data_19), .B(1'h0), .S(RST), .Y(_00617_) );
  \$mux  #( .WIDTH(6) ) _50450_ ( .A(__delay_data_751), .B(6'h00), .S(RST), .Y(_00614_) );
  \$mux  #( .WIDTH(32) ) _50451_ ( .A(_reduceadd_data_17), .B(0), .S(RST), .Y(_00611_) );
  \$mux  #( .WIDTH(1) ) _50452_ ( .A(_greaterthan_data_3), .B(1'h0), .S(RST), .Y(_00610_) );
  \$mux  #( .WIDTH(66) ) _50453_ ( .A(_28509_), .B(66'h00000000000000000), .S(RST), .Y(_01882_) );
  \$mux  #( .WIDTH(6) ) _50454_ ( .A(__variable_wdata_1), .B(6'h00), .S(RST), .Y(_00613_) );
  \$mux  #( .WIDTH(33) ) _50455_ ( .A(_29149_), .B(33'h000000000), .S(_acc_0_reduce_reset), .Y(_26636_) );
  \$mux  #( .WIDTH(33) ) _50456_ ( .A(_26636_), .B(33'h000000000), .S(RST), .Y(_01820_) );
  \$mux  #( .WIDTH(1) ) _50457_ ( .A(_06148_), .B(1'h0), .S(RST), .Y(_01822_) );
  \$mux  #( .WIDTH(33) ) _50458_ ( .A(_29148_), .B(33'h000000000), .S(_acc_0_reduce_reset), .Y(_26637_) );
  \$mux  #( .WIDTH(33) ) _50459_ ( .A(_26637_), .B(33'h000000000), .S(RST), .Y(_01837_) );
  \$mux  #( .WIDTH(32) ) _50460_ ( .A(_24290_), .B(__variable_wdata_0), .S(_acc_0_reduce_reset), .Y(_26638_) );
  \$mux  #( .WIDTH(32) ) _50461_ ( .A(__variable_wdata_0), .B(_26638_), .S(_05720_), .Y(_26639_) );
  \$mux  #( .WIDTH(32) ) _50462_ ( .A(_26639_), .B(0), .S(RST), .Y(_01838_) );
  \$mux  #( .WIDTH(6) ) _50463_ ( .A(_28618_), .B(6'h00), .S(RST), .Y(_01807_) );
  \$mux  #( .WIDTH(1) ) _50464_ ( .A(_06163_), .B(1'h0), .S(RST), .Y(_01697_) );
  \$mux  #( .WIDTH(34) ) _50465_ ( .A(_tmp_1018), .B(_28563_), .S(_06683_), .Y(_26640_) );
  \$mux  #( .WIDTH(34) ) _50466_ ( .A(_26640_), .B(_28617_), .S(_06684_), .Y(_26641_) );
  \$mux  #( .WIDTH(34) ) _50467_ ( .A(_26641_), .B(34'h000000000), .S(RST), .Y(_02865_) );
  \$mux  #( .WIDTH(1) ) _50468_ ( .A(_tmp_1017), .B(1'h0), .S(_06681_), .Y(_26642_) );
  \$mux  #( .WIDTH(1) ) _50469_ ( .A(_26642_), .B(_tmp_1016), .S(_06682_), .Y(_26643_) );
  \$mux  #( .WIDTH(1) ) _50470_ ( .A(_26643_), .B(1'h0), .S(RST), .Y(_02864_) );
  \$mux  #( .WIDTH(1) ) _50471_ ( .A(_tmp_1016), .B(1'h0), .S(_06682_), .Y(_26644_) );
  \$mux  #( .WIDTH(1) ) _50472_ ( .A(_26644_), .B(_06099_), .S(_06683_), .Y(_26645_) );
  \$mux  #( .WIDTH(1) ) _50473_ ( .A(_26645_), .B(1'h0), .S(_06684_), .Y(_26646_) );
  \$mux  #( .WIDTH(1) ) _50474_ ( .A(_26646_), .B(1'h1), .S(_06685_), .Y(_26647_) );
  \$mux  #( .WIDTH(1) ) _50475_ ( .A(_26647_), .B(1'h0), .S(RST), .Y(_02863_) );
  \$mux  #( .WIDTH(1) ) _50476_ ( .A(_tmp_1015), .B(1'h0), .S(_06681_), .Y(_26648_) );
  \$mux  #( .WIDTH(1) ) _50477_ ( .A(_26648_), .B(1'h1), .S(_06682_), .Y(_26649_) );
  \$mux  #( .WIDTH(1) ) _50478_ ( .A(_26649_), .B(1'h0), .S(RST), .Y(_02862_) );
  \$mux  #( .WIDTH(1) ) _50479_ ( .A(_tmp_1014), .B(1'h0), .S(_06682_), .Y(_26650_) );
  \$mux  #( .WIDTH(1) ) _50480_ ( .A(_26650_), .B(1'h1), .S(_06683_), .Y(_26651_) );
  \$mux  #( .WIDTH(1) ) _50481_ ( .A(_26651_), .B(1'h1), .S(_06684_), .Y(_26652_) );
  \$mux  #( .WIDTH(1) ) _50482_ ( .A(_26652_), .B(1'h0), .S(RST), .Y(_02861_) );
  \$mux  #( .WIDTH(8) ) _50483_ ( .A(_tmp_1013), .B(8'h00), .S(RST), .Y(_01108_) );
  \$mux  #( .WIDTH(1) ) _50484_ ( .A(_tmp_1012), .B(1'h0), .S(RST), .Y(_01107_) );
  \$mux  #( .WIDTH(1) ) _50485_ ( .A(_tmp_1007), .B(1'h0), .S(_06681_), .Y(_26653_) );
  \$mux  #( .WIDTH(1) ) _50486_ ( .A(_26653_), .B(1'h1), .S(_06682_), .Y(_26654_) );
  \$mux  #( .WIDTH(1) ) _50487_ ( .A(_26654_), .B(1'h0), .S(RST), .Y(_02859_) );
  \$mux  #( .WIDTH(1) ) _50488_ ( .A(_06680_), .B(1'h0), .S(RST), .Y(_01832_) );
  \$mux  #( .WIDTH(9) ) _50489_ ( .A(ram_w8_l2048_id11_3_1_addr), .B(_maxi_write_local_addr[8:0]), .S(_06683_), .Y(_26655_) );
  \$mux  #( .WIDTH(9) ) _50490_ ( .A(_26655_), .B(_24289_[8:0]), .S(_06684_), .Y(_26656_) );
  \$mux  #( .WIDTH(9) ) _50491_ ( .A(_26656_), .B(9'h000), .S(RST), .Y(_03716_) );
  \$mux  #( .WIDTH(1) ) _50492_ ( .A(ram_w8_l2048_id11_3_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id11_3_cond_0_1), .Y(_26657_) );
  \$mux  #( .WIDTH(1) ) _50493_ ( .A(_26657_), .B(1'h1), .S(_06680_), .Y(_26658_) );
  \$mux  #( .WIDTH(1) ) _50494_ ( .A(_26658_), .B(1'h0), .S(RST), .Y(_03715_) );
  \$mux  #( .WIDTH(8) ) _50495_ ( .A(ram_w8_l2048_id11_3_0_wdata), .B(_stream_conv2d_16_sink_37_sink_wdata), .S(_06680_), .Y(_26659_) );
  \$mux  #( .WIDTH(8) ) _50496_ ( .A(_26659_), .B(8'h00), .S(RST), .Y(_03714_) );
  \$mux  #( .WIDTH(9) ) _50497_ ( .A(ram_w8_l2048_id11_3_0_addr), .B(_stream_conv2d_16_sink_37_sink_waddr[10:2]), .S(_06680_), .Y(_26660_) );
  \$mux  #( .WIDTH(9) ) _50498_ ( .A(_26660_), .B(9'h000), .S(RST), .Y(_03713_) );
  \$mux  #( .WIDTH(34) ) _50499_ ( .A(_tmp_1006), .B(_28563_), .S(_06677_), .Y(_26661_) );
  \$mux  #( .WIDTH(34) ) _50500_ ( .A(_26661_), .B(_28616_), .S(_06678_), .Y(_26662_) );
  \$mux  #( .WIDTH(34) ) _50501_ ( .A(_26662_), .B(34'h000000000), .S(RST), .Y(_02858_) );
  \$mux  #( .WIDTH(1) ) _50502_ ( .A(_tmp_1005), .B(1'h0), .S(_06675_), .Y(_26663_) );
  \$mux  #( .WIDTH(1) ) _50503_ ( .A(_26663_), .B(_tmp_1004), .S(_06676_), .Y(_26664_) );
  \$mux  #( .WIDTH(1) ) _50504_ ( .A(_26664_), .B(1'h0), .S(RST), .Y(_02857_) );
  \$mux  #( .WIDTH(1) ) _50505_ ( .A(_tmp_1004), .B(1'h0), .S(_06676_), .Y(_26665_) );
  \$mux  #( .WIDTH(1) ) _50506_ ( .A(_26665_), .B(_06099_), .S(_06677_), .Y(_26666_) );
  \$mux  #( .WIDTH(1) ) _50507_ ( .A(_26666_), .B(1'h0), .S(_06678_), .Y(_26667_) );
  \$mux  #( .WIDTH(1) ) _50508_ ( .A(_26667_), .B(1'h1), .S(_06679_), .Y(_26668_) );
  \$mux  #( .WIDTH(1) ) _50509_ ( .A(_26668_), .B(1'h0), .S(RST), .Y(_02856_) );
  \$mux  #( .WIDTH(1) ) _50510_ ( .A(_tmp_1003), .B(1'h0), .S(_06675_), .Y(_26669_) );
  \$mux  #( .WIDTH(1) ) _50511_ ( .A(_26669_), .B(1'h1), .S(_06676_), .Y(_26670_) );
  \$mux  #( .WIDTH(1) ) _50512_ ( .A(_26670_), .B(1'h0), .S(RST), .Y(_02855_) );
  \$mux  #( .WIDTH(1) ) _50513_ ( .A(_tmp_1002), .B(1'h0), .S(_06676_), .Y(_26671_) );
  \$mux  #( .WIDTH(1) ) _50514_ ( .A(_26671_), .B(1'h1), .S(_06677_), .Y(_26672_) );
  \$mux  #( .WIDTH(1) ) _50515_ ( .A(_26672_), .B(1'h1), .S(_06678_), .Y(_26673_) );
  \$mux  #( .WIDTH(1) ) _50516_ ( .A(_26673_), .B(1'h0), .S(RST), .Y(_02854_) );
  \$mux  #( .WIDTH(8) ) _50517_ ( .A(_tmp_1001), .B(8'h00), .S(RST), .Y(_01106_) );
  \$mux  #( .WIDTH(1) ) _50518_ ( .A(_tmp_1000), .B(1'h0), .S(RST), .Y(_01105_) );
  \$mux  #( .WIDTH(1) ) _50519_ ( .A(_tmp_995), .B(1'h0), .S(_06675_), .Y(_26674_) );
  \$mux  #( .WIDTH(1) ) _50520_ ( .A(_26674_), .B(1'h1), .S(_06676_), .Y(_26675_) );
  \$mux  #( .WIDTH(1) ) _50521_ ( .A(_26675_), .B(1'h0), .S(RST), .Y(_03170_) );
  \$mux  #( .WIDTH(1) ) _50522_ ( .A(_06674_), .B(1'h0), .S(RST), .Y(_01831_) );
  \$mux  #( .WIDTH(9) ) _50523_ ( .A(ram_w8_l2048_id11_2_1_addr), .B(_maxi_write_local_addr[8:0]), .S(_06677_), .Y(_26676_) );
  \$mux  #( .WIDTH(9) ) _50524_ ( .A(_26676_), .B(_24288_[8:0]), .S(_06678_), .Y(_26677_) );
  \$mux  #( .WIDTH(9) ) _50525_ ( .A(_26677_), .B(9'h000), .S(RST), .Y(_03712_) );
  \$mux  #( .WIDTH(1) ) _50526_ ( .A(ram_w8_l2048_id11_2_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id11_2_cond_0_1), .Y(_26678_) );
  \$mux  #( .WIDTH(1) ) _50527_ ( .A(_26678_), .B(1'h1), .S(_06674_), .Y(_26679_) );
  \$mux  #( .WIDTH(1) ) _50528_ ( .A(_26679_), .B(1'h0), .S(RST), .Y(_03711_) );
  \$mux  #( .WIDTH(8) ) _50529_ ( .A(ram_w8_l2048_id11_2_0_wdata), .B(_stream_conv2d_16_sink_37_sink_wdata), .S(_06674_), .Y(_26680_) );
  \$mux  #( .WIDTH(8) ) _50530_ ( .A(_26680_), .B(8'h00), .S(RST), .Y(_03710_) );
  \$mux  #( .WIDTH(9) ) _50531_ ( .A(ram_w8_l2048_id11_2_0_addr), .B(_stream_conv2d_16_sink_37_sink_waddr[10:2]), .S(_06674_), .Y(_26681_) );
  \$mux  #( .WIDTH(9) ) _50532_ ( .A(_26681_), .B(9'h000), .S(RST), .Y(_03709_) );
  \$mux  #( .WIDTH(34) ) _50533_ ( .A(_tmp_994), .B(_28563_), .S(_06671_), .Y(_26682_) );
  \$mux  #( .WIDTH(34) ) _50534_ ( .A(_26682_), .B(_28615_), .S(_06672_), .Y(_26683_) );
  \$mux  #( .WIDTH(34) ) _50535_ ( .A(_26683_), .B(34'h000000000), .S(RST), .Y(_03169_) );
  \$mux  #( .WIDTH(1) ) _50536_ ( .A(_tmp_993), .B(1'h0), .S(_06669_), .Y(_26684_) );
  \$mux  #( .WIDTH(1) ) _50537_ ( .A(_26684_), .B(_tmp_992), .S(_06670_), .Y(_26685_) );
  \$mux  #( .WIDTH(1) ) _50538_ ( .A(_26685_), .B(1'h0), .S(RST), .Y(_03168_) );
  \$mux  #( .WIDTH(1) ) _50539_ ( .A(_tmp_992), .B(1'h0), .S(_06670_), .Y(_26686_) );
  \$mux  #( .WIDTH(1) ) _50540_ ( .A(_26686_), .B(_06099_), .S(_06671_), .Y(_26687_) );
  \$mux  #( .WIDTH(1) ) _50541_ ( .A(_26687_), .B(1'h0), .S(_06672_), .Y(_26688_) );
  \$mux  #( .WIDTH(1) ) _50542_ ( .A(_26688_), .B(1'h1), .S(_06673_), .Y(_26689_) );
  \$mux  #( .WIDTH(1) ) _50543_ ( .A(_26689_), .B(1'h0), .S(RST), .Y(_03167_) );
  \$mux  #( .WIDTH(1) ) _50544_ ( .A(_tmp_991), .B(1'h0), .S(_06669_), .Y(_26690_) );
  \$mux  #( .WIDTH(1) ) _50545_ ( .A(_26690_), .B(1'h1), .S(_06670_), .Y(_26691_) );
  \$mux  #( .WIDTH(1) ) _50546_ ( .A(_26691_), .B(1'h0), .S(RST), .Y(_03166_) );
  \$mux  #( .WIDTH(1) ) _50547_ ( .A(_tmp_990), .B(1'h0), .S(_06670_), .Y(_26692_) );
  \$mux  #( .WIDTH(1) ) _50548_ ( .A(_26692_), .B(1'h1), .S(_06671_), .Y(_26693_) );
  \$mux  #( .WIDTH(1) ) _50549_ ( .A(_26693_), .B(1'h1), .S(_06672_), .Y(_26694_) );
  \$mux  #( .WIDTH(1) ) _50550_ ( .A(_26694_), .B(1'h0), .S(RST), .Y(_03165_) );
  \$mux  #( .WIDTH(8) ) _50551_ ( .A(_tmp_989), .B(8'h00), .S(RST), .Y(_01372_) );
  \$mux  #( .WIDTH(1) ) _50552_ ( .A(_tmp_988), .B(1'h0), .S(RST), .Y(_01371_) );
  \$mux  #( .WIDTH(1) ) _50553_ ( .A(_tmp_983), .B(1'h0), .S(_06669_), .Y(_26695_) );
  \$mux  #( .WIDTH(1) ) _50554_ ( .A(_26695_), .B(1'h1), .S(_06670_), .Y(_26696_) );
  \$mux  #( .WIDTH(1) ) _50555_ ( .A(_26696_), .B(1'h0), .S(RST), .Y(_03164_) );
  \$mux  #( .WIDTH(1) ) _50556_ ( .A(_06668_), .B(1'h0), .S(RST), .Y(_01830_) );
  \$mux  #( .WIDTH(9) ) _50557_ ( .A(ram_w8_l2048_id11_1_1_addr), .B(_maxi_write_local_addr[8:0]), .S(_06671_), .Y(_26697_) );
  \$mux  #( .WIDTH(9) ) _50558_ ( .A(_26697_), .B(_24287_[8:0]), .S(_06672_), .Y(_26698_) );
  \$mux  #( .WIDTH(9) ) _50559_ ( .A(_26698_), .B(9'h000), .S(RST), .Y(_03708_) );
  \$mux  #( .WIDTH(1) ) _50560_ ( .A(ram_w8_l2048_id11_1_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id11_1_cond_0_1), .Y(_26699_) );
  \$mux  #( .WIDTH(1) ) _50561_ ( .A(_26699_), .B(1'h1), .S(_06668_), .Y(_26700_) );
  \$mux  #( .WIDTH(1) ) _50562_ ( .A(_26700_), .B(1'h0), .S(RST), .Y(_03707_) );
  \$mux  #( .WIDTH(8) ) _50563_ ( .A(ram_w8_l2048_id11_1_0_wdata), .B(_stream_conv2d_16_sink_37_sink_wdata), .S(_06668_), .Y(_26701_) );
  \$mux  #( .WIDTH(8) ) _50564_ ( .A(_26701_), .B(8'h00), .S(RST), .Y(_03706_) );
  \$mux  #( .WIDTH(9) ) _50565_ ( .A(ram_w8_l2048_id11_1_0_addr), .B(_stream_conv2d_16_sink_37_sink_waddr[10:2]), .S(_06668_), .Y(_26702_) );
  \$mux  #( .WIDTH(9) ) _50566_ ( .A(_26702_), .B(9'h000), .S(RST), .Y(_03705_) );
  \$mux  #( .WIDTH(1) ) _50567_ ( .A(_dataflow_cat_valid_98), .B(1'h0), .S(_06187_), .Y(_26703_) );
  \$mux  #( .WIDTH(1) ) _50568_ ( .A(_26703_), .B(_06666_), .S(_06667_), .Y(_26704_) );
  \$mux  #( .WIDTH(1) ) _50569_ ( .A(_26704_), .B(1'h0), .S(RST), .Y(_01591_) );
  \$mux  #( .WIDTH(32) ) _50570_ ( .A(_dataflow_cat_data_98), .B({ _tmp_1013, _tmp_1001, _tmp_989, _tmp_977 }), .S(_06667_), .Y(_26705_) );
  \$mux  #( .WIDTH(32) ) _50571_ ( .A(_26705_), .B(0), .S(RST), .Y(_01588_) );
  \$mux  #( .WIDTH(34) ) _50572_ ( .A(_tmp_982), .B(_28563_), .S(_06663_), .Y(_26706_) );
  \$mux  #( .WIDTH(34) ) _50573_ ( .A(_26706_), .B(_28614_), .S(_06664_), .Y(_26707_) );
  \$mux  #( .WIDTH(34) ) _50574_ ( .A(_26707_), .B(34'h000000000), .S(RST), .Y(_03163_) );
  \$mux  #( .WIDTH(1) ) _50575_ ( .A(_tmp_981), .B(1'h0), .S(_06660_), .Y(_26708_) );
  \$mux  #( .WIDTH(1) ) _50576_ ( .A(_26708_), .B(_tmp_980), .S(_06661_), .Y(_26709_) );
  \$mux  #( .WIDTH(1) ) _50577_ ( .A(_26709_), .B(1'h0), .S(RST), .Y(_03162_) );
  \$mux  #( .WIDTH(1) ) _50578_ ( .A(_tmp_980), .B(1'h0), .S(_06661_), .Y(_26710_) );
  \$mux  #( .WIDTH(1) ) _50579_ ( .A(_26710_), .B(_06099_), .S(_06663_), .Y(_26711_) );
  \$mux  #( .WIDTH(1) ) _50580_ ( .A(_26711_), .B(1'h0), .S(_06664_), .Y(_26712_) );
  \$mux  #( .WIDTH(1) ) _50581_ ( .A(_26712_), .B(1'h1), .S(_06665_), .Y(_26713_) );
  \$mux  #( .WIDTH(1) ) _50582_ ( .A(_26713_), .B(1'h0), .S(RST), .Y(_03161_) );
  \$mux  #( .WIDTH(1) ) _50583_ ( .A(_tmp_979), .B(1'h0), .S(_06660_), .Y(_26714_) );
  \$mux  #( .WIDTH(1) ) _50584_ ( .A(_26714_), .B(1'h1), .S(_06661_), .Y(_26715_) );
  \$mux  #( .WIDTH(1) ) _50585_ ( .A(_26715_), .B(1'h0), .S(RST), .Y(_03160_) );
  \$mux  #( .WIDTH(1) ) _50586_ ( .A(_tmp_978), .B(1'h0), .S(_06661_), .Y(_26716_) );
  \$mux  #( .WIDTH(1) ) _50587_ ( .A(_26716_), .B(1'h1), .S(_06663_), .Y(_26717_) );
  \$mux  #( .WIDTH(1) ) _50588_ ( .A(_26717_), .B(1'h1), .S(_06664_), .Y(_26718_) );
  \$mux  #( .WIDTH(1) ) _50589_ ( .A(_26718_), .B(1'h0), .S(RST), .Y(_03159_) );
  \$mux  #( .WIDTH(8) ) _50590_ ( .A(_tmp_977), .B(8'h00), .S(RST), .Y(_01370_) );
  \$mux  #( .WIDTH(1) ) _50591_ ( .A(_tmp_976), .B(1'h0), .S(RST), .Y(_01369_) );
  \$mux  #( .WIDTH(1) ) _50592_ ( .A(_tmp_971), .B(1'h0), .S(_06660_), .Y(_26719_) );
  \$mux  #( .WIDTH(1) ) _50593_ ( .A(_26719_), .B(1'h1), .S(_06661_), .Y(_26720_) );
  \$mux  #( .WIDTH(1) ) _50594_ ( .A(_26720_), .B(1'h0), .S(RST), .Y(_03158_) );
  \$mux  #( .WIDTH(1) ) _50595_ ( .A(_06659_), .B(1'h0), .S(RST), .Y(_01829_) );
  \$mux  #( .WIDTH(9) ) _50596_ ( .A(ram_w8_l2048_id11_0_1_addr), .B(_maxi_write_local_addr[8:0]), .S(_06663_), .Y(_26721_) );
  \$mux  #( .WIDTH(9) ) _50597_ ( .A(_26721_), .B(_24286_[8:0]), .S(_06664_), .Y(_26722_) );
  \$mux  #( .WIDTH(9) ) _50598_ ( .A(_26722_), .B(9'h000), .S(RST), .Y(_03704_) );
  \$mux  #( .WIDTH(1) ) _50599_ ( .A(ram_w8_l2048_id11_0_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id11_0_cond_0_1), .Y(_26723_) );
  \$mux  #( .WIDTH(1) ) _50600_ ( .A(_26723_), .B(1'h1), .S(_06659_), .Y(_26724_) );
  \$mux  #( .WIDTH(1) ) _50601_ ( .A(_26724_), .B(1'h0), .S(RST), .Y(_03703_) );
  \$mux  #( .WIDTH(8) ) _50602_ ( .A(ram_w8_l2048_id11_0_0_wdata), .B(_stream_conv2d_16_sink_37_sink_wdata), .S(_06659_), .Y(_26725_) );
  \$mux  #( .WIDTH(8) ) _50603_ ( .A(_26725_), .B(8'h00), .S(RST), .Y(_03702_) );
  \$mux  #( .WIDTH(9) ) _50604_ ( .A(ram_w8_l2048_id11_0_0_addr), .B(_stream_conv2d_16_sink_37_sink_waddr[10:2]), .S(_06659_), .Y(_26726_) );
  \$mux  #( .WIDTH(9) ) _50605_ ( .A(_26726_), .B(9'h000), .S(RST), .Y(_03701_) );
  \$mux  #( .WIDTH(1) ) _50606_ ( .A(ram_w8_l2048_id10_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26727_) );
  \$mux  #( .WIDTH(1) ) _50607_ ( .A(_26727_), .B(_06133_), .S(_06277_), .Y(_26728_) );
  \$mux  #( .WIDTH(1) ) _50608_ ( .A(_26728_), .B(1'h0), .S(RST), .Y(_03700_) );
  \$mux  #( .WIDTH(8) ) _50609_ ( .A(ram_w8_l2048_id10_3_1_wdata), .B(_dataflow_slice_data_89), .S(_06277_), .Y(_26729_) );
  \$mux  #( .WIDTH(8) ) _50610_ ( .A(_26729_), .B(8'h00), .S(RST), .Y(_03699_) );
  \$mux  #( .WIDTH(9) ) _50611_ ( .A(ram_w8_l2048_id10_3_1_addr), .B(_tmp_452), .S(_06277_), .Y(_26730_) );
  \$mux  #( .WIDTH(9) ) _50612_ ( .A(_26730_), .B(9'h000), .S(RST), .Y(_03698_) );
  \$mux  #( .WIDTH(9) ) _50613_ ( .A(ram_w8_l2048_id10_3_0_addr), .B(_stream_conv2d_16_source_27_source_ram_raddr[10:2]), .S(_tmp_583), .Y(_26731_) );
  \$mux  #( .WIDTH(9) ) _50614_ ( .A(_26731_), .B(9'h000), .S(RST), .Y(_03697_) );
  \$mux  #( .WIDTH(1) ) _50615_ ( .A(ram_w8_l2048_id10_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26732_) );
  \$mux  #( .WIDTH(1) ) _50616_ ( .A(_26732_), .B(_06130_), .S(_06274_), .Y(_26733_) );
  \$mux  #( .WIDTH(1) ) _50617_ ( .A(_26733_), .B(1'h0), .S(RST), .Y(_03696_) );
  \$mux  #( .WIDTH(8) ) _50618_ ( .A(ram_w8_l2048_id10_2_1_wdata), .B(_dataflow_slice_data_86), .S(_06274_), .Y(_26734_) );
  \$mux  #( .WIDTH(8) ) _50619_ ( .A(_26734_), .B(8'h00), .S(RST), .Y(_03695_) );
  \$mux  #( .WIDTH(9) ) _50620_ ( .A(ram_w8_l2048_id10_2_1_addr), .B(_tmp_439), .S(_06274_), .Y(_26735_) );
  \$mux  #( .WIDTH(9) ) _50621_ ( .A(_26735_), .B(9'h000), .S(RST), .Y(_03694_) );
  \$mux  #( .WIDTH(9) ) _50622_ ( .A(ram_w8_l2048_id10_2_0_addr), .B(_stream_conv2d_16_source_27_source_ram_raddr[10:2]), .S(_tmp_583), .Y(_26736_) );
  \$mux  #( .WIDTH(9) ) _50623_ ( .A(_26736_), .B(9'h000), .S(RST), .Y(_03693_) );
  \$mux  #( .WIDTH(1) ) _50624_ ( .A(ram_w8_l2048_id10_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26737_) );
  \$mux  #( .WIDTH(1) ) _50625_ ( .A(_26737_), .B(_06127_), .S(_06271_), .Y(_26738_) );
  \$mux  #( .WIDTH(1) ) _50626_ ( .A(_26738_), .B(1'h0), .S(RST), .Y(_03692_) );
  \$mux  #( .WIDTH(8) ) _50627_ ( .A(ram_w8_l2048_id10_1_1_wdata), .B(_dataflow_slice_data_83), .S(_06271_), .Y(_26739_) );
  \$mux  #( .WIDTH(8) ) _50628_ ( .A(_26739_), .B(8'h00), .S(RST), .Y(_03691_) );
  \$mux  #( .WIDTH(9) ) _50629_ ( .A(ram_w8_l2048_id10_1_1_addr), .B(_tmp_426), .S(_06271_), .Y(_26740_) );
  \$mux  #( .WIDTH(9) ) _50630_ ( .A(_26740_), .B(9'h000), .S(RST), .Y(_03690_) );
  \$mux  #( .WIDTH(9) ) _50631_ ( .A(ram_w8_l2048_id10_1_0_addr), .B(_stream_conv2d_16_source_27_source_ram_raddr[10:2]), .S(_tmp_583), .Y(_26741_) );
  \$mux  #( .WIDTH(9) ) _50632_ ( .A(_26741_), .B(9'h000), .S(RST), .Y(_03689_) );
  \$mux  #( .WIDTH(1) ) _50633_ ( .A(_tmp_583), .B(1'h0), .S(RST), .Y(_01261_) );
  \$mux  #( .WIDTH(1) ) _50634_ ( .A(ram_w8_l2048_id10_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26742_) );
  \$mux  #( .WIDTH(1) ) _50635_ ( .A(_26742_), .B(_06124_), .S(_06268_), .Y(_26743_) );
  \$mux  #( .WIDTH(1) ) _50636_ ( .A(_26743_), .B(1'h0), .S(RST), .Y(_03688_) );
  \$mux  #( .WIDTH(8) ) _50637_ ( .A(ram_w8_l2048_id10_0_1_wdata), .B(_dataflow_slice_data_80), .S(_06268_), .Y(_26744_) );
  \$mux  #( .WIDTH(8) ) _50638_ ( .A(_26744_), .B(8'h00), .S(RST), .Y(_03687_) );
  \$mux  #( .WIDTH(9) ) _50639_ ( .A(ram_w8_l2048_id10_0_1_addr), .B(_tmp_413), .S(_06268_), .Y(_26745_) );
  \$mux  #( .WIDTH(9) ) _50640_ ( .A(_26745_), .B(9'h000), .S(RST), .Y(_03686_) );
  \$mux  #( .WIDTH(9) ) _50641_ ( .A(ram_w8_l2048_id10_0_0_addr), .B(_stream_conv2d_16_source_27_source_ram_raddr[10:2]), .S(_tmp_583), .Y(_26746_) );
  \$mux  #( .WIDTH(9) ) _50642_ ( .A(_26746_), .B(9'h000), .S(RST), .Y(_03685_) );
  \$mux  #( .WIDTH(1) ) _50643_ ( .A(ram_w8_l2048_id9_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26747_) );
  \$mux  #( .WIDTH(1) ) _50644_ ( .A(_26747_), .B(_06135_), .S(_06277_), .Y(_26748_) );
  \$mux  #( .WIDTH(1) ) _50645_ ( .A(_26748_), .B(1'h0), .S(RST), .Y(_03868_) );
  \$mux  #( .WIDTH(8) ) _50646_ ( .A(ram_w8_l2048_id9_3_1_wdata), .B(_dataflow_slice_data_89), .S(_06277_), .Y(_26749_) );
  \$mux  #( .WIDTH(8) ) _50647_ ( .A(_26749_), .B(8'h00), .S(RST), .Y(_03867_) );
  \$mux  #( .WIDTH(9) ) _50648_ ( .A(ram_w8_l2048_id9_3_1_addr), .B(_tmp_451), .S(_06277_), .Y(_26750_) );
  \$mux  #( .WIDTH(9) ) _50649_ ( .A(_26750_), .B(9'h000), .S(RST), .Y(_03866_) );
  \$mux  #( .WIDTH(9) ) _50650_ ( .A(ram_w8_l2048_id9_3_0_addr), .B(_stream_conv2d_16_source_26_source_ram_raddr[10:2]), .S(_tmp_573), .Y(_26751_) );
  \$mux  #( .WIDTH(9) ) _50651_ ( .A(_26751_), .B(9'h000), .S(RST), .Y(_03865_) );
  \$mux  #( .WIDTH(1) ) _50652_ ( .A(ram_w8_l2048_id9_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26752_) );
  \$mux  #( .WIDTH(1) ) _50653_ ( .A(_26752_), .B(_06132_), .S(_06274_), .Y(_26753_) );
  \$mux  #( .WIDTH(1) ) _50654_ ( .A(_26753_), .B(1'h0), .S(RST), .Y(_03864_) );
  \$mux  #( .WIDTH(8) ) _50655_ ( .A(ram_w8_l2048_id9_2_1_wdata), .B(_dataflow_slice_data_86), .S(_06274_), .Y(_26754_) );
  \$mux  #( .WIDTH(8) ) _50656_ ( .A(_26754_), .B(8'h00), .S(RST), .Y(_03863_) );
  \$mux  #( .WIDTH(9) ) _50657_ ( .A(ram_w8_l2048_id9_2_1_addr), .B(_tmp_438), .S(_06274_), .Y(_26755_) );
  \$mux  #( .WIDTH(9) ) _50658_ ( .A(_26755_), .B(9'h000), .S(RST), .Y(_03862_) );
  \$mux  #( .WIDTH(9) ) _50659_ ( .A(ram_w8_l2048_id9_2_0_addr), .B(_stream_conv2d_16_source_26_source_ram_raddr[10:2]), .S(_tmp_573), .Y(_26756_) );
  \$mux  #( .WIDTH(9) ) _50660_ ( .A(_26756_), .B(9'h000), .S(RST), .Y(_03861_) );
  \$mux  #( .WIDTH(1) ) _50661_ ( .A(ram_w8_l2048_id9_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26757_) );
  \$mux  #( .WIDTH(1) ) _50662_ ( .A(_26757_), .B(_06129_), .S(_06271_), .Y(_26758_) );
  \$mux  #( .WIDTH(1) ) _50663_ ( .A(_26758_), .B(1'h0), .S(RST), .Y(_03860_) );
  \$mux  #( .WIDTH(8) ) _50664_ ( .A(ram_w8_l2048_id9_1_1_wdata), .B(_dataflow_slice_data_83), .S(_06271_), .Y(_26759_) );
  \$mux  #( .WIDTH(8) ) _50665_ ( .A(_26759_), .B(8'h00), .S(RST), .Y(_03859_) );
  \$mux  #( .WIDTH(9) ) _50666_ ( .A(ram_w8_l2048_id9_1_1_addr), .B(_tmp_425), .S(_06271_), .Y(_26760_) );
  \$mux  #( .WIDTH(9) ) _50667_ ( .A(_26760_), .B(9'h000), .S(RST), .Y(_03858_) );
  \$mux  #( .WIDTH(9) ) _50668_ ( .A(ram_w8_l2048_id9_1_0_addr), .B(_stream_conv2d_16_source_26_source_ram_raddr[10:2]), .S(_tmp_573), .Y(_26761_) );
  \$mux  #( .WIDTH(9) ) _50669_ ( .A(_26761_), .B(9'h000), .S(RST), .Y(_03857_) );
  \$mux  #( .WIDTH(1) ) _50670_ ( .A(_tmp_573), .B(1'h0), .S(RST), .Y(_01258_) );
  \$mux  #( .WIDTH(1) ) _50671_ ( .A(ram_w8_l2048_id9_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26762_) );
  \$mux  #( .WIDTH(1) ) _50672_ ( .A(_26762_), .B(_06126_), .S(_06268_), .Y(_26763_) );
  \$mux  #( .WIDTH(1) ) _50673_ ( .A(_26763_), .B(1'h0), .S(RST), .Y(_03856_) );
  \$mux  #( .WIDTH(8) ) _50674_ ( .A(ram_w8_l2048_id9_0_1_wdata), .B(_dataflow_slice_data_80), .S(_06268_), .Y(_26764_) );
  \$mux  #( .WIDTH(8) ) _50675_ ( .A(_26764_), .B(8'h00), .S(RST), .Y(_03855_) );
  \$mux  #( .WIDTH(9) ) _50676_ ( .A(ram_w8_l2048_id9_0_1_addr), .B(_tmp_412), .S(_06268_), .Y(_26765_) );
  \$mux  #( .WIDTH(9) ) _50677_ ( .A(_26765_), .B(9'h000), .S(RST), .Y(_03854_) );
  \$mux  #( .WIDTH(9) ) _50678_ ( .A(ram_w8_l2048_id9_0_0_addr), .B(_stream_conv2d_16_source_26_source_ram_raddr[10:2]), .S(_tmp_573), .Y(_26766_) );
  \$mux  #( .WIDTH(9) ) _50679_ ( .A(_26766_), .B(9'h000), .S(RST), .Y(_03853_) );
  \$mux  #( .WIDTH(2) ) _50680_ ( .A(_tmp_456), .B(2'h0), .S(_06652_), .Y(_26767_) );
  \$mux  #( .WIDTH(2) ) _50681_ ( .A(_26767_), .B(_24285_[1:0]), .S(_06653_), .Y(_26768_) );
  \$mux  #( .WIDTH(2) ) _50682_ ( .A(_26768_), .B(2'h0), .S(_06654_), .Y(_26769_) );
  \$mux  #( .WIDTH(2) ) _50683_ ( .A(_26769_), .B(2'h0), .S(RST), .Y(_03137_) );
  \$mux  #( .WIDTH(9) ) _50684_ ( .A(_tmp_449), .B(_28537_[8:0]), .S(_06652_), .Y(_26770_) );
  \$mux  #( .WIDTH(9) ) _50685_ ( .A(_26770_), .B(_tmp_452), .S(_06657_), .Y(_26771_) );
  \$mux  #( .WIDTH(9) ) _50686_ ( .A(_26771_), .B(9'h000), .S(RST), .Y(_03135_) );
  \$mux  #( .WIDTH(9) ) _50687_ ( .A(_tmp_448), .B(_28537_[8:0]), .S(_06652_), .Y(_26772_) );
  \$mux  #( .WIDTH(9) ) _50688_ ( .A(_26772_), .B(_tmp_451), .S(_06656_), .Y(_26773_) );
  \$mux  #( .WIDTH(9) ) _50689_ ( .A(_26773_), .B(9'h000), .S(RST), .Y(_03134_) );
  \$mux  #( .WIDTH(9) ) _50690_ ( .A(_tmp_447), .B(_28537_[8:0]), .S(_06652_), .Y(_26774_) );
  \$mux  #( .WIDTH(9) ) _50691_ ( .A(_26774_), .B(_tmp_450), .S(_06655_), .Y(_26775_) );
  \$mux  #( .WIDTH(9) ) _50692_ ( .A(_26775_), .B(9'h000), .S(RST), .Y(_03133_) );
  \$mux  #( .WIDTH(1) ) _50693_ ( .A(_tmp_446), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26776_) );
  \$mux  #( .WIDTH(1) ) _50694_ ( .A(_26776_), .B(1'h1), .S(_06658_), .Y(_26777_) );
  \$mux  #( .WIDTH(1) ) _50695_ ( .A(_26777_), .B(1'h0), .S(RST), .Y(_03132_) );
  \$mux  #( .WIDTH(34) ) _50696_ ( .A(_tmp_445), .B({ 1'h0, _maxi_read_size }), .S(_06652_), .Y(_26778_) );
  \$mux  #( .WIDTH(34) ) _50697_ ( .A(_26778_), .B(_28613_), .S(_06277_), .Y(_26779_) );
  \$mux  #( .WIDTH(34) ) _50698_ ( .A(_26779_), .B(34'h000000000), .S(RST), .Y(_03131_) );
  \$mux  #( .WIDTH(10) ) _50699_ ( .A(_tmp_444), .B(_28605_[9:0]), .S(_06652_), .Y(_26780_) );
  \$mux  #( .WIDTH(10) ) _50700_ ( .A(_26780_), .B(_28612_[9:0]), .S(_06277_), .Y(_26781_) );
  \$mux  #( .WIDTH(10) ) _50701_ ( .A(_26781_), .B(_28605_[9:0]), .S(_06653_), .Y(_26782_) );
  \$mux  #( .WIDTH(10) ) _50702_ ( .A(_26782_), .B(10'h000), .S(RST), .Y(_03130_) );
  \$mux  #( .WIDTH(1) ) _50703_ ( .A(ram_w8_l2048_id8_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26783_) );
  \$mux  #( .WIDTH(1) ) _50704_ ( .A(_26783_), .B(_06134_), .S(_06277_), .Y(_26784_) );
  \$mux  #( .WIDTH(1) ) _50705_ ( .A(_26784_), .B(1'h0), .S(RST), .Y(_03852_) );
  \$mux  #( .WIDTH(8) ) _50706_ ( .A(ram_w8_l2048_id8_3_1_wdata), .B(_dataflow_slice_data_89), .S(_06277_), .Y(_26785_) );
  \$mux  #( .WIDTH(8) ) _50707_ ( .A(_26785_), .B(8'h00), .S(RST), .Y(_03851_) );
  \$mux  #( .WIDTH(9) ) _50708_ ( .A(ram_w8_l2048_id8_3_1_addr), .B(_tmp_450), .S(_06277_), .Y(_26786_) );
  \$mux  #( .WIDTH(9) ) _50709_ ( .A(_26786_), .B(9'h000), .S(RST), .Y(_03850_) );
  \$mux  #( .WIDTH(9) ) _50710_ ( .A(ram_w8_l2048_id8_3_0_addr), .B(_stream_conv2d_16_source_25_source_ram_raddr[10:2]), .S(_tmp_563), .Y(_26787_) );
  \$mux  #( .WIDTH(9) ) _50711_ ( .A(_26787_), .B(9'h000), .S(RST), .Y(_03849_) );
  \$mux  #( .WIDTH(2) ) _50712_ ( .A(_tmp_443), .B(2'h0), .S(_06645_), .Y(_26788_) );
  \$mux  #( .WIDTH(2) ) _50713_ ( .A(_26788_), .B(_24284_[1:0]), .S(_06646_), .Y(_26789_) );
  \$mux  #( .WIDTH(2) ) _50714_ ( .A(_26789_), .B(2'h0), .S(_06647_), .Y(_26790_) );
  \$mux  #( .WIDTH(2) ) _50715_ ( .A(_26790_), .B(2'h0), .S(RST), .Y(_03129_) );
  \$mux  #( .WIDTH(9) ) _50716_ ( .A(_tmp_436), .B(_28537_[8:0]), .S(_06645_), .Y(_26791_) );
  \$mux  #( .WIDTH(9) ) _50717_ ( .A(_26791_), .B(_tmp_439), .S(_06650_), .Y(_26792_) );
  \$mux  #( .WIDTH(9) ) _50718_ ( .A(_26792_), .B(9'h000), .S(RST), .Y(_03127_) );
  \$mux  #( .WIDTH(9) ) _50719_ ( .A(_tmp_435), .B(_28537_[8:0]), .S(_06645_), .Y(_26793_) );
  \$mux  #( .WIDTH(9) ) _50720_ ( .A(_26793_), .B(_tmp_438), .S(_06649_), .Y(_26794_) );
  \$mux  #( .WIDTH(9) ) _50721_ ( .A(_26794_), .B(9'h000), .S(RST), .Y(_03126_) );
  \$mux  #( .WIDTH(9) ) _50722_ ( .A(_tmp_434), .B(_28537_[8:0]), .S(_06645_), .Y(_26795_) );
  \$mux  #( .WIDTH(9) ) _50723_ ( .A(_26795_), .B(_tmp_437), .S(_06648_), .Y(_26796_) );
  \$mux  #( .WIDTH(9) ) _50724_ ( .A(_26796_), .B(9'h000), .S(RST), .Y(_03125_) );
  \$mux  #( .WIDTH(1) ) _50725_ ( .A(_tmp_433), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26797_) );
  \$mux  #( .WIDTH(1) ) _50726_ ( .A(_26797_), .B(1'h1), .S(_06651_), .Y(_26798_) );
  \$mux  #( .WIDTH(1) ) _50727_ ( .A(_26798_), .B(1'h0), .S(RST), .Y(_03124_) );
  \$mux  #( .WIDTH(34) ) _50728_ ( .A(_tmp_432), .B({ 1'h0, _maxi_read_size }), .S(_06645_), .Y(_26799_) );
  \$mux  #( .WIDTH(34) ) _50729_ ( .A(_26799_), .B(_28611_), .S(_06274_), .Y(_26800_) );
  \$mux  #( .WIDTH(34) ) _50730_ ( .A(_26800_), .B(34'h000000000), .S(RST), .Y(_03123_) );
  \$mux  #( .WIDTH(10) ) _50731_ ( .A(_tmp_431), .B(_28605_[9:0]), .S(_06645_), .Y(_26801_) );
  \$mux  #( .WIDTH(10) ) _50732_ ( .A(_26801_), .B(_28610_[9:0]), .S(_06274_), .Y(_26802_) );
  \$mux  #( .WIDTH(10) ) _50733_ ( .A(_26802_), .B(_28605_[9:0]), .S(_06646_), .Y(_26803_) );
  \$mux  #( .WIDTH(10) ) _50734_ ( .A(_26803_), .B(10'h000), .S(RST), .Y(_03122_) );
  \$mux  #( .WIDTH(1) ) _50735_ ( .A(ram_w8_l2048_id8_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26804_) );
  \$mux  #( .WIDTH(1) ) _50736_ ( .A(_26804_), .B(_06131_), .S(_06274_), .Y(_26805_) );
  \$mux  #( .WIDTH(1) ) _50737_ ( .A(_26805_), .B(1'h0), .S(RST), .Y(_03848_) );
  \$mux  #( .WIDTH(8) ) _50738_ ( .A(ram_w8_l2048_id8_2_1_wdata), .B(_dataflow_slice_data_86), .S(_06274_), .Y(_26806_) );
  \$mux  #( .WIDTH(8) ) _50739_ ( .A(_26806_), .B(8'h00), .S(RST), .Y(_03847_) );
  \$mux  #( .WIDTH(9) ) _50740_ ( .A(ram_w8_l2048_id8_2_1_addr), .B(_tmp_437), .S(_06274_), .Y(_26807_) );
  \$mux  #( .WIDTH(9) ) _50741_ ( .A(_26807_), .B(9'h000), .S(RST), .Y(_03846_) );
  \$mux  #( .WIDTH(9) ) _50742_ ( .A(ram_w8_l2048_id8_2_0_addr), .B(_stream_conv2d_16_source_25_source_ram_raddr[10:2]), .S(_tmp_563), .Y(_26808_) );
  \$mux  #( .WIDTH(9) ) _50743_ ( .A(_26808_), .B(9'h000), .S(RST), .Y(_03845_) );
  \$mux  #( .WIDTH(2) ) _50744_ ( .A(_tmp_430), .B(2'h0), .S(_06638_), .Y(_26809_) );
  \$mux  #( .WIDTH(2) ) _50745_ ( .A(_26809_), .B(_24283_[1:0]), .S(_06639_), .Y(_26810_) );
  \$mux  #( .WIDTH(2) ) _50746_ ( .A(_26810_), .B(2'h0), .S(_06640_), .Y(_26811_) );
  \$mux  #( .WIDTH(2) ) _50747_ ( .A(_26811_), .B(2'h0), .S(RST), .Y(_03121_) );
  \$mux  #( .WIDTH(9) ) _50748_ ( .A(_tmp_423), .B(_28537_[8:0]), .S(_06638_), .Y(_26812_) );
  \$mux  #( .WIDTH(9) ) _50749_ ( .A(_26812_), .B(_tmp_426), .S(_06643_), .Y(_26813_) );
  \$mux  #( .WIDTH(9) ) _50750_ ( .A(_26813_), .B(9'h000), .S(RST), .Y(_03119_) );
  \$mux  #( .WIDTH(9) ) _50751_ ( .A(_tmp_422), .B(_28537_[8:0]), .S(_06638_), .Y(_26814_) );
  \$mux  #( .WIDTH(9) ) _50752_ ( .A(_26814_), .B(_tmp_425), .S(_06642_), .Y(_26815_) );
  \$mux  #( .WIDTH(9) ) _50753_ ( .A(_26815_), .B(9'h000), .S(RST), .Y(_03118_) );
  \$mux  #( .WIDTH(9) ) _50754_ ( .A(_tmp_421), .B(_28537_[8:0]), .S(_06638_), .Y(_26816_) );
  \$mux  #( .WIDTH(9) ) _50755_ ( .A(_26816_), .B(_tmp_424), .S(_06641_), .Y(_26817_) );
  \$mux  #( .WIDTH(9) ) _50756_ ( .A(_26817_), .B(9'h000), .S(RST), .Y(_03117_) );
  \$mux  #( .WIDTH(1) ) _50757_ ( .A(_tmp_420), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26818_) );
  \$mux  #( .WIDTH(1) ) _50758_ ( .A(_26818_), .B(1'h1), .S(_06644_), .Y(_26819_) );
  \$mux  #( .WIDTH(1) ) _50759_ ( .A(_26819_), .B(1'h0), .S(RST), .Y(_03116_) );
  \$mux  #( .WIDTH(34) ) _50760_ ( .A(_tmp_419), .B({ 1'h0, _maxi_read_size }), .S(_06638_), .Y(_26820_) );
  \$mux  #( .WIDTH(34) ) _50761_ ( .A(_26820_), .B(_28609_), .S(_06271_), .Y(_26821_) );
  \$mux  #( .WIDTH(34) ) _50762_ ( .A(_26821_), .B(34'h000000000), .S(RST), .Y(_03114_) );
  \$mux  #( .WIDTH(10) ) _50763_ ( .A(_tmp_418), .B(_28605_[9:0]), .S(_06638_), .Y(_26822_) );
  \$mux  #( .WIDTH(10) ) _50764_ ( .A(_26822_), .B(_28608_[9:0]), .S(_06271_), .Y(_26823_) );
  \$mux  #( .WIDTH(10) ) _50765_ ( .A(_26823_), .B(_28605_[9:0]), .S(_06639_), .Y(_26824_) );
  \$mux  #( .WIDTH(10) ) _50766_ ( .A(_26824_), .B(10'h000), .S(RST), .Y(_03113_) );
  \$mux  #( .WIDTH(1) ) _50767_ ( .A(ram_w8_l2048_id8_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26825_) );
  \$mux  #( .WIDTH(1) ) _50768_ ( .A(_26825_), .B(_06128_), .S(_06271_), .Y(_26826_) );
  \$mux  #( .WIDTH(1) ) _50769_ ( .A(_26826_), .B(1'h0), .S(RST), .Y(_03844_) );
  \$mux  #( .WIDTH(8) ) _50770_ ( .A(ram_w8_l2048_id8_1_1_wdata), .B(_dataflow_slice_data_83), .S(_06271_), .Y(_26827_) );
  \$mux  #( .WIDTH(8) ) _50771_ ( .A(_26827_), .B(8'h00), .S(RST), .Y(_03843_) );
  \$mux  #( .WIDTH(9) ) _50772_ ( .A(ram_w8_l2048_id8_1_1_addr), .B(_tmp_424), .S(_06271_), .Y(_26828_) );
  \$mux  #( .WIDTH(9) ) _50773_ ( .A(_26828_), .B(9'h000), .S(RST), .Y(_03842_) );
  \$mux  #( .WIDTH(9) ) _50774_ ( .A(ram_w8_l2048_id8_1_0_addr), .B(_stream_conv2d_16_source_25_source_ram_raddr[10:2]), .S(_tmp_563), .Y(_26829_) );
  \$mux  #( .WIDTH(9) ) _50775_ ( .A(_26829_), .B(9'h000), .S(RST), .Y(_03841_) );
  \$mux  #( .WIDTH(1) ) _50776_ ( .A(_tmp_563), .B(1'h0), .S(RST), .Y(_01255_) );
  \$mux  #( .WIDTH(2) ) _50777_ ( .A(_tmp_417), .B(2'h0), .S(_06631_), .Y(_26830_) );
  \$mux  #( .WIDTH(2) ) _50778_ ( .A(_26830_), .B(_24282_[1:0]), .S(_06632_), .Y(_26831_) );
  \$mux  #( .WIDTH(2) ) _50779_ ( .A(_26831_), .B(2'h0), .S(_06633_), .Y(_26832_) );
  \$mux  #( .WIDTH(2) ) _50780_ ( .A(_26832_), .B(2'h0), .S(RST), .Y(_03112_) );
  \$mux  #( .WIDTH(9) ) _50781_ ( .A(_tmp_410), .B(_28537_[8:0]), .S(_06631_), .Y(_26833_) );
  \$mux  #( .WIDTH(9) ) _50782_ ( .A(_26833_), .B(_tmp_413), .S(_06636_), .Y(_26834_) );
  \$mux  #( .WIDTH(9) ) _50783_ ( .A(_26834_), .B(9'h000), .S(RST), .Y(_03111_) );
  \$mux  #( .WIDTH(9) ) _50784_ ( .A(_tmp_409), .B(_28537_[8:0]), .S(_06631_), .Y(_26835_) );
  \$mux  #( .WIDTH(9) ) _50785_ ( .A(_26835_), .B(_tmp_412), .S(_06635_), .Y(_26836_) );
  \$mux  #( .WIDTH(9) ) _50786_ ( .A(_26836_), .B(9'h000), .S(RST), .Y(_03109_) );
  \$mux  #( .WIDTH(9) ) _50787_ ( .A(_tmp_408), .B(_28537_[8:0]), .S(_06631_), .Y(_26837_) );
  \$mux  #( .WIDTH(9) ) _50788_ ( .A(_26837_), .B(_tmp_411), .S(_06634_), .Y(_26838_) );
  \$mux  #( .WIDTH(9) ) _50789_ ( .A(_26838_), .B(9'h000), .S(RST), .Y(_03108_) );
  \$mux  #( .WIDTH(1) ) _50790_ ( .A(_tmp_407), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26839_) );
  \$mux  #( .WIDTH(1) ) _50791_ ( .A(_26839_), .B(1'h1), .S(_06637_), .Y(_26840_) );
  \$mux  #( .WIDTH(1) ) _50792_ ( .A(_26840_), .B(1'h0), .S(RST), .Y(_03107_) );
  \$mux  #( .WIDTH(34) ) _50793_ ( .A(_tmp_406), .B({ 1'h0, _maxi_read_size }), .S(_06631_), .Y(_26841_) );
  \$mux  #( .WIDTH(34) ) _50794_ ( .A(_26841_), .B(_28607_), .S(_06268_), .Y(_26842_) );
  \$mux  #( .WIDTH(34) ) _50795_ ( .A(_26842_), .B(34'h000000000), .S(RST), .Y(_03106_) );
  \$mux  #( .WIDTH(10) ) _50796_ ( .A(_tmp_405), .B(_28605_[9:0]), .S(_06631_), .Y(_26843_) );
  \$mux  #( .WIDTH(10) ) _50797_ ( .A(_26843_), .B(_28606_[9:0]), .S(_06268_), .Y(_26844_) );
  \$mux  #( .WIDTH(10) ) _50798_ ( .A(_26844_), .B(_28605_[9:0]), .S(_06632_), .Y(_26845_) );
  \$mux  #( .WIDTH(10) ) _50799_ ( .A(_26845_), .B(10'h000), .S(RST), .Y(_03105_) );
  \$mux  #( .WIDTH(1) ) _50800_ ( .A(ram_w8_l2048_id8_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26846_) );
  \$mux  #( .WIDTH(1) ) _50801_ ( .A(_26846_), .B(_06125_), .S(_06268_), .Y(_26847_) );
  \$mux  #( .WIDTH(1) ) _50802_ ( .A(_26847_), .B(1'h0), .S(RST), .Y(_03840_) );
  \$mux  #( .WIDTH(8) ) _50803_ ( .A(ram_w8_l2048_id8_0_1_wdata), .B(_dataflow_slice_data_80), .S(_06268_), .Y(_26848_) );
  \$mux  #( .WIDTH(8) ) _50804_ ( .A(_26848_), .B(8'h00), .S(RST), .Y(_03839_) );
  \$mux  #( .WIDTH(9) ) _50805_ ( .A(ram_w8_l2048_id8_0_1_addr), .B(_tmp_411), .S(_06268_), .Y(_26849_) );
  \$mux  #( .WIDTH(9) ) _50806_ ( .A(_26849_), .B(9'h000), .S(RST), .Y(_03838_) );
  \$mux  #( .WIDTH(9) ) _50807_ ( .A(ram_w8_l2048_id8_0_0_addr), .B(_stream_conv2d_16_source_25_source_ram_raddr[10:2]), .S(_tmp_563), .Y(_26850_) );
  \$mux  #( .WIDTH(9) ) _50808_ ( .A(_26850_), .B(9'h000), .S(RST), .Y(_03837_) );
  \$mux  #( .WIDTH(1) ) _50809_ ( .A(ram_w8_l2048_id7_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26851_) );
  \$mux  #( .WIDTH(1) ) _50810_ ( .A(_26851_), .B(_06121_), .S(_06265_), .Y(_26852_) );
  \$mux  #( .WIDTH(1) ) _50811_ ( .A(_26852_), .B(1'h0), .S(RST), .Y(_03836_) );
  \$mux  #( .WIDTH(8) ) _50812_ ( .A(ram_w8_l2048_id7_3_1_wdata), .B(_dataflow_slice_data_76), .S(_06265_), .Y(_26853_) );
  \$mux  #( .WIDTH(8) ) _50813_ ( .A(_26853_), .B(8'h00), .S(RST), .Y(_03835_) );
  \$mux  #( .WIDTH(9) ) _50814_ ( .A(ram_w8_l2048_id7_3_1_addr), .B(_tmp_395), .S(_06265_), .Y(_26854_) );
  \$mux  #( .WIDTH(9) ) _50815_ ( .A(_26854_), .B(9'h000), .S(RST), .Y(_03834_) );
  \$mux  #( .WIDTH(9) ) _50816_ ( .A(ram_w8_l2048_id7_3_0_addr), .B(_stream_conv2d_16_source_24_source_ram_raddr[10:2]), .S(_tmp_553), .Y(_26855_) );
  \$mux  #( .WIDTH(9) ) _50817_ ( .A(_26855_), .B(9'h000), .S(RST), .Y(_03833_) );
  \$mux  #( .WIDTH(1) ) _50818_ ( .A(ram_w8_l2048_id7_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26856_) );
  \$mux  #( .WIDTH(1) ) _50819_ ( .A(_26856_), .B(_06118_), .S(_06262_), .Y(_26857_) );
  \$mux  #( .WIDTH(1) ) _50820_ ( .A(_26857_), .B(1'h0), .S(RST), .Y(_03832_) );
  \$mux  #( .WIDTH(8) ) _50821_ ( .A(ram_w8_l2048_id7_2_1_wdata), .B(_dataflow_slice_data_73), .S(_06262_), .Y(_26858_) );
  \$mux  #( .WIDTH(8) ) _50822_ ( .A(_26858_), .B(8'h00), .S(RST), .Y(_03831_) );
  \$mux  #( .WIDTH(9) ) _50823_ ( .A(ram_w8_l2048_id7_2_1_addr), .B(_tmp_382), .S(_06262_), .Y(_26859_) );
  \$mux  #( .WIDTH(9) ) _50824_ ( .A(_26859_), .B(9'h000), .S(RST), .Y(_03830_) );
  \$mux  #( .WIDTH(9) ) _50825_ ( .A(ram_w8_l2048_id7_2_0_addr), .B(_stream_conv2d_16_source_24_source_ram_raddr[10:2]), .S(_tmp_553), .Y(_26860_) );
  \$mux  #( .WIDTH(9) ) _50826_ ( .A(_26860_), .B(9'h000), .S(RST), .Y(_03829_) );
  \$mux  #( .WIDTH(1) ) _50827_ ( .A(ram_w8_l2048_id7_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26861_) );
  \$mux  #( .WIDTH(1) ) _50828_ ( .A(_26861_), .B(_06115_), .S(_06259_), .Y(_26862_) );
  \$mux  #( .WIDTH(1) ) _50829_ ( .A(_26862_), .B(1'h0), .S(RST), .Y(_03828_) );
  \$mux  #( .WIDTH(8) ) _50830_ ( .A(ram_w8_l2048_id7_1_1_wdata), .B(_dataflow_slice_data_70), .S(_06259_), .Y(_26863_) );
  \$mux  #( .WIDTH(8) ) _50831_ ( .A(_26863_), .B(8'h00), .S(RST), .Y(_03827_) );
  \$mux  #( .WIDTH(9) ) _50832_ ( .A(ram_w8_l2048_id7_1_1_addr), .B(_tmp_369), .S(_06259_), .Y(_26864_) );
  \$mux  #( .WIDTH(9) ) _50833_ ( .A(_26864_), .B(9'h000), .S(RST), .Y(_03826_) );
  \$mux  #( .WIDTH(9) ) _50834_ ( .A(ram_w8_l2048_id7_1_0_addr), .B(_stream_conv2d_16_source_24_source_ram_raddr[10:2]), .S(_tmp_553), .Y(_26865_) );
  \$mux  #( .WIDTH(9) ) _50835_ ( .A(_26865_), .B(9'h000), .S(RST), .Y(_03825_) );
  \$mux  #( .WIDTH(1) ) _50836_ ( .A(_tmp_553), .B(1'h0), .S(RST), .Y(_01252_) );
  \$mux  #( .WIDTH(1) ) _50837_ ( .A(ram_w8_l2048_id7_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26866_) );
  \$mux  #( .WIDTH(1) ) _50838_ ( .A(_26866_), .B(_06112_), .S(_06256_), .Y(_26867_) );
  \$mux  #( .WIDTH(1) ) _50839_ ( .A(_26867_), .B(1'h0), .S(RST), .Y(_03824_) );
  \$mux  #( .WIDTH(8) ) _50840_ ( .A(ram_w8_l2048_id7_0_1_wdata), .B(_dataflow_slice_data_67), .S(_06256_), .Y(_26868_) );
  \$mux  #( .WIDTH(8) ) _50841_ ( .A(_26868_), .B(8'h00), .S(RST), .Y(_03823_) );
  \$mux  #( .WIDTH(9) ) _50842_ ( .A(ram_w8_l2048_id7_0_1_addr), .B(_tmp_356), .S(_06256_), .Y(_26869_) );
  \$mux  #( .WIDTH(9) ) _50843_ ( .A(_26869_), .B(9'h000), .S(RST), .Y(_03822_) );
  \$mux  #( .WIDTH(9) ) _50844_ ( .A(ram_w8_l2048_id7_0_0_addr), .B(_stream_conv2d_16_source_24_source_ram_raddr[10:2]), .S(_tmp_553), .Y(_26870_) );
  \$mux  #( .WIDTH(9) ) _50845_ ( .A(_26870_), .B(9'h000), .S(RST), .Y(_03821_) );
  \$mux  #( .WIDTH(1) ) _50846_ ( .A(ram_w8_l2048_id6_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26871_) );
  \$mux  #( .WIDTH(1) ) _50847_ ( .A(_26871_), .B(_06123_), .S(_06265_), .Y(_26872_) );
  \$mux  #( .WIDTH(1) ) _50848_ ( .A(_26872_), .B(1'h0), .S(RST), .Y(_03820_) );
  \$mux  #( .WIDTH(8) ) _50849_ ( .A(ram_w8_l2048_id6_3_1_wdata), .B(_dataflow_slice_data_76), .S(_06265_), .Y(_26873_) );
  \$mux  #( .WIDTH(8) ) _50850_ ( .A(_26873_), .B(8'h00), .S(RST), .Y(_03819_) );
  \$mux  #( .WIDTH(9) ) _50851_ ( .A(ram_w8_l2048_id6_3_1_addr), .B(_tmp_394), .S(_06265_), .Y(_26874_) );
  \$mux  #( .WIDTH(9) ) _50852_ ( .A(_26874_), .B(9'h000), .S(RST), .Y(_03818_) );
  \$mux  #( .WIDTH(9) ) _50853_ ( .A(ram_w8_l2048_id6_3_0_addr), .B(_stream_conv2d_16_source_23_source_ram_raddr[10:2]), .S(_tmp_543), .Y(_26875_) );
  \$mux  #( .WIDTH(9) ) _50854_ ( .A(_26875_), .B(9'h000), .S(RST), .Y(_03817_) );
  \$mux  #( .WIDTH(1) ) _50855_ ( .A(ram_w8_l2048_id6_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26876_) );
  \$mux  #( .WIDTH(1) ) _50856_ ( .A(_26876_), .B(_06120_), .S(_06262_), .Y(_26877_) );
  \$mux  #( .WIDTH(1) ) _50857_ ( .A(_26877_), .B(1'h0), .S(RST), .Y(_03816_) );
  \$mux  #( .WIDTH(8) ) _50858_ ( .A(ram_w8_l2048_id6_2_1_wdata), .B(_dataflow_slice_data_73), .S(_06262_), .Y(_26878_) );
  \$mux  #( .WIDTH(8) ) _50859_ ( .A(_26878_), .B(8'h00), .S(RST), .Y(_03815_) );
  \$mux  #( .WIDTH(9) ) _50860_ ( .A(ram_w8_l2048_id6_2_1_addr), .B(_tmp_381), .S(_06262_), .Y(_26879_) );
  \$mux  #( .WIDTH(9) ) _50861_ ( .A(_26879_), .B(9'h000), .S(RST), .Y(_03814_) );
  \$mux  #( .WIDTH(9) ) _50862_ ( .A(ram_w8_l2048_id6_2_0_addr), .B(_stream_conv2d_16_source_23_source_ram_raddr[10:2]), .S(_tmp_543), .Y(_26880_) );
  \$mux  #( .WIDTH(9) ) _50863_ ( .A(_26880_), .B(9'h000), .S(RST), .Y(_03813_) );
  \$mux  #( .WIDTH(1) ) _50864_ ( .A(ram_w8_l2048_id6_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26881_) );
  \$mux  #( .WIDTH(1) ) _50865_ ( .A(_26881_), .B(_06117_), .S(_06259_), .Y(_26882_) );
  \$mux  #( .WIDTH(1) ) _50866_ ( .A(_26882_), .B(1'h0), .S(RST), .Y(_03812_) );
  \$mux  #( .WIDTH(8) ) _50867_ ( .A(ram_w8_l2048_id6_1_1_wdata), .B(_dataflow_slice_data_70), .S(_06259_), .Y(_26883_) );
  \$mux  #( .WIDTH(8) ) _50868_ ( .A(_26883_), .B(8'h00), .S(RST), .Y(_03811_) );
  \$mux  #( .WIDTH(9) ) _50869_ ( .A(ram_w8_l2048_id6_1_1_addr), .B(_tmp_368), .S(_06259_), .Y(_26884_) );
  \$mux  #( .WIDTH(9) ) _50870_ ( .A(_26884_), .B(9'h000), .S(RST), .Y(_03810_) );
  \$mux  #( .WIDTH(9) ) _50871_ ( .A(ram_w8_l2048_id6_1_0_addr), .B(_stream_conv2d_16_source_23_source_ram_raddr[10:2]), .S(_tmp_543), .Y(_26885_) );
  \$mux  #( .WIDTH(9) ) _50872_ ( .A(_26885_), .B(9'h000), .S(RST), .Y(_03809_) );
  \$mux  #( .WIDTH(1) ) _50873_ ( .A(_tmp_543), .B(1'h0), .S(RST), .Y(_01249_) );
  \$mux  #( .WIDTH(1) ) _50874_ ( .A(ram_w8_l2048_id6_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26886_) );
  \$mux  #( .WIDTH(1) ) _50875_ ( .A(_26886_), .B(_06114_), .S(_06256_), .Y(_26887_) );
  \$mux  #( .WIDTH(1) ) _50876_ ( .A(_26887_), .B(1'h0), .S(RST), .Y(_03808_) );
  \$mux  #( .WIDTH(8) ) _50877_ ( .A(ram_w8_l2048_id6_0_1_wdata), .B(_dataflow_slice_data_67), .S(_06256_), .Y(_26888_) );
  \$mux  #( .WIDTH(8) ) _50878_ ( .A(_26888_), .B(8'h00), .S(RST), .Y(_03807_) );
  \$mux  #( .WIDTH(9) ) _50879_ ( .A(ram_w8_l2048_id6_0_1_addr), .B(_tmp_355), .S(_06256_), .Y(_26889_) );
  \$mux  #( .WIDTH(9) ) _50880_ ( .A(_26889_), .B(9'h000), .S(RST), .Y(_03806_) );
  \$mux  #( .WIDTH(9) ) _50881_ ( .A(ram_w8_l2048_id6_0_0_addr), .B(_stream_conv2d_16_source_23_source_ram_raddr[10:2]), .S(_tmp_543), .Y(_26890_) );
  \$mux  #( .WIDTH(9) ) _50882_ ( .A(_26890_), .B(9'h000), .S(RST), .Y(_03805_) );
  \$mux  #( .WIDTH(2) ) _50883_ ( .A(_tmp_399), .B(2'h0), .S(_06623_), .Y(_26891_) );
  \$mux  #( .WIDTH(2) ) _50884_ ( .A(_26891_), .B(_24281_[1:0]), .S(_06624_), .Y(_26892_) );
  \$mux  #( .WIDTH(2) ) _50885_ ( .A(_26892_), .B(2'h0), .S(_06625_), .Y(_26893_) );
  \$mux  #( .WIDTH(2) ) _50886_ ( .A(_26893_), .B(2'h0), .S(RST), .Y(_03102_) );
  \$mux  #( .WIDTH(9) ) _50887_ ( .A(_tmp_392), .B(_28537_[8:0]), .S(_06623_), .Y(_26894_) );
  \$mux  #( .WIDTH(9) ) _50888_ ( .A(_26894_), .B(_tmp_395), .S(_06628_), .Y(_26895_) );
  \$mux  #( .WIDTH(9) ) _50889_ ( .A(_26895_), .B(9'h000), .S(RST), .Y(_03101_) );
  \$mux  #( .WIDTH(9) ) _50890_ ( .A(_tmp_391), .B(_28537_[8:0]), .S(_06623_), .Y(_26896_) );
  \$mux  #( .WIDTH(9) ) _50891_ ( .A(_26896_), .B(_tmp_394), .S(_06627_), .Y(_26897_) );
  \$mux  #( .WIDTH(9) ) _50892_ ( .A(_26897_), .B(9'h000), .S(RST), .Y(_03100_) );
  \$mux  #( .WIDTH(9) ) _50893_ ( .A(_tmp_390), .B(_28537_[8:0]), .S(_06623_), .Y(_26898_) );
  \$mux  #( .WIDTH(9) ) _50894_ ( .A(_26898_), .B(_tmp_393), .S(_06626_), .Y(_26899_) );
  \$mux  #( .WIDTH(9) ) _50895_ ( .A(_26899_), .B(9'h000), .S(RST), .Y(_03099_) );
  \$mux  #( .WIDTH(1) ) _50896_ ( .A(_tmp_389), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26900_) );
  \$mux  #( .WIDTH(1) ) _50897_ ( .A(_26900_), .B(1'h1), .S(_06629_), .Y(_26901_) );
  \$mux  #( .WIDTH(1) ) _50898_ ( .A(_26901_), .B(1'h0), .S(RST), .Y(_03097_) );
  \$mux  #( .WIDTH(34) ) _50899_ ( .A(_tmp_388), .B({ 1'h0, _maxi_read_size }), .S(_06623_), .Y(_26902_) );
  \$mux  #( .WIDTH(34) ) _50900_ ( .A(_26902_), .B(_28604_), .S(_06265_), .Y(_26903_) );
  \$mux  #( .WIDTH(34) ) _50901_ ( .A(_26903_), .B(34'h000000000), .S(RST), .Y(_03096_) );
  \$mux  #( .WIDTH(10) ) _50902_ ( .A(_tmp_387), .B(_28596_[9:0]), .S(_06623_), .Y(_26904_) );
  \$mux  #( .WIDTH(10) ) _50903_ ( .A(_26904_), .B(_28603_[9:0]), .S(_06265_), .Y(_26905_) );
  \$mux  #( .WIDTH(10) ) _50904_ ( .A(_26905_), .B(_28596_[9:0]), .S(_06624_), .Y(_26906_) );
  \$mux  #( .WIDTH(10) ) _50905_ ( .A(_26906_), .B(10'h000), .S(RST), .Y(_03095_) );
  \$mux  #( .WIDTH(1) ) _50906_ ( .A(ram_w8_l2048_id5_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26907_) );
  \$mux  #( .WIDTH(1) ) _50907_ ( .A(_26907_), .B(_06122_), .S(_06265_), .Y(_26908_) );
  \$mux  #( .WIDTH(1) ) _50908_ ( .A(_26908_), .B(1'h0), .S(RST), .Y(_03804_) );
  \$mux  #( .WIDTH(8) ) _50909_ ( .A(ram_w8_l2048_id5_3_1_wdata), .B(_dataflow_slice_data_76), .S(_06265_), .Y(_26909_) );
  \$mux  #( .WIDTH(8) ) _50910_ ( .A(_26909_), .B(8'h00), .S(RST), .Y(_03803_) );
  \$mux  #( .WIDTH(9) ) _50911_ ( .A(ram_w8_l2048_id5_3_1_addr), .B(_tmp_393), .S(_06265_), .Y(_26910_) );
  \$mux  #( .WIDTH(9) ) _50912_ ( .A(_26910_), .B(9'h000), .S(RST), .Y(_03802_) );
  \$mux  #( .WIDTH(9) ) _50913_ ( .A(ram_w8_l2048_id5_3_0_addr), .B(_stream_conv2d_16_source_22_source_ram_raddr[10:2]), .S(_tmp_533), .Y(_26911_) );
  \$mux  #( .WIDTH(9) ) _50914_ ( .A(_26911_), .B(9'h000), .S(RST), .Y(_03801_) );
  \$mux  #( .WIDTH(2) ) _50915_ ( .A(_tmp_386), .B(2'h0), .S(_06616_), .Y(_26912_) );
  \$mux  #( .WIDTH(2) ) _50916_ ( .A(_26912_), .B(_24280_[1:0]), .S(_06617_), .Y(_26913_) );
  \$mux  #( .WIDTH(2) ) _50917_ ( .A(_26913_), .B(2'h0), .S(_06618_), .Y(_26914_) );
  \$mux  #( .WIDTH(2) ) _50918_ ( .A(_26914_), .B(2'h0), .S(RST), .Y(_03094_) );
  \$mux  #( .WIDTH(9) ) _50919_ ( .A(_tmp_379), .B(_28537_[8:0]), .S(_06616_), .Y(_26915_) );
  \$mux  #( .WIDTH(9) ) _50920_ ( .A(_26915_), .B(_tmp_382), .S(_06621_), .Y(_26916_) );
  \$mux  #( .WIDTH(9) ) _50921_ ( .A(_26916_), .B(9'h000), .S(RST), .Y(_03093_) );
  \$mux  #( .WIDTH(9) ) _50922_ ( .A(_tmp_378), .B(_28537_[8:0]), .S(_06616_), .Y(_26917_) );
  \$mux  #( .WIDTH(9) ) _50923_ ( .A(_26917_), .B(_tmp_381), .S(_06620_), .Y(_26918_) );
  \$mux  #( .WIDTH(9) ) _50924_ ( .A(_26918_), .B(9'h000), .S(RST), .Y(_03092_) );
  \$mux  #( .WIDTH(9) ) _50925_ ( .A(_tmp_377), .B(_28537_[8:0]), .S(_06616_), .Y(_26919_) );
  \$mux  #( .WIDTH(9) ) _50926_ ( .A(_26919_), .B(_tmp_380), .S(_06619_), .Y(_26920_) );
  \$mux  #( .WIDTH(9) ) _50927_ ( .A(_26920_), .B(9'h000), .S(RST), .Y(_03091_) );
  \$mux  #( .WIDTH(1) ) _50928_ ( .A(_tmp_376), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26921_) );
  \$mux  #( .WIDTH(1) ) _50929_ ( .A(_26921_), .B(1'h1), .S(_06622_), .Y(_26922_) );
  \$mux  #( .WIDTH(1) ) _50930_ ( .A(_26922_), .B(1'h0), .S(RST), .Y(_03090_) );
  \$mux  #( .WIDTH(34) ) _50931_ ( .A(_tmp_375), .B({ 1'h0, _maxi_read_size }), .S(_06616_), .Y(_26923_) );
  \$mux  #( .WIDTH(34) ) _50932_ ( .A(_26923_), .B(_28602_), .S(_06262_), .Y(_26924_) );
  \$mux  #( .WIDTH(34) ) _50933_ ( .A(_26924_), .B(34'h000000000), .S(RST), .Y(_03089_) );
  \$mux  #( .WIDTH(10) ) _50934_ ( .A(_tmp_374), .B(_28596_[9:0]), .S(_06616_), .Y(_26925_) );
  \$mux  #( .WIDTH(10) ) _50935_ ( .A(_26925_), .B(_28601_[9:0]), .S(_06262_), .Y(_26926_) );
  \$mux  #( .WIDTH(10) ) _50936_ ( .A(_26926_), .B(_28596_[9:0]), .S(_06617_), .Y(_26927_) );
  \$mux  #( .WIDTH(10) ) _50937_ ( .A(_26927_), .B(10'h000), .S(RST), .Y(_03088_) );
  \$mux  #( .WIDTH(1) ) _50938_ ( .A(ram_w8_l2048_id5_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26928_) );
  \$mux  #( .WIDTH(1) ) _50939_ ( .A(_26928_), .B(_06119_), .S(_06262_), .Y(_26929_) );
  \$mux  #( .WIDTH(1) ) _50940_ ( .A(_26929_), .B(1'h0), .S(RST), .Y(_03800_) );
  \$mux  #( .WIDTH(8) ) _50941_ ( .A(ram_w8_l2048_id5_2_1_wdata), .B(_dataflow_slice_data_73), .S(_06262_), .Y(_26930_) );
  \$mux  #( .WIDTH(8) ) _50942_ ( .A(_26930_), .B(8'h00), .S(RST), .Y(_03799_) );
  \$mux  #( .WIDTH(9) ) _50943_ ( .A(ram_w8_l2048_id5_2_1_addr), .B(_tmp_380), .S(_06262_), .Y(_26931_) );
  \$mux  #( .WIDTH(9) ) _50944_ ( .A(_26931_), .B(9'h000), .S(RST), .Y(_03798_) );
  \$mux  #( .WIDTH(9) ) _50945_ ( .A(ram_w8_l2048_id5_2_0_addr), .B(_stream_conv2d_16_source_22_source_ram_raddr[10:2]), .S(_tmp_533), .Y(_26932_) );
  \$mux  #( .WIDTH(9) ) _50946_ ( .A(_26932_), .B(9'h000), .S(RST), .Y(_03797_) );
  \$mux  #( .WIDTH(2) ) _50947_ ( .A(_tmp_373), .B(2'h0), .S(_06609_), .Y(_26933_) );
  \$mux  #( .WIDTH(2) ) _50948_ ( .A(_26933_), .B(_24279_[1:0]), .S(_06610_), .Y(_26934_) );
  \$mux  #( .WIDTH(2) ) _50949_ ( .A(_26934_), .B(2'h0), .S(_06611_), .Y(_26935_) );
  \$mux  #( .WIDTH(2) ) _50950_ ( .A(_26935_), .B(2'h0), .S(RST), .Y(_03087_) );
  \$mux  #( .WIDTH(9) ) _50951_ ( .A(_tmp_366), .B(_28537_[8:0]), .S(_06609_), .Y(_26936_) );
  \$mux  #( .WIDTH(9) ) _50952_ ( .A(_26936_), .B(_tmp_369), .S(_06614_), .Y(_26937_) );
  \$mux  #( .WIDTH(9) ) _50953_ ( .A(_26937_), .B(9'h000), .S(RST), .Y(_03086_) );
  \$mux  #( .WIDTH(9) ) _50954_ ( .A(_tmp_365), .B(_28537_[8:0]), .S(_06609_), .Y(_26938_) );
  \$mux  #( .WIDTH(9) ) _50955_ ( .A(_26938_), .B(_tmp_368), .S(_06613_), .Y(_26939_) );
  \$mux  #( .WIDTH(9) ) _50956_ ( .A(_26939_), .B(9'h000), .S(RST), .Y(_03085_) );
  \$mux  #( .WIDTH(9) ) _50957_ ( .A(_tmp_364), .B(_28537_[8:0]), .S(_06609_), .Y(_26940_) );
  \$mux  #( .WIDTH(9) ) _50958_ ( .A(_26940_), .B(_tmp_367), .S(_06612_), .Y(_26941_) );
  \$mux  #( .WIDTH(9) ) _50959_ ( .A(_26941_), .B(9'h000), .S(RST), .Y(_03084_) );
  \$mux  #( .WIDTH(1) ) _50960_ ( .A(_tmp_363), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26942_) );
  \$mux  #( .WIDTH(1) ) _50961_ ( .A(_26942_), .B(1'h1), .S(_06615_), .Y(_26943_) );
  \$mux  #( .WIDTH(1) ) _50962_ ( .A(_26943_), .B(1'h0), .S(RST), .Y(_03083_) );
  \$mux  #( .WIDTH(34) ) _50963_ ( .A(_tmp_362), .B({ 1'h0, _maxi_read_size }), .S(_06609_), .Y(_26944_) );
  \$mux  #( .WIDTH(34) ) _50964_ ( .A(_26944_), .B(_28600_), .S(_06259_), .Y(_26945_) );
  \$mux  #( .WIDTH(34) ) _50965_ ( .A(_26945_), .B(34'h000000000), .S(RST), .Y(_03082_) );
  \$mux  #( .WIDTH(10) ) _50966_ ( .A(_tmp_361), .B(_28596_[9:0]), .S(_06609_), .Y(_26946_) );
  \$mux  #( .WIDTH(10) ) _50967_ ( .A(_26946_), .B(_28599_[9:0]), .S(_06259_), .Y(_26947_) );
  \$mux  #( .WIDTH(10) ) _50968_ ( .A(_26947_), .B(_28596_[9:0]), .S(_06610_), .Y(_26948_) );
  \$mux  #( .WIDTH(10) ) _50969_ ( .A(_26948_), .B(10'h000), .S(RST), .Y(_03081_) );
  \$mux  #( .WIDTH(1) ) _50970_ ( .A(ram_w8_l2048_id5_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26949_) );
  \$mux  #( .WIDTH(1) ) _50971_ ( .A(_26949_), .B(_06116_), .S(_06259_), .Y(_26950_) );
  \$mux  #( .WIDTH(1) ) _50972_ ( .A(_26950_), .B(1'h0), .S(RST), .Y(_03796_) );
  \$mux  #( .WIDTH(8) ) _50973_ ( .A(ram_w8_l2048_id5_1_1_wdata), .B(_dataflow_slice_data_70), .S(_06259_), .Y(_26951_) );
  \$mux  #( .WIDTH(8) ) _50974_ ( .A(_26951_), .B(8'h00), .S(RST), .Y(_03795_) );
  \$mux  #( .WIDTH(9) ) _50975_ ( .A(ram_w8_l2048_id5_1_1_addr), .B(_tmp_367), .S(_06259_), .Y(_26952_) );
  \$mux  #( .WIDTH(9) ) _50976_ ( .A(_26952_), .B(9'h000), .S(RST), .Y(_03794_) );
  \$mux  #( .WIDTH(9) ) _50977_ ( .A(ram_w8_l2048_id5_1_0_addr), .B(_stream_conv2d_16_source_22_source_ram_raddr[10:2]), .S(_tmp_533), .Y(_26953_) );
  \$mux  #( .WIDTH(9) ) _50978_ ( .A(_26953_), .B(9'h000), .S(RST), .Y(_03793_) );
  \$mux  #( .WIDTH(1) ) _50979_ ( .A(_tmp_533), .B(1'h0), .S(RST), .Y(_01246_) );
  \$mux  #( .WIDTH(2) ) _50980_ ( .A(_tmp_360), .B(2'h0), .S(_06602_), .Y(_26954_) );
  \$mux  #( .WIDTH(2) ) _50981_ ( .A(_26954_), .B(_24278_[1:0]), .S(_06603_), .Y(_26955_) );
  \$mux  #( .WIDTH(2) ) _50982_ ( .A(_26955_), .B(2'h0), .S(_06604_), .Y(_26956_) );
  \$mux  #( .WIDTH(2) ) _50983_ ( .A(_26956_), .B(2'h0), .S(RST), .Y(_03080_) );
  \$mux  #( .WIDTH(9) ) _50984_ ( .A(_tmp_353), .B(_28537_[8:0]), .S(_06602_), .Y(_26957_) );
  \$mux  #( .WIDTH(9) ) _50985_ ( .A(_26957_), .B(_tmp_356), .S(_06607_), .Y(_26958_) );
  \$mux  #( .WIDTH(9) ) _50986_ ( .A(_26958_), .B(9'h000), .S(RST), .Y(_03079_) );
  \$mux  #( .WIDTH(9) ) _50987_ ( .A(_tmp_352), .B(_28537_[8:0]), .S(_06602_), .Y(_26959_) );
  \$mux  #( .WIDTH(9) ) _50988_ ( .A(_26959_), .B(_tmp_355), .S(_06606_), .Y(_26960_) );
  \$mux  #( .WIDTH(9) ) _50989_ ( .A(_26960_), .B(9'h000), .S(RST), .Y(_03078_) );
  \$mux  #( .WIDTH(9) ) _50990_ ( .A(_tmp_351), .B(_28537_[8:0]), .S(_06602_), .Y(_26961_) );
  \$mux  #( .WIDTH(9) ) _50991_ ( .A(_26961_), .B(_tmp_354), .S(_06605_), .Y(_26962_) );
  \$mux  #( .WIDTH(9) ) _50992_ ( .A(_26962_), .B(9'h000), .S(RST), .Y(_03077_) );
  \$mux  #( .WIDTH(1) ) _50993_ ( .A(_tmp_350), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26963_) );
  \$mux  #( .WIDTH(1) ) _50994_ ( .A(_26963_), .B(1'h1), .S(_06608_), .Y(_26964_) );
  \$mux  #( .WIDTH(1) ) _50995_ ( .A(_26964_), .B(1'h0), .S(RST), .Y(_03076_) );
  \$mux  #( .WIDTH(34) ) _50996_ ( .A(_tmp_349), .B({ 1'h0, _maxi_read_size }), .S(_06602_), .Y(_26965_) );
  \$mux  #( .WIDTH(34) ) _50997_ ( .A(_26965_), .B(_28598_), .S(_06256_), .Y(_26966_) );
  \$mux  #( .WIDTH(34) ) _50998_ ( .A(_26966_), .B(34'h000000000), .S(RST), .Y(_03075_) );
  \$mux  #( .WIDTH(10) ) _50999_ ( .A(_tmp_348), .B(_28596_[9:0]), .S(_06602_), .Y(_26967_) );
  \$mux  #( .WIDTH(10) ) _51000_ ( .A(_26967_), .B(_28597_[9:0]), .S(_06256_), .Y(_26968_) );
  \$mux  #( .WIDTH(10) ) _51001_ ( .A(_26968_), .B(_28596_[9:0]), .S(_06603_), .Y(_26969_) );
  \$mux  #( .WIDTH(10) ) _51002_ ( .A(_26969_), .B(10'h000), .S(RST), .Y(_03074_) );
  \$mux  #( .WIDTH(1) ) _51003_ ( .A(ram_w8_l2048_id5_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26970_) );
  \$mux  #( .WIDTH(1) ) _51004_ ( .A(_26970_), .B(_06113_), .S(_06256_), .Y(_26971_) );
  \$mux  #( .WIDTH(1) ) _51005_ ( .A(_26971_), .B(1'h0), .S(RST), .Y(_03792_) );
  \$mux  #( .WIDTH(8) ) _51006_ ( .A(ram_w8_l2048_id5_0_1_wdata), .B(_dataflow_slice_data_67), .S(_06256_), .Y(_26972_) );
  \$mux  #( .WIDTH(8) ) _51007_ ( .A(_26972_), .B(8'h00), .S(RST), .Y(_03791_) );
  \$mux  #( .WIDTH(9) ) _51008_ ( .A(ram_w8_l2048_id5_0_1_addr), .B(_tmp_354), .S(_06256_), .Y(_26973_) );
  \$mux  #( .WIDTH(9) ) _51009_ ( .A(_26973_), .B(9'h000), .S(RST), .Y(_03790_) );
  \$mux  #( .WIDTH(9) ) _51010_ ( .A(ram_w8_l2048_id5_0_0_addr), .B(_stream_conv2d_16_source_22_source_ram_raddr[10:2]), .S(_tmp_533), .Y(_26974_) );
  \$mux  #( .WIDTH(9) ) _51011_ ( .A(_26974_), .B(9'h000), .S(RST), .Y(_03789_) );
  \$mux  #( .WIDTH(1) ) _51012_ ( .A(ram_w8_l2048_id4_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26975_) );
  \$mux  #( .WIDTH(1) ) _51013_ ( .A(_26975_), .B(_06109_), .S(_06253_), .Y(_26976_) );
  \$mux  #( .WIDTH(1) ) _51014_ ( .A(_26976_), .B(1'h0), .S(RST), .Y(_03788_) );
  \$mux  #( .WIDTH(8) ) _51015_ ( .A(ram_w8_l2048_id4_3_1_wdata), .B(_dataflow_slice_data_63), .S(_06253_), .Y(_26977_) );
  \$mux  #( .WIDTH(8) ) _51016_ ( .A(_26977_), .B(8'h00), .S(RST), .Y(_03787_) );
  \$mux  #( .WIDTH(9) ) _51017_ ( .A(ram_w8_l2048_id4_3_1_addr), .B(_tmp_338), .S(_06253_), .Y(_26978_) );
  \$mux  #( .WIDTH(9) ) _51018_ ( .A(_26978_), .B(9'h000), .S(RST), .Y(_03786_) );
  \$mux  #( .WIDTH(9) ) _51019_ ( .A(ram_w8_l2048_id4_3_0_addr), .B(_stream_conv2d_16_source_21_source_ram_raddr[10:2]), .S(_tmp_523), .Y(_26979_) );
  \$mux  #( .WIDTH(9) ) _51020_ ( .A(_26979_), .B(9'h000), .S(RST), .Y(_03785_) );
  \$mux  #( .WIDTH(1) ) _51021_ ( .A(ram_w8_l2048_id4_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26980_) );
  \$mux  #( .WIDTH(1) ) _51022_ ( .A(_26980_), .B(_06106_), .S(_06250_), .Y(_26981_) );
  \$mux  #( .WIDTH(1) ) _51023_ ( .A(_26981_), .B(1'h0), .S(RST), .Y(_03784_) );
  \$mux  #( .WIDTH(8) ) _51024_ ( .A(ram_w8_l2048_id4_2_1_wdata), .B(_dataflow_slice_data_60), .S(_06250_), .Y(_26982_) );
  \$mux  #( .WIDTH(8) ) _51025_ ( .A(_26982_), .B(8'h00), .S(RST), .Y(_03783_) );
  \$mux  #( .WIDTH(9) ) _51026_ ( .A(ram_w8_l2048_id4_2_1_addr), .B(_tmp_325), .S(_06250_), .Y(_26983_) );
  \$mux  #( .WIDTH(9) ) _51027_ ( .A(_26983_), .B(9'h000), .S(RST), .Y(_03782_) );
  \$mux  #( .WIDTH(9) ) _51028_ ( .A(ram_w8_l2048_id4_2_0_addr), .B(_stream_conv2d_16_source_21_source_ram_raddr[10:2]), .S(_tmp_523), .Y(_26984_) );
  \$mux  #( .WIDTH(9) ) _51029_ ( .A(_26984_), .B(9'h000), .S(RST), .Y(_03781_) );
  \$mux  #( .WIDTH(1) ) _51030_ ( .A(ram_w8_l2048_id4_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26985_) );
  \$mux  #( .WIDTH(1) ) _51031_ ( .A(_26985_), .B(_06103_), .S(_06247_), .Y(_26986_) );
  \$mux  #( .WIDTH(1) ) _51032_ ( .A(_26986_), .B(1'h0), .S(RST), .Y(_03780_) );
  \$mux  #( .WIDTH(8) ) _51033_ ( .A(ram_w8_l2048_id4_1_1_wdata), .B(_dataflow_slice_data_57), .S(_06247_), .Y(_26987_) );
  \$mux  #( .WIDTH(8) ) _51034_ ( .A(_26987_), .B(8'h00), .S(RST), .Y(_03779_) );
  \$mux  #( .WIDTH(9) ) _51035_ ( .A(ram_w8_l2048_id4_1_1_addr), .B(_tmp_312), .S(_06247_), .Y(_26988_) );
  \$mux  #( .WIDTH(9) ) _51036_ ( .A(_26988_), .B(9'h000), .S(RST), .Y(_03778_) );
  \$mux  #( .WIDTH(9) ) _51037_ ( .A(ram_w8_l2048_id4_1_0_addr), .B(_stream_conv2d_16_source_21_source_ram_raddr[10:2]), .S(_tmp_523), .Y(_26989_) );
  \$mux  #( .WIDTH(9) ) _51038_ ( .A(_26989_), .B(9'h000), .S(RST), .Y(_03777_) );
  \$mux  #( .WIDTH(1) ) _51039_ ( .A(_tmp_523), .B(1'h0), .S(RST), .Y(_01243_) );
  \$mux  #( .WIDTH(1) ) _51040_ ( .A(ram_w8_l2048_id4_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26990_) );
  \$mux  #( .WIDTH(1) ) _51041_ ( .A(_26990_), .B(_06100_), .S(_06244_), .Y(_26991_) );
  \$mux  #( .WIDTH(1) ) _51042_ ( .A(_26991_), .B(1'h0), .S(RST), .Y(_03776_) );
  \$mux  #( .WIDTH(8) ) _51043_ ( .A(ram_w8_l2048_id4_0_1_wdata), .B(_dataflow_slice_data_54), .S(_06244_), .Y(_26992_) );
  \$mux  #( .WIDTH(8) ) _51044_ ( .A(_26992_), .B(8'h00), .S(RST), .Y(_03775_) );
  \$mux  #( .WIDTH(9) ) _51045_ ( .A(ram_w8_l2048_id4_0_1_addr), .B(_tmp_299), .S(_06244_), .Y(_26993_) );
  \$mux  #( .WIDTH(9) ) _51046_ ( .A(_26993_), .B(9'h000), .S(RST), .Y(_03774_) );
  \$mux  #( .WIDTH(9) ) _51047_ ( .A(ram_w8_l2048_id4_0_0_addr), .B(_stream_conv2d_16_source_21_source_ram_raddr[10:2]), .S(_tmp_523), .Y(_26994_) );
  \$mux  #( .WIDTH(9) ) _51048_ ( .A(_26994_), .B(9'h000), .S(RST), .Y(_03773_) );
  \$mux  #( .WIDTH(1) ) _51049_ ( .A(_tmp_1162), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26995_) );
  \$mux  #( .WIDTH(1) ) _51050_ ( .A(_26995_), .B(1'h1), .S(_06600_), .Y(_26996_) );
  \$mux  #( .WIDTH(1) ) _51051_ ( .A(_26996_), .B(1'h0), .S(RST), .Y(_02935_) );
  \$mux  #( .WIDTH(34) ) _51052_ ( .A(_tmp_1161), .B({ 1'h0, _maxi_read_size }), .S(_06599_), .Y(_26997_) );
  \$mux  #( .WIDTH(34) ) _51053_ ( .A(_26997_), .B(_28595_), .S(_06325_), .Y(_26998_) );
  \$mux  #( .WIDTH(34) ) _51054_ ( .A(_26998_), .B(34'h000000000), .S(RST), .Y(_02934_) );
  \$mux  #( .WIDTH(1) ) _51055_ ( .A(ram_w8_l2048_id3_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_26999_) );
  \$mux  #( .WIDTH(1) ) _51056_ ( .A(_26999_), .B(_06111_), .S(_06253_), .Y(_27000_) );
  \$mux  #( .WIDTH(1) ) _51057_ ( .A(_27000_), .B(1'h1), .S(_06325_), .Y(_27001_) );
  \$mux  #( .WIDTH(1) ) _51058_ ( .A(_27001_), .B(1'h0), .S(RST), .Y(_03772_) );
  \$mux  #( .WIDTH(8) ) _51059_ ( .A(ram_w8_l2048_id3_3_1_wdata), .B(_dataflow_slice_data_63), .S(_06253_), .Y(_27002_) );
  \$mux  #( .WIDTH(8) ) _51060_ ( .A(_27002_), .B(_dataflow_slice_data_158), .S(_06325_), .Y(_27003_) );
  \$mux  #( .WIDTH(8) ) _51061_ ( .A(_27003_), .B(8'h00), .S(RST), .Y(_03771_) );
  \$mux  #( .WIDTH(9) ) _51062_ ( .A(ram_w8_l2048_id3_3_1_addr), .B(_tmp_337), .S(_06253_), .Y(_27004_) );
  \$mux  #( .WIDTH(9) ) _51063_ ( .A(_27004_), .B(_28537_[8:0]), .S(_06599_), .Y(_27005_) );
  \$mux  #( .WIDTH(9) ) _51064_ ( .A(_27005_), .B(_24277_[8:0]), .S(_06325_), .Y(_27006_) );
  \$mux  #( .WIDTH(9) ) _51065_ ( .A(_27006_), .B(9'h000), .S(RST), .Y(_03770_) );
  \$mux  #( .WIDTH(9) ) _51066_ ( .A(ram_w8_l2048_id3_3_0_addr), .B(_stream_conv2d_16_source_20_source_ram_raddr[10:2]), .S(_tmp_513), .Y(_27007_) );
  \$mux  #( .WIDTH(9) ) _51067_ ( .A(_27007_), .B(_stream_matmul_29_source_19_source_ram_raddr[10:2]), .S(_tmp_1209), .Y(_27008_) );
  \$mux  #( .WIDTH(9) ) _51068_ ( .A(_27008_), .B(9'h000), .S(RST), .Y(_03769_) );
  \$mux  #( .WIDTH(1) ) _51069_ ( .A(_tmp_1160), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27009_) );
  \$mux  #( .WIDTH(1) ) _51070_ ( .A(_27009_), .B(1'h1), .S(_06598_), .Y(_27010_) );
  \$mux  #( .WIDTH(1) ) _51071_ ( .A(_27010_), .B(1'h0), .S(RST), .Y(_02933_) );
  \$mux  #( .WIDTH(34) ) _51072_ ( .A(_tmp_1159), .B({ 1'h0, _maxi_read_size }), .S(_06597_), .Y(_27011_) );
  \$mux  #( .WIDTH(34) ) _51073_ ( .A(_27011_), .B(_28594_), .S(_06322_), .Y(_27012_) );
  \$mux  #( .WIDTH(34) ) _51074_ ( .A(_27012_), .B(34'h000000000), .S(RST), .Y(_02932_) );
  \$mux  #( .WIDTH(1) ) _51075_ ( .A(ram_w8_l2048_id3_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27013_) );
  \$mux  #( .WIDTH(1) ) _51076_ ( .A(_27013_), .B(_06108_), .S(_06250_), .Y(_27014_) );
  \$mux  #( .WIDTH(1) ) _51077_ ( .A(_27014_), .B(1'h1), .S(_06322_), .Y(_27015_) );
  \$mux  #( .WIDTH(1) ) _51078_ ( .A(_27015_), .B(1'h0), .S(RST), .Y(_03768_) );
  \$mux  #( .WIDTH(8) ) _51079_ ( .A(ram_w8_l2048_id3_2_1_wdata), .B(_dataflow_slice_data_60), .S(_06250_), .Y(_27016_) );
  \$mux  #( .WIDTH(8) ) _51080_ ( .A(_27016_), .B(_dataflow_slice_data_155), .S(_06322_), .Y(_27017_) );
  \$mux  #( .WIDTH(8) ) _51081_ ( .A(_27017_), .B(8'h00), .S(RST), .Y(_03767_) );
  \$mux  #( .WIDTH(9) ) _51082_ ( .A(ram_w8_l2048_id3_2_1_addr), .B(_tmp_324), .S(_06250_), .Y(_27018_) );
  \$mux  #( .WIDTH(9) ) _51083_ ( .A(_27018_), .B(_28537_[8:0]), .S(_06597_), .Y(_27019_) );
  \$mux  #( .WIDTH(9) ) _51084_ ( .A(_27019_), .B(_24276_[8:0]), .S(_06322_), .Y(_27020_) );
  \$mux  #( .WIDTH(9) ) _51085_ ( .A(_27020_), .B(9'h000), .S(RST), .Y(_03766_) );
  \$mux  #( .WIDTH(9) ) _51086_ ( .A(ram_w8_l2048_id3_2_0_addr), .B(_stream_conv2d_16_source_20_source_ram_raddr[10:2]), .S(_tmp_513), .Y(_27021_) );
  \$mux  #( .WIDTH(9) ) _51087_ ( .A(_27021_), .B(_stream_matmul_29_source_19_source_ram_raddr[10:2]), .S(_tmp_1209), .Y(_27022_) );
  \$mux  #( .WIDTH(9) ) _51088_ ( .A(_27022_), .B(9'h000), .S(RST), .Y(_03765_) );
  \$mux  #( .WIDTH(1) ) _51089_ ( .A(_tmp_1158), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27023_) );
  \$mux  #( .WIDTH(1) ) _51090_ ( .A(_27023_), .B(1'h1), .S(_06596_), .Y(_27024_) );
  \$mux  #( .WIDTH(1) ) _51091_ ( .A(_27024_), .B(1'h0), .S(RST), .Y(_02931_) );
  \$mux  #( .WIDTH(34) ) _51092_ ( .A(_tmp_1157), .B({ 1'h0, _maxi_read_size }), .S(_06595_), .Y(_27025_) );
  \$mux  #( .WIDTH(34) ) _51093_ ( .A(_27025_), .B(_28593_), .S(_06319_), .Y(_27026_) );
  \$mux  #( .WIDTH(34) ) _51094_ ( .A(_27026_), .B(34'h000000000), .S(RST), .Y(_02930_) );
  \$mux  #( .WIDTH(1) ) _51095_ ( .A(ram_w8_l2048_id3_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27027_) );
  \$mux  #( .WIDTH(1) ) _51096_ ( .A(_27027_), .B(_06105_), .S(_06247_), .Y(_27028_) );
  \$mux  #( .WIDTH(1) ) _51097_ ( .A(_27028_), .B(1'h1), .S(_06319_), .Y(_27029_) );
  \$mux  #( .WIDTH(1) ) _51098_ ( .A(_27029_), .B(1'h0), .S(RST), .Y(_03764_) );
  \$mux  #( .WIDTH(8) ) _51099_ ( .A(ram_w8_l2048_id3_1_1_wdata), .B(_dataflow_slice_data_57), .S(_06247_), .Y(_27030_) );
  \$mux  #( .WIDTH(8) ) _51100_ ( .A(_27030_), .B(_dataflow_slice_data_152), .S(_06319_), .Y(_27031_) );
  \$mux  #( .WIDTH(8) ) _51101_ ( .A(_27031_), .B(8'h00), .S(RST), .Y(_03763_) );
  \$mux  #( .WIDTH(9) ) _51102_ ( .A(ram_w8_l2048_id3_1_1_addr), .B(_tmp_311), .S(_06247_), .Y(_27032_) );
  \$mux  #( .WIDTH(9) ) _51103_ ( .A(_27032_), .B(_28537_[8:0]), .S(_06595_), .Y(_27033_) );
  \$mux  #( .WIDTH(9) ) _51104_ ( .A(_27033_), .B(_24275_[8:0]), .S(_06319_), .Y(_27034_) );
  \$mux  #( .WIDTH(9) ) _51105_ ( .A(_27034_), .B(9'h000), .S(RST), .Y(_03762_) );
  \$mux  #( .WIDTH(9) ) _51106_ ( .A(ram_w8_l2048_id3_1_0_addr), .B(_stream_conv2d_16_source_20_source_ram_raddr[10:2]), .S(_tmp_513), .Y(_27035_) );
  \$mux  #( .WIDTH(9) ) _51107_ ( .A(_27035_), .B(_stream_matmul_29_source_19_source_ram_raddr[10:2]), .S(_tmp_1209), .Y(_27036_) );
  \$mux  #( .WIDTH(9) ) _51108_ ( .A(_27036_), .B(9'h000), .S(RST), .Y(_03761_) );
  \$mux  #( .WIDTH(1) ) _51109_ ( .A(_tmp_1209), .B(1'h0), .S(RST), .Y(_01147_) );
  \$mux  #( .WIDTH(1) ) _51110_ ( .A(_tmp_1156), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27037_) );
  \$mux  #( .WIDTH(1) ) _51111_ ( .A(_27037_), .B(1'h1), .S(_06594_), .Y(_27038_) );
  \$mux  #( .WIDTH(1) ) _51112_ ( .A(_27038_), .B(1'h0), .S(RST), .Y(_02929_) );
  \$mux  #( .WIDTH(34) ) _51113_ ( .A(_tmp_1155), .B({ 1'h0, _maxi_read_size }), .S(_06593_), .Y(_27039_) );
  \$mux  #( .WIDTH(34) ) _51114_ ( .A(_27039_), .B(_28592_), .S(_06316_), .Y(_27040_) );
  \$mux  #( .WIDTH(34) ) _51115_ ( .A(_27040_), .B(34'h000000000), .S(RST), .Y(_02928_) );
  \$mux  #( .WIDTH(1) ) _51116_ ( .A(_tmp_513), .B(1'h0), .S(RST), .Y(_01240_) );
  \$mux  #( .WIDTH(1) ) _51117_ ( .A(ram_w8_l2048_id3_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27041_) );
  \$mux  #( .WIDTH(1) ) _51118_ ( .A(_27041_), .B(_06102_), .S(_06244_), .Y(_27042_) );
  \$mux  #( .WIDTH(1) ) _51119_ ( .A(_27042_), .B(1'h1), .S(_06316_), .Y(_27043_) );
  \$mux  #( .WIDTH(1) ) _51120_ ( .A(_27043_), .B(1'h0), .S(RST), .Y(_03760_) );
  \$mux  #( .WIDTH(8) ) _51121_ ( .A(ram_w8_l2048_id3_0_1_wdata), .B(_dataflow_slice_data_54), .S(_06244_), .Y(_27044_) );
  \$mux  #( .WIDTH(8) ) _51122_ ( .A(_27044_), .B(_dataflow_slice_data_149), .S(_06316_), .Y(_27045_) );
  \$mux  #( .WIDTH(8) ) _51123_ ( .A(_27045_), .B(8'h00), .S(RST), .Y(_03759_) );
  \$mux  #( .WIDTH(9) ) _51124_ ( .A(ram_w8_l2048_id3_0_1_addr), .B(_tmp_298), .S(_06244_), .Y(_27046_) );
  \$mux  #( .WIDTH(9) ) _51125_ ( .A(_27046_), .B(_28537_[8:0]), .S(_06593_), .Y(_27047_) );
  \$mux  #( .WIDTH(9) ) _51126_ ( .A(_27047_), .B(_24274_[8:0]), .S(_06316_), .Y(_27048_) );
  \$mux  #( .WIDTH(9) ) _51127_ ( .A(_27048_), .B(9'h000), .S(RST), .Y(_03758_) );
  \$mux  #( .WIDTH(9) ) _51128_ ( .A(ram_w8_l2048_id3_0_0_addr), .B(_stream_conv2d_16_source_20_source_ram_raddr[10:2]), .S(_tmp_513), .Y(_27049_) );
  \$mux  #( .WIDTH(9) ) _51129_ ( .A(_27049_), .B(_stream_matmul_29_source_19_source_ram_raddr[10:2]), .S(_tmp_1209), .Y(_27050_) );
  \$mux  #( .WIDTH(9) ) _51130_ ( .A(_27050_), .B(9'h000), .S(RST), .Y(_03757_) );
  \$mux  #( .WIDTH(1) ) _51131_ ( .A(_tmp_1131), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27051_) );
  \$mux  #( .WIDTH(1) ) _51132_ ( .A(_27051_), .B(1'h1), .S(_06591_), .Y(_27052_) );
  \$mux  #( .WIDTH(1) ) _51133_ ( .A(_27052_), .B(1'h0), .S(RST), .Y(_02911_) );
  \$mux  #( .WIDTH(34) ) _51134_ ( .A(_tmp_1130), .B({ 1'h0, _maxi_read_size }), .S(_06590_), .Y(_27053_) );
  \$mux  #( .WIDTH(34) ) _51135_ ( .A(_27053_), .B(_28591_), .S(_06289_), .Y(_27054_) );
  \$mux  #( .WIDTH(34) ) _51136_ ( .A(_27054_), .B(34'h000000000), .S(RST), .Y(_02910_) );
  \$mux  #( .WIDTH(2) ) _51137_ ( .A(_tmp_342), .B(2'h0), .S(_06583_), .Y(_27055_) );
  \$mux  #( .WIDTH(2) ) _51138_ ( .A(_27055_), .B(_24272_[1:0]), .S(_06584_), .Y(_27056_) );
  \$mux  #( .WIDTH(2) ) _51139_ ( .A(_27056_), .B(2'h0), .S(_06585_), .Y(_27057_) );
  \$mux  #( .WIDTH(2) ) _51140_ ( .A(_27057_), .B(2'h0), .S(RST), .Y(_03073_) );
  \$mux  #( .WIDTH(9) ) _51141_ ( .A(_tmp_335), .B(_28537_[8:0]), .S(_06583_), .Y(_27058_) );
  \$mux  #( .WIDTH(9) ) _51142_ ( .A(_27058_), .B(_tmp_338), .S(_06588_), .Y(_27059_) );
  \$mux  #( .WIDTH(9) ) _51143_ ( .A(_27059_), .B(9'h000), .S(RST), .Y(_03072_) );
  \$mux  #( .WIDTH(9) ) _51144_ ( .A(_tmp_334), .B(_28537_[8:0]), .S(_06583_), .Y(_27060_) );
  \$mux  #( .WIDTH(9) ) _51145_ ( .A(_27060_), .B(_tmp_337), .S(_06587_), .Y(_27061_) );
  \$mux  #( .WIDTH(9) ) _51146_ ( .A(_27061_), .B(9'h000), .S(RST), .Y(_03071_) );
  \$mux  #( .WIDTH(9) ) _51147_ ( .A(_tmp_333), .B(_28537_[8:0]), .S(_06583_), .Y(_27062_) );
  \$mux  #( .WIDTH(9) ) _51148_ ( .A(_27062_), .B(_tmp_336), .S(_06586_), .Y(_27063_) );
  \$mux  #( .WIDTH(9) ) _51149_ ( .A(_27063_), .B(9'h000), .S(RST), .Y(_03070_) );
  \$mux  #( .WIDTH(1) ) _51150_ ( .A(_tmp_332), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27064_) );
  \$mux  #( .WIDTH(1) ) _51151_ ( .A(_27064_), .B(1'h1), .S(_06589_), .Y(_27065_) );
  \$mux  #( .WIDTH(1) ) _51152_ ( .A(_27065_), .B(1'h0), .S(RST), .Y(_03069_) );
  \$mux  #( .WIDTH(34) ) _51153_ ( .A(_tmp_331), .B({ 1'h0, _maxi_read_size }), .S(_06583_), .Y(_27066_) );
  \$mux  #( .WIDTH(34) ) _51154_ ( .A(_27066_), .B(_28590_), .S(_06253_), .Y(_27067_) );
  \$mux  #( .WIDTH(34) ) _51155_ ( .A(_27067_), .B(34'h000000000), .S(RST), .Y(_03068_) );
  \$mux  #( .WIDTH(10) ) _51156_ ( .A(_tmp_330), .B(_28579_[9:0]), .S(_06583_), .Y(_27068_) );
  \$mux  #( .WIDTH(10) ) _51157_ ( .A(_27068_), .B(_28589_[9:0]), .S(_06253_), .Y(_27069_) );
  \$mux  #( .WIDTH(10) ) _51158_ ( .A(_27069_), .B(_28579_[9:0]), .S(_06584_), .Y(_27070_) );
  \$mux  #( .WIDTH(10) ) _51159_ ( .A(_27070_), .B(10'h000), .S(RST), .Y(_03067_) );
  \$mux  #( .WIDTH(1) ) _51160_ ( .A(ram_w8_l2048_id2_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27071_) );
  \$mux  #( .WIDTH(1) ) _51161_ ( .A(_27071_), .B(_06110_), .S(_06253_), .Y(_27072_) );
  \$mux  #( .WIDTH(1) ) _51162_ ( .A(_27072_), .B(1'h1), .S(_06289_), .Y(_27073_) );
  \$mux  #( .WIDTH(1) ) _51163_ ( .A(_27073_), .B(1'h0), .S(RST), .Y(_03756_) );
  \$mux  #( .WIDTH(8) ) _51164_ ( .A(ram_w8_l2048_id2_3_1_wdata), .B(_dataflow_slice_data_63), .S(_06253_), .Y(_27074_) );
  \$mux  #( .WIDTH(8) ) _51165_ ( .A(_27074_), .B(_dataflow_slice_data_120), .S(_06289_), .Y(_27075_) );
  \$mux  #( .WIDTH(8) ) _51166_ ( .A(_27075_), .B(8'h00), .S(RST), .Y(_03755_) );
  \$mux  #( .WIDTH(9) ) _51167_ ( .A(ram_w8_l2048_id2_3_1_addr), .B(_tmp_336), .S(_06253_), .Y(_27076_) );
  \$mux  #( .WIDTH(9) ) _51168_ ( .A(_27076_), .B(_28537_[8:0]), .S(_06590_), .Y(_27077_) );
  \$mux  #( .WIDTH(9) ) _51169_ ( .A(_27077_), .B(_24273_[8:0]), .S(_06289_), .Y(_27078_) );
  \$mux  #( .WIDTH(9) ) _51170_ ( .A(_27078_), .B(9'h000), .S(RST), .Y(_03754_) );
  \$mux  #( .WIDTH(9) ) _51171_ ( .A(ram_w8_l2048_id2_3_0_addr), .B(_stream_conv2d_16_source_19_source_ram_raddr[10:2]), .S(_tmp_503), .Y(_27079_) );
  \$mux  #( .WIDTH(9) ) _51172_ ( .A(_27079_), .B(_stream_matmul_29_source_6_source_ram_raddr[10:2]), .S(_tmp_1178), .Y(_27080_) );
  \$mux  #( .WIDTH(9) ) _51173_ ( .A(_27080_), .B(9'h000), .S(RST), .Y(_03753_) );
  \$mux  #( .WIDTH(1) ) _51174_ ( .A(_tmp_1129), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27081_) );
  \$mux  #( .WIDTH(1) ) _51175_ ( .A(_27081_), .B(1'h1), .S(_06582_), .Y(_27082_) );
  \$mux  #( .WIDTH(1) ) _51176_ ( .A(_27082_), .B(1'h0), .S(RST), .Y(_02909_) );
  \$mux  #( .WIDTH(34) ) _51177_ ( .A(_tmp_1128), .B({ 1'h0, _maxi_read_size }), .S(_06581_), .Y(_27083_) );
  \$mux  #( .WIDTH(34) ) _51178_ ( .A(_27083_), .B(_28588_), .S(_06286_), .Y(_27084_) );
  \$mux  #( .WIDTH(34) ) _51179_ ( .A(_27084_), .B(34'h000000000), .S(RST), .Y(_02908_) );
  \$mux  #( .WIDTH(2) ) _51180_ ( .A(_tmp_329), .B(2'h0), .S(_06574_), .Y(_27085_) );
  \$mux  #( .WIDTH(2) ) _51181_ ( .A(_27085_), .B(_24270_[1:0]), .S(_06575_), .Y(_27086_) );
  \$mux  #( .WIDTH(2) ) _51182_ ( .A(_27086_), .B(2'h0), .S(_06576_), .Y(_27087_) );
  \$mux  #( .WIDTH(2) ) _51183_ ( .A(_27087_), .B(2'h0), .S(RST), .Y(_03065_) );
  \$mux  #( .WIDTH(9) ) _51184_ ( .A(_tmp_322), .B(_28537_[8:0]), .S(_06574_), .Y(_27088_) );
  \$mux  #( .WIDTH(9) ) _51185_ ( .A(_27088_), .B(_tmp_325), .S(_06579_), .Y(_27089_) );
  \$mux  #( .WIDTH(9) ) _51186_ ( .A(_27089_), .B(9'h000), .S(RST), .Y(_03064_) );
  \$mux  #( .WIDTH(9) ) _51187_ ( .A(_tmp_321), .B(_28537_[8:0]), .S(_06574_), .Y(_27090_) );
  \$mux  #( .WIDTH(9) ) _51188_ ( .A(_27090_), .B(_tmp_324), .S(_06578_), .Y(_27091_) );
  \$mux  #( .WIDTH(9) ) _51189_ ( .A(_27091_), .B(9'h000), .S(RST), .Y(_03063_) );
  \$mux  #( .WIDTH(9) ) _51190_ ( .A(_tmp_320), .B(_28537_[8:0]), .S(_06574_), .Y(_27092_) );
  \$mux  #( .WIDTH(9) ) _51191_ ( .A(_27092_), .B(_tmp_323), .S(_06577_), .Y(_27093_) );
  \$mux  #( .WIDTH(9) ) _51192_ ( .A(_27093_), .B(9'h000), .S(RST), .Y(_03062_) );
  \$mux  #( .WIDTH(1) ) _51193_ ( .A(_tmp_319), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27094_) );
  \$mux  #( .WIDTH(1) ) _51194_ ( .A(_27094_), .B(1'h1), .S(_06580_), .Y(_27095_) );
  \$mux  #( .WIDTH(1) ) _51195_ ( .A(_27095_), .B(1'h0), .S(RST), .Y(_03060_) );
  \$mux  #( .WIDTH(34) ) _51196_ ( .A(_tmp_318), .B({ 1'h0, _maxi_read_size }), .S(_06574_), .Y(_27096_) );
  \$mux  #( .WIDTH(34) ) _51197_ ( .A(_27096_), .B(_28587_), .S(_06250_), .Y(_27097_) );
  \$mux  #( .WIDTH(34) ) _51198_ ( .A(_27097_), .B(34'h000000000), .S(RST), .Y(_03059_) );
  \$mux  #( .WIDTH(10) ) _51199_ ( .A(_tmp_317), .B(_28579_[9:0]), .S(_06574_), .Y(_27098_) );
  \$mux  #( .WIDTH(10) ) _51200_ ( .A(_27098_), .B(_28586_[9:0]), .S(_06250_), .Y(_27099_) );
  \$mux  #( .WIDTH(10) ) _51201_ ( .A(_27099_), .B(_28579_[9:0]), .S(_06575_), .Y(_27100_) );
  \$mux  #( .WIDTH(10) ) _51202_ ( .A(_27100_), .B(10'h000), .S(RST), .Y(_03058_) );
  \$mux  #( .WIDTH(1) ) _51203_ ( .A(ram_w8_l2048_id2_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27101_) );
  \$mux  #( .WIDTH(1) ) _51204_ ( .A(_27101_), .B(_06107_), .S(_06250_), .Y(_27102_) );
  \$mux  #( .WIDTH(1) ) _51205_ ( .A(_27102_), .B(1'h1), .S(_06286_), .Y(_27103_) );
  \$mux  #( .WIDTH(1) ) _51206_ ( .A(_27103_), .B(1'h0), .S(RST), .Y(_03752_) );
  \$mux  #( .WIDTH(8) ) _51207_ ( .A(ram_w8_l2048_id2_2_1_wdata), .B(_dataflow_slice_data_60), .S(_06250_), .Y(_27104_) );
  \$mux  #( .WIDTH(8) ) _51208_ ( .A(_27104_), .B(_dataflow_slice_data_117), .S(_06286_), .Y(_27105_) );
  \$mux  #( .WIDTH(8) ) _51209_ ( .A(_27105_), .B(8'h00), .S(RST), .Y(_03751_) );
  \$mux  #( .WIDTH(9) ) _51210_ ( .A(ram_w8_l2048_id2_2_1_addr), .B(_tmp_323), .S(_06250_), .Y(_27106_) );
  \$mux  #( .WIDTH(9) ) _51211_ ( .A(_27106_), .B(_28537_[8:0]), .S(_06581_), .Y(_27107_) );
  \$mux  #( .WIDTH(9) ) _51212_ ( .A(_27107_), .B(_24271_[8:0]), .S(_06286_), .Y(_27108_) );
  \$mux  #( .WIDTH(9) ) _51213_ ( .A(_27108_), .B(9'h000), .S(RST), .Y(_03750_) );
  \$mux  #( .WIDTH(9) ) _51214_ ( .A(ram_w8_l2048_id2_2_0_addr), .B(_stream_conv2d_16_source_19_source_ram_raddr[10:2]), .S(_tmp_503), .Y(_27109_) );
  \$mux  #( .WIDTH(9) ) _51215_ ( .A(_27109_), .B(_stream_matmul_29_source_6_source_ram_raddr[10:2]), .S(_tmp_1178), .Y(_27110_) );
  \$mux  #( .WIDTH(9) ) _51216_ ( .A(_27110_), .B(9'h000), .S(RST), .Y(_03749_) );
  \$mux  #( .WIDTH(1) ) _51217_ ( .A(_tmp_1127), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27111_) );
  \$mux  #( .WIDTH(1) ) _51218_ ( .A(_27111_), .B(1'h1), .S(_06573_), .Y(_27112_) );
  \$mux  #( .WIDTH(1) ) _51219_ ( .A(_27112_), .B(1'h0), .S(RST), .Y(_02907_) );
  \$mux  #( .WIDTH(34) ) _51220_ ( .A(_tmp_1126), .B({ 1'h0, _maxi_read_size }), .S(_06572_), .Y(_27113_) );
  \$mux  #( .WIDTH(34) ) _51221_ ( .A(_27113_), .B(_28585_), .S(_06283_), .Y(_27114_) );
  \$mux  #( .WIDTH(34) ) _51222_ ( .A(_27114_), .B(34'h000000000), .S(RST), .Y(_02906_) );
  \$mux  #( .WIDTH(2) ) _51223_ ( .A(_tmp_316), .B(2'h0), .S(_06565_), .Y(_27115_) );
  \$mux  #( .WIDTH(2) ) _51224_ ( .A(_27115_), .B(_24268_[1:0]), .S(_06566_), .Y(_27116_) );
  \$mux  #( .WIDTH(2) ) _51225_ ( .A(_27116_), .B(2'h0), .S(_06567_), .Y(_27117_) );
  \$mux  #( .WIDTH(2) ) _51226_ ( .A(_27117_), .B(2'h0), .S(RST), .Y(_03057_) );
  \$mux  #( .WIDTH(9) ) _51227_ ( .A(_tmp_309), .B(_28537_[8:0]), .S(_06565_), .Y(_27118_) );
  \$mux  #( .WIDTH(9) ) _51228_ ( .A(_27118_), .B(_tmp_312), .S(_06570_), .Y(_27119_) );
  \$mux  #( .WIDTH(9) ) _51229_ ( .A(_27119_), .B(9'h000), .S(RST), .Y(_03055_) );
  \$mux  #( .WIDTH(9) ) _51230_ ( .A(_tmp_308), .B(_28537_[8:0]), .S(_06565_), .Y(_27120_) );
  \$mux  #( .WIDTH(9) ) _51231_ ( .A(_27120_), .B(_tmp_311), .S(_06569_), .Y(_27121_) );
  \$mux  #( .WIDTH(9) ) _51232_ ( .A(_27121_), .B(9'h000), .S(RST), .Y(_03054_) );
  \$mux  #( .WIDTH(9) ) _51233_ ( .A(_tmp_307), .B(_28537_[8:0]), .S(_06565_), .Y(_27122_) );
  \$mux  #( .WIDTH(9) ) _51234_ ( .A(_27122_), .B(_tmp_310), .S(_06568_), .Y(_27123_) );
  \$mux  #( .WIDTH(9) ) _51235_ ( .A(_27123_), .B(9'h000), .S(RST), .Y(_03053_) );
  \$mux  #( .WIDTH(1) ) _51236_ ( .A(_tmp_306), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27124_) );
  \$mux  #( .WIDTH(1) ) _51237_ ( .A(_27124_), .B(1'h1), .S(_06571_), .Y(_27125_) );
  \$mux  #( .WIDTH(1) ) _51238_ ( .A(_27125_), .B(1'h0), .S(RST), .Y(_03052_) );
  \$mux  #( .WIDTH(34) ) _51239_ ( .A(_tmp_305), .B({ 1'h0, _maxi_read_size }), .S(_06565_), .Y(_27126_) );
  \$mux  #( .WIDTH(34) ) _51240_ ( .A(_27126_), .B(_28584_), .S(_06247_), .Y(_27127_) );
  \$mux  #( .WIDTH(34) ) _51241_ ( .A(_27127_), .B(34'h000000000), .S(RST), .Y(_03051_) );
  \$mux  #( .WIDTH(10) ) _51242_ ( .A(_tmp_304), .B(_28579_[9:0]), .S(_06565_), .Y(_27128_) );
  \$mux  #( .WIDTH(10) ) _51243_ ( .A(_27128_), .B(_28583_[9:0]), .S(_06247_), .Y(_27129_) );
  \$mux  #( .WIDTH(10) ) _51244_ ( .A(_27129_), .B(_28579_[9:0]), .S(_06566_), .Y(_27130_) );
  \$mux  #( .WIDTH(10) ) _51245_ ( .A(_27130_), .B(10'h000), .S(RST), .Y(_03050_) );
  \$mux  #( .WIDTH(1) ) _51246_ ( .A(ram_w8_l2048_id2_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27131_) );
  \$mux  #( .WIDTH(1) ) _51247_ ( .A(_27131_), .B(_06104_), .S(_06247_), .Y(_27132_) );
  \$mux  #( .WIDTH(1) ) _51248_ ( .A(_27132_), .B(1'h1), .S(_06283_), .Y(_27133_) );
  \$mux  #( .WIDTH(1) ) _51249_ ( .A(_27133_), .B(1'h0), .S(RST), .Y(_03748_) );
  \$mux  #( .WIDTH(8) ) _51250_ ( .A(ram_w8_l2048_id2_1_1_wdata), .B(_dataflow_slice_data_57), .S(_06247_), .Y(_27134_) );
  \$mux  #( .WIDTH(8) ) _51251_ ( .A(_27134_), .B(_dataflow_slice_data_114), .S(_06283_), .Y(_27135_) );
  \$mux  #( .WIDTH(8) ) _51252_ ( .A(_27135_), .B(8'h00), .S(RST), .Y(_03747_) );
  \$mux  #( .WIDTH(9) ) _51253_ ( .A(ram_w8_l2048_id2_1_1_addr), .B(_tmp_310), .S(_06247_), .Y(_27136_) );
  \$mux  #( .WIDTH(9) ) _51254_ ( .A(_27136_), .B(_28537_[8:0]), .S(_06572_), .Y(_27137_) );
  \$mux  #( .WIDTH(9) ) _51255_ ( .A(_27137_), .B(_24269_[8:0]), .S(_06283_), .Y(_27138_) );
  \$mux  #( .WIDTH(9) ) _51256_ ( .A(_27138_), .B(9'h000), .S(RST), .Y(_03746_) );
  \$mux  #( .WIDTH(9) ) _51257_ ( .A(ram_w8_l2048_id2_1_0_addr), .B(_stream_conv2d_16_source_19_source_ram_raddr[10:2]), .S(_tmp_503), .Y(_27139_) );
  \$mux  #( .WIDTH(9) ) _51258_ ( .A(_27139_), .B(_stream_matmul_29_source_6_source_ram_raddr[10:2]), .S(_tmp_1178), .Y(_27140_) );
  \$mux  #( .WIDTH(9) ) _51259_ ( .A(_27140_), .B(9'h000), .S(RST), .Y(_03745_) );
  \$mux  #( .WIDTH(1) ) _51260_ ( .A(_tmp_1178), .B(1'h0), .S(RST), .Y(_01141_) );
  \$mux  #( .WIDTH(1) ) _51261_ ( .A(_tmp_1125), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27141_) );
  \$mux  #( .WIDTH(1) ) _51262_ ( .A(_27141_), .B(1'h1), .S(_06564_), .Y(_27142_) );
  \$mux  #( .WIDTH(1) ) _51263_ ( .A(_27142_), .B(1'h0), .S(RST), .Y(_02905_) );
  \$mux  #( .WIDTH(34) ) _51264_ ( .A(_tmp_1124), .B({ 1'h0, _maxi_read_size }), .S(_06563_), .Y(_27143_) );
  \$mux  #( .WIDTH(34) ) _51265_ ( .A(_27143_), .B(_28582_), .S(_06280_), .Y(_27144_) );
  \$mux  #( .WIDTH(34) ) _51266_ ( .A(_27144_), .B(34'h000000000), .S(RST), .Y(_02904_) );
  \$mux  #( .WIDTH(1) ) _51267_ ( .A(_tmp_503), .B(1'h0), .S(RST), .Y(_01237_) );
  \$mux  #( .WIDTH(2) ) _51268_ ( .A(_tmp_303), .B(2'h0), .S(_06555_), .Y(_27145_) );
  \$mux  #( .WIDTH(2) ) _51269_ ( .A(_27145_), .B(_24266_[1:0]), .S(_06556_), .Y(_27146_) );
  \$mux  #( .WIDTH(2) ) _51270_ ( .A(_27146_), .B(2'h0), .S(_06557_), .Y(_27147_) );
  \$mux  #( .WIDTH(2) ) _51271_ ( .A(_27147_), .B(2'h0), .S(RST), .Y(_03049_) );
  \$mux  #( .WIDTH(9) ) _51272_ ( .A(_tmp_296), .B(_28537_[8:0]), .S(_06555_), .Y(_27148_) );
  \$mux  #( .WIDTH(9) ) _51273_ ( .A(_27148_), .B(_tmp_299), .S(_06560_), .Y(_27149_) );
  \$mux  #( .WIDTH(9) ) _51274_ ( .A(_27149_), .B(9'h000), .S(RST), .Y(_03046_) );
  \$mux  #( .WIDTH(9) ) _51275_ ( .A(_tmp_295), .B(_28537_[8:0]), .S(_06555_), .Y(_27150_) );
  \$mux  #( .WIDTH(9) ) _51276_ ( .A(_27150_), .B(_tmp_298), .S(_06559_), .Y(_27151_) );
  \$mux  #( .WIDTH(9) ) _51277_ ( .A(_27151_), .B(9'h000), .S(RST), .Y(_03045_) );
  \$mux  #( .WIDTH(9) ) _51278_ ( .A(_tmp_294), .B(_28537_[8:0]), .S(_06555_), .Y(_27152_) );
  \$mux  #( .WIDTH(9) ) _51279_ ( .A(_27152_), .B(_tmp_297), .S(_06558_), .Y(_27153_) );
  \$mux  #( .WIDTH(9) ) _51280_ ( .A(_27153_), .B(9'h000), .S(RST), .Y(_03044_) );
  \$mux  #( .WIDTH(1) ) _51281_ ( .A(_tmp_293), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27154_) );
  \$mux  #( .WIDTH(1) ) _51282_ ( .A(_27154_), .B(1'h1), .S(_06561_), .Y(_27155_) );
  \$mux  #( .WIDTH(1) ) _51283_ ( .A(_27155_), .B(1'h0), .S(RST), .Y(_03043_) );
  \$mux  #( .WIDTH(34) ) _51284_ ( .A(_tmp_292), .B({ 1'h0, _maxi_read_size }), .S(_06555_), .Y(_27156_) );
  \$mux  #( .WIDTH(34) ) _51285_ ( .A(_27156_), .B(_28581_), .S(_06244_), .Y(_27157_) );
  \$mux  #( .WIDTH(34) ) _51286_ ( .A(_27157_), .B(34'h000000000), .S(RST), .Y(_03042_) );
  \$mux  #( .WIDTH(10) ) _51287_ ( .A(_tmp_291), .B(_28579_[9:0]), .S(_06555_), .Y(_27158_) );
  \$mux  #( .WIDTH(10) ) _51288_ ( .A(_27158_), .B(_28580_[9:0]), .S(_06244_), .Y(_27159_) );
  \$mux  #( .WIDTH(10) ) _51289_ ( .A(_27159_), .B(_28579_[9:0]), .S(_06556_), .Y(_27160_) );
  \$mux  #( .WIDTH(10) ) _51290_ ( .A(_27160_), .B(10'h000), .S(RST), .Y(_03041_) );
  \$mux  #( .WIDTH(1) ) _51291_ ( .A(ram_w8_l2048_id2_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27161_) );
  \$mux  #( .WIDTH(1) ) _51292_ ( .A(_27161_), .B(_06101_), .S(_06244_), .Y(_27162_) );
  \$mux  #( .WIDTH(1) ) _51293_ ( .A(_27162_), .B(1'h1), .S(_06280_), .Y(_27163_) );
  \$mux  #( .WIDTH(1) ) _51294_ ( .A(_27163_), .B(1'h0), .S(RST), .Y(_03744_) );
  \$mux  #( .WIDTH(8) ) _51295_ ( .A(ram_w8_l2048_id2_0_1_wdata), .B(_dataflow_slice_data_54), .S(_06244_), .Y(_27164_) );
  \$mux  #( .WIDTH(8) ) _51296_ ( .A(_27164_), .B(_dataflow_slice_data_111), .S(_06280_), .Y(_27165_) );
  \$mux  #( .WIDTH(8) ) _51297_ ( .A(_27165_), .B(8'h00), .S(RST), .Y(_03743_) );
  \$mux  #( .WIDTH(9) ) _51298_ ( .A(ram_w8_l2048_id2_0_1_addr), .B(_tmp_297), .S(_06244_), .Y(_27166_) );
  \$mux  #( .WIDTH(9) ) _51299_ ( .A(_27166_), .B(_28537_[8:0]), .S(_06563_), .Y(_27167_) );
  \$mux  #( .WIDTH(9) ) _51300_ ( .A(_27167_), .B(_24267_[8:0]), .S(_06280_), .Y(_27168_) );
  \$mux  #( .WIDTH(9) ) _51301_ ( .A(_27168_), .B(9'h000), .S(RST), .Y(_03742_) );
  \$mux  #( .WIDTH(9) ) _51302_ ( .A(ram_w8_l2048_id2_0_0_addr), .B(_stream_conv2d_16_source_19_source_ram_raddr[10:2]), .S(_tmp_503), .Y(_27169_) );
  \$mux  #( .WIDTH(9) ) _51303_ ( .A(_27169_), .B(_stream_matmul_29_source_6_source_ram_raddr[10:2]), .S(_tmp_1178), .Y(_27170_) );
  \$mux  #( .WIDTH(9) ) _51304_ ( .A(_27170_), .B(9'h000), .S(RST), .Y(_03741_) );
  \$mux  #( .WIDTH(34) ) _51305_ ( .A(_tmp_1356), .B(_28563_), .S(_06551_), .Y(_27171_) );
  \$mux  #( .WIDTH(34) ) _51306_ ( .A(_27171_), .B(_28578_), .S(_06552_), .Y(_27172_) );
  \$mux  #( .WIDTH(34) ) _51307_ ( .A(_27172_), .B(34'h000000000), .S(RST), .Y(_02965_) );
  \$mux  #( .WIDTH(1) ) _51308_ ( .A(_tmp_1355), .B(1'h0), .S(_06549_), .Y(_27173_) );
  \$mux  #( .WIDTH(1) ) _51309_ ( .A(_27173_), .B(_tmp_1354), .S(_06550_), .Y(_27174_) );
  \$mux  #( .WIDTH(1) ) _51310_ ( .A(_27174_), .B(1'h0), .S(RST), .Y(_02964_) );
  \$mux  #( .WIDTH(1) ) _51311_ ( .A(_tmp_1354), .B(1'h0), .S(_06550_), .Y(_27175_) );
  \$mux  #( .WIDTH(1) ) _51312_ ( .A(_27175_), .B(_06099_), .S(_06551_), .Y(_27176_) );
  \$mux  #( .WIDTH(1) ) _51313_ ( .A(_27176_), .B(1'h0), .S(_06552_), .Y(_27177_) );
  \$mux  #( .WIDTH(1) ) _51314_ ( .A(_27177_), .B(1'h1), .S(_06553_), .Y(_27178_) );
  \$mux  #( .WIDTH(1) ) _51315_ ( .A(_27178_), .B(1'h0), .S(RST), .Y(_02963_) );
  \$mux  #( .WIDTH(1) ) _51316_ ( .A(_tmp_1353), .B(1'h0), .S(_06549_), .Y(_27179_) );
  \$mux  #( .WIDTH(1) ) _51317_ ( .A(_27179_), .B(1'h1), .S(_06550_), .Y(_27180_) );
  \$mux  #( .WIDTH(1) ) _51318_ ( .A(_27180_), .B(1'h0), .S(RST), .Y(_02962_) );
  \$mux  #( .WIDTH(1) ) _51319_ ( .A(_tmp_1352), .B(1'h0), .S(_06550_), .Y(_27181_) );
  \$mux  #( .WIDTH(1) ) _51320_ ( .A(_27181_), .B(1'h1), .S(_06551_), .Y(_27182_) );
  \$mux  #( .WIDTH(1) ) _51321_ ( .A(_27182_), .B(1'h1), .S(_06552_), .Y(_27183_) );
  \$mux  #( .WIDTH(1) ) _51322_ ( .A(_27183_), .B(1'h0), .S(RST), .Y(_02961_) );
  \$mux  #( .WIDTH(8) ) _51323_ ( .A(_tmp_1351), .B(8'h00), .S(RST), .Y(_01228_) );
  \$mux  #( .WIDTH(1) ) _51324_ ( .A(_tmp_1350), .B(1'h0), .S(RST), .Y(_01227_) );
  \$mux  #( .WIDTH(1) ) _51325_ ( .A(_tmp_1345), .B(1'h0), .S(_06549_), .Y(_27184_) );
  \$mux  #( .WIDTH(1) ) _51326_ ( .A(_27184_), .B(1'h1), .S(_06550_), .Y(_27185_) );
  \$mux  #( .WIDTH(1) ) _51327_ ( .A(_27185_), .B(1'h0), .S(RST), .Y(_02959_) );
  \$mux  #( .WIDTH(1) ) _51328_ ( .A(_06548_), .B(1'h0), .S(RST), .Y(_01836_) );
  \$mux  #( .WIDTH(1) ) _51329_ ( .A(_tmp_19), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27186_) );
  \$mux  #( .WIDTH(1) ) _51330_ ( .A(_27186_), .B(1'h1), .S(_06547_), .Y(_27187_) );
  \$mux  #( .WIDTH(1) ) _51331_ ( .A(_27187_), .B(1'h0), .S(RST), .Y(_03002_) );
  \$mux  #( .WIDTH(34) ) _51332_ ( .A(_tmp_18), .B({ 1'h0, _maxi_read_size }), .S(_06546_), .Y(_27188_) );
  \$mux  #( .WIDTH(34) ) _51333_ ( .A(_27188_), .B(_28577_), .S(_06205_), .Y(_27189_) );
  \$mux  #( .WIDTH(34) ) _51334_ ( .A(_27189_), .B(34'h000000000), .S(RST), .Y(_02993_) );
  \$mux  #( .WIDTH(1) ) _51335_ ( .A(ram_w8_l2048_id1_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27190_) );
  \$mux  #( .WIDTH(1) ) _51336_ ( .A(_27190_), .B(1'h1), .S(_06205_), .Y(_27191_) );
  \$mux  #( .WIDTH(1) ) _51337_ ( .A(_27191_), .B(1'h0), .S(RST), .Y(_03740_) );
  \$mux  #( .WIDTH(8) ) _51338_ ( .A(ram_w8_l2048_id1_3_1_wdata), .B(_dataflow_slice_data_12), .S(_06205_), .Y(_27192_) );
  \$mux  #( .WIDTH(8) ) _51339_ ( .A(_27192_), .B(8'h00), .S(RST), .Y(_03739_) );
  \$mux  #( .WIDTH(9) ) _51340_ ( .A(ram_w8_l2048_id1_3_1_addr), .B(_28537_[8:0]), .S(_06546_), .Y(_27193_) );
  \$mux  #( .WIDTH(9) ) _51341_ ( .A(_27193_), .B(_24264_[8:0]), .S(_06205_), .Y(_27194_) );
  \$mux  #( .WIDTH(9) ) _51342_ ( .A(_27194_), .B(_maxi_write_local_addr[8:0]), .S(_06551_), .Y(_27195_) );
  \$mux  #( .WIDTH(9) ) _51343_ ( .A(_27195_), .B(_24265_[8:0]), .S(_06552_), .Y(_27196_) );
  \$mux  #( .WIDTH(9) ) _51344_ ( .A(_27196_), .B(9'h000), .S(RST), .Y(_03738_) );
  \$mux  #( .WIDTH(1) ) _51345_ ( .A(ram_w8_l2048_id1_3_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id1_3_cond_5_1), .Y(_27197_) );
  \$mux  #( .WIDTH(1) ) _51346_ ( .A(_27197_), .B(1'h1), .S(_06548_), .Y(_27198_) );
  \$mux  #( .WIDTH(1) ) _51347_ ( .A(_27198_), .B(1'h0), .S(RST), .Y(_03737_) );
  \$mux  #( .WIDTH(8) ) _51348_ ( .A(ram_w8_l2048_id1_3_0_wdata), .B(_stream_matmul_29_sink_21_sink_wdata), .S(_06548_), .Y(_27199_) );
  \$mux  #( .WIDTH(8) ) _51349_ ( .A(_27199_), .B(8'h00), .S(RST), .Y(_03736_) );
  \$mux  #( .WIDTH(9) ) _51350_ ( .A(ram_w8_l2048_id1_3_0_addr), .B(_stream_conv2d_16_source_6_source_ram_raddr[10:2]), .S(_tmp_472), .Y(_27200_) );
  \$mux  #( .WIDTH(9) ) _51351_ ( .A(_27200_), .B(_stream_max_pool_serial_18_source_1_source_ram_raddr[10:2]), .S(_tmp_1035), .Y(_27201_) );
  \$mux  #( .WIDTH(9) ) _51352_ ( .A(_27201_), .B(_stream_matmul_29_sink_21_sink_waddr[10:2]), .S(_06548_), .Y(_27202_) );
  \$mux  #( .WIDTH(9) ) _51353_ ( .A(_27202_), .B(9'h000), .S(RST), .Y(_03735_) );
  \$mux  #( .WIDTH(34) ) _51354_ ( .A(_tmp_1344), .B(_28563_), .S(_06543_), .Y(_27203_) );
  \$mux  #( .WIDTH(34) ) _51355_ ( .A(_27203_), .B(_28576_), .S(_06544_), .Y(_27204_) );
  \$mux  #( .WIDTH(34) ) _51356_ ( .A(_27204_), .B(34'h000000000), .S(RST), .Y(_02958_) );
  \$mux  #( .WIDTH(1) ) _51357_ ( .A(_tmp_1343), .B(1'h0), .S(_06541_), .Y(_27205_) );
  \$mux  #( .WIDTH(1) ) _51358_ ( .A(_27205_), .B(_tmp_1342), .S(_06542_), .Y(_27206_) );
  \$mux  #( .WIDTH(1) ) _51359_ ( .A(_27206_), .B(1'h0), .S(RST), .Y(_02957_) );
  \$mux  #( .WIDTH(1) ) _51360_ ( .A(_tmp_1342), .B(1'h0), .S(_06542_), .Y(_27207_) );
  \$mux  #( .WIDTH(1) ) _51361_ ( .A(_27207_), .B(_06099_), .S(_06543_), .Y(_27208_) );
  \$mux  #( .WIDTH(1) ) _51362_ ( .A(_27208_), .B(1'h0), .S(_06544_), .Y(_27209_) );
  \$mux  #( .WIDTH(1) ) _51363_ ( .A(_27209_), .B(1'h1), .S(_06545_), .Y(_27210_) );
  \$mux  #( .WIDTH(1) ) _51364_ ( .A(_27210_), .B(1'h0), .S(RST), .Y(_02956_) );
  \$mux  #( .WIDTH(1) ) _51365_ ( .A(_tmp_1341), .B(1'h0), .S(_06541_), .Y(_27211_) );
  \$mux  #( .WIDTH(1) ) _51366_ ( .A(_27211_), .B(1'h1), .S(_06542_), .Y(_27212_) );
  \$mux  #( .WIDTH(1) ) _51367_ ( .A(_27212_), .B(1'h0), .S(RST), .Y(_02955_) );
  \$mux  #( .WIDTH(1) ) _51368_ ( .A(_tmp_1340), .B(1'h0), .S(_06542_), .Y(_27213_) );
  \$mux  #( .WIDTH(1) ) _51369_ ( .A(_27213_), .B(1'h1), .S(_06543_), .Y(_27214_) );
  \$mux  #( .WIDTH(1) ) _51370_ ( .A(_27214_), .B(1'h1), .S(_06544_), .Y(_27215_) );
  \$mux  #( .WIDTH(1) ) _51371_ ( .A(_27215_), .B(1'h0), .S(RST), .Y(_02954_) );
  \$mux  #( .WIDTH(8) ) _51372_ ( .A(_tmp_1339), .B(8'h00), .S(RST), .Y(_01226_) );
  \$mux  #( .WIDTH(1) ) _51373_ ( .A(_tmp_1338), .B(1'h0), .S(RST), .Y(_01225_) );
  \$mux  #( .WIDTH(1) ) _51374_ ( .A(_tmp_1333), .B(1'h0), .S(_06541_), .Y(_27216_) );
  \$mux  #( .WIDTH(1) ) _51375_ ( .A(_27216_), .B(1'h1), .S(_06542_), .Y(_27217_) );
  \$mux  #( .WIDTH(1) ) _51376_ ( .A(_27217_), .B(1'h0), .S(RST), .Y(_02952_) );
  \$mux  #( .WIDTH(1) ) _51377_ ( .A(_06540_), .B(1'h0), .S(RST), .Y(_01835_) );
  \$mux  #( .WIDTH(1) ) _51378_ ( .A(_tmp_17), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27218_) );
  \$mux  #( .WIDTH(1) ) _51379_ ( .A(_27218_), .B(1'h1), .S(_06539_), .Y(_27219_) );
  \$mux  #( .WIDTH(1) ) _51380_ ( .A(_27219_), .B(1'h0), .S(RST), .Y(_02992_) );
  \$mux  #( .WIDTH(34) ) _51381_ ( .A(_tmp_16), .B({ 1'h0, _maxi_read_size }), .S(_06538_), .Y(_27220_) );
  \$mux  #( .WIDTH(34) ) _51382_ ( .A(_27220_), .B(_28575_), .S(_06202_), .Y(_27221_) );
  \$mux  #( .WIDTH(34) ) _51383_ ( .A(_27221_), .B(34'h000000000), .S(RST), .Y(_02987_) );
  \$mux  #( .WIDTH(1) ) _51384_ ( .A(ram_w8_l2048_id1_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27222_) );
  \$mux  #( .WIDTH(1) ) _51385_ ( .A(_27222_), .B(1'h1), .S(_06202_), .Y(_27223_) );
  \$mux  #( .WIDTH(1) ) _51386_ ( .A(_27223_), .B(1'h0), .S(RST), .Y(_03734_) );
  \$mux  #( .WIDTH(8) ) _51387_ ( .A(ram_w8_l2048_id1_2_1_wdata), .B(_dataflow_slice_data_9), .S(_06202_), .Y(_27224_) );
  \$mux  #( .WIDTH(8) ) _51388_ ( .A(_27224_), .B(8'h00), .S(RST), .Y(_03733_) );
  \$mux  #( .WIDTH(9) ) _51389_ ( .A(ram_w8_l2048_id1_2_1_addr), .B(_28537_[8:0]), .S(_06538_), .Y(_27225_) );
  \$mux  #( .WIDTH(9) ) _51390_ ( .A(_27225_), .B(_24262_[8:0]), .S(_06202_), .Y(_27226_) );
  \$mux  #( .WIDTH(9) ) _51391_ ( .A(_27226_), .B(_maxi_write_local_addr[8:0]), .S(_06543_), .Y(_27227_) );
  \$mux  #( .WIDTH(9) ) _51392_ ( .A(_27227_), .B(_24263_[8:0]), .S(_06544_), .Y(_27228_) );
  \$mux  #( .WIDTH(9) ) _51393_ ( .A(_27228_), .B(9'h000), .S(RST), .Y(_03732_) );
  \$mux  #( .WIDTH(1) ) _51394_ ( .A(ram_w8_l2048_id1_2_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id1_2_cond_5_1), .Y(_27229_) );
  \$mux  #( .WIDTH(1) ) _51395_ ( .A(_27229_), .B(1'h1), .S(_06540_), .Y(_27230_) );
  \$mux  #( .WIDTH(1) ) _51396_ ( .A(_27230_), .B(1'h0), .S(RST), .Y(_03731_) );
  \$mux  #( .WIDTH(8) ) _51397_ ( .A(ram_w8_l2048_id1_2_0_wdata), .B(_stream_matmul_29_sink_21_sink_wdata), .S(_06540_), .Y(_27231_) );
  \$mux  #( .WIDTH(8) ) _51398_ ( .A(_27231_), .B(8'h00), .S(RST), .Y(_03730_) );
  \$mux  #( .WIDTH(9) ) _51399_ ( .A(ram_w8_l2048_id1_2_0_addr), .B(_stream_conv2d_16_source_6_source_ram_raddr[10:2]), .S(_tmp_472), .Y(_27232_) );
  \$mux  #( .WIDTH(9) ) _51400_ ( .A(_27232_), .B(_stream_max_pool_serial_18_source_1_source_ram_raddr[10:2]), .S(_tmp_1035), .Y(_27233_) );
  \$mux  #( .WIDTH(9) ) _51401_ ( .A(_27233_), .B(_stream_matmul_29_sink_21_sink_waddr[10:2]), .S(_06540_), .Y(_27234_) );
  \$mux  #( .WIDTH(9) ) _51402_ ( .A(_27234_), .B(9'h000), .S(RST), .Y(_03729_) );
  \$mux  #( .WIDTH(34) ) _51403_ ( .A(_tmp_1332), .B(_28563_), .S(_06535_), .Y(_27235_) );
  \$mux  #( .WIDTH(34) ) _51404_ ( .A(_27235_), .B(_28574_), .S(_06536_), .Y(_27236_) );
  \$mux  #( .WIDTH(34) ) _51405_ ( .A(_27236_), .B(34'h000000000), .S(RST), .Y(_02951_) );
  \$mux  #( .WIDTH(1) ) _51406_ ( .A(_tmp_1331), .B(1'h0), .S(_06533_), .Y(_27237_) );
  \$mux  #( .WIDTH(1) ) _51407_ ( .A(_27237_), .B(_tmp_1330), .S(_06534_), .Y(_27238_) );
  \$mux  #( .WIDTH(1) ) _51408_ ( .A(_27238_), .B(1'h0), .S(RST), .Y(_02950_) );
  \$mux  #( .WIDTH(1) ) _51409_ ( .A(_tmp_1330), .B(1'h0), .S(_06534_), .Y(_27239_) );
  \$mux  #( .WIDTH(1) ) _51410_ ( .A(_27239_), .B(_06099_), .S(_06535_), .Y(_27240_) );
  \$mux  #( .WIDTH(1) ) _51411_ ( .A(_27240_), .B(1'h0), .S(_06536_), .Y(_27241_) );
  \$mux  #( .WIDTH(1) ) _51412_ ( .A(_27241_), .B(1'h1), .S(_06537_), .Y(_27242_) );
  \$mux  #( .WIDTH(1) ) _51413_ ( .A(_27242_), .B(1'h0), .S(RST), .Y(_02949_) );
  \$mux  #( .WIDTH(1) ) _51414_ ( .A(_tmp_1329), .B(1'h0), .S(_06533_), .Y(_27243_) );
  \$mux  #( .WIDTH(1) ) _51415_ ( .A(_27243_), .B(1'h1), .S(_06534_), .Y(_27244_) );
  \$mux  #( .WIDTH(1) ) _51416_ ( .A(_27244_), .B(1'h0), .S(RST), .Y(_02947_) );
  \$mux  #( .WIDTH(1) ) _51417_ ( .A(_tmp_1328), .B(1'h0), .S(_06534_), .Y(_27245_) );
  \$mux  #( .WIDTH(1) ) _51418_ ( .A(_27245_), .B(1'h1), .S(_06535_), .Y(_27246_) );
  \$mux  #( .WIDTH(1) ) _51419_ ( .A(_27246_), .B(1'h1), .S(_06536_), .Y(_27247_) );
  \$mux  #( .WIDTH(1) ) _51420_ ( .A(_27247_), .B(1'h0), .S(RST), .Y(_02946_) );
  \$mux  #( .WIDTH(8) ) _51421_ ( .A(_tmp_1327), .B(8'h00), .S(RST), .Y(_01224_) );
  \$mux  #( .WIDTH(1) ) _51422_ ( .A(_tmp_1326), .B(1'h0), .S(RST), .Y(_01223_) );
  \$mux  #( .WIDTH(1) ) _51423_ ( .A(_tmp_1321), .B(1'h0), .S(_06533_), .Y(_27248_) );
  \$mux  #( .WIDTH(1) ) _51424_ ( .A(_27248_), .B(1'h1), .S(_06534_), .Y(_27249_) );
  \$mux  #( .WIDTH(1) ) _51425_ ( .A(_27249_), .B(1'h0), .S(RST), .Y(_02945_) );
  \$mux  #( .WIDTH(1) ) _51426_ ( .A(_06532_), .B(1'h0), .S(RST), .Y(_01834_) );
  \$mux  #( .WIDTH(1) ) _51427_ ( .A(_tmp_15), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27250_) );
  \$mux  #( .WIDTH(1) ) _51428_ ( .A(_27250_), .B(1'h1), .S(_06531_), .Y(_27251_) );
  \$mux  #( .WIDTH(1) ) _51429_ ( .A(_27251_), .B(1'h0), .S(RST), .Y(_02977_) );
  \$mux  #( .WIDTH(34) ) _51430_ ( .A(_tmp_14), .B({ 1'h0, _maxi_read_size }), .S(_06530_), .Y(_27252_) );
  \$mux  #( .WIDTH(34) ) _51431_ ( .A(_27252_), .B(_28573_), .S(_06199_), .Y(_27253_) );
  \$mux  #( .WIDTH(34) ) _51432_ ( .A(_27253_), .B(34'h000000000), .S(RST), .Y(_02976_) );
  \$mux  #( .WIDTH(1) ) _51433_ ( .A(ram_w8_l2048_id1_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27254_) );
  \$mux  #( .WIDTH(1) ) _51434_ ( .A(_27254_), .B(1'h1), .S(_06199_), .Y(_27255_) );
  \$mux  #( .WIDTH(1) ) _51435_ ( .A(_27255_), .B(1'h0), .S(RST), .Y(_03728_) );
  \$mux  #( .WIDTH(8) ) _51436_ ( .A(ram_w8_l2048_id1_1_1_wdata), .B(_dataflow_slice_data_6), .S(_06199_), .Y(_27256_) );
  \$mux  #( .WIDTH(8) ) _51437_ ( .A(_27256_), .B(8'h00), .S(RST), .Y(_03727_) );
  \$mux  #( .WIDTH(9) ) _51438_ ( .A(ram_w8_l2048_id1_1_1_addr), .B(_28537_[8:0]), .S(_06530_), .Y(_27257_) );
  \$mux  #( .WIDTH(9) ) _51439_ ( .A(_27257_), .B(_24260_[8:0]), .S(_06199_), .Y(_27258_) );
  \$mux  #( .WIDTH(9) ) _51440_ ( .A(_27258_), .B(_maxi_write_local_addr[8:0]), .S(_06535_), .Y(_27259_) );
  \$mux  #( .WIDTH(9) ) _51441_ ( .A(_27259_), .B(_24261_[8:0]), .S(_06536_), .Y(_27260_) );
  \$mux  #( .WIDTH(9) ) _51442_ ( .A(_27260_), .B(9'h000), .S(RST), .Y(_03726_) );
  \$mux  #( .WIDTH(1) ) _51443_ ( .A(ram_w8_l2048_id1_1_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id1_1_cond_5_1), .Y(_27261_) );
  \$mux  #( .WIDTH(1) ) _51444_ ( .A(_27261_), .B(1'h1), .S(_06532_), .Y(_27262_) );
  \$mux  #( .WIDTH(1) ) _51445_ ( .A(_27262_), .B(1'h0), .S(RST), .Y(_03725_) );
  \$mux  #( .WIDTH(8) ) _51446_ ( .A(ram_w8_l2048_id1_1_0_wdata), .B(_stream_matmul_29_sink_21_sink_wdata), .S(_06532_), .Y(_27263_) );
  \$mux  #( .WIDTH(8) ) _51447_ ( .A(_27263_), .B(8'h00), .S(RST), .Y(_03724_) );
  \$mux  #( .WIDTH(9) ) _51448_ ( .A(ram_w8_l2048_id1_1_0_addr), .B(_stream_conv2d_16_source_6_source_ram_raddr[10:2]), .S(_tmp_472), .Y(_27264_) );
  \$mux  #( .WIDTH(9) ) _51449_ ( .A(_27264_), .B(_stream_max_pool_serial_18_source_1_source_ram_raddr[10:2]), .S(_tmp_1035), .Y(_27265_) );
  \$mux  #( .WIDTH(9) ) _51450_ ( .A(_27265_), .B(_stream_matmul_29_sink_21_sink_waddr[10:2]), .S(_06532_), .Y(_27266_) );
  \$mux  #( .WIDTH(9) ) _51451_ ( .A(_27266_), .B(9'h000), .S(RST), .Y(_03723_) );
  \$mux  #( .WIDTH(1) ) _51452_ ( .A(_dataflow_cat_valid_167), .B(1'h0), .S(_06192_), .Y(_27267_) );
  \$mux  #( .WIDTH(1) ) _51453_ ( .A(_27267_), .B(_06528_), .S(_06529_), .Y(_27268_) );
  \$mux  #( .WIDTH(1) ) _51454_ ( .A(_27268_), .B(1'h0), .S(RST), .Y(_01590_) );
  \$mux  #( .WIDTH(32) ) _51455_ ( .A(_dataflow_cat_data_167), .B({ _tmp_1351, _tmp_1339, _tmp_1327, _tmp_1315 }), .S(_06529_), .Y(_27269_) );
  \$mux  #( .WIDTH(32) ) _51456_ ( .A(_27269_), .B(0), .S(RST), .Y(_01587_) );
  \$mux  #( .WIDTH(34) ) _51457_ ( .A(_tmp_1320), .B(_28563_), .S(_06525_), .Y(_27270_) );
  \$mux  #( .WIDTH(34) ) _51458_ ( .A(_27270_), .B(_28572_), .S(_06526_), .Y(_27271_) );
  \$mux  #( .WIDTH(34) ) _51459_ ( .A(_27271_), .B(34'h000000000), .S(RST), .Y(_02944_) );
  \$mux  #( .WIDTH(1) ) _51460_ ( .A(_tmp_1319), .B(1'h0), .S(_06522_), .Y(_27272_) );
  \$mux  #( .WIDTH(1) ) _51461_ ( .A(_27272_), .B(_tmp_1318), .S(_06523_), .Y(_27273_) );
  \$mux  #( .WIDTH(1) ) _51462_ ( .A(_27273_), .B(1'h0), .S(RST), .Y(_02942_) );
  \$mux  #( .WIDTH(1) ) _51463_ ( .A(_tmp_1318), .B(1'h0), .S(_06523_), .Y(_27274_) );
  \$mux  #( .WIDTH(1) ) _51464_ ( .A(_27274_), .B(_06099_), .S(_06525_), .Y(_27275_) );
  \$mux  #( .WIDTH(1) ) _51465_ ( .A(_27275_), .B(1'h0), .S(_06526_), .Y(_27276_) );
  \$mux  #( .WIDTH(1) ) _51466_ ( .A(_27276_), .B(1'h1), .S(_06527_), .Y(_27277_) );
  \$mux  #( .WIDTH(1) ) _51467_ ( .A(_27277_), .B(1'h0), .S(RST), .Y(_02941_) );
  \$mux  #( .WIDTH(1) ) _51468_ ( .A(_tmp_1317), .B(1'h0), .S(_06522_), .Y(_27278_) );
  \$mux  #( .WIDTH(1) ) _51469_ ( .A(_27278_), .B(1'h1), .S(_06523_), .Y(_27279_) );
  \$mux  #( .WIDTH(1) ) _51470_ ( .A(_27279_), .B(1'h0), .S(RST), .Y(_02940_) );
  \$mux  #( .WIDTH(1) ) _51471_ ( .A(_tmp_1316), .B(1'h0), .S(_06523_), .Y(_27280_) );
  \$mux  #( .WIDTH(1) ) _51472_ ( .A(_27280_), .B(1'h1), .S(_06525_), .Y(_27281_) );
  \$mux  #( .WIDTH(1) ) _51473_ ( .A(_27281_), .B(1'h1), .S(_06526_), .Y(_27282_) );
  \$mux  #( .WIDTH(1) ) _51474_ ( .A(_27282_), .B(1'h0), .S(RST), .Y(_02939_) );
  \$mux  #( .WIDTH(8) ) _51475_ ( .A(_tmp_1315), .B(8'h00), .S(RST), .Y(_01222_) );
  \$mux  #( .WIDTH(1) ) _51476_ ( .A(_tmp_1314), .B(1'h0), .S(RST), .Y(_01221_) );
  \$mux  #( .WIDTH(1) ) _51477_ ( .A(_tmp_1309), .B(1'h0), .S(_06522_), .Y(_27283_) );
  \$mux  #( .WIDTH(1) ) _51478_ ( .A(_27283_), .B(1'h1), .S(_06523_), .Y(_27284_) );
  \$mux  #( .WIDTH(1) ) _51479_ ( .A(_27284_), .B(1'h0), .S(RST), .Y(_02937_) );
  \$mux  #( .WIDTH(1) ) _51480_ ( .A(_06521_), .B(1'h0), .S(RST), .Y(_01833_) );
  \$mux  #( .WIDTH(1) ) _51481_ ( .A(_tmp_1035), .B(1'h0), .S(RST), .Y(_01111_) );
  \$mux  #( .WIDTH(1) ) _51482_ ( .A(_tmp_472), .B(1'h0), .S(RST), .Y(_01231_) );
  \$mux  #( .WIDTH(1) ) _51483_ ( .A(_tmp_13), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27285_) );
  \$mux  #( .WIDTH(1) ) _51484_ ( .A(_27285_), .B(1'h1), .S(_06520_), .Y(_27286_) );
  \$mux  #( .WIDTH(1) ) _51485_ ( .A(_27286_), .B(1'h0), .S(RST), .Y(_02972_) );
  \$mux  #( .WIDTH(34) ) _51486_ ( .A(_tmp_12), .B({ 1'h0, _maxi_read_size }), .S(_06519_), .Y(_27287_) );
  \$mux  #( .WIDTH(34) ) _51487_ ( .A(_27287_), .B(_28571_), .S(_06196_), .Y(_27288_) );
  \$mux  #( .WIDTH(34) ) _51488_ ( .A(_27288_), .B(34'h000000000), .S(RST), .Y(_02936_) );
  \$mux  #( .WIDTH(1) ) _51489_ ( .A(ram_w8_l2048_id1_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27289_) );
  \$mux  #( .WIDTH(1) ) _51490_ ( .A(_27289_), .B(1'h1), .S(_06196_), .Y(_27290_) );
  \$mux  #( .WIDTH(1) ) _51491_ ( .A(_27290_), .B(1'h0), .S(RST), .Y(_03722_) );
  \$mux  #( .WIDTH(8) ) _51492_ ( .A(ram_w8_l2048_id1_0_1_wdata), .B(_dataflow_slice_data_3), .S(_06196_), .Y(_27291_) );
  \$mux  #( .WIDTH(8) ) _51493_ ( .A(_27291_), .B(8'h00), .S(RST), .Y(_03721_) );
  \$mux  #( .WIDTH(9) ) _51494_ ( .A(ram_w8_l2048_id1_0_1_addr), .B(_28537_[8:0]), .S(_06519_), .Y(_27292_) );
  \$mux  #( .WIDTH(9) ) _51495_ ( .A(_27292_), .B(_24258_[8:0]), .S(_06196_), .Y(_27293_) );
  \$mux  #( .WIDTH(9) ) _51496_ ( .A(_27293_), .B(_maxi_write_local_addr[8:0]), .S(_06525_), .Y(_27294_) );
  \$mux  #( .WIDTH(9) ) _51497_ ( .A(_27294_), .B(_24259_[8:0]), .S(_06526_), .Y(_27295_) );
  \$mux  #( .WIDTH(9) ) _51498_ ( .A(_27295_), .B(9'h000), .S(RST), .Y(_03720_) );
  \$mux  #( .WIDTH(1) ) _51499_ ( .A(ram_w8_l2048_id1_0_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id1_0_cond_5_1), .Y(_27296_) );
  \$mux  #( .WIDTH(1) ) _51500_ ( .A(_27296_), .B(1'h1), .S(_06521_), .Y(_27297_) );
  \$mux  #( .WIDTH(1) ) _51501_ ( .A(_27297_), .B(1'h0), .S(RST), .Y(_03719_) );
  \$mux  #( .WIDTH(8) ) _51502_ ( .A(ram_w8_l2048_id1_0_0_wdata), .B(_stream_matmul_29_sink_21_sink_wdata), .S(_06521_), .Y(_27298_) );
  \$mux  #( .WIDTH(8) ) _51503_ ( .A(_27298_), .B(8'h00), .S(RST), .Y(_03718_) );
  \$mux  #( .WIDTH(9) ) _51504_ ( .A(ram_w8_l2048_id1_0_0_addr), .B(_stream_conv2d_16_source_6_source_ram_raddr[10:2]), .S(_tmp_472), .Y(_27299_) );
  \$mux  #( .WIDTH(9) ) _51505_ ( .A(_27299_), .B(_stream_max_pool_serial_18_source_1_source_ram_raddr[10:2]), .S(_tmp_1035), .Y(_27300_) );
  \$mux  #( .WIDTH(9) ) _51506_ ( .A(_27300_), .B(_stream_matmul_29_sink_21_sink_waddr[10:2]), .S(_06521_), .Y(_27301_) );
  \$mux  #( .WIDTH(9) ) _51507_ ( .A(_27301_), .B(9'h000), .S(RST), .Y(_03717_) );
  \$mux  #( .WIDTH(34) ) _51508_ ( .A(_tmp_1119), .B(_28563_), .S(_06515_), .Y(_27302_) );
  \$mux  #( .WIDTH(34) ) _51509_ ( .A(_27302_), .B(_28570_), .S(_06516_), .Y(_27303_) );
  \$mux  #( .WIDTH(34) ) _51510_ ( .A(_27303_), .B(34'h000000000), .S(RST), .Y(_02901_) );
  \$mux  #( .WIDTH(1) ) _51511_ ( .A(_tmp_1118), .B(1'h0), .S(_06513_), .Y(_27304_) );
  \$mux  #( .WIDTH(1) ) _51512_ ( .A(_27304_), .B(_tmp_1117), .S(_06514_), .Y(_27305_) );
  \$mux  #( .WIDTH(1) ) _51513_ ( .A(_27305_), .B(1'h0), .S(RST), .Y(_02900_) );
  \$mux  #( .WIDTH(1) ) _51514_ ( .A(_tmp_1117), .B(1'h0), .S(_06514_), .Y(_27306_) );
  \$mux  #( .WIDTH(1) ) _51515_ ( .A(_27306_), .B(_06099_), .S(_06515_), .Y(_27307_) );
  \$mux  #( .WIDTH(1) ) _51516_ ( .A(_27307_), .B(1'h0), .S(_06516_), .Y(_27308_) );
  \$mux  #( .WIDTH(1) ) _51517_ ( .A(_27308_), .B(1'h1), .S(_06517_), .Y(_27309_) );
  \$mux  #( .WIDTH(1) ) _51518_ ( .A(_27309_), .B(1'h0), .S(RST), .Y(_02899_) );
  \$mux  #( .WIDTH(1) ) _51519_ ( .A(_tmp_1116), .B(1'h0), .S(_06513_), .Y(_27310_) );
  \$mux  #( .WIDTH(1) ) _51520_ ( .A(_27310_), .B(1'h1), .S(_06514_), .Y(_27311_) );
  \$mux  #( .WIDTH(1) ) _51521_ ( .A(_27311_), .B(1'h0), .S(RST), .Y(_02898_) );
  \$mux  #( .WIDTH(1) ) _51522_ ( .A(_tmp_1115), .B(1'h0), .S(_06514_), .Y(_27312_) );
  \$mux  #( .WIDTH(1) ) _51523_ ( .A(_27312_), .B(1'h1), .S(_06515_), .Y(_27313_) );
  \$mux  #( .WIDTH(1) ) _51524_ ( .A(_27313_), .B(1'h1), .S(_06516_), .Y(_27314_) );
  \$mux  #( .WIDTH(1) ) _51525_ ( .A(_27314_), .B(1'h0), .S(RST), .Y(_02897_) );
  \$mux  #( .WIDTH(8) ) _51526_ ( .A(_tmp_1114), .B(8'h00), .S(RST), .Y(_01138_) );
  \$mux  #( .WIDTH(1) ) _51527_ ( .A(_tmp_1113), .B(1'h0), .S(RST), .Y(_01137_) );
  \$mux  #( .WIDTH(1) ) _51528_ ( .A(_tmp_1108), .B(1'h0), .S(_06513_), .Y(_27315_) );
  \$mux  #( .WIDTH(1) ) _51529_ ( .A(_27315_), .B(1'h1), .S(_06514_), .Y(_27316_) );
  \$mux  #( .WIDTH(1) ) _51530_ ( .A(_27316_), .B(1'h0), .S(RST), .Y(_02895_) );
  \$mux  #( .WIDTH(1) ) _51531_ ( .A(_06512_), .B(1'h0), .S(RST), .Y(_01828_) );
  \$mux  #( .WIDTH(1) ) _51532_ ( .A(_tmp_32), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27317_) );
  \$mux  #( .WIDTH(1) ) _51533_ ( .A(_27317_), .B(1'h1), .S(_06511_), .Y(_27318_) );
  \$mux  #( .WIDTH(1) ) _51534_ ( .A(_27318_), .B(1'h0), .S(RST), .Y(_03066_) );
  \$mux  #( .WIDTH(34) ) _51535_ ( .A(_tmp_31), .B({ 1'h0, _maxi_read_size }), .S(_06510_), .Y(_27319_) );
  \$mux  #( .WIDTH(34) ) _51536_ ( .A(_27319_), .B(_28569_), .S(_06217_), .Y(_27320_) );
  \$mux  #( .WIDTH(34) ) _51537_ ( .A(_27320_), .B(34'h000000000), .S(RST), .Y(_03061_) );
  \$mux  #( .WIDTH(1) ) _51538_ ( .A(ram_w8_l2048_id0_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27321_) );
  \$mux  #( .WIDTH(1) ) _51539_ ( .A(_27321_), .B(1'h1), .S(_06217_), .Y(_27322_) );
  \$mux  #( .WIDTH(1) ) _51540_ ( .A(_27322_), .B(1'h0), .S(RST), .Y(_03684_) );
  \$mux  #( .WIDTH(8) ) _51541_ ( .A(ram_w8_l2048_id0_3_1_wdata), .B(_dataflow_slice_data_25), .S(_06217_), .Y(_27323_) );
  \$mux  #( .WIDTH(8) ) _51542_ ( .A(_27323_), .B(8'h00), .S(RST), .Y(_03683_) );
  \$mux  #( .WIDTH(9) ) _51543_ ( .A(ram_w8_l2048_id0_3_1_addr), .B(_28537_[8:0]), .S(_06510_), .Y(_27324_) );
  \$mux  #( .WIDTH(9) ) _51544_ ( .A(_27324_), .B(_24256_[8:0]), .S(_06217_), .Y(_27325_) );
  \$mux  #( .WIDTH(9) ) _51545_ ( .A(_27325_), .B(_maxi_write_local_addr[8:0]), .S(_06515_), .Y(_27326_) );
  \$mux  #( .WIDTH(9) ) _51546_ ( .A(_27326_), .B(_24257_[8:0]), .S(_06516_), .Y(_27327_) );
  \$mux  #( .WIDTH(9) ) _51547_ ( .A(_27327_), .B(9'h000), .S(RST), .Y(_03682_) );
  \$mux  #( .WIDTH(1) ) _51548_ ( .A(ram_w8_l2048_id0_3_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_3_1), .Y(_27328_) );
  \$mux  #( .WIDTH(1) ) _51549_ ( .A(_27328_), .B(1'h1), .S(_06512_), .Y(_27329_) );
  \$mux  #( .WIDTH(1) ) _51550_ ( .A(_27329_), .B(1'h0), .S(RST), .Y(_03681_) );
  \$mux  #( .WIDTH(8) ) _51551_ ( .A(ram_w8_l2048_id0_3_0_wdata), .B(_stream_max_pool_serial_18_sink_3_sink_wdata), .S(_06512_), .Y(_27330_) );
  \$mux  #( .WIDTH(8) ) _51552_ ( .A(_27330_), .B(8'h00), .S(RST), .Y(_03680_) );
  \$mux  #( .WIDTH(9) ) _51553_ ( .A(ram_w8_l2048_id0_3_0_addr), .B(_stream_conv2d_16_source_8_source_ram_raddr[10:2]), .S(_tmp_483), .Y(_27331_) );
  \$mux  #( .WIDTH(9) ) _51554_ ( .A(_27331_), .B(_stream_max_pool_serial_18_sink_3_sink_waddr[10:2]), .S(_06512_), .Y(_27332_) );
  \$mux  #( .WIDTH(9) ) _51555_ ( .A(_27332_), .B(_stream_matmul_29_source_8_source_ram_raddr[10:2]), .S(_tmp_1189), .Y(_27333_) );
  \$mux  #( .WIDTH(9) ) _51556_ ( .A(_27333_), .B(9'h000), .S(RST), .Y(_03679_) );
  \$mux  #( .WIDTH(34) ) _51557_ ( .A(_tmp_1107), .B(_28563_), .S(_06507_), .Y(_27334_) );
  \$mux  #( .WIDTH(34) ) _51558_ ( .A(_27334_), .B(_28568_), .S(_06508_), .Y(_27335_) );
  \$mux  #( .WIDTH(34) ) _51559_ ( .A(_27335_), .B(34'h000000000), .S(RST), .Y(_02894_) );
  \$mux  #( .WIDTH(1) ) _51560_ ( .A(_tmp_1106), .B(1'h0), .S(_06505_), .Y(_27336_) );
  \$mux  #( .WIDTH(1) ) _51561_ ( .A(_27336_), .B(_tmp_1105), .S(_06506_), .Y(_27337_) );
  \$mux  #( .WIDTH(1) ) _51562_ ( .A(_27337_), .B(1'h0), .S(RST), .Y(_02893_) );
  \$mux  #( .WIDTH(1) ) _51563_ ( .A(_tmp_1105), .B(1'h0), .S(_06506_), .Y(_27338_) );
  \$mux  #( .WIDTH(1) ) _51564_ ( .A(_27338_), .B(_06099_), .S(_06507_), .Y(_27339_) );
  \$mux  #( .WIDTH(1) ) _51565_ ( .A(_27339_), .B(1'h0), .S(_06508_), .Y(_27340_) );
  \$mux  #( .WIDTH(1) ) _51566_ ( .A(_27340_), .B(1'h1), .S(_06509_), .Y(_27341_) );
  \$mux  #( .WIDTH(1) ) _51567_ ( .A(_27341_), .B(1'h0), .S(RST), .Y(_02892_) );
  \$mux  #( .WIDTH(1) ) _51568_ ( .A(_tmp_1104), .B(1'h0), .S(_06505_), .Y(_27342_) );
  \$mux  #( .WIDTH(1) ) _51569_ ( .A(_27342_), .B(1'h1), .S(_06506_), .Y(_27343_) );
  \$mux  #( .WIDTH(1) ) _51570_ ( .A(_27343_), .B(1'h0), .S(RST), .Y(_02891_) );
  \$mux  #( .WIDTH(1) ) _51571_ ( .A(_tmp_1103), .B(1'h0), .S(_06506_), .Y(_27344_) );
  \$mux  #( .WIDTH(1) ) _51572_ ( .A(_27344_), .B(1'h1), .S(_06507_), .Y(_27345_) );
  \$mux  #( .WIDTH(1) ) _51573_ ( .A(_27345_), .B(1'h1), .S(_06508_), .Y(_27346_) );
  \$mux  #( .WIDTH(1) ) _51574_ ( .A(_27346_), .B(1'h0), .S(RST), .Y(_02890_) );
  \$mux  #( .WIDTH(8) ) _51575_ ( .A(_tmp_1102), .B(8'h00), .S(RST), .Y(_01136_) );
  \$mux  #( .WIDTH(1) ) _51576_ ( .A(_tmp_1101), .B(1'h0), .S(RST), .Y(_01135_) );
  \$mux  #( .WIDTH(1) ) _51577_ ( .A(_tmp_1096), .B(1'h0), .S(_06505_), .Y(_27347_) );
  \$mux  #( .WIDTH(1) ) _51578_ ( .A(_27347_), .B(1'h1), .S(_06506_), .Y(_27348_) );
  \$mux  #( .WIDTH(1) ) _51579_ ( .A(_27348_), .B(1'h0), .S(RST), .Y(_02888_) );
  \$mux  #( .WIDTH(1) ) _51580_ ( .A(_06504_), .B(1'h0), .S(RST), .Y(_01827_) );
  \$mux  #( .WIDTH(1) ) _51581_ ( .A(_tmp_30), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27349_) );
  \$mux  #( .WIDTH(1) ) _51582_ ( .A(_27349_), .B(1'h1), .S(_06503_), .Y(_27350_) );
  \$mux  #( .WIDTH(1) ) _51583_ ( .A(_27350_), .B(1'h0), .S(RST), .Y(_03056_) );
  \$mux  #( .WIDTH(34) ) _51584_ ( .A(_tmp_29), .B({ 1'h0, _maxi_read_size }), .S(_06502_), .Y(_27351_) );
  \$mux  #( .WIDTH(34) ) _51585_ ( .A(_27351_), .B(_28567_), .S(_06214_), .Y(_27352_) );
  \$mux  #( .WIDTH(34) ) _51586_ ( .A(_27352_), .B(34'h000000000), .S(RST), .Y(_03047_) );
  \$mux  #( .WIDTH(1) ) _51587_ ( .A(ram_w8_l2048_id0_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27353_) );
  \$mux  #( .WIDTH(1) ) _51588_ ( .A(_27353_), .B(1'h1), .S(_06214_), .Y(_27354_) );
  \$mux  #( .WIDTH(1) ) _51589_ ( .A(_27354_), .B(1'h0), .S(RST), .Y(_03678_) );
  \$mux  #( .WIDTH(8) ) _51590_ ( .A(ram_w8_l2048_id0_2_1_wdata), .B(_dataflow_slice_data_22), .S(_06214_), .Y(_27355_) );
  \$mux  #( .WIDTH(8) ) _51591_ ( .A(_27355_), .B(8'h00), .S(RST), .Y(_03677_) );
  \$mux  #( .WIDTH(9) ) _51592_ ( .A(ram_w8_l2048_id0_2_1_addr), .B(_28537_[8:0]), .S(_06502_), .Y(_27356_) );
  \$mux  #( .WIDTH(9) ) _51593_ ( .A(_27356_), .B(_24254_[8:0]), .S(_06214_), .Y(_27357_) );
  \$mux  #( .WIDTH(9) ) _51594_ ( .A(_27357_), .B(_maxi_write_local_addr[8:0]), .S(_06507_), .Y(_27358_) );
  \$mux  #( .WIDTH(9) ) _51595_ ( .A(_27358_), .B(_24255_[8:0]), .S(_06508_), .Y(_27359_) );
  \$mux  #( .WIDTH(9) ) _51596_ ( .A(_27359_), .B(9'h000), .S(RST), .Y(_03676_) );
  \$mux  #( .WIDTH(1) ) _51597_ ( .A(ram_w8_l2048_id0_2_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_2_cond_3_1), .Y(_27360_) );
  \$mux  #( .WIDTH(1) ) _51598_ ( .A(_27360_), .B(1'h1), .S(_06504_), .Y(_27361_) );
  \$mux  #( .WIDTH(1) ) _51599_ ( .A(_27361_), .B(1'h0), .S(RST), .Y(_03675_) );
  \$mux  #( .WIDTH(8) ) _51600_ ( .A(ram_w8_l2048_id0_2_0_wdata), .B(_stream_max_pool_serial_18_sink_3_sink_wdata), .S(_06504_), .Y(_27362_) );
  \$mux  #( .WIDTH(8) ) _51601_ ( .A(_27362_), .B(8'h00), .S(RST), .Y(_03674_) );
  \$mux  #( .WIDTH(9) ) _51602_ ( .A(ram_w8_l2048_id0_2_0_addr), .B(_stream_conv2d_16_source_8_source_ram_raddr[10:2]), .S(_tmp_483), .Y(_27363_) );
  \$mux  #( .WIDTH(9) ) _51603_ ( .A(_27363_), .B(_stream_max_pool_serial_18_sink_3_sink_waddr[10:2]), .S(_06504_), .Y(_27364_) );
  \$mux  #( .WIDTH(9) ) _51604_ ( .A(_27364_), .B(_stream_matmul_29_source_8_source_ram_raddr[10:2]), .S(_tmp_1189), .Y(_27365_) );
  \$mux  #( .WIDTH(9) ) _51605_ ( .A(_27365_), .B(9'h000), .S(RST), .Y(_03673_) );
  \$mux  #( .WIDTH(34) ) _51606_ ( .A(_tmp_1095), .B(_28563_), .S(_06499_), .Y(_27366_) );
  \$mux  #( .WIDTH(34) ) _51607_ ( .A(_27366_), .B(_28566_), .S(_06500_), .Y(_27367_) );
  \$mux  #( .WIDTH(34) ) _51608_ ( .A(_27367_), .B(34'h000000000), .S(RST), .Y(_02887_) );
  \$mux  #( .WIDTH(1) ) _51609_ ( .A(_tmp_1094), .B(1'h0), .S(_06497_), .Y(_27368_) );
  \$mux  #( .WIDTH(1) ) _51610_ ( .A(_27368_), .B(_tmp_1093), .S(_06498_), .Y(_27369_) );
  \$mux  #( .WIDTH(1) ) _51611_ ( .A(_27369_), .B(1'h0), .S(RST), .Y(_02886_) );
  \$mux  #( .WIDTH(1) ) _51612_ ( .A(_tmp_1093), .B(1'h0), .S(_06498_), .Y(_27370_) );
  \$mux  #( .WIDTH(1) ) _51613_ ( .A(_27370_), .B(_06099_), .S(_06499_), .Y(_27371_) );
  \$mux  #( .WIDTH(1) ) _51614_ ( .A(_27371_), .B(1'h0), .S(_06500_), .Y(_27372_) );
  \$mux  #( .WIDTH(1) ) _51615_ ( .A(_27372_), .B(1'h1), .S(_06501_), .Y(_27373_) );
  \$mux  #( .WIDTH(1) ) _51616_ ( .A(_27373_), .B(1'h0), .S(RST), .Y(_02885_) );
  \$mux  #( .WIDTH(1) ) _51617_ ( .A(_tmp_1092), .B(1'h0), .S(_06497_), .Y(_27374_) );
  \$mux  #( .WIDTH(1) ) _51618_ ( .A(_27374_), .B(1'h1), .S(_06498_), .Y(_27375_) );
  \$mux  #( .WIDTH(1) ) _51619_ ( .A(_27375_), .B(1'h0), .S(RST), .Y(_02884_) );
  \$mux  #( .WIDTH(1) ) _51620_ ( .A(_tmp_1091), .B(1'h0), .S(_06498_), .Y(_27376_) );
  \$mux  #( .WIDTH(1) ) _51621_ ( .A(_27376_), .B(1'h1), .S(_06499_), .Y(_27377_) );
  \$mux  #( .WIDTH(1) ) _51622_ ( .A(_27377_), .B(1'h1), .S(_06500_), .Y(_27378_) );
  \$mux  #( .WIDTH(1) ) _51623_ ( .A(_27378_), .B(1'h0), .S(RST), .Y(_02883_) );
  \$mux  #( .WIDTH(8) ) _51624_ ( .A(_tmp_1090), .B(8'h00), .S(RST), .Y(_01134_) );
  \$mux  #( .WIDTH(1) ) _51625_ ( .A(_tmp_1089), .B(1'h0), .S(RST), .Y(_01133_) );
  \$mux  #( .WIDTH(1) ) _51626_ ( .A(_tmp_1084), .B(1'h0), .S(_06497_), .Y(_27379_) );
  \$mux  #( .WIDTH(1) ) _51627_ ( .A(_27379_), .B(1'h1), .S(_06498_), .Y(_27380_) );
  \$mux  #( .WIDTH(1) ) _51628_ ( .A(_27380_), .B(1'h0), .S(RST), .Y(_02881_) );
  \$mux  #( .WIDTH(1) ) _51629_ ( .A(_06496_), .B(1'h0), .S(RST), .Y(_01826_) );
  \$mux  #( .WIDTH(1) ) _51630_ ( .A(_tmp_28), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27381_) );
  \$mux  #( .WIDTH(1) ) _51631_ ( .A(_27381_), .B(1'h1), .S(_06495_), .Y(_27382_) );
  \$mux  #( .WIDTH(1) ) _51632_ ( .A(_27382_), .B(1'h0), .S(RST), .Y(_03040_) );
  \$mux  #( .WIDTH(34) ) _51633_ ( .A(_tmp_27), .B({ 1'h0, _maxi_read_size }), .S(_06494_), .Y(_27383_) );
  \$mux  #( .WIDTH(34) ) _51634_ ( .A(_27383_), .B(_28565_), .S(_06211_), .Y(_27384_) );
  \$mux  #( .WIDTH(34) ) _51635_ ( .A(_27384_), .B(34'h000000000), .S(RST), .Y(_03038_) );
  \$mux  #( .WIDTH(1) ) _51636_ ( .A(ram_w8_l2048_id0_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27385_) );
  \$mux  #( .WIDTH(1) ) _51637_ ( .A(_27385_), .B(1'h1), .S(_06211_), .Y(_27386_) );
  \$mux  #( .WIDTH(1) ) _51638_ ( .A(_27386_), .B(1'h0), .S(RST), .Y(_03672_) );
  \$mux  #( .WIDTH(8) ) _51639_ ( .A(ram_w8_l2048_id0_1_1_wdata), .B(_dataflow_slice_data_19), .S(_06211_), .Y(_27387_) );
  \$mux  #( .WIDTH(8) ) _51640_ ( .A(_27387_), .B(8'h00), .S(RST), .Y(_03671_) );
  \$mux  #( .WIDTH(9) ) _51641_ ( .A(ram_w8_l2048_id0_1_1_addr), .B(_28537_[8:0]), .S(_06494_), .Y(_27388_) );
  \$mux  #( .WIDTH(9) ) _51642_ ( .A(_27388_), .B(_24252_[8:0]), .S(_06211_), .Y(_27389_) );
  \$mux  #( .WIDTH(9) ) _51643_ ( .A(_27389_), .B(_maxi_write_local_addr[8:0]), .S(_06499_), .Y(_27390_) );
  \$mux  #( .WIDTH(9) ) _51644_ ( .A(_27390_), .B(_24253_[8:0]), .S(_06500_), .Y(_27391_) );
  \$mux  #( .WIDTH(9) ) _51645_ ( .A(_27391_), .B(9'h000), .S(RST), .Y(_03670_) );
  \$mux  #( .WIDTH(1) ) _51646_ ( .A(ram_w8_l2048_id0_1_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_1_cond_3_1), .Y(_27392_) );
  \$mux  #( .WIDTH(1) ) _51647_ ( .A(_27392_), .B(1'h1), .S(_06496_), .Y(_27393_) );
  \$mux  #( .WIDTH(1) ) _51648_ ( .A(_27393_), .B(1'h0), .S(RST), .Y(_03669_) );
  \$mux  #( .WIDTH(8) ) _51649_ ( .A(ram_w8_l2048_id0_1_0_wdata), .B(_stream_max_pool_serial_18_sink_3_sink_wdata), .S(_06496_), .Y(_27394_) );
  \$mux  #( .WIDTH(8) ) _51650_ ( .A(_27394_), .B(8'h00), .S(RST), .Y(_03668_) );
  \$mux  #( .WIDTH(9) ) _51651_ ( .A(ram_w8_l2048_id0_1_0_addr), .B(_stream_conv2d_16_source_8_source_ram_raddr[10:2]), .S(_tmp_483), .Y(_27395_) );
  \$mux  #( .WIDTH(9) ) _51652_ ( .A(_27395_), .B(_stream_max_pool_serial_18_sink_3_sink_waddr[10:2]), .S(_06496_), .Y(_27396_) );
  \$mux  #( .WIDTH(9) ) _51653_ ( .A(_27396_), .B(_stream_matmul_29_source_8_source_ram_raddr[10:2]), .S(_tmp_1189), .Y(_27397_) );
  \$mux  #( .WIDTH(9) ) _51654_ ( .A(_27397_), .B(9'h000), .S(RST), .Y(_03667_) );
  \$mux  #( .WIDTH(1) ) _51655_ ( .A(_dataflow_cat_valid_107), .B(1'h0), .S(_06190_), .Y(_27398_) );
  \$mux  #( .WIDTH(1) ) _51656_ ( .A(_27398_), .B(_06492_), .S(_06493_), .Y(_27399_) );
  \$mux  #( .WIDTH(1) ) _51657_ ( .A(_27399_), .B(1'h0), .S(RST), .Y(_01589_) );
  \$mux  #( .WIDTH(32) ) _51658_ ( .A(_dataflow_cat_data_107), .B({ _tmp_1114, _tmp_1102, _tmp_1090, _tmp_1078 }), .S(_06493_), .Y(_27400_) );
  \$mux  #( .WIDTH(32) ) _51659_ ( .A(_27400_), .B(0), .S(RST), .Y(_01586_) );
  \$mux  #( .WIDTH(1) ) _51660_ ( .A(_tmp_1189), .B(1'h0), .S(RST), .Y(_01144_) );
  \$mux  #( .WIDTH(34) ) _51661_ ( .A(_tmp_1083), .B(_28563_), .S(_06489_), .Y(_27401_) );
  \$mux  #( .WIDTH(34) ) _51662_ ( .A(_27401_), .B(_28564_), .S(_06490_), .Y(_27402_) );
  \$mux  #( .WIDTH(34) ) _51663_ ( .A(_27402_), .B(34'h000000000), .S(RST), .Y(_02880_) );
  \$mux  #( .WIDTH(1) ) _51664_ ( .A(_tmp_1082), .B(1'h0), .S(_06486_), .Y(_27403_) );
  \$mux  #( .WIDTH(1) ) _51665_ ( .A(_27403_), .B(_tmp_1081), .S(_06487_), .Y(_27404_) );
  \$mux  #( .WIDTH(1) ) _51666_ ( .A(_27404_), .B(1'h0), .S(RST), .Y(_02879_) );
  \$mux  #( .WIDTH(1) ) _51667_ ( .A(_tmp_1081), .B(1'h0), .S(_06487_), .Y(_27405_) );
  \$mux  #( .WIDTH(1) ) _51668_ ( .A(_27405_), .B(_06099_), .S(_06489_), .Y(_27406_) );
  \$mux  #( .WIDTH(1) ) _51669_ ( .A(_27406_), .B(1'h0), .S(_06490_), .Y(_27407_) );
  \$mux  #( .WIDTH(1) ) _51670_ ( .A(_27407_), .B(1'h1), .S(_06491_), .Y(_27408_) );
  \$mux  #( .WIDTH(1) ) _51671_ ( .A(_27408_), .B(1'h0), .S(RST), .Y(_02878_) );
  \$mux  #( .WIDTH(1) ) _51672_ ( .A(_tmp_1080), .B(1'h0), .S(_06486_), .Y(_27409_) );
  \$mux  #( .WIDTH(1) ) _51673_ ( .A(_27409_), .B(1'h1), .S(_06487_), .Y(_27410_) );
  \$mux  #( .WIDTH(1) ) _51674_ ( .A(_27410_), .B(1'h0), .S(RST), .Y(_02877_) );
  \$mux  #( .WIDTH(1) ) _51675_ ( .A(_tmp_1079), .B(1'h0), .S(_06487_), .Y(_27411_) );
  \$mux  #( .WIDTH(1) ) _51676_ ( .A(_27411_), .B(1'h1), .S(_06489_), .Y(_27412_) );
  \$mux  #( .WIDTH(1) ) _51677_ ( .A(_27412_), .B(1'h1), .S(_06490_), .Y(_27413_) );
  \$mux  #( .WIDTH(1) ) _51678_ ( .A(_27413_), .B(1'h0), .S(RST), .Y(_02875_) );
  \$mux  #( .WIDTH(8) ) _51679_ ( .A(_tmp_1078), .B(8'h00), .S(RST), .Y(_01132_) );
  \$mux  #( .WIDTH(1) ) _51680_ ( .A(_tmp_1077), .B(1'h0), .S(RST), .Y(_01131_) );
  \$mux  #( .WIDTH(1) ) _51681_ ( .A(_tmp_1072), .B(1'h0), .S(_06486_), .Y(_27414_) );
  \$mux  #( .WIDTH(1) ) _51682_ ( .A(_27414_), .B(1'h1), .S(_06487_), .Y(_27415_) );
  \$mux  #( .WIDTH(1) ) _51683_ ( .A(_27415_), .B(1'h0), .S(RST), .Y(_02874_) );
  \$mux  #( .WIDTH(1) ) _51684_ ( .A(_06485_), .B(1'h0), .S(RST), .Y(_01825_) );
  \$mux  #( .WIDTH(1) ) _51685_ ( .A(_tmp_483), .B(1'h0), .S(RST), .Y(_01234_) );
  \$mux  #( .WIDTH(1) ) _51686_ ( .A(_tmp_26), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27416_) );
  \$mux  #( .WIDTH(1) ) _51687_ ( .A(_27416_), .B(1'h1), .S(_06484_), .Y(_27417_) );
  \$mux  #( .WIDTH(1) ) _51688_ ( .A(_27417_), .B(1'h0), .S(RST), .Y(_03037_) );
  \$mux  #( .WIDTH(34) ) _51689_ ( .A(_tmp_25), .B({ 1'h0, _maxi_read_size }), .S(_06483_), .Y(_27418_) );
  \$mux  #( .WIDTH(34) ) _51690_ ( .A(_27418_), .B(_28562_), .S(_06208_), .Y(_27419_) );
  \$mux  #( .WIDTH(34) ) _51691_ ( .A(_27419_), .B(34'h000000000), .S(RST), .Y(_03029_) );
  \$mux  #( .WIDTH(1) ) _51692_ ( .A(ram_w8_l2048_id0_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27420_) );
  \$mux  #( .WIDTH(1) ) _51693_ ( .A(_27420_), .B(1'h1), .S(_06208_), .Y(_27421_) );
  \$mux  #( .WIDTH(1) ) _51694_ ( .A(_27421_), .B(1'h0), .S(RST), .Y(_03666_) );
  \$mux  #( .WIDTH(8) ) _51695_ ( .A(ram_w8_l2048_id0_0_1_wdata), .B(_dataflow_slice_data_16), .S(_06208_), .Y(_27422_) );
  \$mux  #( .WIDTH(8) ) _51696_ ( .A(_27422_), .B(8'h00), .S(RST), .Y(_03665_) );
  \$mux  #( .WIDTH(9) ) _51697_ ( .A(ram_w8_l2048_id0_0_1_addr), .B(_28537_[8:0]), .S(_06483_), .Y(_27423_) );
  \$mux  #( .WIDTH(9) ) _51698_ ( .A(_27423_), .B(_24250_[8:0]), .S(_06208_), .Y(_27424_) );
  \$mux  #( .WIDTH(9) ) _51699_ ( .A(_27424_), .B(_maxi_write_local_addr[8:0]), .S(_06489_), .Y(_27425_) );
  \$mux  #( .WIDTH(9) ) _51700_ ( .A(_27425_), .B(_24251_[8:0]), .S(_06490_), .Y(_27426_) );
  \$mux  #( .WIDTH(9) ) _51701_ ( .A(_27426_), .B(9'h000), .S(RST), .Y(_03664_) );
  \$mux  #( .WIDTH(1) ) _51702_ ( .A(ram_w8_l2048_id0_0_0_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_0_cond_3_1), .Y(_27427_) );
  \$mux  #( .WIDTH(1) ) _51703_ ( .A(_27427_), .B(1'h1), .S(_06485_), .Y(_27428_) );
  \$mux  #( .WIDTH(1) ) _51704_ ( .A(_27428_), .B(1'h0), .S(RST), .Y(_03663_) );
  \$mux  #( .WIDTH(8) ) _51705_ ( .A(ram_w8_l2048_id0_0_0_wdata), .B(_stream_max_pool_serial_18_sink_3_sink_wdata), .S(_06485_), .Y(_27429_) );
  \$mux  #( .WIDTH(8) ) _51706_ ( .A(_27429_), .B(8'h00), .S(RST), .Y(_03662_) );
  \$mux  #( .WIDTH(9) ) _51707_ ( .A(ram_w8_l2048_id0_0_0_addr), .B(_stream_conv2d_16_source_8_source_ram_raddr[10:2]), .S(_tmp_483), .Y(_27430_) );
  \$mux  #( .WIDTH(9) ) _51708_ ( .A(_27430_), .B(_stream_max_pool_serial_18_sink_3_sink_waddr[10:2]), .S(_06485_), .Y(_27431_) );
  \$mux  #( .WIDTH(9) ) _51709_ ( .A(_27431_), .B(_stream_matmul_29_source_8_source_ram_raddr[10:2]), .S(_tmp_1189), .Y(_27432_) );
  \$mux  #( .WIDTH(9) ) _51710_ ( .A(_27432_), .B(9'h000), .S(RST), .Y(_03661_) );
  \$mux  #( .WIDTH(1) ) _51711_ ( .A(ram_w4_l8192_id8_7_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27433_) );
  \$mux  #( .WIDTH(1) ) _51712_ ( .A(_27433_), .B(_06090_), .S(_06241_), .Y(_27434_) );
  \$mux  #( .WIDTH(1) ) _51713_ ( .A(_27434_), .B(1'h0), .S(RST), .Y(_03660_) );
  \$mux  #( .WIDTH(4) ) _51714_ ( .A(ram_w4_l8192_id8_7_1_wdata), .B(_dataflow_slice_data_50), .S(_06241_), .Y(_27435_) );
  \$mux  #( .WIDTH(4) ) _51715_ ( .A(_27435_), .B(4'h0), .S(RST), .Y(_03659_) );
  \$mux  #( .WIDTH(10) ) _51716_ ( .A(ram_w4_l8192_id8_7_1_addr), .B(_tmp_275), .S(_06241_), .Y(_27436_) );
  \$mux  #( .WIDTH(10) ) _51717_ ( .A(_27436_), .B(10'h000), .S(RST), .Y(_03658_) );
  \$mux  #( .WIDTH(10) ) _51718_ ( .A(ram_w4_l8192_id8_7_0_addr), .B(_stream_conv2d_16_source_36_source_ram_raddr[12:3]), .S(_tmp_709), .Y(_27437_) );
  \$mux  #( .WIDTH(10) ) _51719_ ( .A(_27437_), .B(10'h000), .S(RST), .Y(_03657_) );
  \$mux  #( .WIDTH(1) ) _51720_ ( .A(ram_w4_l8192_id8_6_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27438_) );
  \$mux  #( .WIDTH(1) ) _51721_ ( .A(_27438_), .B(_06081_), .S(_06238_), .Y(_27439_) );
  \$mux  #( .WIDTH(1) ) _51722_ ( .A(_27439_), .B(1'h0), .S(RST), .Y(_03656_) );
  \$mux  #( .WIDTH(4) ) _51723_ ( .A(ram_w4_l8192_id8_6_1_wdata), .B(_dataflow_slice_data_47), .S(_06238_), .Y(_27440_) );
  \$mux  #( .WIDTH(4) ) _51724_ ( .A(_27440_), .B(4'h0), .S(RST), .Y(_03655_) );
  \$mux  #( .WIDTH(10) ) _51725_ ( .A(ram_w4_l8192_id8_6_1_addr), .B(_tmp_244), .S(_06238_), .Y(_27441_) );
  \$mux  #( .WIDTH(10) ) _51726_ ( .A(_27441_), .B(10'h000), .S(RST), .Y(_03654_) );
  \$mux  #( .WIDTH(10) ) _51727_ ( .A(ram_w4_l8192_id8_6_0_addr), .B(_stream_conv2d_16_source_36_source_ram_raddr[12:3]), .S(_tmp_709), .Y(_27442_) );
  \$mux  #( .WIDTH(10) ) _51728_ ( .A(_27442_), .B(10'h000), .S(RST), .Y(_03653_) );
  \$mux  #( .WIDTH(1) ) _51729_ ( .A(ram_w4_l8192_id8_5_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27443_) );
  \$mux  #( .WIDTH(1) ) _51730_ ( .A(_27443_), .B(_06072_), .S(_06235_), .Y(_27444_) );
  \$mux  #( .WIDTH(1) ) _51731_ ( .A(_27444_), .B(1'h0), .S(RST), .Y(_03652_) );
  \$mux  #( .WIDTH(4) ) _51732_ ( .A(ram_w4_l8192_id8_5_1_wdata), .B(_dataflow_slice_data_44), .S(_06235_), .Y(_27445_) );
  \$mux  #( .WIDTH(4) ) _51733_ ( .A(_27445_), .B(4'h0), .S(RST), .Y(_03651_) );
  \$mux  #( .WIDTH(10) ) _51734_ ( .A(ram_w4_l8192_id8_5_1_addr), .B(_tmp_213), .S(_06235_), .Y(_27446_) );
  \$mux  #( .WIDTH(10) ) _51735_ ( .A(_27446_), .B(10'h000), .S(RST), .Y(_03650_) );
  \$mux  #( .WIDTH(10) ) _51736_ ( .A(ram_w4_l8192_id8_5_0_addr), .B(_stream_conv2d_16_source_36_source_ram_raddr[12:3]), .S(_tmp_709), .Y(_27447_) );
  \$mux  #( .WIDTH(10) ) _51737_ ( .A(_27447_), .B(10'h000), .S(RST), .Y(_03649_) );
  \$mux  #( .WIDTH(1) ) _51738_ ( .A(ram_w4_l8192_id8_4_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27448_) );
  \$mux  #( .WIDTH(1) ) _51739_ ( .A(_27448_), .B(_06063_), .S(_06232_), .Y(_27449_) );
  \$mux  #( .WIDTH(1) ) _51740_ ( .A(_27449_), .B(1'h0), .S(RST), .Y(_03648_) );
  \$mux  #( .WIDTH(4) ) _51741_ ( .A(ram_w4_l8192_id8_4_1_wdata), .B(_dataflow_slice_data_41), .S(_06232_), .Y(_27450_) );
  \$mux  #( .WIDTH(4) ) _51742_ ( .A(_27450_), .B(4'h0), .S(RST), .Y(_03647_) );
  \$mux  #( .WIDTH(10) ) _51743_ ( .A(ram_w4_l8192_id8_4_1_addr), .B(_tmp_182), .S(_06232_), .Y(_27451_) );
  \$mux  #( .WIDTH(10) ) _51744_ ( .A(_27451_), .B(10'h000), .S(RST), .Y(_03646_) );
  \$mux  #( .WIDTH(10) ) _51745_ ( .A(ram_w4_l8192_id8_4_0_addr), .B(_stream_conv2d_16_source_36_source_ram_raddr[12:3]), .S(_tmp_709), .Y(_27452_) );
  \$mux  #( .WIDTH(10) ) _51746_ ( .A(_27452_), .B(10'h000), .S(RST), .Y(_03645_) );
  \$mux  #( .WIDTH(1) ) _51747_ ( .A(ram_w4_l8192_id8_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27453_) );
  \$mux  #( .WIDTH(1) ) _51748_ ( .A(_27453_), .B(_06054_), .S(_06229_), .Y(_27454_) );
  \$mux  #( .WIDTH(1) ) _51749_ ( .A(_27454_), .B(1'h0), .S(RST), .Y(_03644_) );
  \$mux  #( .WIDTH(4) ) _51750_ ( .A(ram_w4_l8192_id8_3_1_wdata), .B(_dataflow_slice_data_38), .S(_06229_), .Y(_27455_) );
  \$mux  #( .WIDTH(4) ) _51751_ ( .A(_27455_), .B(4'h0), .S(RST), .Y(_03643_) );
  \$mux  #( .WIDTH(10) ) _51752_ ( .A(ram_w4_l8192_id8_3_1_addr), .B(_tmp_151), .S(_06229_), .Y(_27456_) );
  \$mux  #( .WIDTH(10) ) _51753_ ( .A(_27456_), .B(10'h000), .S(RST), .Y(_03642_) );
  \$mux  #( .WIDTH(10) ) _51754_ ( .A(ram_w4_l8192_id8_3_0_addr), .B(_stream_conv2d_16_source_36_source_ram_raddr[12:3]), .S(_tmp_709), .Y(_27457_) );
  \$mux  #( .WIDTH(10) ) _51755_ ( .A(_27457_), .B(10'h000), .S(RST), .Y(_03641_) );
  \$mux  #( .WIDTH(1) ) _51756_ ( .A(ram_w4_l8192_id8_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27458_) );
  \$mux  #( .WIDTH(1) ) _51757_ ( .A(_27458_), .B(_06045_), .S(_06226_), .Y(_27459_) );
  \$mux  #( .WIDTH(1) ) _51758_ ( .A(_27459_), .B(1'h0), .S(RST), .Y(_03640_) );
  \$mux  #( .WIDTH(4) ) _51759_ ( .A(ram_w4_l8192_id8_2_1_wdata), .B(_dataflow_slice_data_35), .S(_06226_), .Y(_27460_) );
  \$mux  #( .WIDTH(4) ) _51760_ ( .A(_27460_), .B(4'h0), .S(RST), .Y(_03639_) );
  \$mux  #( .WIDTH(10) ) _51761_ ( .A(ram_w4_l8192_id8_2_1_addr), .B(_tmp_120), .S(_06226_), .Y(_27461_) );
  \$mux  #( .WIDTH(10) ) _51762_ ( .A(_27461_), .B(10'h000), .S(RST), .Y(_03638_) );
  \$mux  #( .WIDTH(10) ) _51763_ ( .A(ram_w4_l8192_id8_2_0_addr), .B(_stream_conv2d_16_source_36_source_ram_raddr[12:3]), .S(_tmp_709), .Y(_27462_) );
  \$mux  #( .WIDTH(10) ) _51764_ ( .A(_27462_), .B(10'h000), .S(RST), .Y(_03637_) );
  \$mux  #( .WIDTH(1) ) _51765_ ( .A(ram_w4_l8192_id8_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27463_) );
  \$mux  #( .WIDTH(1) ) _51766_ ( .A(_27463_), .B(_06036_), .S(_06223_), .Y(_27464_) );
  \$mux  #( .WIDTH(1) ) _51767_ ( .A(_27464_), .B(1'h0), .S(RST), .Y(_03636_) );
  \$mux  #( .WIDTH(4) ) _51768_ ( .A(ram_w4_l8192_id8_1_1_wdata), .B(_dataflow_slice_data_32), .S(_06223_), .Y(_27465_) );
  \$mux  #( .WIDTH(4) ) _51769_ ( .A(_27465_), .B(4'h0), .S(RST), .Y(_03635_) );
  \$mux  #( .WIDTH(10) ) _51770_ ( .A(ram_w4_l8192_id8_1_1_addr), .B(_tmp_89), .S(_06223_), .Y(_27466_) );
  \$mux  #( .WIDTH(10) ) _51771_ ( .A(_27466_), .B(10'h000), .S(RST), .Y(_03634_) );
  \$mux  #( .WIDTH(10) ) _51772_ ( .A(ram_w4_l8192_id8_1_0_addr), .B(_stream_conv2d_16_source_36_source_ram_raddr[12:3]), .S(_tmp_709), .Y(_27467_) );
  \$mux  #( .WIDTH(10) ) _51773_ ( .A(_27467_), .B(10'h000), .S(RST), .Y(_03633_) );
  \$mux  #( .WIDTH(1) ) _51774_ ( .A(_tmp_709), .B(1'h0), .S(RST), .Y(_01288_) );
  \$mux  #( .WIDTH(1) ) _51775_ ( .A(ram_w4_l8192_id8_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27468_) );
  \$mux  #( .WIDTH(1) ) _51776_ ( .A(_27468_), .B(_06027_), .S(_06220_), .Y(_27469_) );
  \$mux  #( .WIDTH(1) ) _51777_ ( .A(_27469_), .B(1'h0), .S(RST), .Y(_03632_) );
  \$mux  #( .WIDTH(4) ) _51778_ ( .A(ram_w4_l8192_id8_0_1_wdata), .B(_dataflow_slice_data_29), .S(_06220_), .Y(_27470_) );
  \$mux  #( .WIDTH(4) ) _51779_ ( .A(_27470_), .B(4'h0), .S(RST), .Y(_03631_) );
  \$mux  #( .WIDTH(10) ) _51780_ ( .A(ram_w4_l8192_id8_0_1_addr), .B(_tmp_58), .S(_06220_), .Y(_27471_) );
  \$mux  #( .WIDTH(10) ) _51781_ ( .A(_27471_), .B(10'h000), .S(RST), .Y(_03630_) );
  \$mux  #( .WIDTH(10) ) _51782_ ( .A(ram_w4_l8192_id8_0_0_addr), .B(_stream_conv2d_16_source_36_source_ram_raddr[12:3]), .S(_tmp_709), .Y(_27472_) );
  \$mux  #( .WIDTH(10) ) _51783_ ( .A(_27472_), .B(10'h000), .S(RST), .Y(_03629_) );
  \$mux  #( .WIDTH(1) ) _51784_ ( .A(ram_w4_l8192_id7_7_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27473_) );
  \$mux  #( .WIDTH(1) ) _51785_ ( .A(_27473_), .B(_06098_), .S(_06241_), .Y(_27474_) );
  \$mux  #( .WIDTH(1) ) _51786_ ( .A(_27474_), .B(1'h0), .S(RST), .Y(_03628_) );
  \$mux  #( .WIDTH(4) ) _51787_ ( .A(ram_w4_l8192_id7_7_1_wdata), .B(_dataflow_slice_data_50), .S(_06241_), .Y(_27475_) );
  \$mux  #( .WIDTH(4) ) _51788_ ( .A(_27475_), .B(4'h0), .S(RST), .Y(_03627_) );
  \$mux  #( .WIDTH(10) ) _51789_ ( .A(ram_w4_l8192_id7_7_1_addr), .B(_tmp_274), .S(_06241_), .Y(_27476_) );
  \$mux  #( .WIDTH(10) ) _51790_ ( .A(_27476_), .B(10'h000), .S(RST), .Y(_03626_) );
  \$mux  #( .WIDTH(10) ) _51791_ ( .A(ram_w4_l8192_id7_7_0_addr), .B(_stream_conv2d_16_source_35_source_ram_raddr[12:3]), .S(_tmp_695), .Y(_27477_) );
  \$mux  #( .WIDTH(10) ) _51792_ ( .A(_27477_), .B(10'h000), .S(RST), .Y(_03625_) );
  \$mux  #( .WIDTH(1) ) _51793_ ( .A(ram_w4_l8192_id7_6_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27478_) );
  \$mux  #( .WIDTH(1) ) _51794_ ( .A(_27478_), .B(_06089_), .S(_06238_), .Y(_27479_) );
  \$mux  #( .WIDTH(1) ) _51795_ ( .A(_27479_), .B(1'h0), .S(RST), .Y(_03624_) );
  \$mux  #( .WIDTH(4) ) _51796_ ( .A(ram_w4_l8192_id7_6_1_wdata), .B(_dataflow_slice_data_47), .S(_06238_), .Y(_27480_) );
  \$mux  #( .WIDTH(4) ) _51797_ ( .A(_27480_), .B(4'h0), .S(RST), .Y(_03623_) );
  \$mux  #( .WIDTH(10) ) _51798_ ( .A(ram_w4_l8192_id7_6_1_addr), .B(_tmp_243), .S(_06238_), .Y(_27481_) );
  \$mux  #( .WIDTH(10) ) _51799_ ( .A(_27481_), .B(10'h000), .S(RST), .Y(_03622_) );
  \$mux  #( .WIDTH(10) ) _51800_ ( .A(ram_w4_l8192_id7_6_0_addr), .B(_stream_conv2d_16_source_35_source_ram_raddr[12:3]), .S(_tmp_695), .Y(_27482_) );
  \$mux  #( .WIDTH(10) ) _51801_ ( .A(_27482_), .B(10'h000), .S(RST), .Y(_03621_) );
  \$mux  #( .WIDTH(1) ) _51802_ ( .A(ram_w4_l8192_id7_5_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27483_) );
  \$mux  #( .WIDTH(1) ) _51803_ ( .A(_27483_), .B(_06080_), .S(_06235_), .Y(_27484_) );
  \$mux  #( .WIDTH(1) ) _51804_ ( .A(_27484_), .B(1'h0), .S(RST), .Y(_03620_) );
  \$mux  #( .WIDTH(4) ) _51805_ ( .A(ram_w4_l8192_id7_5_1_wdata), .B(_dataflow_slice_data_44), .S(_06235_), .Y(_27485_) );
  \$mux  #( .WIDTH(4) ) _51806_ ( .A(_27485_), .B(4'h0), .S(RST), .Y(_03619_) );
  \$mux  #( .WIDTH(10) ) _51807_ ( .A(ram_w4_l8192_id7_5_1_addr), .B(_tmp_212), .S(_06235_), .Y(_27486_) );
  \$mux  #( .WIDTH(10) ) _51808_ ( .A(_27486_), .B(10'h000), .S(RST), .Y(_03618_) );
  \$mux  #( .WIDTH(10) ) _51809_ ( .A(ram_w4_l8192_id7_5_0_addr), .B(_stream_conv2d_16_source_35_source_ram_raddr[12:3]), .S(_tmp_695), .Y(_27487_) );
  \$mux  #( .WIDTH(10) ) _51810_ ( .A(_27487_), .B(10'h000), .S(RST), .Y(_03617_) );
  \$mux  #( .WIDTH(1) ) _51811_ ( .A(ram_w4_l8192_id7_4_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27488_) );
  \$mux  #( .WIDTH(1) ) _51812_ ( .A(_27488_), .B(_06071_), .S(_06232_), .Y(_27489_) );
  \$mux  #( .WIDTH(1) ) _51813_ ( .A(_27489_), .B(1'h0), .S(RST), .Y(_03616_) );
  \$mux  #( .WIDTH(4) ) _51814_ ( .A(ram_w4_l8192_id7_4_1_wdata), .B(_dataflow_slice_data_41), .S(_06232_), .Y(_27490_) );
  \$mux  #( .WIDTH(4) ) _51815_ ( .A(_27490_), .B(4'h0), .S(RST), .Y(_03615_) );
  \$mux  #( .WIDTH(10) ) _51816_ ( .A(ram_w4_l8192_id7_4_1_addr), .B(_tmp_181), .S(_06232_), .Y(_27491_) );
  \$mux  #( .WIDTH(10) ) _51817_ ( .A(_27491_), .B(10'h000), .S(RST), .Y(_03614_) );
  \$mux  #( .WIDTH(10) ) _51818_ ( .A(ram_w4_l8192_id7_4_0_addr), .B(_stream_conv2d_16_source_35_source_ram_raddr[12:3]), .S(_tmp_695), .Y(_27492_) );
  \$mux  #( .WIDTH(10) ) _51819_ ( .A(_27492_), .B(10'h000), .S(RST), .Y(_03613_) );
  \$mux  #( .WIDTH(1) ) _51820_ ( .A(ram_w4_l8192_id7_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27493_) );
  \$mux  #( .WIDTH(1) ) _51821_ ( .A(_27493_), .B(_06062_), .S(_06229_), .Y(_27494_) );
  \$mux  #( .WIDTH(1) ) _51822_ ( .A(_27494_), .B(1'h0), .S(RST), .Y(_03612_) );
  \$mux  #( .WIDTH(4) ) _51823_ ( .A(ram_w4_l8192_id7_3_1_wdata), .B(_dataflow_slice_data_38), .S(_06229_), .Y(_27495_) );
  \$mux  #( .WIDTH(4) ) _51824_ ( .A(_27495_), .B(4'h0), .S(RST), .Y(_03611_) );
  \$mux  #( .WIDTH(10) ) _51825_ ( .A(ram_w4_l8192_id7_3_1_addr), .B(_tmp_150), .S(_06229_), .Y(_27496_) );
  \$mux  #( .WIDTH(10) ) _51826_ ( .A(_27496_), .B(10'h000), .S(RST), .Y(_03610_) );
  \$mux  #( .WIDTH(10) ) _51827_ ( .A(ram_w4_l8192_id7_3_0_addr), .B(_stream_conv2d_16_source_35_source_ram_raddr[12:3]), .S(_tmp_695), .Y(_27497_) );
  \$mux  #( .WIDTH(10) ) _51828_ ( .A(_27497_), .B(10'h000), .S(RST), .Y(_03609_) );
  \$mux  #( .WIDTH(1) ) _51829_ ( .A(ram_w4_l8192_id7_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27498_) );
  \$mux  #( .WIDTH(1) ) _51830_ ( .A(_27498_), .B(_06053_), .S(_06226_), .Y(_27499_) );
  \$mux  #( .WIDTH(1) ) _51831_ ( .A(_27499_), .B(1'h0), .S(RST), .Y(_03608_) );
  \$mux  #( .WIDTH(4) ) _51832_ ( .A(ram_w4_l8192_id7_2_1_wdata), .B(_dataflow_slice_data_35), .S(_06226_), .Y(_27500_) );
  \$mux  #( .WIDTH(4) ) _51833_ ( .A(_27500_), .B(4'h0), .S(RST), .Y(_03607_) );
  \$mux  #( .WIDTH(10) ) _51834_ ( .A(ram_w4_l8192_id7_2_1_addr), .B(_tmp_119), .S(_06226_), .Y(_27501_) );
  \$mux  #( .WIDTH(10) ) _51835_ ( .A(_27501_), .B(10'h000), .S(RST), .Y(_03606_) );
  \$mux  #( .WIDTH(10) ) _51836_ ( .A(ram_w4_l8192_id7_2_0_addr), .B(_stream_conv2d_16_source_35_source_ram_raddr[12:3]), .S(_tmp_695), .Y(_27502_) );
  \$mux  #( .WIDTH(10) ) _51837_ ( .A(_27502_), .B(10'h000), .S(RST), .Y(_03605_) );
  \$mux  #( .WIDTH(1) ) _51838_ ( .A(ram_w4_l8192_id7_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27503_) );
  \$mux  #( .WIDTH(1) ) _51839_ ( .A(_27503_), .B(_06044_), .S(_06223_), .Y(_27504_) );
  \$mux  #( .WIDTH(1) ) _51840_ ( .A(_27504_), .B(1'h0), .S(RST), .Y(_03604_) );
  \$mux  #( .WIDTH(4) ) _51841_ ( .A(ram_w4_l8192_id7_1_1_wdata), .B(_dataflow_slice_data_32), .S(_06223_), .Y(_27505_) );
  \$mux  #( .WIDTH(4) ) _51842_ ( .A(_27505_), .B(4'h0), .S(RST), .Y(_03603_) );
  \$mux  #( .WIDTH(10) ) _51843_ ( .A(ram_w4_l8192_id7_1_1_addr), .B(_tmp_88), .S(_06223_), .Y(_27506_) );
  \$mux  #( .WIDTH(10) ) _51844_ ( .A(_27506_), .B(10'h000), .S(RST), .Y(_03602_) );
  \$mux  #( .WIDTH(10) ) _51845_ ( .A(ram_w4_l8192_id7_1_0_addr), .B(_stream_conv2d_16_source_35_source_ram_raddr[12:3]), .S(_tmp_695), .Y(_27507_) );
  \$mux  #( .WIDTH(10) ) _51846_ ( .A(_27507_), .B(10'h000), .S(RST), .Y(_03601_) );
  \$mux  #( .WIDTH(1) ) _51847_ ( .A(_tmp_695), .B(1'h0), .S(RST), .Y(_01285_) );
  \$mux  #( .WIDTH(1) ) _51848_ ( .A(ram_w4_l8192_id7_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27508_) );
  \$mux  #( .WIDTH(1) ) _51849_ ( .A(_27508_), .B(_06035_), .S(_06220_), .Y(_27509_) );
  \$mux  #( .WIDTH(1) ) _51850_ ( .A(_27509_), .B(1'h0), .S(RST), .Y(_03600_) );
  \$mux  #( .WIDTH(4) ) _51851_ ( .A(ram_w4_l8192_id7_0_1_wdata), .B(_dataflow_slice_data_29), .S(_06220_), .Y(_27510_) );
  \$mux  #( .WIDTH(4) ) _51852_ ( .A(_27510_), .B(4'h0), .S(RST), .Y(_03599_) );
  \$mux  #( .WIDTH(10) ) _51853_ ( .A(ram_w4_l8192_id7_0_1_addr), .B(_tmp_57), .S(_06220_), .Y(_27511_) );
  \$mux  #( .WIDTH(10) ) _51854_ ( .A(_27511_), .B(10'h000), .S(RST), .Y(_03598_) );
  \$mux  #( .WIDTH(10) ) _51855_ ( .A(ram_w4_l8192_id7_0_0_addr), .B(_stream_conv2d_16_source_35_source_ram_raddr[12:3]), .S(_tmp_695), .Y(_27512_) );
  \$mux  #( .WIDTH(10) ) _51856_ ( .A(_27512_), .B(10'h000), .S(RST), .Y(_03597_) );
  \$mux  #( .WIDTH(1) ) _51857_ ( .A(ram_w4_l8192_id6_7_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27513_) );
  \$mux  #( .WIDTH(1) ) _51858_ ( .A(_27513_), .B(_06097_), .S(_06241_), .Y(_27514_) );
  \$mux  #( .WIDTH(1) ) _51859_ ( .A(_27514_), .B(1'h0), .S(RST), .Y(_03596_) );
  \$mux  #( .WIDTH(4) ) _51860_ ( .A(ram_w4_l8192_id6_7_1_wdata), .B(_dataflow_slice_data_50), .S(_06241_), .Y(_27515_) );
  \$mux  #( .WIDTH(4) ) _51861_ ( .A(_27515_), .B(4'h0), .S(RST), .Y(_03595_) );
  \$mux  #( .WIDTH(10) ) _51862_ ( .A(ram_w4_l8192_id6_7_1_addr), .B(_tmp_273), .S(_06241_), .Y(_27516_) );
  \$mux  #( .WIDTH(10) ) _51863_ ( .A(_27516_), .B(10'h000), .S(RST), .Y(_03594_) );
  \$mux  #( .WIDTH(10) ) _51864_ ( .A(ram_w4_l8192_id6_7_0_addr), .B(_stream_conv2d_16_source_34_source_ram_raddr[12:3]), .S(_tmp_681), .Y(_27517_) );
  \$mux  #( .WIDTH(10) ) _51865_ ( .A(_27517_), .B(10'h000), .S(RST), .Y(_03593_) );
  \$mux  #( .WIDTH(1) ) _51866_ ( .A(ram_w4_l8192_id6_6_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27518_) );
  \$mux  #( .WIDTH(1) ) _51867_ ( .A(_27518_), .B(_06088_), .S(_06238_), .Y(_27519_) );
  \$mux  #( .WIDTH(1) ) _51868_ ( .A(_27519_), .B(1'h0), .S(RST), .Y(_03592_) );
  \$mux  #( .WIDTH(4) ) _51869_ ( .A(ram_w4_l8192_id6_6_1_wdata), .B(_dataflow_slice_data_47), .S(_06238_), .Y(_27520_) );
  \$mux  #( .WIDTH(4) ) _51870_ ( .A(_27520_), .B(4'h0), .S(RST), .Y(_03591_) );
  \$mux  #( .WIDTH(10) ) _51871_ ( .A(ram_w4_l8192_id6_6_1_addr), .B(_tmp_242), .S(_06238_), .Y(_27521_) );
  \$mux  #( .WIDTH(10) ) _51872_ ( .A(_27521_), .B(10'h000), .S(RST), .Y(_03590_) );
  \$mux  #( .WIDTH(10) ) _51873_ ( .A(ram_w4_l8192_id6_6_0_addr), .B(_stream_conv2d_16_source_34_source_ram_raddr[12:3]), .S(_tmp_681), .Y(_27522_) );
  \$mux  #( .WIDTH(10) ) _51874_ ( .A(_27522_), .B(10'h000), .S(RST), .Y(_03589_) );
  \$mux  #( .WIDTH(1) ) _51875_ ( .A(ram_w4_l8192_id6_5_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27523_) );
  \$mux  #( .WIDTH(1) ) _51876_ ( .A(_27523_), .B(_06079_), .S(_06235_), .Y(_27524_) );
  \$mux  #( .WIDTH(1) ) _51877_ ( .A(_27524_), .B(1'h0), .S(RST), .Y(_03588_) );
  \$mux  #( .WIDTH(4) ) _51878_ ( .A(ram_w4_l8192_id6_5_1_wdata), .B(_dataflow_slice_data_44), .S(_06235_), .Y(_27525_) );
  \$mux  #( .WIDTH(4) ) _51879_ ( .A(_27525_), .B(4'h0), .S(RST), .Y(_03587_) );
  \$mux  #( .WIDTH(10) ) _51880_ ( .A(ram_w4_l8192_id6_5_1_addr), .B(_tmp_211), .S(_06235_), .Y(_27526_) );
  \$mux  #( .WIDTH(10) ) _51881_ ( .A(_27526_), .B(10'h000), .S(RST), .Y(_03586_) );
  \$mux  #( .WIDTH(10) ) _51882_ ( .A(ram_w4_l8192_id6_5_0_addr), .B(_stream_conv2d_16_source_34_source_ram_raddr[12:3]), .S(_tmp_681), .Y(_27527_) );
  \$mux  #( .WIDTH(10) ) _51883_ ( .A(_27527_), .B(10'h000), .S(RST), .Y(_03585_) );
  \$mux  #( .WIDTH(1) ) _51884_ ( .A(ram_w4_l8192_id6_4_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27528_) );
  \$mux  #( .WIDTH(1) ) _51885_ ( .A(_27528_), .B(_06070_), .S(_06232_), .Y(_27529_) );
  \$mux  #( .WIDTH(1) ) _51886_ ( .A(_27529_), .B(1'h0), .S(RST), .Y(_03584_) );
  \$mux  #( .WIDTH(4) ) _51887_ ( .A(ram_w4_l8192_id6_4_1_wdata), .B(_dataflow_slice_data_41), .S(_06232_), .Y(_27530_) );
  \$mux  #( .WIDTH(4) ) _51888_ ( .A(_27530_), .B(4'h0), .S(RST), .Y(_03583_) );
  \$mux  #( .WIDTH(10) ) _51889_ ( .A(ram_w4_l8192_id6_4_1_addr), .B(_tmp_180), .S(_06232_), .Y(_27531_) );
  \$mux  #( .WIDTH(10) ) _51890_ ( .A(_27531_), .B(10'h000), .S(RST), .Y(_03582_) );
  \$mux  #( .WIDTH(10) ) _51891_ ( .A(ram_w4_l8192_id6_4_0_addr), .B(_stream_conv2d_16_source_34_source_ram_raddr[12:3]), .S(_tmp_681), .Y(_27532_) );
  \$mux  #( .WIDTH(10) ) _51892_ ( .A(_27532_), .B(10'h000), .S(RST), .Y(_03581_) );
  \$mux  #( .WIDTH(1) ) _51893_ ( .A(ram_w4_l8192_id6_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27533_) );
  \$mux  #( .WIDTH(1) ) _51894_ ( .A(_27533_), .B(_06061_), .S(_06229_), .Y(_27534_) );
  \$mux  #( .WIDTH(1) ) _51895_ ( .A(_27534_), .B(1'h0), .S(RST), .Y(_03580_) );
  \$mux  #( .WIDTH(4) ) _51896_ ( .A(ram_w4_l8192_id6_3_1_wdata), .B(_dataflow_slice_data_38), .S(_06229_), .Y(_27535_) );
  \$mux  #( .WIDTH(4) ) _51897_ ( .A(_27535_), .B(4'h0), .S(RST), .Y(_03579_) );
  \$mux  #( .WIDTH(10) ) _51898_ ( .A(ram_w4_l8192_id6_3_1_addr), .B(_tmp_149), .S(_06229_), .Y(_27536_) );
  \$mux  #( .WIDTH(10) ) _51899_ ( .A(_27536_), .B(10'h000), .S(RST), .Y(_03578_) );
  \$mux  #( .WIDTH(10) ) _51900_ ( .A(ram_w4_l8192_id6_3_0_addr), .B(_stream_conv2d_16_source_34_source_ram_raddr[12:3]), .S(_tmp_681), .Y(_27537_) );
  \$mux  #( .WIDTH(10) ) _51901_ ( .A(_27537_), .B(10'h000), .S(RST), .Y(_03577_) );
  \$mux  #( .WIDTH(1) ) _51902_ ( .A(ram_w4_l8192_id6_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27538_) );
  \$mux  #( .WIDTH(1) ) _51903_ ( .A(_27538_), .B(_06052_), .S(_06226_), .Y(_27539_) );
  \$mux  #( .WIDTH(1) ) _51904_ ( .A(_27539_), .B(1'h0), .S(RST), .Y(_03576_) );
  \$mux  #( .WIDTH(4) ) _51905_ ( .A(ram_w4_l8192_id6_2_1_wdata), .B(_dataflow_slice_data_35), .S(_06226_), .Y(_27540_) );
  \$mux  #( .WIDTH(4) ) _51906_ ( .A(_27540_), .B(4'h0), .S(RST), .Y(_03575_) );
  \$mux  #( .WIDTH(10) ) _51907_ ( .A(ram_w4_l8192_id6_2_1_addr), .B(_tmp_118), .S(_06226_), .Y(_27541_) );
  \$mux  #( .WIDTH(10) ) _51908_ ( .A(_27541_), .B(10'h000), .S(RST), .Y(_03574_) );
  \$mux  #( .WIDTH(10) ) _51909_ ( .A(ram_w4_l8192_id6_2_0_addr), .B(_stream_conv2d_16_source_34_source_ram_raddr[12:3]), .S(_tmp_681), .Y(_27542_) );
  \$mux  #( .WIDTH(10) ) _51910_ ( .A(_27542_), .B(10'h000), .S(RST), .Y(_03573_) );
  \$mux  #( .WIDTH(1) ) _51911_ ( .A(ram_w4_l8192_id6_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27543_) );
  \$mux  #( .WIDTH(1) ) _51912_ ( .A(_27543_), .B(_06043_), .S(_06223_), .Y(_27544_) );
  \$mux  #( .WIDTH(1) ) _51913_ ( .A(_27544_), .B(1'h0), .S(RST), .Y(_03572_) );
  \$mux  #( .WIDTH(4) ) _51914_ ( .A(ram_w4_l8192_id6_1_1_wdata), .B(_dataflow_slice_data_32), .S(_06223_), .Y(_27545_) );
  \$mux  #( .WIDTH(4) ) _51915_ ( .A(_27545_), .B(4'h0), .S(RST), .Y(_03571_) );
  \$mux  #( .WIDTH(10) ) _51916_ ( .A(ram_w4_l8192_id6_1_1_addr), .B(_tmp_87), .S(_06223_), .Y(_27546_) );
  \$mux  #( .WIDTH(10) ) _51917_ ( .A(_27546_), .B(10'h000), .S(RST), .Y(_03570_) );
  \$mux  #( .WIDTH(10) ) _51918_ ( .A(ram_w4_l8192_id6_1_0_addr), .B(_stream_conv2d_16_source_34_source_ram_raddr[12:3]), .S(_tmp_681), .Y(_27547_) );
  \$mux  #( .WIDTH(10) ) _51919_ ( .A(_27547_), .B(10'h000), .S(RST), .Y(_03569_) );
  \$mux  #( .WIDTH(1) ) _51920_ ( .A(_tmp_681), .B(1'h0), .S(RST), .Y(_01282_) );
  \$mux  #( .WIDTH(1) ) _51921_ ( .A(ram_w4_l8192_id6_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27548_) );
  \$mux  #( .WIDTH(1) ) _51922_ ( .A(_27548_), .B(_06034_), .S(_06220_), .Y(_27549_) );
  \$mux  #( .WIDTH(1) ) _51923_ ( .A(_27549_), .B(1'h0), .S(RST), .Y(_03568_) );
  \$mux  #( .WIDTH(4) ) _51924_ ( .A(ram_w4_l8192_id6_0_1_wdata), .B(_dataflow_slice_data_29), .S(_06220_), .Y(_27550_) );
  \$mux  #( .WIDTH(4) ) _51925_ ( .A(_27550_), .B(4'h0), .S(RST), .Y(_03567_) );
  \$mux  #( .WIDTH(10) ) _51926_ ( .A(ram_w4_l8192_id6_0_1_addr), .B(_tmp_56), .S(_06220_), .Y(_27551_) );
  \$mux  #( .WIDTH(10) ) _51927_ ( .A(_27551_), .B(10'h000), .S(RST), .Y(_03566_) );
  \$mux  #( .WIDTH(10) ) _51928_ ( .A(ram_w4_l8192_id6_0_0_addr), .B(_stream_conv2d_16_source_34_source_ram_raddr[12:3]), .S(_tmp_681), .Y(_27552_) );
  \$mux  #( .WIDTH(10) ) _51929_ ( .A(_27552_), .B(10'h000), .S(RST), .Y(_03565_) );
  \$mux  #( .WIDTH(1) ) _51930_ ( .A(ram_w4_l8192_id5_7_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27553_) );
  \$mux  #( .WIDTH(1) ) _51931_ ( .A(_27553_), .B(_06096_), .S(_06241_), .Y(_27554_) );
  \$mux  #( .WIDTH(1) ) _51932_ ( .A(_27554_), .B(1'h0), .S(RST), .Y(_03564_) );
  \$mux  #( .WIDTH(4) ) _51933_ ( .A(ram_w4_l8192_id5_7_1_wdata), .B(_dataflow_slice_data_50), .S(_06241_), .Y(_27555_) );
  \$mux  #( .WIDTH(4) ) _51934_ ( .A(_27555_), .B(4'h0), .S(RST), .Y(_03563_) );
  \$mux  #( .WIDTH(10) ) _51935_ ( .A(ram_w4_l8192_id5_7_1_addr), .B(_tmp_272), .S(_06241_), .Y(_27556_) );
  \$mux  #( .WIDTH(10) ) _51936_ ( .A(_27556_), .B(10'h000), .S(RST), .Y(_03562_) );
  \$mux  #( .WIDTH(10) ) _51937_ ( .A(ram_w4_l8192_id5_7_0_addr), .B(_stream_conv2d_16_source_33_source_ram_raddr[12:3]), .S(_tmp_667), .Y(_27557_) );
  \$mux  #( .WIDTH(10) ) _51938_ ( .A(_27557_), .B(10'h000), .S(RST), .Y(_03561_) );
  \$mux  #( .WIDTH(1) ) _51939_ ( .A(ram_w4_l8192_id5_6_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27558_) );
  \$mux  #( .WIDTH(1) ) _51940_ ( .A(_27558_), .B(_06087_), .S(_06238_), .Y(_27559_) );
  \$mux  #( .WIDTH(1) ) _51941_ ( .A(_27559_), .B(1'h0), .S(RST), .Y(_03560_) );
  \$mux  #( .WIDTH(4) ) _51942_ ( .A(ram_w4_l8192_id5_6_1_wdata), .B(_dataflow_slice_data_47), .S(_06238_), .Y(_27560_) );
  \$mux  #( .WIDTH(4) ) _51943_ ( .A(_27560_), .B(4'h0), .S(RST), .Y(_03559_) );
  \$mux  #( .WIDTH(10) ) _51944_ ( .A(ram_w4_l8192_id5_6_1_addr), .B(_tmp_241), .S(_06238_), .Y(_27561_) );
  \$mux  #( .WIDTH(10) ) _51945_ ( .A(_27561_), .B(10'h000), .S(RST), .Y(_03558_) );
  \$mux  #( .WIDTH(10) ) _51946_ ( .A(ram_w4_l8192_id5_6_0_addr), .B(_stream_conv2d_16_source_33_source_ram_raddr[12:3]), .S(_tmp_667), .Y(_27562_) );
  \$mux  #( .WIDTH(10) ) _51947_ ( .A(_27562_), .B(10'h000), .S(RST), .Y(_03557_) );
  \$mux  #( .WIDTH(1) ) _51948_ ( .A(ram_w4_l8192_id5_5_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27563_) );
  \$mux  #( .WIDTH(1) ) _51949_ ( .A(_27563_), .B(_06078_), .S(_06235_), .Y(_27564_) );
  \$mux  #( .WIDTH(1) ) _51950_ ( .A(_27564_), .B(1'h0), .S(RST), .Y(_03556_) );
  \$mux  #( .WIDTH(4) ) _51951_ ( .A(ram_w4_l8192_id5_5_1_wdata), .B(_dataflow_slice_data_44), .S(_06235_), .Y(_27565_) );
  \$mux  #( .WIDTH(4) ) _51952_ ( .A(_27565_), .B(4'h0), .S(RST), .Y(_03555_) );
  \$mux  #( .WIDTH(10) ) _51953_ ( .A(ram_w4_l8192_id5_5_1_addr), .B(_tmp_210), .S(_06235_), .Y(_27566_) );
  \$mux  #( .WIDTH(10) ) _51954_ ( .A(_27566_), .B(10'h000), .S(RST), .Y(_03554_) );
  \$mux  #( .WIDTH(10) ) _51955_ ( .A(ram_w4_l8192_id5_5_0_addr), .B(_stream_conv2d_16_source_33_source_ram_raddr[12:3]), .S(_tmp_667), .Y(_27567_) );
  \$mux  #( .WIDTH(10) ) _51956_ ( .A(_27567_), .B(10'h000), .S(RST), .Y(_03553_) );
  \$mux  #( .WIDTH(1) ) _51957_ ( .A(ram_w4_l8192_id5_4_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27568_) );
  \$mux  #( .WIDTH(1) ) _51958_ ( .A(_27568_), .B(_06069_), .S(_06232_), .Y(_27569_) );
  \$mux  #( .WIDTH(1) ) _51959_ ( .A(_27569_), .B(1'h0), .S(RST), .Y(_03552_) );
  \$mux  #( .WIDTH(4) ) _51960_ ( .A(ram_w4_l8192_id5_4_1_wdata), .B(_dataflow_slice_data_41), .S(_06232_), .Y(_27570_) );
  \$mux  #( .WIDTH(4) ) _51961_ ( .A(_27570_), .B(4'h0), .S(RST), .Y(_03551_) );
  \$mux  #( .WIDTH(10) ) _51962_ ( .A(ram_w4_l8192_id5_4_1_addr), .B(_tmp_179), .S(_06232_), .Y(_27571_) );
  \$mux  #( .WIDTH(10) ) _51963_ ( .A(_27571_), .B(10'h000), .S(RST), .Y(_03550_) );
  \$mux  #( .WIDTH(10) ) _51964_ ( .A(ram_w4_l8192_id5_4_0_addr), .B(_stream_conv2d_16_source_33_source_ram_raddr[12:3]), .S(_tmp_667), .Y(_27572_) );
  \$mux  #( .WIDTH(10) ) _51965_ ( .A(_27572_), .B(10'h000), .S(RST), .Y(_03549_) );
  \$mux  #( .WIDTH(1) ) _51966_ ( .A(ram_w4_l8192_id5_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27573_) );
  \$mux  #( .WIDTH(1) ) _51967_ ( .A(_27573_), .B(_06060_), .S(_06229_), .Y(_27574_) );
  \$mux  #( .WIDTH(1) ) _51968_ ( .A(_27574_), .B(1'h0), .S(RST), .Y(_03548_) );
  \$mux  #( .WIDTH(4) ) _51969_ ( .A(ram_w4_l8192_id5_3_1_wdata), .B(_dataflow_slice_data_38), .S(_06229_), .Y(_27575_) );
  \$mux  #( .WIDTH(4) ) _51970_ ( .A(_27575_), .B(4'h0), .S(RST), .Y(_03547_) );
  \$mux  #( .WIDTH(10) ) _51971_ ( .A(ram_w4_l8192_id5_3_1_addr), .B(_tmp_148), .S(_06229_), .Y(_27576_) );
  \$mux  #( .WIDTH(10) ) _51972_ ( .A(_27576_), .B(10'h000), .S(RST), .Y(_03546_) );
  \$mux  #( .WIDTH(10) ) _51973_ ( .A(ram_w4_l8192_id5_3_0_addr), .B(_stream_conv2d_16_source_33_source_ram_raddr[12:3]), .S(_tmp_667), .Y(_27577_) );
  \$mux  #( .WIDTH(10) ) _51974_ ( .A(_27577_), .B(10'h000), .S(RST), .Y(_03545_) );
  \$mux  #( .WIDTH(1) ) _51975_ ( .A(ram_w4_l8192_id5_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27578_) );
  \$mux  #( .WIDTH(1) ) _51976_ ( .A(_27578_), .B(_06051_), .S(_06226_), .Y(_27579_) );
  \$mux  #( .WIDTH(1) ) _51977_ ( .A(_27579_), .B(1'h0), .S(RST), .Y(_03544_) );
  \$mux  #( .WIDTH(4) ) _51978_ ( .A(ram_w4_l8192_id5_2_1_wdata), .B(_dataflow_slice_data_35), .S(_06226_), .Y(_27580_) );
  \$mux  #( .WIDTH(4) ) _51979_ ( .A(_27580_), .B(4'h0), .S(RST), .Y(_03543_) );
  \$mux  #( .WIDTH(10) ) _51980_ ( .A(ram_w4_l8192_id5_2_1_addr), .B(_tmp_117), .S(_06226_), .Y(_27581_) );
  \$mux  #( .WIDTH(10) ) _51981_ ( .A(_27581_), .B(10'h000), .S(RST), .Y(_03542_) );
  \$mux  #( .WIDTH(10) ) _51982_ ( .A(ram_w4_l8192_id5_2_0_addr), .B(_stream_conv2d_16_source_33_source_ram_raddr[12:3]), .S(_tmp_667), .Y(_27582_) );
  \$mux  #( .WIDTH(10) ) _51983_ ( .A(_27582_), .B(10'h000), .S(RST), .Y(_03541_) );
  \$mux  #( .WIDTH(1) ) _51984_ ( .A(ram_w4_l8192_id5_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27583_) );
  \$mux  #( .WIDTH(1) ) _51985_ ( .A(_27583_), .B(_06042_), .S(_06223_), .Y(_27584_) );
  \$mux  #( .WIDTH(1) ) _51986_ ( .A(_27584_), .B(1'h0), .S(RST), .Y(_03540_) );
  \$mux  #( .WIDTH(4) ) _51987_ ( .A(ram_w4_l8192_id5_1_1_wdata), .B(_dataflow_slice_data_32), .S(_06223_), .Y(_27585_) );
  \$mux  #( .WIDTH(4) ) _51988_ ( .A(_27585_), .B(4'h0), .S(RST), .Y(_03539_) );
  \$mux  #( .WIDTH(10) ) _51989_ ( .A(ram_w4_l8192_id5_1_1_addr), .B(_tmp_86), .S(_06223_), .Y(_27586_) );
  \$mux  #( .WIDTH(10) ) _51990_ ( .A(_27586_), .B(10'h000), .S(RST), .Y(_03538_) );
  \$mux  #( .WIDTH(10) ) _51991_ ( .A(ram_w4_l8192_id5_1_0_addr), .B(_stream_conv2d_16_source_33_source_ram_raddr[12:3]), .S(_tmp_667), .Y(_27587_) );
  \$mux  #( .WIDTH(10) ) _51992_ ( .A(_27587_), .B(10'h000), .S(RST), .Y(_03537_) );
  \$mux  #( .WIDTH(1) ) _51993_ ( .A(_tmp_667), .B(1'h0), .S(RST), .Y(_01279_) );
  \$mux  #( .WIDTH(1) ) _51994_ ( .A(ram_w4_l8192_id5_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27588_) );
  \$mux  #( .WIDTH(1) ) _51995_ ( .A(_27588_), .B(_06033_), .S(_06220_), .Y(_27589_) );
  \$mux  #( .WIDTH(1) ) _51996_ ( .A(_27589_), .B(1'h0), .S(RST), .Y(_03536_) );
  \$mux  #( .WIDTH(4) ) _51997_ ( .A(ram_w4_l8192_id5_0_1_wdata), .B(_dataflow_slice_data_29), .S(_06220_), .Y(_27590_) );
  \$mux  #( .WIDTH(4) ) _51998_ ( .A(_27590_), .B(4'h0), .S(RST), .Y(_03535_) );
  \$mux  #( .WIDTH(10) ) _51999_ ( .A(ram_w4_l8192_id5_0_1_addr), .B(_tmp_55), .S(_06220_), .Y(_27591_) );
  \$mux  #( .WIDTH(10) ) _52000_ ( .A(_27591_), .B(10'h000), .S(RST), .Y(_03534_) );
  \$mux  #( .WIDTH(10) ) _52001_ ( .A(ram_w4_l8192_id5_0_0_addr), .B(_stream_conv2d_16_source_33_source_ram_raddr[12:3]), .S(_tmp_667), .Y(_27592_) );
  \$mux  #( .WIDTH(10) ) _52002_ ( .A(_27592_), .B(10'h000), .S(RST), .Y(_03533_) );
  \$mux  #( .WIDTH(1) ) _52003_ ( .A(ram_w4_l8192_id4_7_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27593_) );
  \$mux  #( .WIDTH(1) ) _52004_ ( .A(_27593_), .B(_06095_), .S(_06241_), .Y(_27594_) );
  \$mux  #( .WIDTH(1) ) _52005_ ( .A(_27594_), .B(1'h0), .S(RST), .Y(_03532_) );
  \$mux  #( .WIDTH(4) ) _52006_ ( .A(ram_w4_l8192_id4_7_1_wdata), .B(_dataflow_slice_data_50), .S(_06241_), .Y(_27595_) );
  \$mux  #( .WIDTH(4) ) _52007_ ( .A(_27595_), .B(4'h0), .S(RST), .Y(_03531_) );
  \$mux  #( .WIDTH(10) ) _52008_ ( .A(ram_w4_l8192_id4_7_1_addr), .B(_tmp_271), .S(_06241_), .Y(_27596_) );
  \$mux  #( .WIDTH(10) ) _52009_ ( .A(_27596_), .B(10'h000), .S(RST), .Y(_03530_) );
  \$mux  #( .WIDTH(10) ) _52010_ ( .A(ram_w4_l8192_id4_7_0_addr), .B(_stream_conv2d_16_source_32_source_ram_raddr[12:3]), .S(_tmp_653), .Y(_27597_) );
  \$mux  #( .WIDTH(10) ) _52011_ ( .A(_27597_), .B(10'h000), .S(RST), .Y(_03529_) );
  \$mux  #( .WIDTH(1) ) _52012_ ( .A(ram_w4_l8192_id4_6_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27598_) );
  \$mux  #( .WIDTH(1) ) _52013_ ( .A(_27598_), .B(_06086_), .S(_06238_), .Y(_27599_) );
  \$mux  #( .WIDTH(1) ) _52014_ ( .A(_27599_), .B(1'h0), .S(RST), .Y(_03528_) );
  \$mux  #( .WIDTH(4) ) _52015_ ( .A(ram_w4_l8192_id4_6_1_wdata), .B(_dataflow_slice_data_47), .S(_06238_), .Y(_27600_) );
  \$mux  #( .WIDTH(4) ) _52016_ ( .A(_27600_), .B(4'h0), .S(RST), .Y(_03527_) );
  \$mux  #( .WIDTH(10) ) _52017_ ( .A(ram_w4_l8192_id4_6_1_addr), .B(_tmp_240), .S(_06238_), .Y(_27601_) );
  \$mux  #( .WIDTH(10) ) _52018_ ( .A(_27601_), .B(10'h000), .S(RST), .Y(_03526_) );
  \$mux  #( .WIDTH(10) ) _52019_ ( .A(ram_w4_l8192_id4_6_0_addr), .B(_stream_conv2d_16_source_32_source_ram_raddr[12:3]), .S(_tmp_653), .Y(_27602_) );
  \$mux  #( .WIDTH(10) ) _52020_ ( .A(_27602_), .B(10'h000), .S(RST), .Y(_03525_) );
  \$mux  #( .WIDTH(1) ) _52021_ ( .A(ram_w4_l8192_id4_5_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27603_) );
  \$mux  #( .WIDTH(1) ) _52022_ ( .A(_27603_), .B(_06077_), .S(_06235_), .Y(_27604_) );
  \$mux  #( .WIDTH(1) ) _52023_ ( .A(_27604_), .B(1'h0), .S(RST), .Y(_03524_) );
  \$mux  #( .WIDTH(4) ) _52024_ ( .A(ram_w4_l8192_id4_5_1_wdata), .B(_dataflow_slice_data_44), .S(_06235_), .Y(_27605_) );
  \$mux  #( .WIDTH(4) ) _52025_ ( .A(_27605_), .B(4'h0), .S(RST), .Y(_03523_) );
  \$mux  #( .WIDTH(10) ) _52026_ ( .A(ram_w4_l8192_id4_5_1_addr), .B(_tmp_209), .S(_06235_), .Y(_27606_) );
  \$mux  #( .WIDTH(10) ) _52027_ ( .A(_27606_), .B(10'h000), .S(RST), .Y(_03522_) );
  \$mux  #( .WIDTH(10) ) _52028_ ( .A(ram_w4_l8192_id4_5_0_addr), .B(_stream_conv2d_16_source_32_source_ram_raddr[12:3]), .S(_tmp_653), .Y(_27607_) );
  \$mux  #( .WIDTH(10) ) _52029_ ( .A(_27607_), .B(10'h000), .S(RST), .Y(_03521_) );
  \$mux  #( .WIDTH(1) ) _52030_ ( .A(ram_w4_l8192_id4_4_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27608_) );
  \$mux  #( .WIDTH(1) ) _52031_ ( .A(_27608_), .B(_06068_), .S(_06232_), .Y(_27609_) );
  \$mux  #( .WIDTH(1) ) _52032_ ( .A(_27609_), .B(1'h0), .S(RST), .Y(_03520_) );
  \$mux  #( .WIDTH(4) ) _52033_ ( .A(ram_w4_l8192_id4_4_1_wdata), .B(_dataflow_slice_data_41), .S(_06232_), .Y(_27610_) );
  \$mux  #( .WIDTH(4) ) _52034_ ( .A(_27610_), .B(4'h0), .S(RST), .Y(_03519_) );
  \$mux  #( .WIDTH(10) ) _52035_ ( .A(ram_w4_l8192_id4_4_1_addr), .B(_tmp_178), .S(_06232_), .Y(_27611_) );
  \$mux  #( .WIDTH(10) ) _52036_ ( .A(_27611_), .B(10'h000), .S(RST), .Y(_03518_) );
  \$mux  #( .WIDTH(10) ) _52037_ ( .A(ram_w4_l8192_id4_4_0_addr), .B(_stream_conv2d_16_source_32_source_ram_raddr[12:3]), .S(_tmp_653), .Y(_27612_) );
  \$mux  #( .WIDTH(10) ) _52038_ ( .A(_27612_), .B(10'h000), .S(RST), .Y(_03517_) );
  \$mux  #( .WIDTH(1) ) _52039_ ( .A(ram_w4_l8192_id4_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27613_) );
  \$mux  #( .WIDTH(1) ) _52040_ ( .A(_27613_), .B(_06059_), .S(_06229_), .Y(_27614_) );
  \$mux  #( .WIDTH(1) ) _52041_ ( .A(_27614_), .B(1'h0), .S(RST), .Y(_03516_) );
  \$mux  #( .WIDTH(4) ) _52042_ ( .A(ram_w4_l8192_id4_3_1_wdata), .B(_dataflow_slice_data_38), .S(_06229_), .Y(_27615_) );
  \$mux  #( .WIDTH(4) ) _52043_ ( .A(_27615_), .B(4'h0), .S(RST), .Y(_03515_) );
  \$mux  #( .WIDTH(10) ) _52044_ ( .A(ram_w4_l8192_id4_3_1_addr), .B(_tmp_147), .S(_06229_), .Y(_27616_) );
  \$mux  #( .WIDTH(10) ) _52045_ ( .A(_27616_), .B(10'h000), .S(RST), .Y(_03514_) );
  \$mux  #( .WIDTH(10) ) _52046_ ( .A(ram_w4_l8192_id4_3_0_addr), .B(_stream_conv2d_16_source_32_source_ram_raddr[12:3]), .S(_tmp_653), .Y(_27617_) );
  \$mux  #( .WIDTH(10) ) _52047_ ( .A(_27617_), .B(10'h000), .S(RST), .Y(_03513_) );
  \$mux  #( .WIDTH(1) ) _52048_ ( .A(ram_w4_l8192_id4_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27618_) );
  \$mux  #( .WIDTH(1) ) _52049_ ( .A(_27618_), .B(_06050_), .S(_06226_), .Y(_27619_) );
  \$mux  #( .WIDTH(1) ) _52050_ ( .A(_27619_), .B(1'h0), .S(RST), .Y(_03512_) );
  \$mux  #( .WIDTH(4) ) _52051_ ( .A(ram_w4_l8192_id4_2_1_wdata), .B(_dataflow_slice_data_35), .S(_06226_), .Y(_27620_) );
  \$mux  #( .WIDTH(4) ) _52052_ ( .A(_27620_), .B(4'h0), .S(RST), .Y(_03511_) );
  \$mux  #( .WIDTH(10) ) _52053_ ( .A(ram_w4_l8192_id4_2_1_addr), .B(_tmp_116), .S(_06226_), .Y(_27621_) );
  \$mux  #( .WIDTH(10) ) _52054_ ( .A(_27621_), .B(10'h000), .S(RST), .Y(_03510_) );
  \$mux  #( .WIDTH(10) ) _52055_ ( .A(ram_w4_l8192_id4_2_0_addr), .B(_stream_conv2d_16_source_32_source_ram_raddr[12:3]), .S(_tmp_653), .Y(_27622_) );
  \$mux  #( .WIDTH(10) ) _52056_ ( .A(_27622_), .B(10'h000), .S(RST), .Y(_03509_) );
  \$mux  #( .WIDTH(1) ) _52057_ ( .A(ram_w4_l8192_id4_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27623_) );
  \$mux  #( .WIDTH(1) ) _52058_ ( .A(_27623_), .B(_06041_), .S(_06223_), .Y(_27624_) );
  \$mux  #( .WIDTH(1) ) _52059_ ( .A(_27624_), .B(1'h0), .S(RST), .Y(_03508_) );
  \$mux  #( .WIDTH(4) ) _52060_ ( .A(ram_w4_l8192_id4_1_1_wdata), .B(_dataflow_slice_data_32), .S(_06223_), .Y(_27625_) );
  \$mux  #( .WIDTH(4) ) _52061_ ( .A(_27625_), .B(4'h0), .S(RST), .Y(_03507_) );
  \$mux  #( .WIDTH(10) ) _52062_ ( .A(ram_w4_l8192_id4_1_1_addr), .B(_tmp_85), .S(_06223_), .Y(_27626_) );
  \$mux  #( .WIDTH(10) ) _52063_ ( .A(_27626_), .B(10'h000), .S(RST), .Y(_03506_) );
  \$mux  #( .WIDTH(10) ) _52064_ ( .A(ram_w4_l8192_id4_1_0_addr), .B(_stream_conv2d_16_source_32_source_ram_raddr[12:3]), .S(_tmp_653), .Y(_27627_) );
  \$mux  #( .WIDTH(10) ) _52065_ ( .A(_27627_), .B(10'h000), .S(RST), .Y(_03505_) );
  \$mux  #( .WIDTH(1) ) _52066_ ( .A(_tmp_653), .B(1'h0), .S(RST), .Y(_01276_) );
  \$mux  #( .WIDTH(1) ) _52067_ ( .A(ram_w4_l8192_id4_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27628_) );
  \$mux  #( .WIDTH(1) ) _52068_ ( .A(_27628_), .B(_06032_), .S(_06220_), .Y(_27629_) );
  \$mux  #( .WIDTH(1) ) _52069_ ( .A(_27629_), .B(1'h0), .S(RST), .Y(_03504_) );
  \$mux  #( .WIDTH(4) ) _52070_ ( .A(ram_w4_l8192_id4_0_1_wdata), .B(_dataflow_slice_data_29), .S(_06220_), .Y(_27630_) );
  \$mux  #( .WIDTH(4) ) _52071_ ( .A(_27630_), .B(4'h0), .S(RST), .Y(_03503_) );
  \$mux  #( .WIDTH(10) ) _52072_ ( .A(ram_w4_l8192_id4_0_1_addr), .B(_tmp_54), .S(_06220_), .Y(_27631_) );
  \$mux  #( .WIDTH(10) ) _52073_ ( .A(_27631_), .B(10'h000), .S(RST), .Y(_03502_) );
  \$mux  #( .WIDTH(10) ) _52074_ ( .A(ram_w4_l8192_id4_0_0_addr), .B(_stream_conv2d_16_source_32_source_ram_raddr[12:3]), .S(_tmp_653), .Y(_27632_) );
  \$mux  #( .WIDTH(10) ) _52075_ ( .A(_27632_), .B(10'h000), .S(RST), .Y(_03501_) );
  \$mux  #( .WIDTH(1) ) _52076_ ( .A(ram_w4_l8192_id3_7_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27633_) );
  \$mux  #( .WIDTH(1) ) _52077_ ( .A(_27633_), .B(_06094_), .S(_06241_), .Y(_27634_) );
  \$mux  #( .WIDTH(1) ) _52078_ ( .A(_27634_), .B(1'h0), .S(RST), .Y(_03500_) );
  \$mux  #( .WIDTH(4) ) _52079_ ( .A(ram_w4_l8192_id3_7_1_wdata), .B(_dataflow_slice_data_50), .S(_06241_), .Y(_27635_) );
  \$mux  #( .WIDTH(4) ) _52080_ ( .A(_27635_), .B(4'h0), .S(RST), .Y(_03499_) );
  \$mux  #( .WIDTH(10) ) _52081_ ( .A(ram_w4_l8192_id3_7_1_addr), .B(_tmp_270), .S(_06241_), .Y(_27636_) );
  \$mux  #( .WIDTH(10) ) _52082_ ( .A(_27636_), .B(10'h000), .S(RST), .Y(_03498_) );
  \$mux  #( .WIDTH(10) ) _52083_ ( .A(ram_w4_l8192_id3_7_0_addr), .B(_stream_conv2d_16_source_31_source_ram_raddr[12:3]), .S(_tmp_639), .Y(_27637_) );
  \$mux  #( .WIDTH(10) ) _52084_ ( .A(_27637_), .B(10'h000), .S(RST), .Y(_03497_) );
  \$mux  #( .WIDTH(1) ) _52085_ ( .A(ram_w4_l8192_id3_6_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27638_) );
  \$mux  #( .WIDTH(1) ) _52086_ ( .A(_27638_), .B(_06085_), .S(_06238_), .Y(_27639_) );
  \$mux  #( .WIDTH(1) ) _52087_ ( .A(_27639_), .B(1'h0), .S(RST), .Y(_03496_) );
  \$mux  #( .WIDTH(4) ) _52088_ ( .A(ram_w4_l8192_id3_6_1_wdata), .B(_dataflow_slice_data_47), .S(_06238_), .Y(_27640_) );
  \$mux  #( .WIDTH(4) ) _52089_ ( .A(_27640_), .B(4'h0), .S(RST), .Y(_03495_) );
  \$mux  #( .WIDTH(10) ) _52090_ ( .A(ram_w4_l8192_id3_6_1_addr), .B(_tmp_239), .S(_06238_), .Y(_27641_) );
  \$mux  #( .WIDTH(10) ) _52091_ ( .A(_27641_), .B(10'h000), .S(RST), .Y(_03494_) );
  \$mux  #( .WIDTH(10) ) _52092_ ( .A(ram_w4_l8192_id3_6_0_addr), .B(_stream_conv2d_16_source_31_source_ram_raddr[12:3]), .S(_tmp_639), .Y(_27642_) );
  \$mux  #( .WIDTH(10) ) _52093_ ( .A(_27642_), .B(10'h000), .S(RST), .Y(_03493_) );
  \$mux  #( .WIDTH(1) ) _52094_ ( .A(1'h1), .B(1'h0), .S(RST), .Y(_01824_) );
  \$mux  #( .WIDTH(1) ) _52095_ ( .A(ram_w4_l8192_id3_5_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27643_) );
  \$mux  #( .WIDTH(1) ) _52096_ ( .A(_27643_), .B(_06076_), .S(_06235_), .Y(_27644_) );
  \$mux  #( .WIDTH(1) ) _52097_ ( .A(_27644_), .B(1'h0), .S(RST), .Y(_03492_) );
  \$mux  #( .WIDTH(4) ) _52098_ ( .A(ram_w4_l8192_id3_5_1_wdata), .B(_dataflow_slice_data_44), .S(_06235_), .Y(_27645_) );
  \$mux  #( .WIDTH(4) ) _52099_ ( .A(_27645_), .B(4'h0), .S(RST), .Y(_03491_) );
  \$mux  #( .WIDTH(10) ) _52100_ ( .A(ram_w4_l8192_id3_5_1_addr), .B(_tmp_208), .S(_06235_), .Y(_27646_) );
  \$mux  #( .WIDTH(10) ) _52101_ ( .A(_27646_), .B(10'h000), .S(RST), .Y(_03490_) );
  \$mux  #( .WIDTH(10) ) _52102_ ( .A(ram_w4_l8192_id3_5_0_addr), .B(_stream_conv2d_16_source_31_source_ram_raddr[12:3]), .S(_tmp_639), .Y(_27647_) );
  \$mux  #( .WIDTH(10) ) _52103_ ( .A(_27647_), .B(10'h000), .S(RST), .Y(_03489_) );
  \$mux  #( .WIDTH(1) ) _52104_ ( .A(_tmp_639), .B(1'h0), .S(RST), .Y(_01273_) );
  \$mux  #( .WIDTH(1) ) _52105_ ( .A(ram_w4_l8192_id3_4_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27648_) );
  \$mux  #( .WIDTH(1) ) _52106_ ( .A(_27648_), .B(_06067_), .S(_06232_), .Y(_27649_) );
  \$mux  #( .WIDTH(1) ) _52107_ ( .A(_27649_), .B(1'h0), .S(RST), .Y(_03488_) );
  \$mux  #( .WIDTH(4) ) _52108_ ( .A(ram_w4_l8192_id3_4_1_wdata), .B(_dataflow_slice_data_41), .S(_06232_), .Y(_27650_) );
  \$mux  #( .WIDTH(4) ) _52109_ ( .A(_27650_), .B(4'h0), .S(RST), .Y(_03487_) );
  \$mux  #( .WIDTH(10) ) _52110_ ( .A(ram_w4_l8192_id3_4_1_addr), .B(_tmp_177), .S(_06232_), .Y(_27651_) );
  \$mux  #( .WIDTH(10) ) _52111_ ( .A(_27651_), .B(10'h000), .S(RST), .Y(_03486_) );
  \$mux  #( .WIDTH(10) ) _52112_ ( .A(ram_w4_l8192_id3_4_0_addr), .B(_stream_conv2d_16_source_31_source_ram_raddr[12:3]), .S(_tmp_639), .Y(_27652_) );
  \$mux  #( .WIDTH(10) ) _52113_ ( .A(_27652_), .B(10'h000), .S(RST), .Y(_03485_) );
  \$mux  #( .WIDTH(1) ) _52114_ ( .A(ram_w4_l8192_id3_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27653_) );
  \$mux  #( .WIDTH(1) ) _52115_ ( .A(_27653_), .B(_06058_), .S(_06229_), .Y(_27654_) );
  \$mux  #( .WIDTH(1) ) _52116_ ( .A(_27654_), .B(1'h0), .S(RST), .Y(_03484_) );
  \$mux  #( .WIDTH(4) ) _52117_ ( .A(ram_w4_l8192_id3_3_1_wdata), .B(_dataflow_slice_data_38), .S(_06229_), .Y(_27655_) );
  \$mux  #( .WIDTH(4) ) _52118_ ( .A(_27655_), .B(4'h0), .S(RST), .Y(_03483_) );
  \$mux  #( .WIDTH(10) ) _52119_ ( .A(ram_w4_l8192_id3_3_1_addr), .B(_tmp_146), .S(_06229_), .Y(_27656_) );
  \$mux  #( .WIDTH(10) ) _52120_ ( .A(_27656_), .B(10'h000), .S(RST), .Y(_03482_) );
  \$mux  #( .WIDTH(10) ) _52121_ ( .A(ram_w4_l8192_id3_3_0_addr), .B(_stream_conv2d_16_source_31_source_ram_raddr[12:3]), .S(_tmp_639), .Y(_27657_) );
  \$mux  #( .WIDTH(10) ) _52122_ ( .A(_27657_), .B(10'h000), .S(RST), .Y(_03481_) );
  \$mux  #( .WIDTH(1) ) _52123_ ( .A(ram_w4_l8192_id3_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27658_) );
  \$mux  #( .WIDTH(1) ) _52124_ ( .A(_27658_), .B(_06049_), .S(_06226_), .Y(_27659_) );
  \$mux  #( .WIDTH(1) ) _52125_ ( .A(_27659_), .B(1'h0), .S(RST), .Y(_03480_) );
  \$mux  #( .WIDTH(4) ) _52126_ ( .A(ram_w4_l8192_id3_2_1_wdata), .B(_dataflow_slice_data_35), .S(_06226_), .Y(_27660_) );
  \$mux  #( .WIDTH(4) ) _52127_ ( .A(_27660_), .B(4'h0), .S(RST), .Y(_03479_) );
  \$mux  #( .WIDTH(10) ) _52128_ ( .A(ram_w4_l8192_id3_2_1_addr), .B(_tmp_115), .S(_06226_), .Y(_27661_) );
  \$mux  #( .WIDTH(10) ) _52129_ ( .A(_27661_), .B(10'h000), .S(RST), .Y(_03478_) );
  \$mux  #( .WIDTH(10) ) _52130_ ( .A(ram_w4_l8192_id3_2_0_addr), .B(_stream_conv2d_16_source_31_source_ram_raddr[12:3]), .S(_tmp_639), .Y(_27662_) );
  \$mux  #( .WIDTH(10) ) _52131_ ( .A(_27662_), .B(10'h000), .S(RST), .Y(_03477_) );
  \$mux  #( .WIDTH(1) ) _52132_ ( .A(ram_w4_l8192_id3_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27663_) );
  \$mux  #( .WIDTH(1) ) _52133_ ( .A(_27663_), .B(_06040_), .S(_06223_), .Y(_27664_) );
  \$mux  #( .WIDTH(1) ) _52134_ ( .A(_27664_), .B(1'h0), .S(RST), .Y(_03476_) );
  \$mux  #( .WIDTH(4) ) _52135_ ( .A(ram_w4_l8192_id3_1_1_wdata), .B(_dataflow_slice_data_32), .S(_06223_), .Y(_27665_) );
  \$mux  #( .WIDTH(4) ) _52136_ ( .A(_27665_), .B(4'h0), .S(RST), .Y(_03475_) );
  \$mux  #( .WIDTH(10) ) _52137_ ( .A(ram_w4_l8192_id3_1_1_addr), .B(_tmp_84), .S(_06223_), .Y(_27666_) );
  \$mux  #( .WIDTH(10) ) _52138_ ( .A(_27666_), .B(10'h000), .S(RST), .Y(_03474_) );
  \$mux  #( .WIDTH(10) ) _52139_ ( .A(ram_w4_l8192_id3_1_0_addr), .B(_stream_conv2d_16_source_31_source_ram_raddr[12:3]), .S(_tmp_639), .Y(_27667_) );
  \$mux  #( .WIDTH(10) ) _52140_ ( .A(_27667_), .B(10'h000), .S(RST), .Y(_03473_) );
  \$mux  #( .WIDTH(1) ) _52141_ ( .A(ram_w4_l8192_id3_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27668_) );
  \$mux  #( .WIDTH(1) ) _52142_ ( .A(_27668_), .B(_06031_), .S(_06220_), .Y(_27669_) );
  \$mux  #( .WIDTH(1) ) _52143_ ( .A(_27669_), .B(1'h0), .S(RST), .Y(_03472_) );
  \$mux  #( .WIDTH(4) ) _52144_ ( .A(ram_w4_l8192_id3_0_1_wdata), .B(_dataflow_slice_data_29), .S(_06220_), .Y(_27670_) );
  \$mux  #( .WIDTH(4) ) _52145_ ( .A(_27670_), .B(4'h0), .S(RST), .Y(_03471_) );
  \$mux  #( .WIDTH(10) ) _52146_ ( .A(ram_w4_l8192_id3_0_1_addr), .B(_tmp_53), .S(_06220_), .Y(_27671_) );
  \$mux  #( .WIDTH(10) ) _52147_ ( .A(_27671_), .B(10'h000), .S(RST), .Y(_03470_) );
  \$mux  #( .WIDTH(10) ) _52148_ ( .A(ram_w4_l8192_id3_0_0_addr), .B(_stream_conv2d_16_source_31_source_ram_raddr[12:3]), .S(_tmp_639), .Y(_27672_) );
  \$mux  #( .WIDTH(10) ) _52149_ ( .A(_27672_), .B(10'h000), .S(RST), .Y(_03469_) );
  \$mux  #( .WIDTH(1) ) _52150_ ( .A(ram_w4_l8192_id2_7_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27673_) );
  \$mux  #( .WIDTH(1) ) _52151_ ( .A(_27673_), .B(_06093_), .S(_06241_), .Y(_27674_) );
  \$mux  #( .WIDTH(1) ) _52152_ ( .A(_27674_), .B(1'h0), .S(RST), .Y(_03468_) );
  \$mux  #( .WIDTH(4) ) _52153_ ( .A(ram_w4_l8192_id2_7_1_wdata), .B(_dataflow_slice_data_50), .S(_06241_), .Y(_27675_) );
  \$mux  #( .WIDTH(4) ) _52154_ ( .A(_27675_), .B(4'h0), .S(RST), .Y(_03467_) );
  \$mux  #( .WIDTH(10) ) _52155_ ( .A(ram_w4_l8192_id2_7_1_addr), .B(_tmp_269), .S(_06241_), .Y(_27676_) );
  \$mux  #( .WIDTH(10) ) _52156_ ( .A(_27676_), .B(10'h000), .S(RST), .Y(_03466_) );
  \$mux  #( .WIDTH(10) ) _52157_ ( .A(ram_w4_l8192_id2_7_0_addr), .B(_stream_conv2d_16_source_30_source_ram_raddr[12:3]), .S(_tmp_625), .Y(_27677_) );
  \$mux  #( .WIDTH(10) ) _52158_ ( .A(_27677_), .B(10'h000), .S(RST), .Y(_03465_) );
  \$mux  #( .WIDTH(1) ) _52159_ ( .A(ram_w4_l8192_id2_6_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27678_) );
  \$mux  #( .WIDTH(1) ) _52160_ ( .A(_27678_), .B(_06084_), .S(_06238_), .Y(_27679_) );
  \$mux  #( .WIDTH(1) ) _52161_ ( .A(_27679_), .B(1'h0), .S(RST), .Y(_03464_) );
  \$mux  #( .WIDTH(4) ) _52162_ ( .A(ram_w4_l8192_id2_6_1_wdata), .B(_dataflow_slice_data_47), .S(_06238_), .Y(_27680_) );
  \$mux  #( .WIDTH(4) ) _52163_ ( .A(_27680_), .B(4'h0), .S(RST), .Y(_03463_) );
  \$mux  #( .WIDTH(10) ) _52164_ ( .A(ram_w4_l8192_id2_6_1_addr), .B(_tmp_238), .S(_06238_), .Y(_27681_) );
  \$mux  #( .WIDTH(10) ) _52165_ ( .A(_27681_), .B(10'h000), .S(RST), .Y(_03462_) );
  \$mux  #( .WIDTH(10) ) _52166_ ( .A(ram_w4_l8192_id2_6_0_addr), .B(_stream_conv2d_16_source_30_source_ram_raddr[12:3]), .S(_tmp_625), .Y(_27682_) );
  \$mux  #( .WIDTH(10) ) _52167_ ( .A(_27682_), .B(10'h000), .S(RST), .Y(_03461_) );
  \$mux  #( .WIDTH(1) ) _52168_ ( .A(ram_w4_l8192_id2_5_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27683_) );
  \$mux  #( .WIDTH(1) ) _52169_ ( .A(_27683_), .B(_06075_), .S(_06235_), .Y(_27684_) );
  \$mux  #( .WIDTH(1) ) _52170_ ( .A(_27684_), .B(1'h0), .S(RST), .Y(_03460_) );
  \$mux  #( .WIDTH(4) ) _52171_ ( .A(ram_w4_l8192_id2_5_1_wdata), .B(_dataflow_slice_data_44), .S(_06235_), .Y(_27685_) );
  \$mux  #( .WIDTH(4) ) _52172_ ( .A(_27685_), .B(4'h0), .S(RST), .Y(_03459_) );
  \$mux  #( .WIDTH(10) ) _52173_ ( .A(ram_w4_l8192_id2_5_1_addr), .B(_tmp_207), .S(_06235_), .Y(_27686_) );
  \$mux  #( .WIDTH(10) ) _52174_ ( .A(_27686_), .B(10'h000), .S(RST), .Y(_03458_) );
  \$mux  #( .WIDTH(10) ) _52175_ ( .A(ram_w4_l8192_id2_5_0_addr), .B(_stream_conv2d_16_source_30_source_ram_raddr[12:3]), .S(_tmp_625), .Y(_27687_) );
  \$mux  #( .WIDTH(10) ) _52176_ ( .A(_27687_), .B(10'h000), .S(RST), .Y(_03457_) );
  \$mux  #( .WIDTH(1) ) _52177_ ( .A(ram_w4_l8192_id2_4_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27688_) );
  \$mux  #( .WIDTH(1) ) _52178_ ( .A(_27688_), .B(_06066_), .S(_06232_), .Y(_27689_) );
  \$mux  #( .WIDTH(1) ) _52179_ ( .A(_27689_), .B(1'h0), .S(RST), .Y(_03456_) );
  \$mux  #( .WIDTH(4) ) _52180_ ( .A(ram_w4_l8192_id2_4_1_wdata), .B(_dataflow_slice_data_41), .S(_06232_), .Y(_27690_) );
  \$mux  #( .WIDTH(4) ) _52181_ ( .A(_27690_), .B(4'h0), .S(RST), .Y(_03455_) );
  \$mux  #( .WIDTH(10) ) _52182_ ( .A(ram_w4_l8192_id2_4_1_addr), .B(_tmp_176), .S(_06232_), .Y(_27691_) );
  \$mux  #( .WIDTH(10) ) _52183_ ( .A(_27691_), .B(10'h000), .S(RST), .Y(_03454_) );
  \$mux  #( .WIDTH(10) ) _52184_ ( .A(ram_w4_l8192_id2_4_0_addr), .B(_stream_conv2d_16_source_30_source_ram_raddr[12:3]), .S(_tmp_625), .Y(_27692_) );
  \$mux  #( .WIDTH(10) ) _52185_ ( .A(_27692_), .B(10'h000), .S(RST), .Y(_03453_) );
  \$mux  #( .WIDTH(1) ) _52186_ ( .A(ram_w4_l8192_id2_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27693_) );
  \$mux  #( .WIDTH(1) ) _52187_ ( .A(_27693_), .B(_06057_), .S(_06229_), .Y(_27694_) );
  \$mux  #( .WIDTH(1) ) _52188_ ( .A(_27694_), .B(1'h0), .S(RST), .Y(_03452_) );
  \$mux  #( .WIDTH(4) ) _52189_ ( .A(ram_w4_l8192_id2_3_1_wdata), .B(_dataflow_slice_data_38), .S(_06229_), .Y(_27695_) );
  \$mux  #( .WIDTH(4) ) _52190_ ( .A(_27695_), .B(4'h0), .S(RST), .Y(_03451_) );
  \$mux  #( .WIDTH(10) ) _52191_ ( .A(ram_w4_l8192_id2_3_1_addr), .B(_tmp_145), .S(_06229_), .Y(_27696_) );
  \$mux  #( .WIDTH(10) ) _52192_ ( .A(_27696_), .B(10'h000), .S(RST), .Y(_03450_) );
  \$mux  #( .WIDTH(10) ) _52193_ ( .A(ram_w4_l8192_id2_3_0_addr), .B(_stream_conv2d_16_source_30_source_ram_raddr[12:3]), .S(_tmp_625), .Y(_27697_) );
  \$mux  #( .WIDTH(10) ) _52194_ ( .A(_27697_), .B(10'h000), .S(RST), .Y(_03449_) );
  \$mux  #( .WIDTH(1) ) _52195_ ( .A(ram_w4_l8192_id2_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27698_) );
  \$mux  #( .WIDTH(1) ) _52196_ ( .A(_27698_), .B(_06048_), .S(_06226_), .Y(_27699_) );
  \$mux  #( .WIDTH(1) ) _52197_ ( .A(_27699_), .B(1'h0), .S(RST), .Y(_03448_) );
  \$mux  #( .WIDTH(4) ) _52198_ ( .A(ram_w4_l8192_id2_2_1_wdata), .B(_dataflow_slice_data_35), .S(_06226_), .Y(_27700_) );
  \$mux  #( .WIDTH(4) ) _52199_ ( .A(_27700_), .B(4'h0), .S(RST), .Y(_03447_) );
  \$mux  #( .WIDTH(10) ) _52200_ ( .A(ram_w4_l8192_id2_2_1_addr), .B(_tmp_114), .S(_06226_), .Y(_27701_) );
  \$mux  #( .WIDTH(10) ) _52201_ ( .A(_27701_), .B(10'h000), .S(RST), .Y(_03446_) );
  \$mux  #( .WIDTH(10) ) _52202_ ( .A(ram_w4_l8192_id2_2_0_addr), .B(_stream_conv2d_16_source_30_source_ram_raddr[12:3]), .S(_tmp_625), .Y(_27702_) );
  \$mux  #( .WIDTH(10) ) _52203_ ( .A(_27702_), .B(10'h000), .S(RST), .Y(_03445_) );
  \$mux  #( .WIDTH(1) ) _52204_ ( .A(ram_w4_l8192_id2_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27703_) );
  \$mux  #( .WIDTH(1) ) _52205_ ( .A(_27703_), .B(_06039_), .S(_06223_), .Y(_27704_) );
  \$mux  #( .WIDTH(1) ) _52206_ ( .A(_27704_), .B(1'h0), .S(RST), .Y(_03444_) );
  \$mux  #( .WIDTH(4) ) _52207_ ( .A(ram_w4_l8192_id2_1_1_wdata), .B(_dataflow_slice_data_32), .S(_06223_), .Y(_27705_) );
  \$mux  #( .WIDTH(4) ) _52208_ ( .A(_27705_), .B(4'h0), .S(RST), .Y(_03443_) );
  \$mux  #( .WIDTH(10) ) _52209_ ( .A(ram_w4_l8192_id2_1_1_addr), .B(_tmp_83), .S(_06223_), .Y(_27706_) );
  \$mux  #( .WIDTH(10) ) _52210_ ( .A(_27706_), .B(10'h000), .S(RST), .Y(_03442_) );
  \$mux  #( .WIDTH(10) ) _52211_ ( .A(ram_w4_l8192_id2_1_0_addr), .B(_stream_conv2d_16_source_30_source_ram_raddr[12:3]), .S(_tmp_625), .Y(_27707_) );
  \$mux  #( .WIDTH(10) ) _52212_ ( .A(_27707_), .B(10'h000), .S(RST), .Y(_03441_) );
  \$mux  #( .WIDTH(1) ) _52213_ ( .A(ram_w4_l8192_id2_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27708_) );
  \$mux  #( .WIDTH(1) ) _52214_ ( .A(_27708_), .B(_06030_), .S(_06220_), .Y(_27709_) );
  \$mux  #( .WIDTH(1) ) _52215_ ( .A(_27709_), .B(1'h0), .S(RST), .Y(_03440_) );
  \$mux  #( .WIDTH(4) ) _52216_ ( .A(ram_w4_l8192_id2_0_1_wdata), .B(_dataflow_slice_data_29), .S(_06220_), .Y(_27710_) );
  \$mux  #( .WIDTH(4) ) _52217_ ( .A(_27710_), .B(4'h0), .S(RST), .Y(_03439_) );
  \$mux  #( .WIDTH(10) ) _52218_ ( .A(ram_w4_l8192_id2_0_1_addr), .B(_tmp_52), .S(_06220_), .Y(_27711_) );
  \$mux  #( .WIDTH(10) ) _52219_ ( .A(_27711_), .B(10'h000), .S(RST), .Y(_03438_) );
  \$mux  #( .WIDTH(10) ) _52220_ ( .A(ram_w4_l8192_id2_0_0_addr), .B(_stream_conv2d_16_source_30_source_ram_raddr[12:3]), .S(_tmp_625), .Y(_27712_) );
  \$mux  #( .WIDTH(10) ) _52221_ ( .A(_27712_), .B(10'h000), .S(RST), .Y(_03437_) );
  \$mux  #( .WIDTH(1) ) _52222_ ( .A(ram_w4_l8192_id1_7_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27713_) );
  \$mux  #( .WIDTH(1) ) _52223_ ( .A(_27713_), .B(_06092_), .S(_06241_), .Y(_27714_) );
  \$mux  #( .WIDTH(1) ) _52224_ ( .A(_27714_), .B(1'h0), .S(RST), .Y(_03436_) );
  \$mux  #( .WIDTH(4) ) _52225_ ( .A(ram_w4_l8192_id1_7_1_wdata), .B(_dataflow_slice_data_50), .S(_06241_), .Y(_27715_) );
  \$mux  #( .WIDTH(4) ) _52226_ ( .A(_27715_), .B(4'h0), .S(RST), .Y(_03435_) );
  \$mux  #( .WIDTH(10) ) _52227_ ( .A(ram_w4_l8192_id1_7_1_addr), .B(_tmp_268), .S(_06241_), .Y(_27716_) );
  \$mux  #( .WIDTH(10) ) _52228_ ( .A(_27716_), .B(10'h000), .S(RST), .Y(_03434_) );
  \$mux  #( .WIDTH(10) ) _52229_ ( .A(ram_w4_l8192_id1_7_0_addr), .B(_stream_conv2d_16_source_29_source_ram_raddr[12:3]), .S(_tmp_611), .Y(_27717_) );
  \$mux  #( .WIDTH(10) ) _52230_ ( .A(_27717_), .B(10'h000), .S(RST), .Y(_03433_) );
  \$mux  #( .WIDTH(1) ) _52231_ ( .A(ram_w4_l8192_id1_6_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27718_) );
  \$mux  #( .WIDTH(1) ) _52232_ ( .A(_27718_), .B(_06083_), .S(_06238_), .Y(_27719_) );
  \$mux  #( .WIDTH(1) ) _52233_ ( .A(_27719_), .B(1'h0), .S(RST), .Y(_03432_) );
  \$mux  #( .WIDTH(4) ) _52234_ ( .A(ram_w4_l8192_id1_6_1_wdata), .B(_dataflow_slice_data_47), .S(_06238_), .Y(_27720_) );
  \$mux  #( .WIDTH(4) ) _52235_ ( .A(_27720_), .B(4'h0), .S(RST), .Y(_03431_) );
  \$mux  #( .WIDTH(10) ) _52236_ ( .A(ram_w4_l8192_id1_6_1_addr), .B(_tmp_237), .S(_06238_), .Y(_27721_) );
  \$mux  #( .WIDTH(10) ) _52237_ ( .A(_27721_), .B(10'h000), .S(RST), .Y(_03430_) );
  \$mux  #( .WIDTH(10) ) _52238_ ( .A(ram_w4_l8192_id1_6_0_addr), .B(_stream_conv2d_16_source_29_source_ram_raddr[12:3]), .S(_tmp_611), .Y(_27722_) );
  \$mux  #( .WIDTH(10) ) _52239_ ( .A(_27722_), .B(10'h000), .S(RST), .Y(_03429_) );
  \$mux  #( .WIDTH(1) ) _52240_ ( .A(ram_w4_l8192_id1_5_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27723_) );
  \$mux  #( .WIDTH(1) ) _52241_ ( .A(_27723_), .B(_06074_), .S(_06235_), .Y(_27724_) );
  \$mux  #( .WIDTH(1) ) _52242_ ( .A(_27724_), .B(1'h0), .S(RST), .Y(_03428_) );
  \$mux  #( .WIDTH(4) ) _52243_ ( .A(ram_w4_l8192_id1_5_1_wdata), .B(_dataflow_slice_data_44), .S(_06235_), .Y(_27725_) );
  \$mux  #( .WIDTH(4) ) _52244_ ( .A(_27725_), .B(4'h0), .S(RST), .Y(_03427_) );
  \$mux  #( .WIDTH(10) ) _52245_ ( .A(ram_w4_l8192_id1_5_1_addr), .B(_tmp_206), .S(_06235_), .Y(_27726_) );
  \$mux  #( .WIDTH(10) ) _52246_ ( .A(_27726_), .B(10'h000), .S(RST), .Y(_03426_) );
  \$mux  #( .WIDTH(10) ) _52247_ ( .A(ram_w4_l8192_id1_5_0_addr), .B(_stream_conv2d_16_source_29_source_ram_raddr[12:3]), .S(_tmp_611), .Y(_27727_) );
  \$mux  #( .WIDTH(10) ) _52248_ ( .A(_27727_), .B(10'h000), .S(RST), .Y(_03425_) );
  \$mux  #( .WIDTH(1) ) _52249_ ( .A(ram_w4_l8192_id1_4_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27728_) );
  \$mux  #( .WIDTH(1) ) _52250_ ( .A(_27728_), .B(_06065_), .S(_06232_), .Y(_27729_) );
  \$mux  #( .WIDTH(1) ) _52251_ ( .A(_27729_), .B(1'h0), .S(RST), .Y(_03424_) );
  \$mux  #( .WIDTH(4) ) _52252_ ( .A(ram_w4_l8192_id1_4_1_wdata), .B(_dataflow_slice_data_41), .S(_06232_), .Y(_27730_) );
  \$mux  #( .WIDTH(4) ) _52253_ ( .A(_27730_), .B(4'h0), .S(RST), .Y(_03423_) );
  \$mux  #( .WIDTH(10) ) _52254_ ( .A(ram_w4_l8192_id1_4_1_addr), .B(_tmp_175), .S(_06232_), .Y(_27731_) );
  \$mux  #( .WIDTH(10) ) _52255_ ( .A(_27731_), .B(10'h000), .S(RST), .Y(_03422_) );
  \$mux  #( .WIDTH(10) ) _52256_ ( .A(ram_w4_l8192_id1_4_0_addr), .B(_stream_conv2d_16_source_29_source_ram_raddr[12:3]), .S(_tmp_611), .Y(_27732_) );
  \$mux  #( .WIDTH(10) ) _52257_ ( .A(_27732_), .B(10'h000), .S(RST), .Y(_03421_) );
  \$mux  #( .WIDTH(1) ) _52258_ ( .A(ram_w4_l8192_id1_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27733_) );
  \$mux  #( .WIDTH(1) ) _52259_ ( .A(_27733_), .B(_06056_), .S(_06229_), .Y(_27734_) );
  \$mux  #( .WIDTH(1) ) _52260_ ( .A(_27734_), .B(1'h0), .S(RST), .Y(_03420_) );
  \$mux  #( .WIDTH(4) ) _52261_ ( .A(ram_w4_l8192_id1_3_1_wdata), .B(_dataflow_slice_data_38), .S(_06229_), .Y(_27735_) );
  \$mux  #( .WIDTH(4) ) _52262_ ( .A(_27735_), .B(4'h0), .S(RST), .Y(_03419_) );
  \$mux  #( .WIDTH(10) ) _52263_ ( .A(ram_w4_l8192_id1_3_1_addr), .B(_tmp_144), .S(_06229_), .Y(_27736_) );
  \$mux  #( .WIDTH(10) ) _52264_ ( .A(_27736_), .B(10'h000), .S(RST), .Y(_03418_) );
  \$mux  #( .WIDTH(10) ) _52265_ ( .A(ram_w4_l8192_id1_3_0_addr), .B(_stream_conv2d_16_source_29_source_ram_raddr[12:3]), .S(_tmp_611), .Y(_27737_) );
  \$mux  #( .WIDTH(10) ) _52266_ ( .A(_27737_), .B(10'h000), .S(RST), .Y(_03417_) );
  \$mux  #( .WIDTH(1) ) _52267_ ( .A(ram_w4_l8192_id1_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27738_) );
  \$mux  #( .WIDTH(1) ) _52268_ ( .A(_27738_), .B(_06047_), .S(_06226_), .Y(_27739_) );
  \$mux  #( .WIDTH(1) ) _52269_ ( .A(_27739_), .B(1'h0), .S(RST), .Y(_03416_) );
  \$mux  #( .WIDTH(4) ) _52270_ ( .A(ram_w4_l8192_id1_2_1_wdata), .B(_dataflow_slice_data_35), .S(_06226_), .Y(_27740_) );
  \$mux  #( .WIDTH(4) ) _52271_ ( .A(_27740_), .B(4'h0), .S(RST), .Y(_03415_) );
  \$mux  #( .WIDTH(10) ) _52272_ ( .A(ram_w4_l8192_id1_2_1_addr), .B(_tmp_113), .S(_06226_), .Y(_27741_) );
  \$mux  #( .WIDTH(10) ) _52273_ ( .A(_27741_), .B(10'h000), .S(RST), .Y(_03414_) );
  \$mux  #( .WIDTH(10) ) _52274_ ( .A(ram_w4_l8192_id1_2_0_addr), .B(_stream_conv2d_16_source_29_source_ram_raddr[12:3]), .S(_tmp_611), .Y(_27742_) );
  \$mux  #( .WIDTH(10) ) _52275_ ( .A(_27742_), .B(10'h000), .S(RST), .Y(_03413_) );
  \$mux  #( .WIDTH(1) ) _52276_ ( .A(ram_w4_l8192_id1_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27743_) );
  \$mux  #( .WIDTH(1) ) _52277_ ( .A(_27743_), .B(_06038_), .S(_06223_), .Y(_27744_) );
  \$mux  #( .WIDTH(1) ) _52278_ ( .A(_27744_), .B(1'h0), .S(RST), .Y(_03412_) );
  \$mux  #( .WIDTH(4) ) _52279_ ( .A(ram_w4_l8192_id1_1_1_wdata), .B(_dataflow_slice_data_32), .S(_06223_), .Y(_27745_) );
  \$mux  #( .WIDTH(4) ) _52280_ ( .A(_27745_), .B(4'h0), .S(RST), .Y(_03411_) );
  \$mux  #( .WIDTH(10) ) _52281_ ( .A(ram_w4_l8192_id1_1_1_addr), .B(_tmp_82), .S(_06223_), .Y(_27746_) );
  \$mux  #( .WIDTH(10) ) _52282_ ( .A(_27746_), .B(10'h000), .S(RST), .Y(_03410_) );
  \$mux  #( .WIDTH(10) ) _52283_ ( .A(ram_w4_l8192_id1_1_0_addr), .B(_stream_conv2d_16_source_29_source_ram_raddr[12:3]), .S(_tmp_611), .Y(_27747_) );
  \$mux  #( .WIDTH(10) ) _52284_ ( .A(_27747_), .B(10'h000), .S(RST), .Y(_03409_) );
  \$mux  #( .WIDTH(1) ) _52285_ ( .A(ram_w4_l8192_id1_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27748_) );
  \$mux  #( .WIDTH(1) ) _52286_ ( .A(_27748_), .B(_06029_), .S(_06220_), .Y(_27749_) );
  \$mux  #( .WIDTH(1) ) _52287_ ( .A(_27749_), .B(1'h0), .S(RST), .Y(_03408_) );
  \$mux  #( .WIDTH(4) ) _52288_ ( .A(ram_w4_l8192_id1_0_1_wdata), .B(_dataflow_slice_data_29), .S(_06220_), .Y(_27750_) );
  \$mux  #( .WIDTH(4) ) _52289_ ( .A(_27750_), .B(4'h0), .S(RST), .Y(_03407_) );
  \$mux  #( .WIDTH(10) ) _52290_ ( .A(ram_w4_l8192_id1_0_1_addr), .B(_tmp_51), .S(_06220_), .Y(_27751_) );
  \$mux  #( .WIDTH(10) ) _52291_ ( .A(_27751_), .B(10'h000), .S(RST), .Y(_03406_) );
  \$mux  #( .WIDTH(10) ) _52292_ ( .A(ram_w4_l8192_id1_0_0_addr), .B(_stream_conv2d_16_source_29_source_ram_raddr[12:3]), .S(_tmp_611), .Y(_27752_) );
  \$mux  #( .WIDTH(10) ) _52293_ ( .A(_27752_), .B(10'h000), .S(RST), .Y(_03405_) );
  \$mux  #( .WIDTH(1) ) _52294_ ( .A(_tmp_1151), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27753_) );
  \$mux  #( .WIDTH(1) ) _52295_ ( .A(_27753_), .B(1'h1), .S(_06481_), .Y(_27754_) );
  \$mux  #( .WIDTH(1) ) _52296_ ( .A(_27754_), .B(1'h0), .S(RST), .Y(_02927_) );
  \$mux  #( .WIDTH(34) ) _52297_ ( .A(_tmp_1150), .B({ 1'h0, _maxi_read_size }), .S(_06480_), .Y(_27755_) );
  \$mux  #( .WIDTH(34) ) _52298_ ( .A(_27755_), .B(_28561_), .S(_06313_), .Y(_27756_) );
  \$mux  #( .WIDTH(34) ) _52299_ ( .A(_27756_), .B(34'h000000000), .S(RST), .Y(_02926_) );
  \$mux  #( .WIDTH(4) ) _52300_ ( .A(_tmp_285), .B(4'h0), .S(_06467_), .Y(_27757_) );
  \$mux  #( .WIDTH(4) ) _52301_ ( .A(_27757_), .B(_24248_[3:0]), .S(_06468_), .Y(_27758_) );
  \$mux  #( .WIDTH(4) ) _52302_ ( .A(_27758_), .B(4'h0), .S(_06469_), .Y(_27759_) );
  \$mux  #( .WIDTH(4) ) _52303_ ( .A(_27759_), .B(4'h0), .S(RST), .Y(_03039_) );
  \$mux  #( .WIDTH(10) ) _52304_ ( .A(_tmp_266), .B(_28537_[9:0]), .S(_06467_), .Y(_27760_) );
  \$mux  #( .WIDTH(10) ) _52305_ ( .A(_27760_), .B(_tmp_275), .S(_06478_), .Y(_27761_) );
  \$mux  #( .WIDTH(10) ) _52306_ ( .A(_27761_), .B(10'h000), .S(RST), .Y(_03036_) );
  \$mux  #( .WIDTH(10) ) _52307_ ( .A(_tmp_265), .B(_28537_[9:0]), .S(_06467_), .Y(_27762_) );
  \$mux  #( .WIDTH(10) ) _52308_ ( .A(_27762_), .B(_tmp_274), .S(_06477_), .Y(_27763_) );
  \$mux  #( .WIDTH(10) ) _52309_ ( .A(_27763_), .B(10'h000), .S(RST), .Y(_03035_) );
  \$mux  #( .WIDTH(10) ) _52310_ ( .A(_tmp_264), .B(_28537_[9:0]), .S(_06467_), .Y(_27764_) );
  \$mux  #( .WIDTH(10) ) _52311_ ( .A(_27764_), .B(_tmp_273), .S(_06476_), .Y(_27765_) );
  \$mux  #( .WIDTH(10) ) _52312_ ( .A(_27765_), .B(10'h000), .S(RST), .Y(_03034_) );
  \$mux  #( .WIDTH(10) ) _52313_ ( .A(_tmp_263), .B(_28537_[9:0]), .S(_06467_), .Y(_27766_) );
  \$mux  #( .WIDTH(10) ) _52314_ ( .A(_27766_), .B(_tmp_272), .S(_06475_), .Y(_27767_) );
  \$mux  #( .WIDTH(10) ) _52315_ ( .A(_27767_), .B(10'h000), .S(RST), .Y(_03033_) );
  \$mux  #( .WIDTH(10) ) _52316_ ( .A(_tmp_262), .B(_28537_[9:0]), .S(_06467_), .Y(_27768_) );
  \$mux  #( .WIDTH(10) ) _52317_ ( .A(_27768_), .B(_tmp_271), .S(_06474_), .Y(_27769_) );
  \$mux  #( .WIDTH(10) ) _52318_ ( .A(_27769_), .B(10'h000), .S(RST), .Y(_03032_) );
  \$mux  #( .WIDTH(10) ) _52319_ ( .A(_tmp_261), .B(_28537_[9:0]), .S(_06467_), .Y(_27770_) );
  \$mux  #( .WIDTH(10) ) _52320_ ( .A(_27770_), .B(_tmp_270), .S(_06473_), .Y(_27771_) );
  \$mux  #( .WIDTH(10) ) _52321_ ( .A(_27771_), .B(10'h000), .S(RST), .Y(_03031_) );
  \$mux  #( .WIDTH(10) ) _52322_ ( .A(_tmp_260), .B(_28537_[9:0]), .S(_06467_), .Y(_27772_) );
  \$mux  #( .WIDTH(10) ) _52323_ ( .A(_27772_), .B(_tmp_269), .S(_06472_), .Y(_27773_) );
  \$mux  #( .WIDTH(10) ) _52324_ ( .A(_27773_), .B(10'h000), .S(RST), .Y(_03030_) );
  \$mux  #( .WIDTH(10) ) _52325_ ( .A(_tmp_259), .B(_28537_[9:0]), .S(_06467_), .Y(_27774_) );
  \$mux  #( .WIDTH(10) ) _52326_ ( .A(_27774_), .B(_tmp_268), .S(_06471_), .Y(_27775_) );
  \$mux  #( .WIDTH(10) ) _52327_ ( .A(_27775_), .B(10'h000), .S(RST), .Y(_03028_) );
  \$mux  #( .WIDTH(10) ) _52328_ ( .A(_tmp_258), .B(_28537_[9:0]), .S(_06467_), .Y(_27776_) );
  \$mux  #( .WIDTH(10) ) _52329_ ( .A(_27776_), .B(_tmp_267), .S(_06470_), .Y(_27777_) );
  \$mux  #( .WIDTH(10) ) _52330_ ( .A(_27777_), .B(10'h000), .S(RST), .Y(_03027_) );
  \$mux  #( .WIDTH(1) ) _52331_ ( .A(_tmp_257), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27778_) );
  \$mux  #( .WIDTH(1) ) _52332_ ( .A(_27778_), .B(1'h1), .S(_06479_), .Y(_27779_) );
  \$mux  #( .WIDTH(1) ) _52333_ ( .A(_27779_), .B(1'h0), .S(RST), .Y(_03026_) );
  \$mux  #( .WIDTH(34) ) _52334_ ( .A(_tmp_256), .B({ 1'h0, _maxi_read_size }), .S(_06467_), .Y(_27780_) );
  \$mux  #( .WIDTH(34) ) _52335_ ( .A(_27780_), .B(_28560_), .S(_06241_), .Y(_27781_) );
  \$mux  #( .WIDTH(34) ) _52336_ ( .A(_27781_), .B(34'h000000000), .S(RST), .Y(_03025_) );
  \$mux  #( .WIDTH(11) ) _52337_ ( .A(_tmp_255), .B(_28536_[10:0]), .S(_06467_), .Y(_27782_) );
  \$mux  #( .WIDTH(11) ) _52338_ ( .A(_27782_), .B(_28559_[10:0]), .S(_06241_), .Y(_27783_) );
  \$mux  #( .WIDTH(11) ) _52339_ ( .A(_27783_), .B(_28536_[10:0]), .S(_06468_), .Y(_27784_) );
  \$mux  #( .WIDTH(11) ) _52340_ ( .A(_27784_), .B(11'h000), .S(RST), .Y(_03024_) );
  \$mux  #( .WIDTH(1) ) _52341_ ( .A(ram_w4_l8192_id0_7_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27785_) );
  \$mux  #( .WIDTH(1) ) _52342_ ( .A(_27785_), .B(_06091_), .S(_06241_), .Y(_27786_) );
  \$mux  #( .WIDTH(1) ) _52343_ ( .A(_27786_), .B(1'h1), .S(_06313_), .Y(_27787_) );
  \$mux  #( .WIDTH(1) ) _52344_ ( .A(_27787_), .B(1'h0), .S(RST), .Y(_03404_) );
  \$mux  #( .WIDTH(4) ) _52345_ ( .A(ram_w4_l8192_id0_7_1_wdata), .B(_dataflow_slice_data_50), .S(_06241_), .Y(_27788_) );
  \$mux  #( .WIDTH(4) ) _52346_ ( .A(_27788_), .B(_dataflow_slice_data_145), .S(_06313_), .Y(_27789_) );
  \$mux  #( .WIDTH(4) ) _52347_ ( .A(_27789_), .B(4'h0), .S(RST), .Y(_03403_) );
  \$mux  #( .WIDTH(10) ) _52348_ ( .A(ram_w4_l8192_id0_7_1_addr), .B(_tmp_267), .S(_06241_), .Y(_27790_) );
  \$mux  #( .WIDTH(10) ) _52349_ ( .A(_27790_), .B(_28537_[9:0]), .S(_06480_), .Y(_27791_) );
  \$mux  #( .WIDTH(10) ) _52350_ ( .A(_27791_), .B(_24249_[9:0]), .S(_06313_), .Y(_27792_) );
  \$mux  #( .WIDTH(10) ) _52351_ ( .A(_27792_), .B(10'h000), .S(RST), .Y(_03402_) );
  \$mux  #( .WIDTH(10) ) _52352_ ( .A(ram_w4_l8192_id0_7_0_addr), .B(_stream_conv2d_16_source_28_source_ram_raddr[12:3]), .S(_tmp_597), .Y(_27793_) );
  \$mux  #( .WIDTH(10) ) _52353_ ( .A(_27793_), .B(_stream_matmul_29_source_20_source_ram_raddr[12:3]), .S(_tmp_1223), .Y(_27794_) );
  \$mux  #( .WIDTH(10) ) _52354_ ( .A(_27794_), .B(10'h000), .S(RST), .Y(_03401_) );
  \$mux  #( .WIDTH(1) ) _52355_ ( .A(_tmp_1149), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27795_) );
  \$mux  #( .WIDTH(1) ) _52356_ ( .A(_27795_), .B(1'h1), .S(_06466_), .Y(_27796_) );
  \$mux  #( .WIDTH(1) ) _52357_ ( .A(_27796_), .B(1'h0), .S(RST), .Y(_02925_) );
  \$mux  #( .WIDTH(34) ) _52358_ ( .A(_tmp_1148), .B({ 1'h0, _maxi_read_size }), .S(_06465_), .Y(_27797_) );
  \$mux  #( .WIDTH(34) ) _52359_ ( .A(_27797_), .B(_28558_), .S(_06310_), .Y(_27798_) );
  \$mux  #( .WIDTH(34) ) _52360_ ( .A(_27798_), .B(34'h000000000), .S(RST), .Y(_02924_) );
  \$mux  #( .WIDTH(4) ) _52361_ ( .A(_tmp_254), .B(4'h0), .S(_06452_), .Y(_27799_) );
  \$mux  #( .WIDTH(4) ) _52362_ ( .A(_27799_), .B(_24246_[3:0]), .S(_06453_), .Y(_27800_) );
  \$mux  #( .WIDTH(4) ) _52363_ ( .A(_27800_), .B(4'h0), .S(_06454_), .Y(_27801_) );
  \$mux  #( .WIDTH(4) ) _52364_ ( .A(_27801_), .B(4'h0), .S(RST), .Y(_03023_) );
  \$mux  #( .WIDTH(10) ) _52365_ ( .A(_tmp_235), .B(_28537_[9:0]), .S(_06452_), .Y(_27802_) );
  \$mux  #( .WIDTH(10) ) _52366_ ( .A(_27802_), .B(_tmp_244), .S(_06463_), .Y(_27803_) );
  \$mux  #( .WIDTH(10) ) _52367_ ( .A(_27803_), .B(10'h000), .S(RST), .Y(_03022_) );
  \$mux  #( .WIDTH(10) ) _52368_ ( .A(_tmp_234), .B(_28537_[9:0]), .S(_06452_), .Y(_27804_) );
  \$mux  #( .WIDTH(10) ) _52369_ ( .A(_27804_), .B(_tmp_243), .S(_06462_), .Y(_27805_) );
  \$mux  #( .WIDTH(10) ) _52370_ ( .A(_27805_), .B(10'h000), .S(RST), .Y(_03021_) );
  \$mux  #( .WIDTH(10) ) _52371_ ( .A(_tmp_233), .B(_28537_[9:0]), .S(_06452_), .Y(_27806_) );
  \$mux  #( .WIDTH(10) ) _52372_ ( .A(_27806_), .B(_tmp_242), .S(_06461_), .Y(_27807_) );
  \$mux  #( .WIDTH(10) ) _52373_ ( .A(_27807_), .B(10'h000), .S(RST), .Y(_03020_) );
  \$mux  #( .WIDTH(10) ) _52374_ ( .A(_tmp_232), .B(_28537_[9:0]), .S(_06452_), .Y(_27808_) );
  \$mux  #( .WIDTH(10) ) _52375_ ( .A(_27808_), .B(_tmp_241), .S(_06460_), .Y(_27809_) );
  \$mux  #( .WIDTH(10) ) _52376_ ( .A(_27809_), .B(10'h000), .S(RST), .Y(_03019_) );
  \$mux  #( .WIDTH(10) ) _52377_ ( .A(_tmp_231), .B(_28537_[9:0]), .S(_06452_), .Y(_27810_) );
  \$mux  #( .WIDTH(10) ) _52378_ ( .A(_27810_), .B(_tmp_240), .S(_06459_), .Y(_27811_) );
  \$mux  #( .WIDTH(10) ) _52379_ ( .A(_27811_), .B(10'h000), .S(RST), .Y(_03018_) );
  \$mux  #( .WIDTH(10) ) _52380_ ( .A(_tmp_230), .B(_28537_[9:0]), .S(_06452_), .Y(_27812_) );
  \$mux  #( .WIDTH(10) ) _52381_ ( .A(_27812_), .B(_tmp_239), .S(_06458_), .Y(_27813_) );
  \$mux  #( .WIDTH(10) ) _52382_ ( .A(_27813_), .B(10'h000), .S(RST), .Y(_03017_) );
  \$mux  #( .WIDTH(10) ) _52383_ ( .A(_tmp_229), .B(_28537_[9:0]), .S(_06452_), .Y(_27814_) );
  \$mux  #( .WIDTH(10) ) _52384_ ( .A(_27814_), .B(_tmp_238), .S(_06457_), .Y(_27815_) );
  \$mux  #( .WIDTH(10) ) _52385_ ( .A(_27815_), .B(10'h000), .S(RST), .Y(_03016_) );
  \$mux  #( .WIDTH(10) ) _52386_ ( .A(_tmp_228), .B(_28537_[9:0]), .S(_06452_), .Y(_27816_) );
  \$mux  #( .WIDTH(10) ) _52387_ ( .A(_27816_), .B(_tmp_237), .S(_06456_), .Y(_27817_) );
  \$mux  #( .WIDTH(10) ) _52388_ ( .A(_27817_), .B(10'h000), .S(RST), .Y(_03015_) );
  \$mux  #( .WIDTH(10) ) _52389_ ( .A(_tmp_227), .B(_28537_[9:0]), .S(_06452_), .Y(_27818_) );
  \$mux  #( .WIDTH(10) ) _52390_ ( .A(_27818_), .B(_tmp_236), .S(_06455_), .Y(_27819_) );
  \$mux  #( .WIDTH(10) ) _52391_ ( .A(_27819_), .B(10'h000), .S(RST), .Y(_03014_) );
  \$mux  #( .WIDTH(1) ) _52392_ ( .A(_tmp_226), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27820_) );
  \$mux  #( .WIDTH(1) ) _52393_ ( .A(_27820_), .B(1'h1), .S(_06464_), .Y(_27821_) );
  \$mux  #( .WIDTH(1) ) _52394_ ( .A(_27821_), .B(1'h0), .S(RST), .Y(_03013_) );
  \$mux  #( .WIDTH(34) ) _52395_ ( .A(_tmp_225), .B({ 1'h0, _maxi_read_size }), .S(_06452_), .Y(_27822_) );
  \$mux  #( .WIDTH(34) ) _52396_ ( .A(_27822_), .B(_28557_), .S(_06238_), .Y(_27823_) );
  \$mux  #( .WIDTH(34) ) _52397_ ( .A(_27823_), .B(34'h000000000), .S(RST), .Y(_03012_) );
  \$mux  #( .WIDTH(11) ) _52398_ ( .A(_tmp_224), .B(_28536_[10:0]), .S(_06452_), .Y(_27824_) );
  \$mux  #( .WIDTH(11) ) _52399_ ( .A(_27824_), .B(_28556_[10:0]), .S(_06238_), .Y(_27825_) );
  \$mux  #( .WIDTH(11) ) _52400_ ( .A(_27825_), .B(_28536_[10:0]), .S(_06453_), .Y(_27826_) );
  \$mux  #( .WIDTH(11) ) _52401_ ( .A(_27826_), .B(11'h000), .S(RST), .Y(_03011_) );
  \$mux  #( .WIDTH(1) ) _52402_ ( .A(ram_w4_l8192_id0_6_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27827_) );
  \$mux  #( .WIDTH(1) ) _52403_ ( .A(_27827_), .B(_06082_), .S(_06238_), .Y(_27828_) );
  \$mux  #( .WIDTH(1) ) _52404_ ( .A(_27828_), .B(1'h1), .S(_06310_), .Y(_27829_) );
  \$mux  #( .WIDTH(1) ) _52405_ ( .A(_27829_), .B(1'h0), .S(RST), .Y(_03400_) );
  \$mux  #( .WIDTH(4) ) _52406_ ( .A(ram_w4_l8192_id0_6_1_wdata), .B(_dataflow_slice_data_47), .S(_06238_), .Y(_27830_) );
  \$mux  #( .WIDTH(4) ) _52407_ ( .A(_27830_), .B(_dataflow_slice_data_142), .S(_06310_), .Y(_27831_) );
  \$mux  #( .WIDTH(4) ) _52408_ ( .A(_27831_), .B(4'h0), .S(RST), .Y(_03399_) );
  \$mux  #( .WIDTH(10) ) _52409_ ( .A(ram_w4_l8192_id0_6_1_addr), .B(_tmp_236), .S(_06238_), .Y(_27832_) );
  \$mux  #( .WIDTH(10) ) _52410_ ( .A(_27832_), .B(_28537_[9:0]), .S(_06465_), .Y(_27833_) );
  \$mux  #( .WIDTH(10) ) _52411_ ( .A(_27833_), .B(_24247_[9:0]), .S(_06310_), .Y(_27834_) );
  \$mux  #( .WIDTH(10) ) _52412_ ( .A(_27834_), .B(10'h000), .S(RST), .Y(_03398_) );
  \$mux  #( .WIDTH(10) ) _52413_ ( .A(ram_w4_l8192_id0_6_0_addr), .B(_stream_conv2d_16_source_28_source_ram_raddr[12:3]), .S(_tmp_597), .Y(_27835_) );
  \$mux  #( .WIDTH(10) ) _52414_ ( .A(_27835_), .B(_stream_matmul_29_source_20_source_ram_raddr[12:3]), .S(_tmp_1223), .Y(_27836_) );
  \$mux  #( .WIDTH(10) ) _52415_ ( .A(_27836_), .B(10'h000), .S(RST), .Y(_03397_) );
  \$mux  #( .WIDTH(1) ) _52416_ ( .A(_tmp_1147), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27837_) );
  \$mux  #( .WIDTH(1) ) _52417_ ( .A(_27837_), .B(1'h1), .S(_06451_), .Y(_27838_) );
  \$mux  #( .WIDTH(1) ) _52418_ ( .A(_27838_), .B(1'h0), .S(RST), .Y(_02923_) );
  \$mux  #( .WIDTH(34) ) _52419_ ( .A(_tmp_1146), .B({ 1'h0, _maxi_read_size }), .S(_06450_), .Y(_27839_) );
  \$mux  #( .WIDTH(34) ) _52420_ ( .A(_27839_), .B(_28555_), .S(_06307_), .Y(_27840_) );
  \$mux  #( .WIDTH(34) ) _52421_ ( .A(_27840_), .B(34'h000000000), .S(RST), .Y(_02922_) );
  \$mux  #( .WIDTH(4) ) _52422_ ( .A(_tmp_223), .B(4'h0), .S(_06437_), .Y(_27841_) );
  \$mux  #( .WIDTH(4) ) _52423_ ( .A(_27841_), .B(_24244_[3:0]), .S(_06438_), .Y(_27842_) );
  \$mux  #( .WIDTH(4) ) _52424_ ( .A(_27842_), .B(4'h0), .S(_06439_), .Y(_27843_) );
  \$mux  #( .WIDTH(4) ) _52425_ ( .A(_27843_), .B(4'h0), .S(RST), .Y(_03010_) );
  \$mux  #( .WIDTH(10) ) _52426_ ( .A(_tmp_204), .B(_28537_[9:0]), .S(_06437_), .Y(_27844_) );
  \$mux  #( .WIDTH(10) ) _52427_ ( .A(_27844_), .B(_tmp_213), .S(_06448_), .Y(_27845_) );
  \$mux  #( .WIDTH(10) ) _52428_ ( .A(_27845_), .B(10'h000), .S(RST), .Y(_03008_) );
  \$mux  #( .WIDTH(10) ) _52429_ ( .A(_tmp_203), .B(_28537_[9:0]), .S(_06437_), .Y(_27846_) );
  \$mux  #( .WIDTH(10) ) _52430_ ( .A(_27846_), .B(_tmp_212), .S(_06447_), .Y(_27847_) );
  \$mux  #( .WIDTH(10) ) _52431_ ( .A(_27847_), .B(10'h000), .S(RST), .Y(_03007_) );
  \$mux  #( .WIDTH(10) ) _52432_ ( .A(_tmp_202), .B(_28537_[9:0]), .S(_06437_), .Y(_27848_) );
  \$mux  #( .WIDTH(10) ) _52433_ ( .A(_27848_), .B(_tmp_211), .S(_06446_), .Y(_27849_) );
  \$mux  #( .WIDTH(10) ) _52434_ ( .A(_27849_), .B(10'h000), .S(RST), .Y(_03006_) );
  \$mux  #( .WIDTH(10) ) _52435_ ( .A(_tmp_201), .B(_28537_[9:0]), .S(_06437_), .Y(_27850_) );
  \$mux  #( .WIDTH(10) ) _52436_ ( .A(_27850_), .B(_tmp_210), .S(_06445_), .Y(_27851_) );
  \$mux  #( .WIDTH(10) ) _52437_ ( .A(_27851_), .B(10'h000), .S(RST), .Y(_03005_) );
  \$mux  #( .WIDTH(10) ) _52438_ ( .A(_tmp_200), .B(_28537_[9:0]), .S(_06437_), .Y(_27852_) );
  \$mux  #( .WIDTH(10) ) _52439_ ( .A(_27852_), .B(_tmp_209), .S(_06444_), .Y(_27853_) );
  \$mux  #( .WIDTH(10) ) _52440_ ( .A(_27853_), .B(10'h000), .S(RST), .Y(_03004_) );
  \$mux  #( .WIDTH(10) ) _52441_ ( .A(_tmp_199), .B(_28537_[9:0]), .S(_06437_), .Y(_27854_) );
  \$mux  #( .WIDTH(10) ) _52442_ ( .A(_27854_), .B(_tmp_208), .S(_06443_), .Y(_27855_) );
  \$mux  #( .WIDTH(10) ) _52443_ ( .A(_27855_), .B(10'h000), .S(RST), .Y(_03001_) );
  \$mux  #( .WIDTH(10) ) _52444_ ( .A(_tmp_198), .B(_28537_[9:0]), .S(_06437_), .Y(_27856_) );
  \$mux  #( .WIDTH(10) ) _52445_ ( .A(_27856_), .B(_tmp_207), .S(_06442_), .Y(_27857_) );
  \$mux  #( .WIDTH(10) ) _52446_ ( .A(_27857_), .B(10'h000), .S(RST), .Y(_03000_) );
  \$mux  #( .WIDTH(10) ) _52447_ ( .A(_tmp_197), .B(_28537_[9:0]), .S(_06437_), .Y(_27858_) );
  \$mux  #( .WIDTH(10) ) _52448_ ( .A(_27858_), .B(_tmp_206), .S(_06441_), .Y(_27859_) );
  \$mux  #( .WIDTH(10) ) _52449_ ( .A(_27859_), .B(10'h000), .S(RST), .Y(_02999_) );
  \$mux  #( .WIDTH(10) ) _52450_ ( .A(_tmp_196), .B(_28537_[9:0]), .S(_06437_), .Y(_27860_) );
  \$mux  #( .WIDTH(10) ) _52451_ ( .A(_27860_), .B(_tmp_205), .S(_06440_), .Y(_27861_) );
  \$mux  #( .WIDTH(10) ) _52452_ ( .A(_27861_), .B(10'h000), .S(RST), .Y(_02998_) );
  \$mux  #( .WIDTH(1) ) _52453_ ( .A(_tmp_195), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27862_) );
  \$mux  #( .WIDTH(1) ) _52454_ ( .A(_27862_), .B(1'h1), .S(_06449_), .Y(_27863_) );
  \$mux  #( .WIDTH(1) ) _52455_ ( .A(_27863_), .B(1'h0), .S(RST), .Y(_02997_) );
  \$mux  #( .WIDTH(34) ) _52456_ ( .A(_tmp_194), .B({ 1'h0, _maxi_read_size }), .S(_06437_), .Y(_27864_) );
  \$mux  #( .WIDTH(34) ) _52457_ ( .A(_27864_), .B(_28554_), .S(_06235_), .Y(_27865_) );
  \$mux  #( .WIDTH(34) ) _52458_ ( .A(_27865_), .B(34'h000000000), .S(RST), .Y(_02996_) );
  \$mux  #( .WIDTH(11) ) _52459_ ( .A(_tmp_193), .B(_28536_[10:0]), .S(_06437_), .Y(_27866_) );
  \$mux  #( .WIDTH(11) ) _52460_ ( .A(_27866_), .B(_28553_[10:0]), .S(_06235_), .Y(_27867_) );
  \$mux  #( .WIDTH(11) ) _52461_ ( .A(_27867_), .B(_28536_[10:0]), .S(_06438_), .Y(_27868_) );
  \$mux  #( .WIDTH(11) ) _52462_ ( .A(_27868_), .B(11'h000), .S(RST), .Y(_02995_) );
  \$mux  #( .WIDTH(1) ) _52463_ ( .A(ram_w4_l8192_id0_5_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27869_) );
  \$mux  #( .WIDTH(1) ) _52464_ ( .A(_27869_), .B(_06073_), .S(_06235_), .Y(_27870_) );
  \$mux  #( .WIDTH(1) ) _52465_ ( .A(_27870_), .B(1'h1), .S(_06307_), .Y(_27871_) );
  \$mux  #( .WIDTH(1) ) _52466_ ( .A(_27871_), .B(1'h0), .S(RST), .Y(_03396_) );
  \$mux  #( .WIDTH(4) ) _52467_ ( .A(ram_w4_l8192_id0_5_1_wdata), .B(_dataflow_slice_data_44), .S(_06235_), .Y(_27872_) );
  \$mux  #( .WIDTH(4) ) _52468_ ( .A(_27872_), .B(_dataflow_slice_data_139), .S(_06307_), .Y(_27873_) );
  \$mux  #( .WIDTH(4) ) _52469_ ( .A(_27873_), .B(4'h0), .S(RST), .Y(_03395_) );
  \$mux  #( .WIDTH(10) ) _52470_ ( .A(ram_w4_l8192_id0_5_1_addr), .B(_tmp_205), .S(_06235_), .Y(_27874_) );
  \$mux  #( .WIDTH(10) ) _52471_ ( .A(_27874_), .B(_28537_[9:0]), .S(_06450_), .Y(_27875_) );
  \$mux  #( .WIDTH(10) ) _52472_ ( .A(_27875_), .B(_24245_[9:0]), .S(_06307_), .Y(_27876_) );
  \$mux  #( .WIDTH(10) ) _52473_ ( .A(_27876_), .B(10'h000), .S(RST), .Y(_03394_) );
  \$mux  #( .WIDTH(10) ) _52474_ ( .A(ram_w4_l8192_id0_5_0_addr), .B(_stream_conv2d_16_source_28_source_ram_raddr[12:3]), .S(_tmp_597), .Y(_27877_) );
  \$mux  #( .WIDTH(10) ) _52475_ ( .A(_27877_), .B(_stream_matmul_29_source_20_source_ram_raddr[12:3]), .S(_tmp_1223), .Y(_27878_) );
  \$mux  #( .WIDTH(10) ) _52476_ ( .A(_27878_), .B(10'h000), .S(RST), .Y(_03393_) );
  \$mux  #( .WIDTH(1) ) _52477_ ( .A(_tmp_1145), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27879_) );
  \$mux  #( .WIDTH(1) ) _52478_ ( .A(_27879_), .B(1'h1), .S(_06436_), .Y(_27880_) );
  \$mux  #( .WIDTH(1) ) _52479_ ( .A(_27880_), .B(1'h0), .S(RST), .Y(_02921_) );
  \$mux  #( .WIDTH(34) ) _52480_ ( .A(_tmp_1144), .B({ 1'h0, _maxi_read_size }), .S(_06435_), .Y(_27881_) );
  \$mux  #( .WIDTH(34) ) _52481_ ( .A(_27881_), .B(_28552_), .S(_06304_), .Y(_27882_) );
  \$mux  #( .WIDTH(34) ) _52482_ ( .A(_27882_), .B(34'h000000000), .S(RST), .Y(_02920_) );
  \$mux  #( .WIDTH(4) ) _52483_ ( .A(_tmp_192), .B(4'h0), .S(_06422_), .Y(_27883_) );
  \$mux  #( .WIDTH(4) ) _52484_ ( .A(_27883_), .B(_24242_[3:0]), .S(_06423_), .Y(_27884_) );
  \$mux  #( .WIDTH(4) ) _52485_ ( .A(_27884_), .B(4'h0), .S(_06424_), .Y(_27885_) );
  \$mux  #( .WIDTH(4) ) _52486_ ( .A(_27885_), .B(4'h0), .S(RST), .Y(_02994_) );
  \$mux  #( .WIDTH(10) ) _52487_ ( .A(_tmp_173), .B(_28537_[9:0]), .S(_06422_), .Y(_27886_) );
  \$mux  #( .WIDTH(10) ) _52488_ ( .A(_27886_), .B(_tmp_182), .S(_06433_), .Y(_27887_) );
  \$mux  #( .WIDTH(10) ) _52489_ ( .A(_27887_), .B(10'h000), .S(RST), .Y(_02991_) );
  \$mux  #( .WIDTH(10) ) _52490_ ( .A(_tmp_172), .B(_28537_[9:0]), .S(_06422_), .Y(_27888_) );
  \$mux  #( .WIDTH(10) ) _52491_ ( .A(_27888_), .B(_tmp_181), .S(_06432_), .Y(_27889_) );
  \$mux  #( .WIDTH(10) ) _52492_ ( .A(_27889_), .B(10'h000), .S(RST), .Y(_02990_) );
  \$mux  #( .WIDTH(10) ) _52493_ ( .A(_tmp_171), .B(_28537_[9:0]), .S(_06422_), .Y(_27890_) );
  \$mux  #( .WIDTH(10) ) _52494_ ( .A(_27890_), .B(_tmp_180), .S(_06431_), .Y(_27891_) );
  \$mux  #( .WIDTH(10) ) _52495_ ( .A(_27891_), .B(10'h000), .S(RST), .Y(_02989_) );
  \$mux  #( .WIDTH(10) ) _52496_ ( .A(_tmp_170), .B(_28537_[9:0]), .S(_06422_), .Y(_27892_) );
  \$mux  #( .WIDTH(10) ) _52497_ ( .A(_27892_), .B(_tmp_179), .S(_06430_), .Y(_27893_) );
  \$mux  #( .WIDTH(10) ) _52498_ ( .A(_27893_), .B(10'h000), .S(RST), .Y(_02988_) );
  \$mux  #( .WIDTH(10) ) _52499_ ( .A(_tmp_169), .B(_28537_[9:0]), .S(_06422_), .Y(_27894_) );
  \$mux  #( .WIDTH(10) ) _52500_ ( .A(_27894_), .B(_tmp_178), .S(_06429_), .Y(_27895_) );
  \$mux  #( .WIDTH(10) ) _52501_ ( .A(_27895_), .B(10'h000), .S(RST), .Y(_02986_) );
  \$mux  #( .WIDTH(10) ) _52502_ ( .A(_tmp_168), .B(_28537_[9:0]), .S(_06422_), .Y(_27896_) );
  \$mux  #( .WIDTH(10) ) _52503_ ( .A(_27896_), .B(_tmp_177), .S(_06428_), .Y(_27897_) );
  \$mux  #( .WIDTH(10) ) _52504_ ( .A(_27897_), .B(10'h000), .S(RST), .Y(_02985_) );
  \$mux  #( .WIDTH(10) ) _52505_ ( .A(_tmp_167), .B(_28537_[9:0]), .S(_06422_), .Y(_27898_) );
  \$mux  #( .WIDTH(10) ) _52506_ ( .A(_27898_), .B(_tmp_176), .S(_06427_), .Y(_27899_) );
  \$mux  #( .WIDTH(10) ) _52507_ ( .A(_27899_), .B(10'h000), .S(RST), .Y(_02984_) );
  \$mux  #( .WIDTH(10) ) _52508_ ( .A(_tmp_166), .B(_28537_[9:0]), .S(_06422_), .Y(_27900_) );
  \$mux  #( .WIDTH(10) ) _52509_ ( .A(_27900_), .B(_tmp_175), .S(_06426_), .Y(_27901_) );
  \$mux  #( .WIDTH(10) ) _52510_ ( .A(_27901_), .B(10'h000), .S(RST), .Y(_02983_) );
  \$mux  #( .WIDTH(10) ) _52511_ ( .A(_tmp_165), .B(_28537_[9:0]), .S(_06422_), .Y(_27902_) );
  \$mux  #( .WIDTH(10) ) _52512_ ( .A(_27902_), .B(_tmp_174), .S(_06425_), .Y(_27903_) );
  \$mux  #( .WIDTH(10) ) _52513_ ( .A(_27903_), .B(10'h000), .S(RST), .Y(_02982_) );
  \$mux  #( .WIDTH(1) ) _52514_ ( .A(_tmp_164), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27904_) );
  \$mux  #( .WIDTH(1) ) _52515_ ( .A(_27904_), .B(1'h1), .S(_06434_), .Y(_27905_) );
  \$mux  #( .WIDTH(1) ) _52516_ ( .A(_27905_), .B(1'h0), .S(RST), .Y(_02981_) );
  \$mux  #( .WIDTH(34) ) _52517_ ( .A(_tmp_163), .B({ 1'h0, _maxi_read_size }), .S(_06422_), .Y(_27906_) );
  \$mux  #( .WIDTH(34) ) _52518_ ( .A(_27906_), .B(_28551_), .S(_06232_), .Y(_27907_) );
  \$mux  #( .WIDTH(34) ) _52519_ ( .A(_27907_), .B(34'h000000000), .S(RST), .Y(_02980_) );
  \$mux  #( .WIDTH(11) ) _52520_ ( .A(_tmp_162), .B(_28536_[10:0]), .S(_06422_), .Y(_27908_) );
  \$mux  #( .WIDTH(11) ) _52521_ ( .A(_27908_), .B(_28550_[10:0]), .S(_06232_), .Y(_27909_) );
  \$mux  #( .WIDTH(11) ) _52522_ ( .A(_27909_), .B(_28536_[10:0]), .S(_06423_), .Y(_27910_) );
  \$mux  #( .WIDTH(11) ) _52523_ ( .A(_27910_), .B(11'h000), .S(RST), .Y(_02979_) );
  \$mux  #( .WIDTH(1) ) _52524_ ( .A(ram_w4_l8192_id0_4_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27911_) );
  \$mux  #( .WIDTH(1) ) _52525_ ( .A(_27911_), .B(_06064_), .S(_06232_), .Y(_27912_) );
  \$mux  #( .WIDTH(1) ) _52526_ ( .A(_27912_), .B(1'h1), .S(_06304_), .Y(_27913_) );
  \$mux  #( .WIDTH(1) ) _52527_ ( .A(_27913_), .B(1'h0), .S(RST), .Y(_03392_) );
  \$mux  #( .WIDTH(4) ) _52528_ ( .A(ram_w4_l8192_id0_4_1_wdata), .B(_dataflow_slice_data_41), .S(_06232_), .Y(_27914_) );
  \$mux  #( .WIDTH(4) ) _52529_ ( .A(_27914_), .B(_dataflow_slice_data_136), .S(_06304_), .Y(_27915_) );
  \$mux  #( .WIDTH(4) ) _52530_ ( .A(_27915_), .B(4'h0), .S(RST), .Y(_03391_) );
  \$mux  #( .WIDTH(10) ) _52531_ ( .A(ram_w4_l8192_id0_4_1_addr), .B(_tmp_174), .S(_06232_), .Y(_27916_) );
  \$mux  #( .WIDTH(10) ) _52532_ ( .A(_27916_), .B(_28537_[9:0]), .S(_06435_), .Y(_27917_) );
  \$mux  #( .WIDTH(10) ) _52533_ ( .A(_27917_), .B(_24243_[9:0]), .S(_06304_), .Y(_27918_) );
  \$mux  #( .WIDTH(10) ) _52534_ ( .A(_27918_), .B(10'h000), .S(RST), .Y(_03390_) );
  \$mux  #( .WIDTH(10) ) _52535_ ( .A(ram_w4_l8192_id0_4_0_addr), .B(_stream_conv2d_16_source_28_source_ram_raddr[12:3]), .S(_tmp_597), .Y(_27919_) );
  \$mux  #( .WIDTH(10) ) _52536_ ( .A(_27919_), .B(_stream_matmul_29_source_20_source_ram_raddr[12:3]), .S(_tmp_1223), .Y(_27920_) );
  \$mux  #( .WIDTH(10) ) _52537_ ( .A(_27920_), .B(10'h000), .S(RST), .Y(_03389_) );
  \$mux  #( .WIDTH(1) ) _52538_ ( .A(_tmp_1143), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27921_) );
  \$mux  #( .WIDTH(1) ) _52539_ ( .A(_27921_), .B(1'h1), .S(_06421_), .Y(_27922_) );
  \$mux  #( .WIDTH(1) ) _52540_ ( .A(_27922_), .B(1'h0), .S(RST), .Y(_02919_) );
  \$mux  #( .WIDTH(34) ) _52541_ ( .A(_tmp_1142), .B({ 1'h0, _maxi_read_size }), .S(_06420_), .Y(_27923_) );
  \$mux  #( .WIDTH(34) ) _52542_ ( .A(_27923_), .B(_28549_), .S(_06301_), .Y(_27924_) );
  \$mux  #( .WIDTH(34) ) _52543_ ( .A(_27924_), .B(34'h000000000), .S(RST), .Y(_02918_) );
  \$mux  #( .WIDTH(4) ) _52544_ ( .A(_tmp_161), .B(4'h0), .S(_06407_), .Y(_27925_) );
  \$mux  #( .WIDTH(4) ) _52545_ ( .A(_27925_), .B(_24240_[3:0]), .S(_06408_), .Y(_27926_) );
  \$mux  #( .WIDTH(4) ) _52546_ ( .A(_27926_), .B(4'h0), .S(_06409_), .Y(_27927_) );
  \$mux  #( .WIDTH(4) ) _52547_ ( .A(_27927_), .B(4'h0), .S(RST), .Y(_02978_) );
  \$mux  #( .WIDTH(10) ) _52548_ ( .A(_tmp_142), .B(_28537_[9:0]), .S(_06407_), .Y(_27928_) );
  \$mux  #( .WIDTH(10) ) _52549_ ( .A(_27928_), .B(_tmp_151), .S(_06418_), .Y(_27929_) );
  \$mux  #( .WIDTH(10) ) _52550_ ( .A(_27929_), .B(10'h000), .S(RST), .Y(_02975_) );
  \$mux  #( .WIDTH(10) ) _52551_ ( .A(_tmp_141), .B(_28537_[9:0]), .S(_06407_), .Y(_27930_) );
  \$mux  #( .WIDTH(10) ) _52552_ ( .A(_27930_), .B(_tmp_150), .S(_06417_), .Y(_27931_) );
  \$mux  #( .WIDTH(10) ) _52553_ ( .A(_27931_), .B(10'h000), .S(RST), .Y(_02974_) );
  \$mux  #( .WIDTH(10) ) _52554_ ( .A(_tmp_140), .B(_28537_[9:0]), .S(_06407_), .Y(_27932_) );
  \$mux  #( .WIDTH(10) ) _52555_ ( .A(_27932_), .B(_tmp_149), .S(_06416_), .Y(_27933_) );
  \$mux  #( .WIDTH(10) ) _52556_ ( .A(_27933_), .B(10'h000), .S(RST), .Y(_02973_) );
  \$mux  #( .WIDTH(10) ) _52557_ ( .A(_tmp_139), .B(_28537_[9:0]), .S(_06407_), .Y(_27934_) );
  \$mux  #( .WIDTH(10) ) _52558_ ( .A(_27934_), .B(_tmp_148), .S(_06415_), .Y(_27935_) );
  \$mux  #( .WIDTH(10) ) _52559_ ( .A(_27935_), .B(10'h000), .S(RST), .Y(_02971_) );
  \$mux  #( .WIDTH(10) ) _52560_ ( .A(_tmp_138), .B(_28537_[9:0]), .S(_06407_), .Y(_27936_) );
  \$mux  #( .WIDTH(10) ) _52561_ ( .A(_27936_), .B(_tmp_147), .S(_06414_), .Y(_27937_) );
  \$mux  #( .WIDTH(10) ) _52562_ ( .A(_27937_), .B(10'h000), .S(RST), .Y(_02970_) );
  \$mux  #( .WIDTH(10) ) _52563_ ( .A(_tmp_137), .B(_28537_[9:0]), .S(_06407_), .Y(_27938_) );
  \$mux  #( .WIDTH(10) ) _52564_ ( .A(_27938_), .B(_tmp_146), .S(_06413_), .Y(_27939_) );
  \$mux  #( .WIDTH(10) ) _52565_ ( .A(_27939_), .B(10'h000), .S(RST), .Y(_02969_) );
  \$mux  #( .WIDTH(10) ) _52566_ ( .A(_tmp_136), .B(_28537_[9:0]), .S(_06407_), .Y(_27940_) );
  \$mux  #( .WIDTH(10) ) _52567_ ( .A(_27940_), .B(_tmp_145), .S(_06412_), .Y(_27941_) );
  \$mux  #( .WIDTH(10) ) _52568_ ( .A(_27941_), .B(10'h000), .S(RST), .Y(_02968_) );
  \$mux  #( .WIDTH(10) ) _52569_ ( .A(_tmp_135), .B(_28537_[9:0]), .S(_06407_), .Y(_27942_) );
  \$mux  #( .WIDTH(10) ) _52570_ ( .A(_27942_), .B(_tmp_144), .S(_06411_), .Y(_27943_) );
  \$mux  #( .WIDTH(10) ) _52571_ ( .A(_27943_), .B(10'h000), .S(RST), .Y(_02967_) );
  \$mux  #( .WIDTH(10) ) _52572_ ( .A(_tmp_134), .B(_28537_[9:0]), .S(_06407_), .Y(_27944_) );
  \$mux  #( .WIDTH(10) ) _52573_ ( .A(_27944_), .B(_tmp_143), .S(_06410_), .Y(_27945_) );
  \$mux  #( .WIDTH(10) ) _52574_ ( .A(_27945_), .B(10'h000), .S(RST), .Y(_02960_) );
  \$mux  #( .WIDTH(1) ) _52575_ ( .A(_tmp_133), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27946_) );
  \$mux  #( .WIDTH(1) ) _52576_ ( .A(_27946_), .B(1'h1), .S(_06419_), .Y(_27947_) );
  \$mux  #( .WIDTH(1) ) _52577_ ( .A(_27947_), .B(1'h0), .S(RST), .Y(_02953_) );
  \$mux  #( .WIDTH(34) ) _52578_ ( .A(_tmp_132), .B({ 1'h0, _maxi_read_size }), .S(_06407_), .Y(_27948_) );
  \$mux  #( .WIDTH(34) ) _52579_ ( .A(_27948_), .B(_28548_), .S(_06229_), .Y(_27949_) );
  \$mux  #( .WIDTH(34) ) _52580_ ( .A(_27949_), .B(34'h000000000), .S(RST), .Y(_02948_) );
  \$mux  #( .WIDTH(11) ) _52581_ ( .A(_tmp_131), .B(_28536_[10:0]), .S(_06407_), .Y(_27950_) );
  \$mux  #( .WIDTH(11) ) _52582_ ( .A(_27950_), .B(_28547_[10:0]), .S(_06229_), .Y(_27951_) );
  \$mux  #( .WIDTH(11) ) _52583_ ( .A(_27951_), .B(_28536_[10:0]), .S(_06408_), .Y(_27952_) );
  \$mux  #( .WIDTH(11) ) _52584_ ( .A(_27952_), .B(11'h000), .S(RST), .Y(_02943_) );
  \$mux  #( .WIDTH(1) ) _52585_ ( .A(ram_w4_l8192_id0_3_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27953_) );
  \$mux  #( .WIDTH(1) ) _52586_ ( .A(_27953_), .B(_06055_), .S(_06229_), .Y(_27954_) );
  \$mux  #( .WIDTH(1) ) _52587_ ( .A(_27954_), .B(1'h1), .S(_06301_), .Y(_27955_) );
  \$mux  #( .WIDTH(1) ) _52588_ ( .A(_27955_), .B(1'h0), .S(RST), .Y(_03388_) );
  \$mux  #( .WIDTH(4) ) _52589_ ( .A(ram_w4_l8192_id0_3_1_wdata), .B(_dataflow_slice_data_38), .S(_06229_), .Y(_27956_) );
  \$mux  #( .WIDTH(4) ) _52590_ ( .A(_27956_), .B(_dataflow_slice_data_133), .S(_06301_), .Y(_27957_) );
  \$mux  #( .WIDTH(4) ) _52591_ ( .A(_27957_), .B(4'h0), .S(RST), .Y(_03387_) );
  \$mux  #( .WIDTH(10) ) _52592_ ( .A(ram_w4_l8192_id0_3_1_addr), .B(_tmp_143), .S(_06229_), .Y(_27958_) );
  \$mux  #( .WIDTH(10) ) _52593_ ( .A(_27958_), .B(_28537_[9:0]), .S(_06420_), .Y(_27959_) );
  \$mux  #( .WIDTH(10) ) _52594_ ( .A(_27959_), .B(_24241_[9:0]), .S(_06301_), .Y(_27960_) );
  \$mux  #( .WIDTH(10) ) _52595_ ( .A(_27960_), .B(10'h000), .S(RST), .Y(_03386_) );
  \$mux  #( .WIDTH(10) ) _52596_ ( .A(ram_w4_l8192_id0_3_0_addr), .B(_stream_conv2d_16_source_28_source_ram_raddr[12:3]), .S(_tmp_597), .Y(_27961_) );
  \$mux  #( .WIDTH(10) ) _52597_ ( .A(_27961_), .B(_stream_matmul_29_source_20_source_ram_raddr[12:3]), .S(_tmp_1223), .Y(_27962_) );
  \$mux  #( .WIDTH(10) ) _52598_ ( .A(_27962_), .B(10'h000), .S(RST), .Y(_03385_) );
  \$mux  #( .WIDTH(1) ) _52599_ ( .A(_tmp_1141), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27963_) );
  \$mux  #( .WIDTH(1) ) _52600_ ( .A(_27963_), .B(1'h1), .S(_06406_), .Y(_27964_) );
  \$mux  #( .WIDTH(1) ) _52601_ ( .A(_27964_), .B(1'h0), .S(RST), .Y(_02917_) );
  \$mux  #( .WIDTH(34) ) _52602_ ( .A(_tmp_1140), .B({ 1'h0, _maxi_read_size }), .S(_06405_), .Y(_27965_) );
  \$mux  #( .WIDTH(34) ) _52603_ ( .A(_27965_), .B(_28546_), .S(_06298_), .Y(_27966_) );
  \$mux  #( .WIDTH(34) ) _52604_ ( .A(_27966_), .B(34'h000000000), .S(RST), .Y(_02916_) );
  \$mux  #( .WIDTH(4) ) _52605_ ( .A(_tmp_130), .B(4'h0), .S(_06392_), .Y(_27967_) );
  \$mux  #( .WIDTH(4) ) _52606_ ( .A(_27967_), .B(_24238_[3:0]), .S(_06393_), .Y(_27968_) );
  \$mux  #( .WIDTH(4) ) _52607_ ( .A(_27968_), .B(4'h0), .S(_06394_), .Y(_27969_) );
  \$mux  #( .WIDTH(4) ) _52608_ ( .A(_27969_), .B(4'h0), .S(RST), .Y(_02938_) );
  \$mux  #( .WIDTH(10) ) _52609_ ( .A(_tmp_111), .B(_28537_[9:0]), .S(_06392_), .Y(_27970_) );
  \$mux  #( .WIDTH(10) ) _52610_ ( .A(_27970_), .B(_tmp_120), .S(_06403_), .Y(_27971_) );
  \$mux  #( .WIDTH(10) ) _52611_ ( .A(_27971_), .B(10'h000), .S(RST), .Y(_02902_) );
  \$mux  #( .WIDTH(10) ) _52612_ ( .A(_tmp_110), .B(_28537_[9:0]), .S(_06392_), .Y(_27972_) );
  \$mux  #( .WIDTH(10) ) _52613_ ( .A(_27972_), .B(_tmp_119), .S(_06402_), .Y(_27973_) );
  \$mux  #( .WIDTH(10) ) _52614_ ( .A(_27973_), .B(10'h000), .S(RST), .Y(_02896_) );
  \$mux  #( .WIDTH(10) ) _52615_ ( .A(_tmp_109), .B(_28537_[9:0]), .S(_06392_), .Y(_27974_) );
  \$mux  #( .WIDTH(10) ) _52616_ ( .A(_27974_), .B(_tmp_118), .S(_06401_), .Y(_27975_) );
  \$mux  #( .WIDTH(10) ) _52617_ ( .A(_27975_), .B(10'h000), .S(RST), .Y(_02889_) );
  \$mux  #( .WIDTH(10) ) _52618_ ( .A(_tmp_108), .B(_28537_[9:0]), .S(_06392_), .Y(_27976_) );
  \$mux  #( .WIDTH(10) ) _52619_ ( .A(_27976_), .B(_tmp_117), .S(_06400_), .Y(_27977_) );
  \$mux  #( .WIDTH(10) ) _52620_ ( .A(_27977_), .B(10'h000), .S(RST), .Y(_02882_) );
  \$mux  #( .WIDTH(10) ) _52621_ ( .A(_tmp_107), .B(_28537_[9:0]), .S(_06392_), .Y(_27978_) );
  \$mux  #( .WIDTH(10) ) _52622_ ( .A(_27978_), .B(_tmp_116), .S(_06399_), .Y(_27979_) );
  \$mux  #( .WIDTH(10) ) _52623_ ( .A(_27979_), .B(10'h000), .S(RST), .Y(_02876_) );
  \$mux  #( .WIDTH(10) ) _52624_ ( .A(_tmp_106), .B(_28537_[9:0]), .S(_06392_), .Y(_27980_) );
  \$mux  #( .WIDTH(10) ) _52625_ ( .A(_27980_), .B(_tmp_115), .S(_06398_), .Y(_27981_) );
  \$mux  #( .WIDTH(10) ) _52626_ ( .A(_27981_), .B(10'h000), .S(RST), .Y(_02873_) );
  \$mux  #( .WIDTH(10) ) _52627_ ( .A(_tmp_105), .B(_28537_[9:0]), .S(_06392_), .Y(_27982_) );
  \$mux  #( .WIDTH(10) ) _52628_ ( .A(_27982_), .B(_tmp_114), .S(_06397_), .Y(_27983_) );
  \$mux  #( .WIDTH(10) ) _52629_ ( .A(_27983_), .B(10'h000), .S(RST), .Y(_02872_) );
  \$mux  #( .WIDTH(10) ) _52630_ ( .A(_tmp_104), .B(_28537_[9:0]), .S(_06392_), .Y(_27984_) );
  \$mux  #( .WIDTH(10) ) _52631_ ( .A(_27984_), .B(_tmp_113), .S(_06396_), .Y(_27985_) );
  \$mux  #( .WIDTH(10) ) _52632_ ( .A(_27985_), .B(10'h000), .S(RST), .Y(_02871_) );
  \$mux  #( .WIDTH(10) ) _52633_ ( .A(_tmp_103), .B(_28537_[9:0]), .S(_06392_), .Y(_27986_) );
  \$mux  #( .WIDTH(10) ) _52634_ ( .A(_27986_), .B(_tmp_112), .S(_06395_), .Y(_27987_) );
  \$mux  #( .WIDTH(10) ) _52635_ ( .A(_27987_), .B(10'h000), .S(RST), .Y(_02870_) );
  \$mux  #( .WIDTH(1) ) _52636_ ( .A(_tmp_102), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27988_) );
  \$mux  #( .WIDTH(1) ) _52637_ ( .A(_27988_), .B(1'h1), .S(_06404_), .Y(_27989_) );
  \$mux  #( .WIDTH(1) ) _52638_ ( .A(_27989_), .B(1'h0), .S(RST), .Y(_02869_) );
  \$mux  #( .WIDTH(34) ) _52639_ ( .A(_tmp_101), .B({ 1'h0, _maxi_read_size }), .S(_06392_), .Y(_27990_) );
  \$mux  #( .WIDTH(34) ) _52640_ ( .A(_27990_), .B(_28545_), .S(_06226_), .Y(_27991_) );
  \$mux  #( .WIDTH(34) ) _52641_ ( .A(_27991_), .B(34'h000000000), .S(RST), .Y(_02867_) );
  \$mux  #( .WIDTH(11) ) _52642_ ( .A(_tmp_100), .B(_28536_[10:0]), .S(_06392_), .Y(_27992_) );
  \$mux  #( .WIDTH(11) ) _52643_ ( .A(_27992_), .B(_28544_[10:0]), .S(_06226_), .Y(_27993_) );
  \$mux  #( .WIDTH(11) ) _52644_ ( .A(_27993_), .B(_28536_[10:0]), .S(_06393_), .Y(_27994_) );
  \$mux  #( .WIDTH(11) ) _52645_ ( .A(_27994_), .B(11'h000), .S(RST), .Y(_02860_) );
  \$mux  #( .WIDTH(1) ) _52646_ ( .A(ram_w4_l8192_id0_2_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_27995_) );
  \$mux  #( .WIDTH(1) ) _52647_ ( .A(_27995_), .B(_06046_), .S(_06226_), .Y(_27996_) );
  \$mux  #( .WIDTH(1) ) _52648_ ( .A(_27996_), .B(1'h1), .S(_06298_), .Y(_27997_) );
  \$mux  #( .WIDTH(1) ) _52649_ ( .A(_27997_), .B(1'h0), .S(RST), .Y(_03384_) );
  \$mux  #( .WIDTH(4) ) _52650_ ( .A(ram_w4_l8192_id0_2_1_wdata), .B(_dataflow_slice_data_35), .S(_06226_), .Y(_27998_) );
  \$mux  #( .WIDTH(4) ) _52651_ ( .A(_27998_), .B(_dataflow_slice_data_130), .S(_06298_), .Y(_27999_) );
  \$mux  #( .WIDTH(4) ) _52652_ ( .A(_27999_), .B(4'h0), .S(RST), .Y(_03383_) );
  \$mux  #( .WIDTH(10) ) _52653_ ( .A(ram_w4_l8192_id0_2_1_addr), .B(_tmp_112), .S(_06226_), .Y(_28000_) );
  \$mux  #( .WIDTH(10) ) _52654_ ( .A(_28000_), .B(_28537_[9:0]), .S(_06405_), .Y(_28001_) );
  \$mux  #( .WIDTH(10) ) _52655_ ( .A(_28001_), .B(_24239_[9:0]), .S(_06298_), .Y(_28002_) );
  \$mux  #( .WIDTH(10) ) _52656_ ( .A(_28002_), .B(10'h000), .S(RST), .Y(_03382_) );
  \$mux  #( .WIDTH(10) ) _52657_ ( .A(ram_w4_l8192_id0_2_0_addr), .B(_stream_conv2d_16_source_28_source_ram_raddr[12:3]), .S(_tmp_597), .Y(_28003_) );
  \$mux  #( .WIDTH(10) ) _52658_ ( .A(_28003_), .B(_stream_matmul_29_source_20_source_ram_raddr[12:3]), .S(_tmp_1223), .Y(_28004_) );
  \$mux  #( .WIDTH(10) ) _52659_ ( .A(_28004_), .B(10'h000), .S(RST), .Y(_03381_) );
  \$mux  #( .WIDTH(1) ) _52660_ ( .A(_tmp_1139), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_28005_) );
  \$mux  #( .WIDTH(1) ) _52661_ ( .A(_28005_), .B(1'h1), .S(_06391_), .Y(_28006_) );
  \$mux  #( .WIDTH(1) ) _52662_ ( .A(_28006_), .B(1'h0), .S(RST), .Y(_02915_) );
  \$mux  #( .WIDTH(34) ) _52663_ ( .A(_tmp_1138), .B({ 1'h0, _maxi_read_size }), .S(_06390_), .Y(_28007_) );
  \$mux  #( .WIDTH(34) ) _52664_ ( .A(_28007_), .B(_28543_), .S(_06295_), .Y(_28008_) );
  \$mux  #( .WIDTH(34) ) _52665_ ( .A(_28008_), .B(34'h000000000), .S(RST), .Y(_02914_) );
  \$mux  #( .WIDTH(4) ) _52666_ ( .A(_tmp_99), .B(4'h0), .S(_06377_), .Y(_28009_) );
  \$mux  #( .WIDTH(4) ) _52667_ ( .A(_28009_), .B(_24236_[3:0]), .S(_06378_), .Y(_28010_) );
  \$mux  #( .WIDTH(4) ) _52668_ ( .A(_28010_), .B(4'h0), .S(_06379_), .Y(_28011_) );
  \$mux  #( .WIDTH(4) ) _52669_ ( .A(_28011_), .B(4'h0), .S(RST), .Y(_03171_) );
  \$mux  #( .WIDTH(10) ) _52670_ ( .A(_tmp_80), .B(_28537_[9:0]), .S(_06377_), .Y(_28012_) );
  \$mux  #( .WIDTH(10) ) _52671_ ( .A(_28012_), .B(_tmp_89), .S(_06388_), .Y(_28013_) );
  \$mux  #( .WIDTH(10) ) _52672_ ( .A(_28013_), .B(10'h000), .S(RST), .Y(_03157_) );
  \$mux  #( .WIDTH(10) ) _52673_ ( .A(_tmp_79), .B(_28537_[9:0]), .S(_06377_), .Y(_28014_) );
  \$mux  #( .WIDTH(10) ) _52674_ ( .A(_28014_), .B(_tmp_88), .S(_06387_), .Y(_28015_) );
  \$mux  #( .WIDTH(10) ) _52675_ ( .A(_28015_), .B(10'h000), .S(RST), .Y(_03156_) );
  \$mux  #( .WIDTH(10) ) _52676_ ( .A(_tmp_78), .B(_28537_[9:0]), .S(_06377_), .Y(_28016_) );
  \$mux  #( .WIDTH(10) ) _52677_ ( .A(_28016_), .B(_tmp_87), .S(_06386_), .Y(_28017_) );
  \$mux  #( .WIDTH(10) ) _52678_ ( .A(_28017_), .B(10'h000), .S(RST), .Y(_03155_) );
  \$mux  #( .WIDTH(10) ) _52679_ ( .A(_tmp_77), .B(_28537_[9:0]), .S(_06377_), .Y(_28018_) );
  \$mux  #( .WIDTH(10) ) _52680_ ( .A(_28018_), .B(_tmp_86), .S(_06385_), .Y(_28019_) );
  \$mux  #( .WIDTH(10) ) _52681_ ( .A(_28019_), .B(10'h000), .S(RST), .Y(_03154_) );
  \$mux  #( .WIDTH(10) ) _52682_ ( .A(_tmp_76), .B(_28537_[9:0]), .S(_06377_), .Y(_28020_) );
  \$mux  #( .WIDTH(10) ) _52683_ ( .A(_28020_), .B(_tmp_85), .S(_06384_), .Y(_28021_) );
  \$mux  #( .WIDTH(10) ) _52684_ ( .A(_28021_), .B(10'h000), .S(RST), .Y(_03153_) );
  \$mux  #( .WIDTH(10) ) _52685_ ( .A(_tmp_75), .B(_28537_[9:0]), .S(_06377_), .Y(_28022_) );
  \$mux  #( .WIDTH(10) ) _52686_ ( .A(_28022_), .B(_tmp_84), .S(_06383_), .Y(_28023_) );
  \$mux  #( .WIDTH(10) ) _52687_ ( .A(_28023_), .B(10'h000), .S(RST), .Y(_03152_) );
  \$mux  #( .WIDTH(10) ) _52688_ ( .A(_tmp_74), .B(_28537_[9:0]), .S(_06377_), .Y(_28024_) );
  \$mux  #( .WIDTH(10) ) _52689_ ( .A(_28024_), .B(_tmp_83), .S(_06382_), .Y(_28025_) );
  \$mux  #( .WIDTH(10) ) _52690_ ( .A(_28025_), .B(10'h000), .S(RST), .Y(_03151_) );
  \$mux  #( .WIDTH(10) ) _52691_ ( .A(_tmp_73), .B(_28537_[9:0]), .S(_06377_), .Y(_28026_) );
  \$mux  #( .WIDTH(10) ) _52692_ ( .A(_28026_), .B(_tmp_82), .S(_06381_), .Y(_28027_) );
  \$mux  #( .WIDTH(10) ) _52693_ ( .A(_28027_), .B(10'h000), .S(RST), .Y(_03150_) );
  \$mux  #( .WIDTH(10) ) _52694_ ( .A(_tmp_72), .B(_28537_[9:0]), .S(_06377_), .Y(_28028_) );
  \$mux  #( .WIDTH(10) ) _52695_ ( .A(_28028_), .B(_tmp_81), .S(_06380_), .Y(_28029_) );
  \$mux  #( .WIDTH(10) ) _52696_ ( .A(_28029_), .B(10'h000), .S(RST), .Y(_03149_) );
  \$mux  #( .WIDTH(1) ) _52697_ ( .A(_tmp_71), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_28030_) );
  \$mux  #( .WIDTH(1) ) _52698_ ( .A(_28030_), .B(1'h1), .S(_06389_), .Y(_28031_) );
  \$mux  #( .WIDTH(1) ) _52699_ ( .A(_28031_), .B(1'h0), .S(RST), .Y(_03148_) );
  \$mux  #( .WIDTH(34) ) _52700_ ( .A(_tmp_70), .B({ 1'h0, _maxi_read_size }), .S(_06377_), .Y(_28032_) );
  \$mux  #( .WIDTH(34) ) _52701_ ( .A(_28032_), .B(_28542_), .S(_06223_), .Y(_28033_) );
  \$mux  #( .WIDTH(34) ) _52702_ ( .A(_28033_), .B(34'h000000000), .S(RST), .Y(_03147_) );
  \$mux  #( .WIDTH(11) ) _52703_ ( .A(_tmp_69), .B(_28536_[10:0]), .S(_06377_), .Y(_28034_) );
  \$mux  #( .WIDTH(11) ) _52704_ ( .A(_28034_), .B(_28541_[10:0]), .S(_06223_), .Y(_28035_) );
  \$mux  #( .WIDTH(11) ) _52705_ ( .A(_28035_), .B(_28536_[10:0]), .S(_06378_), .Y(_28036_) );
  \$mux  #( .WIDTH(11) ) _52706_ ( .A(_28036_), .B(11'h000), .S(RST), .Y(_03146_) );
  \$mux  #( .WIDTH(1) ) _52707_ ( .A(ram_w4_l8192_id0_1_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_28037_) );
  \$mux  #( .WIDTH(1) ) _52708_ ( .A(_28037_), .B(_06037_), .S(_06223_), .Y(_28038_) );
  \$mux  #( .WIDTH(1) ) _52709_ ( .A(_28038_), .B(1'h1), .S(_06295_), .Y(_28039_) );
  \$mux  #( .WIDTH(1) ) _52710_ ( .A(_28039_), .B(1'h0), .S(RST), .Y(_03380_) );
  \$mux  #( .WIDTH(4) ) _52711_ ( .A(ram_w4_l8192_id0_1_1_wdata), .B(_dataflow_slice_data_32), .S(_06223_), .Y(_28040_) );
  \$mux  #( .WIDTH(4) ) _52712_ ( .A(_28040_), .B(_dataflow_slice_data_127), .S(_06295_), .Y(_28041_) );
  \$mux  #( .WIDTH(4) ) _52713_ ( .A(_28041_), .B(4'h0), .S(RST), .Y(_03379_) );
  \$mux  #( .WIDTH(10) ) _52714_ ( .A(ram_w4_l8192_id0_1_1_addr), .B(_tmp_81), .S(_06223_), .Y(_28042_) );
  \$mux  #( .WIDTH(10) ) _52715_ ( .A(_28042_), .B(_28537_[9:0]), .S(_06390_), .Y(_28043_) );
  \$mux  #( .WIDTH(10) ) _52716_ ( .A(_28043_), .B(_24237_[9:0]), .S(_06295_), .Y(_28044_) );
  \$mux  #( .WIDTH(10) ) _52717_ ( .A(_28044_), .B(10'h000), .S(RST), .Y(_03378_) );
  \$mux  #( .WIDTH(10) ) _52718_ ( .A(ram_w4_l8192_id0_1_0_addr), .B(_stream_conv2d_16_source_28_source_ram_raddr[12:3]), .S(_tmp_597), .Y(_28045_) );
  \$mux  #( .WIDTH(10) ) _52719_ ( .A(_28045_), .B(_stream_matmul_29_source_20_source_ram_raddr[12:3]), .S(_tmp_1223), .Y(_28046_) );
  \$mux  #( .WIDTH(10) ) _52720_ ( .A(_28046_), .B(10'h000), .S(RST), .Y(_03377_) );
  \$mux  #( .WIDTH(1) ) _52721_ ( .A(_tmp_1137), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_28047_) );
  \$mux  #( .WIDTH(1) ) _52722_ ( .A(_28047_), .B(1'h1), .S(_06376_), .Y(_28048_) );
  \$mux  #( .WIDTH(1) ) _52723_ ( .A(_28048_), .B(1'h0), .S(RST), .Y(_02913_) );
  \$mux  #( .WIDTH(34) ) _52724_ ( .A(_tmp_1136), .B({ 1'h0, _maxi_read_size }), .S(_06375_), .Y(_28049_) );
  \$mux  #( .WIDTH(34) ) _52725_ ( .A(_28049_), .B(_28540_), .S(_06292_), .Y(_28050_) );
  \$mux  #( .WIDTH(34) ) _52726_ ( .A(_28050_), .B(34'h000000000), .S(RST), .Y(_02912_) );
  \$mux  #( .WIDTH(4) ) _52727_ ( .A(_tmp_68), .B(4'h0), .S(_06361_), .Y(_28051_) );
  \$mux  #( .WIDTH(4) ) _52728_ ( .A(_28051_), .B(_24234_[3:0]), .S(_06362_), .Y(_28052_) );
  \$mux  #( .WIDTH(4) ) _52729_ ( .A(_28052_), .B(4'h0), .S(_06363_), .Y(_28053_) );
  \$mux  #( .WIDTH(4) ) _52730_ ( .A(_28053_), .B(4'h0), .S(RST), .Y(_03145_) );
  \$mux  #( .WIDTH(10) ) _52731_ ( .A(_tmp_49), .B(_28537_[9:0]), .S(_06361_), .Y(_28054_) );
  \$mux  #( .WIDTH(10) ) _52732_ ( .A(_28054_), .B(_tmp_58), .S(_06372_), .Y(_28055_) );
  \$mux  #( .WIDTH(10) ) _52733_ ( .A(_28055_), .B(10'h000), .S(RST), .Y(_03142_) );
  \$mux  #( .WIDTH(10) ) _52734_ ( .A(_tmp_48), .B(_28537_[9:0]), .S(_06361_), .Y(_28056_) );
  \$mux  #( .WIDTH(10) ) _52735_ ( .A(_28056_), .B(_tmp_57), .S(_06371_), .Y(_28057_) );
  \$mux  #( .WIDTH(10) ) _52736_ ( .A(_28057_), .B(10'h000), .S(RST), .Y(_03141_) );
  \$mux  #( .WIDTH(10) ) _52737_ ( .A(_tmp_47), .B(_28537_[9:0]), .S(_06361_), .Y(_28058_) );
  \$mux  #( .WIDTH(10) ) _52738_ ( .A(_28058_), .B(_tmp_56), .S(_06370_), .Y(_28059_) );
  \$mux  #( .WIDTH(10) ) _52739_ ( .A(_28059_), .B(10'h000), .S(RST), .Y(_03140_) );
  \$mux  #( .WIDTH(10) ) _52740_ ( .A(_tmp_46), .B(_28537_[9:0]), .S(_06361_), .Y(_28060_) );
  \$mux  #( .WIDTH(10) ) _52741_ ( .A(_28060_), .B(_tmp_55), .S(_06369_), .Y(_28061_) );
  \$mux  #( .WIDTH(10) ) _52742_ ( .A(_28061_), .B(10'h000), .S(RST), .Y(_03139_) );
  \$mux  #( .WIDTH(10) ) _52743_ ( .A(_tmp_45), .B(_28537_[9:0]), .S(_06361_), .Y(_28062_) );
  \$mux  #( .WIDTH(10) ) _52744_ ( .A(_28062_), .B(_tmp_54), .S(_06368_), .Y(_28063_) );
  \$mux  #( .WIDTH(10) ) _52745_ ( .A(_28063_), .B(10'h000), .S(RST), .Y(_03138_) );
  \$mux  #( .WIDTH(10) ) _52746_ ( .A(_tmp_44), .B(_28537_[9:0]), .S(_06361_), .Y(_28064_) );
  \$mux  #( .WIDTH(10) ) _52747_ ( .A(_28064_), .B(_tmp_53), .S(_06367_), .Y(_28065_) );
  \$mux  #( .WIDTH(10) ) _52748_ ( .A(_28065_), .B(10'h000), .S(RST), .Y(_03136_) );
  \$mux  #( .WIDTH(10) ) _52749_ ( .A(_tmp_43), .B(_28537_[9:0]), .S(_06361_), .Y(_28066_) );
  \$mux  #( .WIDTH(10) ) _52750_ ( .A(_28066_), .B(_tmp_52), .S(_06366_), .Y(_28067_) );
  \$mux  #( .WIDTH(10) ) _52751_ ( .A(_28067_), .B(10'h000), .S(RST), .Y(_03128_) );
  \$mux  #( .WIDTH(10) ) _52752_ ( .A(_tmp_42), .B(_28537_[9:0]), .S(_06361_), .Y(_28068_) );
  \$mux  #( .WIDTH(10) ) _52753_ ( .A(_28068_), .B(_tmp_51), .S(_06365_), .Y(_28069_) );
  \$mux  #( .WIDTH(10) ) _52754_ ( .A(_28069_), .B(10'h000), .S(RST), .Y(_03120_) );
  \$mux  #( .WIDTH(10) ) _52755_ ( .A(_tmp_41), .B(_28537_[9:0]), .S(_06361_), .Y(_28070_) );
  \$mux  #( .WIDTH(10) ) _52756_ ( .A(_28070_), .B(_tmp_50), .S(_06364_), .Y(_28071_) );
  \$mux  #( .WIDTH(10) ) _52757_ ( .A(_28071_), .B(10'h000), .S(RST), .Y(_03115_) );
  \$mux  #( .WIDTH(1) ) _52758_ ( .A(_tmp_40), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_28072_) );
  \$mux  #( .WIDTH(1) ) _52759_ ( .A(_28072_), .B(1'h1), .S(_06373_), .Y(_28073_) );
  \$mux  #( .WIDTH(1) ) _52760_ ( .A(_28073_), .B(1'h0), .S(RST), .Y(_03110_) );
  \$mux  #( .WIDTH(34) ) _52761_ ( .A(_tmp_39), .B({ 1'h0, _maxi_read_size }), .S(_06361_), .Y(_28074_) );
  \$mux  #( .WIDTH(34) ) _52762_ ( .A(_28074_), .B(_28539_), .S(_06220_), .Y(_28075_) );
  \$mux  #( .WIDTH(34) ) _52763_ ( .A(_28075_), .B(34'h000000000), .S(RST), .Y(_03103_) );
  \$mux  #( .WIDTH(11) ) _52764_ ( .A(_tmp_38), .B(_28536_[10:0]), .S(_06361_), .Y(_28076_) );
  \$mux  #( .WIDTH(11) ) _52765_ ( .A(_28076_), .B(_28538_[10:0]), .S(_06220_), .Y(_28077_) );
  \$mux  #( .WIDTH(11) ) _52766_ ( .A(_28077_), .B(_28536_[10:0]), .S(_06362_), .Y(_28078_) );
  \$mux  #( .WIDTH(11) ) _52767_ ( .A(_28078_), .B(11'h000), .S(RST), .Y(_03098_) );
  \$mux  #( .WIDTH(1) ) _52768_ ( .A(ram_w4_l8192_id0_0_1_wenable), .B(1'h0), .S(_ram_w8_l2048_id0_3_cond_0_1), .Y(_28079_) );
  \$mux  #( .WIDTH(1) ) _52769_ ( .A(_28079_), .B(_06028_), .S(_06220_), .Y(_28080_) );
  \$mux  #( .WIDTH(1) ) _52770_ ( .A(_28080_), .B(1'h1), .S(_06292_), .Y(_28081_) );
  \$mux  #( .WIDTH(1) ) _52771_ ( .A(_28081_), .B(1'h0), .S(RST), .Y(_03376_) );
  \$mux  #( .WIDTH(4) ) _52772_ ( .A(ram_w4_l8192_id0_0_1_wdata), .B(_dataflow_slice_data_29), .S(_06220_), .Y(_28082_) );
  \$mux  #( .WIDTH(4) ) _52773_ ( .A(_28082_), .B(_dataflow_slice_data_124), .S(_06292_), .Y(_28083_) );
  \$mux  #( .WIDTH(4) ) _52774_ ( .A(_28083_), .B(4'h0), .S(RST), .Y(_03375_) );
  \$mux  #( .WIDTH(10) ) _52775_ ( .A(ram_w4_l8192_id0_0_1_addr), .B(_tmp_50), .S(_06220_), .Y(_28084_) );
  \$mux  #( .WIDTH(10) ) _52776_ ( .A(_28084_), .B(_28537_[9:0]), .S(_06375_), .Y(_28085_) );
  \$mux  #( .WIDTH(10) ) _52777_ ( .A(_28085_), .B(_24235_[9:0]), .S(_06292_), .Y(_28086_) );
  \$mux  #( .WIDTH(10) ) _52778_ ( .A(_28086_), .B(10'h000), .S(RST), .Y(_03374_) );
  \$mux  #( .WIDTH(10) ) _52779_ ( .A(ram_w4_l8192_id0_0_0_addr), .B(_stream_conv2d_16_source_28_source_ram_raddr[12:3]), .S(_tmp_597), .Y(_28087_) );
  \$mux  #( .WIDTH(10) ) _52780_ ( .A(_28087_), .B(_stream_matmul_29_source_20_source_ram_raddr[12:3]), .S(_tmp_1223), .Y(_28088_) );
  \$mux  #( .WIDTH(10) ) _52781_ ( .A(_28088_), .B(10'h000), .S(RST), .Y(_03373_) );
  \$mux  #( .WIDTH(4) ) _52782_ ( .A(_tmp_5), .B(_tmp_0[5:2]), .S(_06878_), .Y(_28089_) );
  \$mux  #( .WIDTH(4) ) _52783_ ( .A(_28089_), .B(_tmp_5), .S(_05688_), .Y(_28090_) );
  \$mux  #( .WIDTH(4) ) _52784_ ( .A(_28090_), .B(_tmp_5), .S(_RESETN_inv_2), .Y(_03144_) );
  \$mux  #( .WIDTH(32) ) _52785_ ( .A(_saxi_register_fsm), .B(0), .S(_06877_), .Y({ _23883_, _23882_, _23880_, _23879_, _23878_, _23877_, _23876_, _23875_, _23874_, _23873_, _23872_, _23871_, _23869_, _23868_, _23867_, _23866_, _23865_, _23864_, _23863_, _23862_, _23861_, _23860_, _23890_, _23889_, _23888_, _23887_, _23886_, _23885_, _23884_, _23881_, _23870_, _23859_ }) );
  \$mux  #( .WIDTH(32) ) _52786_ ( .A(_saxi_register_fsm), .B(1), .S(_tmp_2), .Y(_28092_) );
  \$mux  #( .WIDTH(32) ) _52787_ ( .A(_28092_), .B(2), .S(_tmp_1), .Y({ _23915_, _23914_, _23912_, _23911_, _23910_, _23909_, _23908_, _23907_, _23906_, _23905_, _23904_, _23903_, _23901_, _23900_, _23899_, _23898_, _23897_, _23896_, _23895_, _23894_, _23893_, _23892_, _23922_, _23921_, _23920_, _23919_, _23918_, _23917_, _23916_, _23913_, _23902_, _23891_ }) );
  \$mux  #( .WIDTH(32) ) _52788_ ( .A(_28091_), .B(0), .S(_RESETN_inv_2), .Y(_01869_) );
  \$mux  #( .WIDTH(1) ) _52789_ ( .A(1'h1), .B(1'h0), .S(_RESETN_inv_2), .Y(_01704_) );
  \$mux  #( .WIDTH(1) ) _52790_ ( .A(saxi_arvalid), .B(1'h0), .S(_RESETN_inv_2), .Y(_03143_) );
  \$mux  #( .WIDTH(1) ) _52791_ ( .A(saxi_awvalid), .B(1'h0), .S(_RESETN_inv_2), .Y(_03104_) );
  \$mux  #( .WIDTH(1) ) _52792_ ( .A(1'h0), .B(1'h1), .S(_06329_), .Y(_28093_) );
  \$mux  #( .WIDTH(1) ) _52793_ ( .A(_28093_), .B(1'h0), .S(_06328_), .Y(_28094_) );
  \$mux  #( .WIDTH(1) ) _52794_ ( .A(_28094_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03048_) );
  \$mux  #( .WIDTH(1) ) _52795_ ( .A(1'h0), .B(1'h1), .S(_06328_), .Y(_28095_) );
  \$mux  #( .WIDTH(1) ) _52796_ ( .A(_28095_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03003_) );
  \$mux  #( .WIDTH(6) ) _52797_ ( .A(_tmp_0), .B(saxi_araddr), .S(_06329_), .Y(_28096_) );
  \$mux  #( .WIDTH(6) ) _52798_ ( .A(_28096_), .B(saxi_awaddr), .S(_06328_), .Y(_28097_) );
  \$mux  #( .WIDTH(6) ) _52799_ ( .A(_28097_), .B(6'h00), .S(_RESETN_inv_2), .Y(_02853_) );
  \$mux  #( .WIDTH(1) ) _52800_ ( .A(_saxi_flag_13), .B(1'h0), .S(_06345_), .Y(_28098_) );
  \$mux  #( .WIDTH(1) ) _52801_ ( .A(_28098_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01845_) );
  \$mux  #( .WIDTH(1) ) _52802_ ( .A(_saxi_flag_12), .B(1'h0), .S(_06344_), .Y(_28099_) );
  \$mux  #( .WIDTH(1) ) _52803_ ( .A(_28099_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01844_) );
  \$mux  #( .WIDTH(1) ) _52804_ ( .A(_saxi_flag_11), .B(1'h0), .S(_06343_), .Y(_28100_) );
  \$mux  #( .WIDTH(1) ) _52805_ ( .A(_28100_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01843_) );
  \$mux  #( .WIDTH(1) ) _52806_ ( .A(_saxi_flag_10), .B(1'h0), .S(_06342_), .Y(_28101_) );
  \$mux  #( .WIDTH(1) ) _52807_ ( .A(_28101_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01842_) );
  \$mux  #( .WIDTH(1) ) _52808_ ( .A(_saxi_flag_9), .B(1'h0), .S(_06341_), .Y(_28102_) );
  \$mux  #( .WIDTH(1) ) _52809_ ( .A(_28102_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01854_) );
  \$mux  #( .WIDTH(1) ) _52810_ ( .A(_saxi_flag_8), .B(1'h0), .S(_06340_), .Y(_28103_) );
  \$mux  #( .WIDTH(1) ) _52811_ ( .A(_28103_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01853_) );
  \$mux  #( .WIDTH(1) ) _52812_ ( .A(_saxi_flag_7), .B(1'h0), .S(_06339_), .Y(_28104_) );
  \$mux  #( .WIDTH(1) ) _52813_ ( .A(_28104_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01852_) );
  \$mux  #( .WIDTH(1) ) _52814_ ( .A(_saxi_flag_6), .B(1'h0), .S(_06338_), .Y(_28105_) );
  \$mux  #( .WIDTH(1) ) _52815_ ( .A(_28105_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01851_) );
  \$mux  #( .WIDTH(1) ) _52816_ ( .A(_saxi_flag_5), .B(1'h0), .S(_06337_), .Y(_28106_) );
  \$mux  #( .WIDTH(1) ) _52817_ ( .A(1'h0), .B(_28106_), .S(_05743_), .Y(_28107_) );
  \$mux  #( .WIDTH(1) ) _52818_ ( .A(1'h0), .B(_28107_), .S(_06022_), .Y(_28108_) );
  \$mux  #( .WIDTH(1) ) _52819_ ( .A(_28108_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01850_) );
  \$mux  #( .WIDTH(1) ) _52820_ ( .A(_saxi_flag_4), .B(1'h0), .S(_06336_), .Y(_28109_) );
  \$mux  #( .WIDTH(1) ) _52821_ ( .A(1'h0), .B(_28109_), .S(_05742_), .Y(_28110_) );
  \$mux  #( .WIDTH(1) ) _52822_ ( .A(_28110_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01849_) );
  \$mux  #( .WIDTH(1) ) _52823_ ( .A(_saxi_flag_3), .B(1'h0), .S(_06335_), .Y(_28111_) );
  \$mux  #( .WIDTH(1) ) _52824_ ( .A(_28111_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01848_) );
  \$mux  #( .WIDTH(1) ) _52825_ ( .A(_saxi_flag_2), .B(1'h0), .S(_06334_), .Y(_28112_) );
  \$mux  #( .WIDTH(1) ) _52826_ ( .A(_28112_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01847_) );
  \$mux  #( .WIDTH(1) ) _52827_ ( .A(_saxi_flag_1), .B(1'h0), .S(_06333_), .Y(_28113_) );
  \$mux  #( .WIDTH(1) ) _52828_ ( .A(_28113_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01846_) );
  \$mux  #( .WIDTH(1) ) _52829_ ( .A(_saxi_flag_0), .B(1'h0), .S(_06332_), .Y(_28114_) );
  \$mux  #( .WIDTH(1) ) _52830_ ( .A(_28114_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01841_) );
  \$mux  #( .WIDTH(32) ) _52831_ ( .A(_saxi_register_13), .B(_tmp_8), .S(_06345_), .Y(_28115_) );
  \$mux  #( .WIDTH(32) ) _52832_ ( .A(_28115_), .B(saxi_wdata), .S(_06359_), .Y(_28116_) );
  \$mux  #( .WIDTH(32) ) _52833_ ( .A(_28116_), .B(4160), .S(_RESETN_inv_2), .Y(_01859_) );
  \$mux  #( .WIDTH(32) ) _52834_ ( .A(_saxi_register_12), .B(_tmp_8), .S(_06344_), .Y(_28117_) );
  \$mux  #( .WIDTH(32) ) _52835_ ( .A(_28117_), .B(saxi_wdata), .S(_06358_), .Y(_28118_) );
  \$mux  #( .WIDTH(32) ) _52836_ ( .A(_28118_), .B(64), .S(_RESETN_inv_2), .Y(_01858_) );
  \$mux  #( .WIDTH(32) ) _52837_ ( .A(_saxi_register_11), .B(_tmp_8), .S(_06343_), .Y(_28119_) );
  \$mux  #( .WIDTH(32) ) _52838_ ( .A(_28119_), .B(saxi_wdata), .S(_06357_), .Y(_28120_) );
  \$mux  #( .WIDTH(32) ) _52839_ ( .A(_28120_), .B(0), .S(_RESETN_inv_2), .Y(_01857_) );
  \$mux  #( .WIDTH(32) ) _52840_ ( .A(_saxi_register_10), .B(_tmp_8), .S(_06342_), .Y(_28121_) );
  \$mux  #( .WIDTH(32) ) _52841_ ( .A(_28121_), .B(saxi_wdata), .S(_06356_), .Y(_28122_) );
  \$mux  #( .WIDTH(32) ) _52842_ ( .A(_28122_), .B(165376), .S(_RESETN_inv_2), .Y(_01856_) );
  \$mux  #( .WIDTH(32) ) _52843_ ( .A(_saxi_register_9), .B(_tmp_8), .S(_06341_), .Y(_28123_) );
  \$mux  #( .WIDTH(32) ) _52844_ ( .A(_28123_), .B(saxi_wdata), .S(_06355_), .Y(_28124_) );
  \$mux  #( .WIDTH(32) ) _52845_ ( .A(_28124_), .B(0), .S(_RESETN_inv_2), .Y(_01868_) );
  \$mux  #( .WIDTH(32) ) _52846_ ( .A(_saxi_register_8), .B(_tmp_8), .S(_06340_), .Y(_28125_) );
  \$mux  #( .WIDTH(32) ) _52847_ ( .A(_28125_), .B(saxi_wdata), .S(_06354_), .Y(_28126_) );
  \$mux  #( .WIDTH(32) ) _52848_ ( .A(_28126_), .B(0), .S(_RESETN_inv_2), .Y(_01867_) );
  \$mux  #( .WIDTH(32) ) _52849_ ( .A(_saxi_register_7), .B(_tmp_8), .S(_06339_), .Y(_28127_) );
  \$mux  #( .WIDTH(32) ) _52850_ ( .A(_28127_), .B(saxi_wdata), .S(_06353_), .Y(_28128_) );
  \$mux  #( .WIDTH(32) ) _52851_ ( .A(0), .B(_28128_), .S(_05684_), .Y(_28129_) );
  \$mux  #( .WIDTH(32) ) _52852_ ( .A(_28129_), .B(0), .S(_RESETN_inv_2), .Y(_01866_) );
  \$mux  #( .WIDTH(32) ) _52853_ ( .A(_saxi_register_6), .B(_tmp_8), .S(_06338_), .Y(_28130_) );
  \$mux  #( .WIDTH(32) ) _52854_ ( .A(_28130_), .B(saxi_wdata), .S(_06352_), .Y(_28131_) );
  \$mux  #( .WIDTH(32) ) _52855_ ( .A(0), .B(_28131_), .S(_05684_), .Y(_28132_) );
  \$mux  #( .WIDTH(32) ) _52856_ ( .A(_28132_), .B(0), .S(_RESETN_inv_2), .Y(_01865_) );
  \$mux  #( .WIDTH(32) ) _52857_ ( .A(_saxi_register_5), .B(_tmp_8), .S(_06337_), .Y(_28133_) );
  \$mux  #( .WIDTH(32) ) _52858_ ( .A(_28133_), .B(saxi_wdata), .S(_06351_), .Y(_28134_) );
  \$mux  #( .WIDTH(32) ) _52859_ ( .A(0), .B(_28134_), .S(_05684_), .Y(_28135_) );
  \$mux  #( .WIDTH(32) ) _52860_ ( .A(1), .B(_28135_), .S(_05743_), .Y(_28136_) );
  \$mux  #( .WIDTH(32) ) _52861_ ( .A(0), .B(_28136_), .S(_06022_), .Y(_28137_) );
  \$mux  #( .WIDTH(32) ) _52862_ ( .A(_28137_), .B(0), .S(_RESETN_inv_2), .Y(_01864_) );
  \$mux  #( .WIDTH(32) ) _52863_ ( .A(_saxi_register_4), .B(_tmp_8), .S(_06336_), .Y(_28138_) );
  \$mux  #( .WIDTH(32) ) _52864_ ( .A(_28138_), .B(saxi_wdata), .S(_06350_), .Y(_28139_) );
  \$mux  #( .WIDTH(32) ) _52865_ ( .A(0), .B(_28139_), .S(_05742_), .Y(_28140_) );
  \$mux  #( .WIDTH(32) ) _52866_ ( .A(_28140_), .B(0), .S(_RESETN_inv_2), .Y(_01863_) );
  \$mux  #( .WIDTH(32) ) _52867_ ( .A(_saxi_register_3), .B(_tmp_8), .S(_06335_), .Y(_28141_) );
  \$mux  #( .WIDTH(32) ) _52868_ ( .A(_28141_), .B(saxi_wdata), .S(_06349_), .Y(_28142_) );
  \$mux  #( .WIDTH(32) ) _52869_ ( .A(_28142_), .B(0), .S(_RESETN_inv_2), .Y(_01862_) );
  \$mux  #( .WIDTH(32) ) _52870_ ( .A(_saxi_register_2), .B(_tmp_8), .S(_06334_), .Y(_28143_) );
  \$mux  #( .WIDTH(32) ) _52871_ ( .A(_28143_), .B(saxi_wdata), .S(_06348_), .Y(_28144_) );
  \$mux  #( .WIDTH(32) ) _52872_ ( .A(_28144_), .B(0), .S(_RESETN_inv_2), .Y(_01861_) );
  \$mux  #( .WIDTH(32) ) _52873_ ( .A(_saxi_register_1), .B(_tmp_8), .S(_06333_), .Y(_28145_) );
  \$mux  #( .WIDTH(32) ) _52874_ ( .A(_28145_), .B(saxi_wdata), .S(_06347_), .Y(_28146_) );
  \$mux  #( .WIDTH(32) ) _52875_ ( .A(_28146_), .B(0), .S(_RESETN_inv_2), .Y(_01860_) );
  \$mux  #( .WIDTH(32) ) _52876_ ( .A(_saxi_register_0), .B(_tmp_8), .S(_06332_), .Y(_28147_) );
  \$mux  #( .WIDTH(32) ) _52877_ ( .A(_28147_), .B(saxi_wdata), .S(_06346_), .Y(_28148_) );
  \$mux  #( .WIDTH(32) ) _52878_ ( .A(_28148_), .B(0), .S(_RESETN_inv_2), .Y(_01855_) );
  \$mux  #( .WIDTH(1) ) _52879_ ( .A(saxi_rvalid), .B(1'h0), .S(_saxi_cond_0_1), .Y(_28149_) );
  \$mux  #( .WIDTH(1) ) _52880_ ( .A(_28149_), .B(1'h1), .S(_06330_), .Y(_28150_) );
  \$mux  #( .WIDTH(1) ) _52881_ ( .A(_28150_), .B(saxi_rvalid), .S(_06331_), .Y(_28151_) );
  \$mux  #( .WIDTH(1) ) _52882_ ( .A(_28151_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03875_) );
  \$mux  #( .WIDTH(32) ) _52883_ ( .A(saxi_rdata), .B(_tmp_6), .S(_06330_), .Y(_28152_) );
  \$mux  #( .WIDTH(32) ) _52884_ ( .A(_28152_), .B(0), .S(_RESETN_inv_2), .Y(_03874_) );
  \$mux  #( .WIDTH(1) ) _52885_ ( .A(saxi_bvalid), .B(1'h0), .S(_06326_), .Y(_28153_) );
  \$mux  #( .WIDTH(1) ) _52886_ ( .A(_28153_), .B(1'h1), .S(_06327_), .Y(_28154_) );
  \$mux  #( .WIDTH(1) ) _52887_ ( .A(_28154_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03873_) );
  \$mux  #( .WIDTH(1) ) _52888_ ( .A(_dataflow_slice_valid_158), .B(1'h0), .S(_06325_), .Y(_28155_) );
  \$mux  #( .WIDTH(1) ) _52889_ ( .A(_28155_), .B(_wvalid_1154), .S(_06323_), .Y(_28156_) );
  \$mux  #( .WIDTH(1) ) _52890_ ( .A(_28156_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01652_) );
  \$mux  #( .WIDTH(8) ) _52891_ ( .A(_dataflow_slice_data_158), .B(_wdata_1153[31:24]), .S(_06324_), .Y(_28157_) );
  \$mux  #( .WIDTH(8) ) _52892_ ( .A(_28157_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01608_) );
  \$mux  #( .WIDTH(1) ) _52893_ ( .A(_dataflow_slice_valid_155), .B(1'h0), .S(_06322_), .Y(_28158_) );
  \$mux  #( .WIDTH(1) ) _52894_ ( .A(_28158_), .B(_wvalid_1154), .S(_06320_), .Y(_28159_) );
  \$mux  #( .WIDTH(1) ) _52895_ ( .A(_28159_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01651_) );
  \$mux  #( .WIDTH(8) ) _52896_ ( .A(_dataflow_slice_data_155), .B(_wdata_1153[23:16]), .S(_06321_), .Y(_28160_) );
  \$mux  #( .WIDTH(8) ) _52897_ ( .A(_28160_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01607_) );
  \$mux  #( .WIDTH(1) ) _52898_ ( .A(_dataflow_slice_valid_152), .B(1'h0), .S(_06319_), .Y(_28161_) );
  \$mux  #( .WIDTH(1) ) _52899_ ( .A(_28161_), .B(_wvalid_1154), .S(_06317_), .Y(_28162_) );
  \$mux  #( .WIDTH(1) ) _52900_ ( .A(_28162_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01650_) );
  \$mux  #( .WIDTH(8) ) _52901_ ( .A(_dataflow_slice_data_152), .B(_wdata_1153[15:8]), .S(_06318_), .Y(_28163_) );
  \$mux  #( .WIDTH(8) ) _52902_ ( .A(_28163_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01606_) );
  \$mux  #( .WIDTH(1) ) _52903_ ( .A(_dataflow_slice_valid_149), .B(1'h0), .S(_06316_), .Y(_28164_) );
  \$mux  #( .WIDTH(1) ) _52904_ ( .A(_28164_), .B(_wvalid_1154), .S(_06314_), .Y(_28165_) );
  \$mux  #( .WIDTH(1) ) _52905_ ( .A(_28165_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01649_) );
  \$mux  #( .WIDTH(8) ) _52906_ ( .A(_dataflow_slice_data_149), .B(_wdata_1153[7:0]), .S(_06315_), .Y(_28166_) );
  \$mux  #( .WIDTH(8) ) _52907_ ( .A(_28166_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01605_) );
  \$mux  #( .WIDTH(1) ) _52908_ ( .A(_dataflow_slice_valid_145), .B(1'h0), .S(_06313_), .Y(_28167_) );
  \$mux  #( .WIDTH(1) ) _52909_ ( .A(_28167_), .B(_wvalid_1135), .S(_06311_), .Y(_28168_) );
  \$mux  #( .WIDTH(1) ) _52910_ ( .A(_28168_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01648_) );
  \$mux  #( .WIDTH(4) ) _52911_ ( .A(_dataflow_slice_data_145), .B(_wdata_1134[31:28]), .S(_06312_), .Y(_28169_) );
  \$mux  #( .WIDTH(4) ) _52912_ ( .A(_28169_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01604_) );
  \$mux  #( .WIDTH(1) ) _52913_ ( .A(_dataflow_slice_valid_142), .B(1'h0), .S(_06310_), .Y(_28170_) );
  \$mux  #( .WIDTH(1) ) _52914_ ( .A(_28170_), .B(_wvalid_1135), .S(_06308_), .Y(_28171_) );
  \$mux  #( .WIDTH(1) ) _52915_ ( .A(_28171_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01647_) );
  \$mux  #( .WIDTH(4) ) _52916_ ( .A(_dataflow_slice_data_142), .B(_wdata_1134[27:24]), .S(_06309_), .Y(_28172_) );
  \$mux  #( .WIDTH(4) ) _52917_ ( .A(_28172_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01603_) );
  \$mux  #( .WIDTH(1) ) _52918_ ( .A(_dataflow_slice_valid_139), .B(1'h0), .S(_06307_), .Y(_28173_) );
  \$mux  #( .WIDTH(1) ) _52919_ ( .A(_28173_), .B(_wvalid_1135), .S(_06305_), .Y(_28174_) );
  \$mux  #( .WIDTH(1) ) _52920_ ( .A(_28174_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01646_) );
  \$mux  #( .WIDTH(4) ) _52921_ ( .A(_dataflow_slice_data_139), .B(_wdata_1134[23:20]), .S(_06306_), .Y(_28175_) );
  \$mux  #( .WIDTH(4) ) _52922_ ( .A(_28175_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01602_) );
  \$mux  #( .WIDTH(1) ) _52923_ ( .A(_dataflow_slice_valid_136), .B(1'h0), .S(_06304_), .Y(_28176_) );
  \$mux  #( .WIDTH(1) ) _52924_ ( .A(_28176_), .B(_wvalid_1135), .S(_06302_), .Y(_28177_) );
  \$mux  #( .WIDTH(1) ) _52925_ ( .A(_28177_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01645_) );
  \$mux  #( .WIDTH(4) ) _52926_ ( .A(_dataflow_slice_data_136), .B(_wdata_1134[19:16]), .S(_06303_), .Y(_28178_) );
  \$mux  #( .WIDTH(4) ) _52927_ ( .A(_28178_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01601_) );
  \$mux  #( .WIDTH(1) ) _52928_ ( .A(_dataflow_slice_valid_133), .B(1'h0), .S(_06301_), .Y(_28179_) );
  \$mux  #( .WIDTH(1) ) _52929_ ( .A(_28179_), .B(_wvalid_1135), .S(_06299_), .Y(_28180_) );
  \$mux  #( .WIDTH(1) ) _52930_ ( .A(_28180_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01644_) );
  \$mux  #( .WIDTH(4) ) _52931_ ( .A(_dataflow_slice_data_133), .B(_wdata_1134[15:12]), .S(_06300_), .Y(_28181_) );
  \$mux  #( .WIDTH(4) ) _52932_ ( .A(_28181_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01600_) );
  \$mux  #( .WIDTH(1) ) _52933_ ( .A(_dataflow_slice_valid_130), .B(1'h0), .S(_06298_), .Y(_28182_) );
  \$mux  #( .WIDTH(1) ) _52934_ ( .A(_28182_), .B(_wvalid_1135), .S(_06296_), .Y(_28183_) );
  \$mux  #( .WIDTH(1) ) _52935_ ( .A(_28183_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01643_) );
  \$mux  #( .WIDTH(4) ) _52936_ ( .A(_dataflow_slice_data_130), .B(_wdata_1134[11:8]), .S(_06297_), .Y(_28184_) );
  \$mux  #( .WIDTH(4) ) _52937_ ( .A(_28184_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01599_) );
  \$mux  #( .WIDTH(1) ) _52938_ ( .A(_dataflow_slice_valid_127), .B(1'h0), .S(_06295_), .Y(_28185_) );
  \$mux  #( .WIDTH(1) ) _52939_ ( .A(_28185_), .B(_wvalid_1135), .S(_06293_), .Y(_28186_) );
  \$mux  #( .WIDTH(1) ) _52940_ ( .A(_28186_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01641_) );
  \$mux  #( .WIDTH(4) ) _52941_ ( .A(_dataflow_slice_data_127), .B(_wdata_1134[7:4]), .S(_06294_), .Y(_28187_) );
  \$mux  #( .WIDTH(4) ) _52942_ ( .A(_28187_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01597_) );
  \$mux  #( .WIDTH(1) ) _52943_ ( .A(_dataflow_slice_valid_124), .B(1'h0), .S(_06292_), .Y(_28188_) );
  \$mux  #( .WIDTH(1) ) _52944_ ( .A(_28188_), .B(_wvalid_1135), .S(_06290_), .Y(_28189_) );
  \$mux  #( .WIDTH(1) ) _52945_ ( .A(_28189_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01640_) );
  \$mux  #( .WIDTH(4) ) _52946_ ( .A(_dataflow_slice_data_124), .B(_wdata_1134[3:0]), .S(_06291_), .Y(_28190_) );
  \$mux  #( .WIDTH(4) ) _52947_ ( .A(_28190_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01596_) );
  \$mux  #( .WIDTH(1) ) _52948_ ( .A(_dataflow_slice_valid_120), .B(1'h0), .S(_06289_), .Y(_28191_) );
  \$mux  #( .WIDTH(1) ) _52949_ ( .A(_28191_), .B(_wvalid_1123), .S(_06287_), .Y(_28192_) );
  \$mux  #( .WIDTH(1) ) _52950_ ( .A(_28192_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01639_) );
  \$mux  #( .WIDTH(8) ) _52951_ ( .A(_dataflow_slice_data_120), .B(_wdata_1122[31:24]), .S(_06288_), .Y(_28193_) );
  \$mux  #( .WIDTH(8) ) _52952_ ( .A(_28193_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01595_) );
  \$mux  #( .WIDTH(1) ) _52953_ ( .A(_dataflow_slice_valid_117), .B(1'h0), .S(_06286_), .Y(_28194_) );
  \$mux  #( .WIDTH(1) ) _52954_ ( .A(_28194_), .B(_wvalid_1123), .S(_06284_), .Y(_28195_) );
  \$mux  #( .WIDTH(1) ) _52955_ ( .A(_28195_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01638_) );
  \$mux  #( .WIDTH(8) ) _52956_ ( .A(_dataflow_slice_data_117), .B(_wdata_1122[23:16]), .S(_06285_), .Y(_28196_) );
  \$mux  #( .WIDTH(8) ) _52957_ ( .A(_28196_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01594_) );
  \$mux  #( .WIDTH(1) ) _52958_ ( .A(_dataflow_slice_valid_114), .B(1'h0), .S(_06283_), .Y(_28197_) );
  \$mux  #( .WIDTH(1) ) _52959_ ( .A(_28197_), .B(_wvalid_1123), .S(_06281_), .Y(_28198_) );
  \$mux  #( .WIDTH(1) ) _52960_ ( .A(_28198_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01637_) );
  \$mux  #( .WIDTH(8) ) _52961_ ( .A(_dataflow_slice_data_114), .B(_wdata_1122[15:8]), .S(_06282_), .Y(_28199_) );
  \$mux  #( .WIDTH(8) ) _52962_ ( .A(_28199_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01593_) );
  \$mux  #( .WIDTH(1) ) _52963_ ( .A(_dataflow_slice_valid_111), .B(1'h0), .S(_06280_), .Y(_28200_) );
  \$mux  #( .WIDTH(1) ) _52964_ ( .A(_28200_), .B(_wvalid_1123), .S(_06278_), .Y(_28201_) );
  \$mux  #( .WIDTH(1) ) _52965_ ( .A(_28201_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01636_) );
  \$mux  #( .WIDTH(8) ) _52966_ ( .A(_dataflow_slice_data_111), .B(_wdata_1122[7:0]), .S(_06279_), .Y(_28202_) );
  \$mux  #( .WIDTH(8) ) _52967_ ( .A(_28202_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01592_) );
  \$mux  #( .WIDTH(1) ) _52968_ ( .A(_dataflow_slice_valid_89), .B(1'h0), .S(_06277_), .Y(_28203_) );
  \$mux  #( .WIDTH(1) ) _52969_ ( .A(_28203_), .B(_wvalid_404), .S(_06275_), .Y(_28204_) );
  \$mux  #( .WIDTH(1) ) _52970_ ( .A(_28204_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01678_) );
  \$mux  #( .WIDTH(8) ) _52971_ ( .A(_dataflow_slice_data_89), .B(_wdata_403[31:24]), .S(_06276_), .Y(_28205_) );
  \$mux  #( .WIDTH(8) ) _52972_ ( .A(_28205_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01634_) );
  \$mux  #( .WIDTH(1) ) _52973_ ( .A(_dataflow_slice_valid_86), .B(1'h0), .S(_06274_), .Y(_28206_) );
  \$mux  #( .WIDTH(1) ) _52974_ ( .A(_28206_), .B(_wvalid_404), .S(_06272_), .Y(_28207_) );
  \$mux  #( .WIDTH(1) ) _52975_ ( .A(_28207_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01677_) );
  \$mux  #( .WIDTH(8) ) _52976_ ( .A(_dataflow_slice_data_86), .B(_wdata_403[23:16]), .S(_06273_), .Y(_28208_) );
  \$mux  #( .WIDTH(8) ) _52977_ ( .A(_28208_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01633_) );
  \$mux  #( .WIDTH(1) ) _52978_ ( .A(_dataflow_slice_valid_83), .B(1'h0), .S(_06271_), .Y(_28209_) );
  \$mux  #( .WIDTH(1) ) _52979_ ( .A(_28209_), .B(_wvalid_404), .S(_06269_), .Y(_28210_) );
  \$mux  #( .WIDTH(1) ) _52980_ ( .A(_28210_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01676_) );
  \$mux  #( .WIDTH(8) ) _52981_ ( .A(_dataflow_slice_data_83), .B(_wdata_403[15:8]), .S(_06270_), .Y(_28211_) );
  \$mux  #( .WIDTH(8) ) _52982_ ( .A(_28211_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01632_) );
  \$mux  #( .WIDTH(1) ) _52983_ ( .A(_dataflow_slice_valid_80), .B(1'h0), .S(_06268_), .Y(_28212_) );
  \$mux  #( .WIDTH(1) ) _52984_ ( .A(_28212_), .B(_wvalid_404), .S(_06266_), .Y(_28213_) );
  \$mux  #( .WIDTH(1) ) _52985_ ( .A(_28213_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01675_) );
  \$mux  #( .WIDTH(8) ) _52986_ ( .A(_dataflow_slice_data_80), .B(_wdata_403[7:0]), .S(_06267_), .Y(_28214_) );
  \$mux  #( .WIDTH(8) ) _52987_ ( .A(_28214_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01631_) );
  \$mux  #( .WIDTH(1) ) _52988_ ( .A(_dataflow_slice_valid_76), .B(1'h0), .S(_06265_), .Y(_28215_) );
  \$mux  #( .WIDTH(1) ) _52989_ ( .A(_28215_), .B(_wvalid_347), .S(_06263_), .Y(_28216_) );
  \$mux  #( .WIDTH(1) ) _52990_ ( .A(_28216_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01674_) );
  \$mux  #( .WIDTH(8) ) _52991_ ( .A(_dataflow_slice_data_76), .B(_wdata_346[31:24]), .S(_06264_), .Y(_28217_) );
  \$mux  #( .WIDTH(8) ) _52992_ ( .A(_28217_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01630_) );
  \$mux  #( .WIDTH(1) ) _52993_ ( .A(_dataflow_slice_valid_73), .B(1'h0), .S(_06262_), .Y(_28218_) );
  \$mux  #( .WIDTH(1) ) _52994_ ( .A(_28218_), .B(_wvalid_347), .S(_06260_), .Y(_28219_) );
  \$mux  #( .WIDTH(1) ) _52995_ ( .A(_28219_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01673_) );
  \$mux  #( .WIDTH(8) ) _52996_ ( .A(_dataflow_slice_data_73), .B(_wdata_346[23:16]), .S(_06261_), .Y(_28220_) );
  \$mux  #( .WIDTH(8) ) _52997_ ( .A(_28220_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01629_) );
  \$mux  #( .WIDTH(1) ) _52998_ ( .A(_dataflow_slice_valid_70), .B(1'h0), .S(_06259_), .Y(_28221_) );
  \$mux  #( .WIDTH(1) ) _52999_ ( .A(_28221_), .B(_wvalid_347), .S(_06257_), .Y(_28222_) );
  \$mux  #( .WIDTH(1) ) _53000_ ( .A(_28222_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01672_) );
  \$mux  #( .WIDTH(8) ) _53001_ ( .A(_dataflow_slice_data_70), .B(_wdata_346[15:8]), .S(_06258_), .Y(_28223_) );
  \$mux  #( .WIDTH(8) ) _53002_ ( .A(_28223_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01628_) );
  \$mux  #( .WIDTH(1) ) _53003_ ( .A(_dataflow_slice_valid_67), .B(1'h0), .S(_06256_), .Y(_28224_) );
  \$mux  #( .WIDTH(1) ) _53004_ ( .A(_28224_), .B(_wvalid_347), .S(_06254_), .Y(_28225_) );
  \$mux  #( .WIDTH(1) ) _53005_ ( .A(_28225_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01670_) );
  \$mux  #( .WIDTH(8) ) _53006_ ( .A(_dataflow_slice_data_67), .B(_wdata_346[7:0]), .S(_06255_), .Y(_28226_) );
  \$mux  #( .WIDTH(8) ) _53007_ ( .A(_28226_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01626_) );
  \$mux  #( .WIDTH(1) ) _53008_ ( .A(_dataflow_slice_valid_63), .B(1'h0), .S(_06253_), .Y(_28227_) );
  \$mux  #( .WIDTH(1) ) _53009_ ( .A(_28227_), .B(_wvalid_290), .S(_06251_), .Y(_28228_) );
  \$mux  #( .WIDTH(1) ) _53010_ ( .A(_28228_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01669_) );
  \$mux  #( .WIDTH(8) ) _53011_ ( .A(_dataflow_slice_data_63), .B(_wdata_289[31:24]), .S(_06252_), .Y(_28229_) );
  \$mux  #( .WIDTH(8) ) _53012_ ( .A(_28229_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01625_) );
  \$mux  #( .WIDTH(1) ) _53013_ ( .A(_dataflow_slice_valid_60), .B(1'h0), .S(_06250_), .Y(_28230_) );
  \$mux  #( .WIDTH(1) ) _53014_ ( .A(_28230_), .B(_wvalid_290), .S(_06248_), .Y(_28231_) );
  \$mux  #( .WIDTH(1) ) _53015_ ( .A(_28231_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01668_) );
  \$mux  #( .WIDTH(8) ) _53016_ ( .A(_dataflow_slice_data_60), .B(_wdata_289[23:16]), .S(_06249_), .Y(_28232_) );
  \$mux  #( .WIDTH(8) ) _53017_ ( .A(_28232_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01624_) );
  \$mux  #( .WIDTH(1) ) _53018_ ( .A(_dataflow_slice_valid_57), .B(1'h0), .S(_06247_), .Y(_28233_) );
  \$mux  #( .WIDTH(1) ) _53019_ ( .A(_28233_), .B(_wvalid_290), .S(_06245_), .Y(_28234_) );
  \$mux  #( .WIDTH(1) ) _53020_ ( .A(_28234_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01667_) );
  \$mux  #( .WIDTH(8) ) _53021_ ( .A(_dataflow_slice_data_57), .B(_wdata_289[15:8]), .S(_06246_), .Y(_28235_) );
  \$mux  #( .WIDTH(8) ) _53022_ ( .A(_28235_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01623_) );
  \$mux  #( .WIDTH(1) ) _53023_ ( .A(_dataflow_slice_valid_54), .B(1'h0), .S(_06244_), .Y(_28236_) );
  \$mux  #( .WIDTH(1) ) _53024_ ( .A(_28236_), .B(_wvalid_290), .S(_06242_), .Y(_28237_) );
  \$mux  #( .WIDTH(1) ) _53025_ ( .A(_28237_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01666_) );
  \$mux  #( .WIDTH(8) ) _53026_ ( .A(_dataflow_slice_data_54), .B(_wdata_289[7:0]), .S(_06243_), .Y(_28238_) );
  \$mux  #( .WIDTH(8) ) _53027_ ( .A(_28238_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01622_) );
  \$mux  #( .WIDTH(1) ) _53028_ ( .A(_dataflow_slice_valid_50), .B(1'h0), .S(_06241_), .Y(_28239_) );
  \$mux  #( .WIDTH(1) ) _53029_ ( .A(_28239_), .B(_wvalid_37), .S(_06239_), .Y(_28240_) );
  \$mux  #( .WIDTH(1) ) _53030_ ( .A(_28240_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01665_) );
  \$mux  #( .WIDTH(4) ) _53031_ ( .A(_dataflow_slice_data_50), .B(_wdata_36[31:28]), .S(_06240_), .Y(_28241_) );
  \$mux  #( .WIDTH(4) ) _53032_ ( .A(_28241_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01621_) );
  \$mux  #( .WIDTH(1) ) _53033_ ( .A(_dataflow_slice_valid_47), .B(1'h0), .S(_06238_), .Y(_28242_) );
  \$mux  #( .WIDTH(1) ) _53034_ ( .A(_28242_), .B(_wvalid_37), .S(_06236_), .Y(_28243_) );
  \$mux  #( .WIDTH(1) ) _53035_ ( .A(_28243_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01664_) );
  \$mux  #( .WIDTH(4) ) _53036_ ( .A(_dataflow_slice_data_47), .B(_wdata_36[27:24]), .S(_06237_), .Y(_28244_) );
  \$mux  #( .WIDTH(4) ) _53037_ ( .A(_28244_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01620_) );
  \$mux  #( .WIDTH(1) ) _53038_ ( .A(_dataflow_slice_valid_44), .B(1'h0), .S(_06235_), .Y(_28245_) );
  \$mux  #( .WIDTH(1) ) _53039_ ( .A(_28245_), .B(_wvalid_37), .S(_06233_), .Y(_28246_) );
  \$mux  #( .WIDTH(1) ) _53040_ ( .A(_28246_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01663_) );
  \$mux  #( .WIDTH(4) ) _53041_ ( .A(_dataflow_slice_data_44), .B(_wdata_36[23:20]), .S(_06234_), .Y(_28247_) );
  \$mux  #( .WIDTH(4) ) _53042_ ( .A(_28247_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01619_) );
  \$mux  #( .WIDTH(1) ) _53043_ ( .A(_dataflow_slice_valid_41), .B(1'h0), .S(_06232_), .Y(_28248_) );
  \$mux  #( .WIDTH(1) ) _53044_ ( .A(_28248_), .B(_wvalid_37), .S(_06230_), .Y(_28249_) );
  \$mux  #( .WIDTH(1) ) _53045_ ( .A(_28249_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01662_) );
  \$mux  #( .WIDTH(4) ) _53046_ ( .A(_dataflow_slice_data_41), .B(_wdata_36[19:16]), .S(_06231_), .Y(_28250_) );
  \$mux  #( .WIDTH(4) ) _53047_ ( .A(_28250_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01618_) );
  \$mux  #( .WIDTH(1) ) _53048_ ( .A(_dataflow_slice_valid_38), .B(1'h0), .S(_06229_), .Y(_28251_) );
  \$mux  #( .WIDTH(1) ) _53049_ ( .A(_28251_), .B(_wvalid_37), .S(_06227_), .Y(_28252_) );
  \$mux  #( .WIDTH(1) ) _53050_ ( .A(_28252_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01660_) );
  \$mux  #( .WIDTH(4) ) _53051_ ( .A(_dataflow_slice_data_38), .B(_wdata_36[15:12]), .S(_06228_), .Y(_28253_) );
  \$mux  #( .WIDTH(4) ) _53052_ ( .A(_28253_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01616_) );
  \$mux  #( .WIDTH(1) ) _53053_ ( .A(_dataflow_slice_valid_35), .B(1'h0), .S(_06226_), .Y(_28254_) );
  \$mux  #( .WIDTH(1) ) _53054_ ( .A(_28254_), .B(_wvalid_37), .S(_06224_), .Y(_28255_) );
  \$mux  #( .WIDTH(1) ) _53055_ ( .A(_28255_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01659_) );
  \$mux  #( .WIDTH(4) ) _53056_ ( .A(_dataflow_slice_data_35), .B(_wdata_36[11:8]), .S(_06225_), .Y(_28256_) );
  \$mux  #( .WIDTH(4) ) _53057_ ( .A(_28256_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01615_) );
  \$mux  #( .WIDTH(1) ) _53058_ ( .A(_dataflow_slice_valid_32), .B(1'h0), .S(_06223_), .Y(_28257_) );
  \$mux  #( .WIDTH(1) ) _53059_ ( .A(_28257_), .B(_wvalid_37), .S(_06221_), .Y(_28258_) );
  \$mux  #( .WIDTH(1) ) _53060_ ( .A(_28258_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01658_) );
  \$mux  #( .WIDTH(4) ) _53061_ ( .A(_dataflow_slice_data_32), .B(_wdata_36[7:4]), .S(_06222_), .Y(_28259_) );
  \$mux  #( .WIDTH(4) ) _53062_ ( .A(_28259_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01614_) );
  \$mux  #( .WIDTH(1) ) _53063_ ( .A(_dataflow_slice_valid_29), .B(1'h0), .S(_06220_), .Y(_28260_) );
  \$mux  #( .WIDTH(1) ) _53064_ ( .A(_28260_), .B(_wvalid_37), .S(_06218_), .Y(_28261_) );
  \$mux  #( .WIDTH(1) ) _53065_ ( .A(_28261_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01657_) );
  \$mux  #( .WIDTH(4) ) _53066_ ( .A(_dataflow_slice_data_29), .B(_wdata_36[3:0]), .S(_06219_), .Y(_28262_) );
  \$mux  #( .WIDTH(4) ) _53067_ ( .A(_28262_), .B(4'h0), .S(_RESETN_inv_2), .Y(_01613_) );
  \$mux  #( .WIDTH(1) ) _53068_ ( .A(_dataflow_slice_valid_25), .B(1'h0), .S(_06217_), .Y(_28263_) );
  \$mux  #( .WIDTH(1) ) _53069_ ( .A(_28263_), .B(_wvalid_24), .S(_06215_), .Y(_28264_) );
  \$mux  #( .WIDTH(1) ) _53070_ ( .A(_28264_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01656_) );
  \$mux  #( .WIDTH(8) ) _53071_ ( .A(_dataflow_slice_data_25), .B(_wdata_23[31:24]), .S(_06216_), .Y(_28265_) );
  \$mux  #( .WIDTH(8) ) _53072_ ( .A(_28265_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01612_) );
  \$mux  #( .WIDTH(1) ) _53073_ ( .A(_dataflow_slice_valid_22), .B(1'h0), .S(_06214_), .Y(_28266_) );
  \$mux  #( .WIDTH(1) ) _53074_ ( .A(_28266_), .B(_wvalid_24), .S(_06212_), .Y(_28267_) );
  \$mux  #( .WIDTH(1) ) _53075_ ( .A(_28267_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01655_) );
  \$mux  #( .WIDTH(8) ) _53076_ ( .A(_dataflow_slice_data_22), .B(_wdata_23[23:16]), .S(_06213_), .Y(_28268_) );
  \$mux  #( .WIDTH(8) ) _53077_ ( .A(_28268_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01611_) );
  \$mux  #( .WIDTH(1) ) _53078_ ( .A(_dataflow_slice_valid_19), .B(1'h0), .S(_06211_), .Y(_28269_) );
  \$mux  #( .WIDTH(1) ) _53079_ ( .A(_28269_), .B(_wvalid_24), .S(_06209_), .Y(_28270_) );
  \$mux  #( .WIDTH(1) ) _53080_ ( .A(_28270_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01654_) );
  \$mux  #( .WIDTH(8) ) _53081_ ( .A(_dataflow_slice_data_19), .B(_wdata_23[15:8]), .S(_06210_), .Y(_28271_) );
  \$mux  #( .WIDTH(8) ) _53082_ ( .A(_28271_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01610_) );
  \$mux  #( .WIDTH(1) ) _53083_ ( .A(_dataflow_slice_valid_16), .B(1'h0), .S(_06208_), .Y(_28272_) );
  \$mux  #( .WIDTH(1) ) _53084_ ( .A(_28272_), .B(_wvalid_24), .S(_06206_), .Y(_28273_) );
  \$mux  #( .WIDTH(1) ) _53085_ ( .A(_28273_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01653_) );
  \$mux  #( .WIDTH(8) ) _53086_ ( .A(_dataflow_slice_data_16), .B(_wdata_23[7:0]), .S(_06207_), .Y(_28274_) );
  \$mux  #( .WIDTH(8) ) _53087_ ( .A(_28274_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01609_) );
  \$mux  #( .WIDTH(1) ) _53088_ ( .A(_dataflow_slice_valid_12), .B(1'h0), .S(_06205_), .Y(_28275_) );
  \$mux  #( .WIDTH(1) ) _53089_ ( .A(_28275_), .B(_wvalid_11), .S(_06203_), .Y(_28276_) );
  \$mux  #( .WIDTH(1) ) _53090_ ( .A(_28276_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01642_) );
  \$mux  #( .WIDTH(8) ) _53091_ ( .A(_dataflow_slice_data_12), .B(_wdata_10[31:24]), .S(_06204_), .Y(_28277_) );
  \$mux  #( .WIDTH(8) ) _53092_ ( .A(_28277_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01598_) );
  \$mux  #( .WIDTH(1) ) _53093_ ( .A(_dataflow_slice_valid_9), .B(1'h0), .S(_06202_), .Y(_28278_) );
  \$mux  #( .WIDTH(1) ) _53094_ ( .A(_28278_), .B(_wvalid_11), .S(_06200_), .Y(_28279_) );
  \$mux  #( .WIDTH(1) ) _53095_ ( .A(_28279_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01679_) );
  \$mux  #( .WIDTH(8) ) _53096_ ( .A(_dataflow_slice_data_9), .B(_wdata_10[23:16]), .S(_06201_), .Y(_28280_) );
  \$mux  #( .WIDTH(8) ) _53097_ ( .A(_28280_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01635_) );
  \$mux  #( .WIDTH(1) ) _53098_ ( .A(_dataflow_slice_valid_6), .B(1'h0), .S(_06199_), .Y(_28281_) );
  \$mux  #( .WIDTH(1) ) _53099_ ( .A(_28281_), .B(_wvalid_11), .S(_06197_), .Y(_28282_) );
  \$mux  #( .WIDTH(1) ) _53100_ ( .A(_28282_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01671_) );
  \$mux  #( .WIDTH(8) ) _53101_ ( .A(_dataflow_slice_data_6), .B(_wdata_10[15:8]), .S(_06198_), .Y(_28283_) );
  \$mux  #( .WIDTH(8) ) _53102_ ( .A(_28283_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01627_) );
  \$mux  #( .WIDTH(1) ) _53103_ ( .A(_dataflow_slice_valid_3), .B(1'h0), .S(_06196_), .Y(_28284_) );
  \$mux  #( .WIDTH(1) ) _53104_ ( .A(_28284_), .B(_wvalid_11), .S(_06194_), .Y(_28285_) );
  \$mux  #( .WIDTH(1) ) _53105_ ( .A(_28285_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01661_) );
  \$mux  #( .WIDTH(8) ) _53106_ ( .A(_dataflow_slice_data_3), .B(_wdata_10[7:0]), .S(_06195_), .Y(_28286_) );
  \$mux  #( .WIDTH(8) ) _53107_ ( .A(_28286_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01617_) );
  \$mux  #( .WIDTH(1) ) _53108_ ( .A(_tmp_1357), .B(1'h0), .S(_saxi_cond_0_1), .Y(_28287_) );
  \$mux  #( .WIDTH(1) ) _53109_ ( .A(_28287_), .B(1'h1), .S(_06193_), .Y(_28288_) );
  \$mux  #( .WIDTH(1) ) _53110_ ( .A(_28288_), .B(_tmp_1357), .S(_06189_), .Y(_28289_) );
  \$mux  #( .WIDTH(1) ) _53111_ ( .A(_28289_), .B(1'h0), .S(_RESETN_inv_2), .Y(_02966_) );
  \$mux  #( .WIDTH(32) ) _53112_ ( .A(_maxi_ram_w8_l2048_id1_1_write_local_stride), .B(1), .S(axim_flag_1308), .Y(_28290_) );
  \$mux  #( .WIDTH(32) ) _53113_ ( .A(_28290_), .B(0), .S(_RESETN_inv_2), .Y(_01744_) );
  \$mux  #( .WIDTH(33) ) _53114_ ( .A(_maxi_ram_w8_l2048_id1_1_write_size), .B(_24233_), .S(axim_flag_1308), .Y(_28291_) );
  \$mux  #( .WIDTH(33) ) _53115_ ( .A(_28291_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01746_) );
  \$mux  #( .WIDTH(32) ) _53116_ ( .A(_maxi_ram_w8_l2048_id1_1_write_global_addr), .B(_24232_), .S(axim_flag_1308), .Y(_28292_) );
  \$mux  #( .WIDTH(32) ) _53117_ ( .A(_28292_), .B(0), .S(_RESETN_inv_2), .Y(_01742_) );
  \$mux  #( .WIDTH(32) ) _53118_ ( .A(_maxi_ram_w8_l2048_id1_1_write_local_addr), .B({ 2'h0, _24231_[31:2] }), .S(axim_flag_1308), .Y(_28293_) );
  \$mux  #( .WIDTH(32) ) _53119_ ( .A(_28293_), .B(0), .S(_RESETN_inv_2), .Y(_01743_) );
  \$mux  #( .WIDTH(8) ) _53120_ ( .A(_maxi_ram_w8_l2048_id1_1_write_op_sel), .B(8'h03), .S(axim_flag_1308), .Y(_28294_) );
  \$mux  #( .WIDTH(8) ) _53121_ ( .A(_28294_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01745_) );
  \$mux  #( .WIDTH(1) ) _53122_ ( .A(1'h0), .B(1'h1), .S(axim_flag_1308), .Y(_28295_) );
  \$mux  #( .WIDTH(1) ) _53123_ ( .A(_28295_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01747_) );
  \$mux  #( .WIDTH(32) ) _53124_ ( .A(_maxi_ram_w8_l2048_id3_1_read_local_stride), .B(1), .S(axim_flag_1152), .Y(_28296_) );
  \$mux  #( .WIDTH(32) ) _53125_ ( .A(_28296_), .B(0), .S(_RESETN_inv_2), .Y(_01762_) );
  \$mux  #( .WIDTH(33) ) _53126_ ( .A(_maxi_ram_w8_l2048_id3_1_read_size), .B(_24230_), .S(axim_flag_1152), .Y(_28297_) );
  \$mux  #( .WIDTH(33) ) _53127_ ( .A(_28297_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01764_) );
  \$mux  #( .WIDTH(32) ) _53128_ ( .A(_maxi_ram_w8_l2048_id3_1_read_global_addr), .B(matmul_29_mux_act_gaddr_0), .S(axim_flag_1152), .Y(_28298_) );
  \$mux  #( .WIDTH(32) ) _53129_ ( .A(_28298_), .B(0), .S(_RESETN_inv_2), .Y(_01760_) );
  \$mux  #( .WIDTH(32) ) _53130_ ( .A(_maxi_ram_w8_l2048_id3_1_read_local_addr), .B({ 2'h0, matmul_29_act_page_dma_offset_0[31:2] }), .S(axim_flag_1152), .Y(_28299_) );
  \$mux  #( .WIDTH(32) ) _53131_ ( .A(_28299_), .B(0), .S(_RESETN_inv_2), .Y(_01761_) );
  \$mux  #( .WIDTH(8) ) _53132_ ( .A(_maxi_ram_w8_l2048_id3_1_read_op_sel), .B(8'h09), .S(axim_flag_1152), .Y(_28300_) );
  \$mux  #( .WIDTH(8) ) _53133_ ( .A(_28300_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01763_) );
  \$mux  #( .WIDTH(1) ) _53134_ ( .A(1'h0), .B(1'h1), .S(axim_flag_1152), .Y(_28301_) );
  \$mux  #( .WIDTH(1) ) _53135_ ( .A(_28301_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01765_) );
  \$mux  #( .WIDTH(32) ) _53136_ ( .A(_maxi_ram_w4_l8192_id0_1_read_local_stride), .B(1), .S(axim_flag_1133), .Y(_28302_) );
  \$mux  #( .WIDTH(32) ) _53137_ ( .A(_28302_), .B(0), .S(_RESETN_inv_2), .Y(_01708_) );
  \$mux  #( .WIDTH(33) ) _53138_ ( .A(_maxi_ram_w4_l8192_id0_1_read_size), .B(_24229_), .S(axim_flag_1133), .Y(_28303_) );
  \$mux  #( .WIDTH(33) ) _53139_ ( .A(_28303_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01710_) );
  \$mux  #( .WIDTH(32) ) _53140_ ( .A(_maxi_ram_w4_l8192_id0_1_read_global_addr), .B(_24228_), .S(axim_flag_1133), .Y(_28304_) );
  \$mux  #( .WIDTH(32) ) _53141_ ( .A(_28304_), .B(0), .S(_RESETN_inv_2), .Y(_01706_) );
  \$mux  #( .WIDTH(32) ) _53142_ ( .A(_maxi_ram_w4_l8192_id0_1_read_local_addr), .B({ 3'h0, matmul_29_filter_page_dma_offset[31:3] }), .S(axim_flag_1133), .Y(_28305_) );
  \$mux  #( .WIDTH(32) ) _53143_ ( .A(_28305_), .B(0), .S(_RESETN_inv_2), .Y(_01707_) );
  \$mux  #( .WIDTH(8) ) _53144_ ( .A(_maxi_ram_w4_l8192_id0_1_read_op_sel), .B(8'h08), .S(axim_flag_1133), .Y(_28306_) );
  \$mux  #( .WIDTH(8) ) _53145_ ( .A(_28306_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01709_) );
  \$mux  #( .WIDTH(1) ) _53146_ ( .A(1'h0), .B(1'h1), .S(axim_flag_1133), .Y(_28307_) );
  \$mux  #( .WIDTH(1) ) _53147_ ( .A(_28307_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01711_) );
  \$mux  #( .WIDTH(32) ) _53148_ ( .A(_maxi_ram_w8_l2048_id2_1_read_local_stride), .B(1), .S(axim_flag_1121), .Y(_28308_) );
  \$mux  #( .WIDTH(32) ) _53149_ ( .A(_28308_), .B(0), .S(_RESETN_inv_2), .Y(_01750_) );
  \$mux  #( .WIDTH(33) ) _53150_ ( .A(_maxi_ram_w8_l2048_id2_1_read_size), .B(_24227_), .S(axim_flag_1121), .Y(_28309_) );
  \$mux  #( .WIDTH(33) ) _53151_ ( .A(_28309_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01752_) );
  \$mux  #( .WIDTH(32) ) _53152_ ( .A(_maxi_ram_w8_l2048_id2_1_read_global_addr), .B(matmul_29_arg_objaddr_2), .S(axim_flag_1121), .Y(_28310_) );
  \$mux  #( .WIDTH(32) ) _53153_ ( .A(_28310_), .B(0), .S(_RESETN_inv_2), .Y(_01748_) );
  \$mux  #( .WIDTH(32) ) _53154_ ( .A(_maxi_ram_w8_l2048_id2_1_read_local_addr), .B(0), .S(axim_flag_1121), .Y(_28311_) );
  \$mux  #( .WIDTH(32) ) _53155_ ( .A(_28311_), .B(0), .S(_RESETN_inv_2), .Y(_01749_) );
  \$mux  #( .WIDTH(8) ) _53156_ ( .A(_maxi_ram_w8_l2048_id2_1_read_op_sel), .B(8'h07), .S(axim_flag_1121), .Y(_28312_) );
  \$mux  #( .WIDTH(8) ) _53157_ ( .A(_28312_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01751_) );
  \$mux  #( .WIDTH(1) ) _53158_ ( .A(1'h0), .B(1'h1), .S(axim_flag_1121), .Y(_28313_) );
  \$mux  #( .WIDTH(1) ) _53159_ ( .A(_28313_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01753_) );
  \$mux  #( .WIDTH(1) ) _53160_ ( .A(_tmp_1120), .B(1'h0), .S(_saxi_cond_0_1), .Y(_28314_) );
  \$mux  #( .WIDTH(1) ) _53161_ ( .A(_28314_), .B(1'h1), .S(_06191_), .Y(_28315_) );
  \$mux  #( .WIDTH(1) ) _53162_ ( .A(_28315_), .B(_tmp_1120), .S(_06189_), .Y(_28316_) );
  \$mux  #( .WIDTH(1) ) _53163_ ( .A(_28316_), .B(1'h0), .S(_RESETN_inv_2), .Y(_02903_) );
  \$mux  #( .WIDTH(32) ) _53164_ ( .A(_maxi_ram_w8_l2048_id0_1_write_local_stride), .B(1), .S(axim_flag_1071), .Y(_28317_) );
  \$mux  #( .WIDTH(32) ) _53165_ ( .A(_28317_), .B(0), .S(_RESETN_inv_2), .Y(_01726_) );
  \$mux  #( .WIDTH(33) ) _53166_ ( .A(_maxi_ram_w8_l2048_id0_1_write_size), .B(33'h000000040), .S(axim_flag_1071), .Y(_28318_) );
  \$mux  #( .WIDTH(33) ) _53167_ ( .A(_28318_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01728_) );
  \$mux  #( .WIDTH(32) ) _53168_ ( .A(_maxi_ram_w8_l2048_id0_1_write_global_addr), .B(_24226_), .S(axim_flag_1071), .Y(_28319_) );
  \$mux  #( .WIDTH(32) ) _53169_ ( .A(_28319_), .B(0), .S(_RESETN_inv_2), .Y(_01724_) );
  \$mux  #( .WIDTH(32) ) _53170_ ( .A(_maxi_ram_w8_l2048_id0_1_write_local_addr), .B({ 2'h0, max_pool_serial_18_out_page_dma_offset[31:2] }), .S(axim_flag_1071), .Y(_28320_) );
  \$mux  #( .WIDTH(32) ) _53171_ ( .A(_28320_), .B(0), .S(_RESETN_inv_2), .Y(_01725_) );
  \$mux  #( .WIDTH(8) ) _53172_ ( .A(_maxi_ram_w8_l2048_id0_1_write_op_sel), .B(8'h02), .S(axim_flag_1071), .Y(_28321_) );
  \$mux  #( .WIDTH(8) ) _53173_ ( .A(_28321_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01727_) );
  \$mux  #( .WIDTH(1) ) _53174_ ( .A(1'h0), .B(1'h1), .S(axim_flag_1071), .Y(_28322_) );
  \$mux  #( .WIDTH(1) ) _53175_ ( .A(_28322_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01729_) );
  \$mux  #( .WIDTH(1) ) _53176_ ( .A(_tmp_1020), .B(1'h0), .S(_saxi_cond_0_1), .Y(_28323_) );
  \$mux  #( .WIDTH(1) ) _53177_ ( .A(_28323_), .B(1'h1), .S(_06188_), .Y(_28324_) );
  \$mux  #( .WIDTH(1) ) _53178_ ( .A(_28324_), .B(_tmp_1020), .S(_06189_), .Y(_28325_) );
  \$mux  #( .WIDTH(1) ) _53179_ ( .A(_28325_), .B(1'h0), .S(_RESETN_inv_2), .Y(_02868_) );
  \$mux  #( .WIDTH(9) ) _53180_ ( .A(_tmp_1019), .B(_maxi_write_cur_size[8:0]), .S(_06184_), .Y(_28326_) );
  \$mux  #( .WIDTH(9) ) _53181_ ( .A(_28326_), .B(_28535_[8:0]), .S(_06187_), .Y(_28327_) );
  \$mux  #( .WIDTH(9) ) _53182_ ( .A(_28327_), .B(_28535_[8:0]), .S(_06190_), .Y(_28328_) );
  \$mux  #( .WIDTH(9) ) _53183_ ( .A(_28328_), .B(_28535_[8:0]), .S(_06192_), .Y(_28329_) );
  \$mux  #( .WIDTH(9) ) _53184_ ( .A(_28329_), .B(9'h000), .S(_RESETN_inv_2), .Y(_02866_) );
  \$mux  #( .WIDTH(32) ) _53185_ ( .A(_maxi_ram_w8_l2048_id11_1_write_local_stride), .B(1), .S(axim_flag_970), .Y(_28330_) );
  \$mux  #( .WIDTH(32) ) _53186_ ( .A(_28330_), .B(0), .S(_RESETN_inv_2), .Y(_01732_) );
  \$mux  #( .WIDTH(33) ) _53187_ ( .A(_maxi_ram_w8_l2048_id11_1_write_size), .B(_24221_), .S(axim_flag_970), .Y(_28331_) );
  \$mux  #( .WIDTH(33) ) _53188_ ( .A(_28331_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01734_) );
  \$mux  #( .WIDTH(32) ) _53189_ ( .A(_maxi_ram_w8_l2048_id11_1_write_global_addr), .B(_24220_), .S(axim_flag_970), .Y(_28332_) );
  \$mux  #( .WIDTH(32) ) _53190_ ( .A(_28332_), .B(0), .S(_RESETN_inv_2), .Y(_01730_) );
  \$mux  #( .WIDTH(32) ) _53191_ ( .A(_maxi_ram_w8_l2048_id11_1_write_local_addr), .B({ 2'h0, _24219_[31:2] }), .S(axim_flag_970), .Y(_28333_) );
  \$mux  #( .WIDTH(32) ) _53192_ ( .A(_28333_), .B(0), .S(_RESETN_inv_2), .Y(_01731_) );
  \$mux  #( .WIDTH(8) ) _53193_ ( .A(_maxi_ram_w8_l2048_id11_1_write_op_sel), .B(8'h01), .S(axim_flag_970), .Y(_28334_) );
  \$mux  #( .WIDTH(8) ) _53194_ ( .A(_28334_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01733_) );
  \$mux  #( .WIDTH(1) ) _53195_ ( .A(1'h0), .B(1'h1), .S(axim_flag_970), .Y(_28335_) );
  \$mux  #( .WIDTH(1) ) _53196_ ( .A(_28335_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01735_) );
  \$mux  #( .WIDTH(32) ) _53197_ ( .A(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_stride), .B(1), .S(axim_flag_402), .Y(_28336_) );
  \$mux  #( .WIDTH(32) ) _53198_ ( .A(_28336_), .B(0), .S(_RESETN_inv_2), .Y(_01774_) );
  \$mux  #( .WIDTH(33) ) _53199_ ( .A(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_size), .B(_24218_), .S(axim_flag_402), .Y(_28337_) );
  \$mux  #( .WIDTH(33) ) _53200_ ( .A(_28337_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01776_) );
  \$mux  #( .WIDTH(32) ) _53201_ ( .A(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_global_addr), .B(conv2d_16_mux_act_gaddr_2), .S(axim_flag_402), .Y(_28338_) );
  \$mux  #( .WIDTH(32) ) _53202_ ( .A(_28338_), .B(0), .S(_RESETN_inv_2), .Y(_01772_) );
  \$mux  #( .WIDTH(32) ) _53203_ ( .A(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_addr), .B({ 2'h0, conv2d_16_act_page_dma_offset_2[31:2] }), .S(axim_flag_402), .Y(_28339_) );
  \$mux  #( .WIDTH(32) ) _53204_ ( .A(_28339_), .B(0), .S(_RESETN_inv_2), .Y(_01773_) );
  \$mux  #( .WIDTH(8) ) _53205_ ( .A(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_op_sel), .B(8'h06), .S(axim_flag_402), .Y(_28340_) );
  \$mux  #( .WIDTH(8) ) _53206_ ( .A(_28340_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01775_) );
  \$mux  #( .WIDTH(1) ) _53207_ ( .A(1'h0), .B(1'h1), .S(axim_flag_402), .Y(_28341_) );
  \$mux  #( .WIDTH(1) ) _53208_ ( .A(_28341_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01777_) );
  \$mux  #( .WIDTH(32) ) _53209_ ( .A(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_stride), .B(1), .S(axim_flag_345), .Y(_28342_) );
  \$mux  #( .WIDTH(32) ) _53210_ ( .A(_28342_), .B(0), .S(_RESETN_inv_2), .Y(_01768_) );
  \$mux  #( .WIDTH(33) ) _53211_ ( .A(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_size), .B(_24218_), .S(axim_flag_345), .Y(_28343_) );
  \$mux  #( .WIDTH(33) ) _53212_ ( .A(_28343_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01770_) );
  \$mux  #( .WIDTH(32) ) _53213_ ( .A(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_global_addr), .B(conv2d_16_mux_act_gaddr_1), .S(axim_flag_345), .Y(_28344_) );
  \$mux  #( .WIDTH(32) ) _53214_ ( .A(_28344_), .B(0), .S(_RESETN_inv_2), .Y(_01766_) );
  \$mux  #( .WIDTH(32) ) _53215_ ( .A(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_addr), .B({ 2'h0, conv2d_16_act_page_dma_offset_1[31:2] }), .S(axim_flag_345), .Y(_28345_) );
  \$mux  #( .WIDTH(32) ) _53216_ ( .A(_28345_), .B(0), .S(_RESETN_inv_2), .Y(_01767_) );
  \$mux  #( .WIDTH(8) ) _53217_ ( .A(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_op_sel), .B(8'h05), .S(axim_flag_345), .Y(_28346_) );
  \$mux  #( .WIDTH(8) ) _53218_ ( .A(_28346_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01769_) );
  \$mux  #( .WIDTH(1) ) _53219_ ( .A(1'h0), .B(1'h1), .S(axim_flag_345), .Y(_28347_) );
  \$mux  #( .WIDTH(1) ) _53220_ ( .A(_28347_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01771_) );
  \$mux  #( .WIDTH(32) ) _53221_ ( .A(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_stride), .B(1), .S(axim_flag_288), .Y(_28348_) );
  \$mux  #( .WIDTH(32) ) _53222_ ( .A(_28348_), .B(0), .S(_RESETN_inv_2), .Y(_01756_) );
  \$mux  #( .WIDTH(33) ) _53223_ ( .A(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_size), .B(_24218_), .S(axim_flag_288), .Y(_28349_) );
  \$mux  #( .WIDTH(33) ) _53224_ ( .A(_28349_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01758_) );
  \$mux  #( .WIDTH(32) ) _53225_ ( .A(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_global_addr), .B(conv2d_16_mux_act_gaddr_0), .S(axim_flag_288), .Y(_28350_) );
  \$mux  #( .WIDTH(32) ) _53226_ ( .A(_28350_), .B(0), .S(_RESETN_inv_2), .Y(_01754_) );
  \$mux  #( .WIDTH(32) ) _53227_ ( .A(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_addr), .B({ 2'h0, conv2d_16_act_page_dma_offset_0[31:2] }), .S(axim_flag_288), .Y(_28351_) );
  \$mux  #( .WIDTH(32) ) _53228_ ( .A(_28351_), .B(0), .S(_RESETN_inv_2), .Y(_01755_) );
  \$mux  #( .WIDTH(8) ) _53229_ ( .A(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_op_sel), .B(8'h04), .S(axim_flag_288), .Y(_28352_) );
  \$mux  #( .WIDTH(8) ) _53230_ ( .A(_28352_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01757_) );
  \$mux  #( .WIDTH(1) ) _53231_ ( .A(1'h0), .B(1'h1), .S(axim_flag_288), .Y(_28353_) );
  \$mux  #( .WIDTH(1) ) _53232_ ( .A(_28353_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01759_) );
  \$mux  #( .WIDTH(32) ) _53233_ ( .A(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_stride), .B(1), .S(axim_flag_35), .Y(_28354_) );
  \$mux  #( .WIDTH(32) ) _53234_ ( .A(_28354_), .B(0), .S(_RESETN_inv_2), .Y(_01714_) );
  \$mux  #( .WIDTH(33) ) _53235_ ( .A(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_size), .B(_24217_), .S(axim_flag_35), .Y(_28355_) );
  \$mux  #( .WIDTH(33) ) _53236_ ( .A(_28355_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01716_) );
  \$mux  #( .WIDTH(32) ) _53237_ ( .A(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_global_addr), .B(_24216_), .S(axim_flag_35), .Y(_28356_) );
  \$mux  #( .WIDTH(32) ) _53238_ ( .A(_28356_), .B(0), .S(_RESETN_inv_2), .Y(_01712_) );
  \$mux  #( .WIDTH(32) ) _53239_ ( .A(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_addr), .B({ 3'h0, conv2d_16_filter_page_dma_offset[31:3] }), .S(axim_flag_35), .Y(_28357_) );
  \$mux  #( .WIDTH(32) ) _53240_ ( .A(_28357_), .B(0), .S(_RESETN_inv_2), .Y(_01713_) );
  \$mux  #( .WIDTH(8) ) _53241_ ( .A(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_op_sel), .B(8'h03), .S(axim_flag_35), .Y(_28358_) );
  \$mux  #( .WIDTH(8) ) _53242_ ( .A(_28358_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01715_) );
  \$mux  #( .WIDTH(1) ) _53243_ ( .A(1'h0), .B(1'h1), .S(axim_flag_35), .Y(_28359_) );
  \$mux  #( .WIDTH(1) ) _53244_ ( .A(_28359_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01717_) );
  \$mux  #( .WIDTH(32) ) _53245_ ( .A(_maxi_ram_w8_l2048_id0_1_read_local_stride), .B(1), .S(axim_flag_22), .Y(_28360_) );
  \$mux  #( .WIDTH(32) ) _53246_ ( .A(_28360_), .B(1), .S(axim_flag_1132), .Y(_28361_) );
  \$mux  #( .WIDTH(32) ) _53247_ ( .A(_28361_), .B(0), .S(_RESETN_inv_2), .Y(_01720_) );
  \$mux  #( .WIDTH(33) ) _53248_ ( .A(_maxi_ram_w8_l2048_id0_1_read_size), .B(33'h000000001), .S(axim_flag_22), .Y(_28362_) );
  \$mux  #( .WIDTH(33) ) _53249_ ( .A(_28362_), .B(33'h000000001), .S(axim_flag_1132), .Y(_28363_) );
  \$mux  #( .WIDTH(33) ) _53250_ ( .A(_28363_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01722_) );
  \$mux  #( .WIDTH(32) ) _53251_ ( .A(_maxi_ram_w8_l2048_id0_1_read_global_addr), .B(conv2d_16_arg_objaddr_3), .S(axim_flag_22), .Y(_28364_) );
  \$mux  #( .WIDTH(32) ) _53252_ ( .A(_28364_), .B(matmul_29_arg_objaddr_3), .S(axim_flag_1132), .Y(_28365_) );
  \$mux  #( .WIDTH(32) ) _53253_ ( .A(_28365_), .B(0), .S(_RESETN_inv_2), .Y(_01718_) );
  \$mux  #( .WIDTH(32) ) _53254_ ( .A(_maxi_ram_w8_l2048_id0_1_read_local_addr), .B(0), .S(axim_flag_22), .Y(_28366_) );
  \$mux  #( .WIDTH(32) ) _53255_ ( .A(_28366_), .B(0), .S(axim_flag_1132), .Y(_28367_) );
  \$mux  #( .WIDTH(32) ) _53256_ ( .A(_28367_), .B(0), .S(_RESETN_inv_2), .Y(_01719_) );
  \$mux  #( .WIDTH(8) ) _53257_ ( .A(_maxi_ram_w8_l2048_id0_1_read_op_sel), .B(8'h02), .S(axim_flag_22), .Y(_28368_) );
  \$mux  #( .WIDTH(8) ) _53258_ ( .A(_28368_), .B(8'h02), .S(axim_flag_1132), .Y(_28369_) );
  \$mux  #( .WIDTH(8) ) _53259_ ( .A(_28369_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01721_) );
  \$mux  #( .WIDTH(1) ) _53260_ ( .A(1'h0), .B(1'h1), .S(axim_flag_22), .Y(_28370_) );
  \$mux  #( .WIDTH(1) ) _53261_ ( .A(_28370_), .B(1'h1), .S(axim_flag_1132), .Y(_28371_) );
  \$mux  #( .WIDTH(1) ) _53262_ ( .A(_28371_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01723_) );
  \$mux  #( .WIDTH(9) ) _53263_ ( .A(_tmp_20), .B(_maxi_read_cur_size[8:0]), .S(_06181_), .Y(_28372_) );
  \$mux  #( .WIDTH(9) ) _53264_ ( .A(_28372_), .B(_28533_[8:0]), .S(_06183_), .Y(_28373_) );
  \$mux  #( .WIDTH(9) ) _53265_ ( .A(_28373_), .B(9'h000), .S(_RESETN_inv_2), .Y(_03009_) );
  \$mux  #( .WIDTH(32) ) _53266_ ( .A(_maxi_ram_w8_l2048_id1_1_read_local_stride), .B(1), .S(axim_flag_9), .Y(_28374_) );
  \$mux  #( .WIDTH(32) ) _53267_ ( .A(_28374_), .B(1), .S(axim_flag_1022), .Y(_28375_) );
  \$mux  #( .WIDTH(32) ) _53268_ ( .A(_28375_), .B(1), .S(axim_flag_1023), .Y(_28376_) );
  \$mux  #( .WIDTH(32) ) _53269_ ( .A(_28376_), .B(0), .S(_RESETN_inv_2), .Y(_01738_) );
  \$mux  #( .WIDTH(33) ) _53270_ ( .A(_maxi_ram_w8_l2048_id1_1_read_size), .B(_24215_), .S(axim_flag_9), .Y(_28377_) );
  \$mux  #( .WIDTH(33) ) _53271_ ( .A(_28377_), .B(33'h000000080), .S(axim_flag_1022), .Y(_28378_) );
  \$mux  #( .WIDTH(33) ) _53272_ ( .A(_28378_), .B(33'h000000080), .S(axim_flag_1023), .Y(_28379_) );
  \$mux  #( .WIDTH(33) ) _53273_ ( .A(_28379_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01740_) );
  \$mux  #( .WIDTH(32) ) _53274_ ( .A(_maxi_ram_w8_l2048_id1_1_read_global_addr), .B(conv2d_16_arg_objaddr_2), .S(axim_flag_9), .Y(_28380_) );
  \$mux  #( .WIDTH(32) ) _53275_ ( .A(_28380_), .B(_24222_), .S(axim_flag_1022), .Y(_28381_) );
  \$mux  #( .WIDTH(32) ) _53276_ ( .A(_28381_), .B(_24225_), .S(axim_flag_1023), .Y(_28382_) );
  \$mux  #( .WIDTH(32) ) _53277_ ( .A(_28382_), .B(0), .S(_RESETN_inv_2), .Y(_01736_) );
  \$mux  #( .WIDTH(32) ) _53278_ ( .A(_maxi_ram_w8_l2048_id1_1_read_local_addr), .B(0), .S(axim_flag_9), .Y(_28383_) );
  \$mux  #( .WIDTH(32) ) _53279_ ( .A(_28383_), .B({ 2'h0, max_pool_serial_18_act_page_dma_offset[31:2] }), .S(axim_flag_1022), .Y(_28384_) );
  \$mux  #( .WIDTH(32) ) _53280_ ( .A(_28384_), .B({ 2'h0, _24223_[31:2] }), .S(axim_flag_1023), .Y(_28385_) );
  \$mux  #( .WIDTH(32) ) _53281_ ( .A(_28385_), .B(0), .S(_RESETN_inv_2), .Y(_01737_) );
  \$mux  #( .WIDTH(8) ) _53282_ ( .A(_maxi_ram_w8_l2048_id1_1_read_op_sel), .B(8'h01), .S(axim_flag_9), .Y(_28386_) );
  \$mux  #( .WIDTH(8) ) _53283_ ( .A(_28386_), .B(8'h01), .S(axim_flag_1022), .Y(_28387_) );
  \$mux  #( .WIDTH(8) ) _53284_ ( .A(_28387_), .B(8'h01), .S(axim_flag_1023), .Y(_28388_) );
  \$mux  #( .WIDTH(8) ) _53285_ ( .A(_28388_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01739_) );
  \$mux  #( .WIDTH(1) ) _53286_ ( .A(1'h0), .B(1'h1), .S(axim_flag_9), .Y(_28389_) );
  \$mux  #( .WIDTH(1) ) _53287_ ( .A(_28389_), .B(1'h1), .S(axim_flag_1022), .Y(_28390_) );
  \$mux  #( .WIDTH(1) ) _53288_ ( .A(_28390_), .B(1'h1), .S(axim_flag_1023), .Y(_28391_) );
  \$mux  #( .WIDTH(1) ) _53289_ ( .A(_28391_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01741_) );
  \$mux  #( .WIDTH(32) ) _53290_ ( .A(_saxi_register_9), .B(0), .S(_RESETN_inv_2), .Y(_01705_) );
  \$mux  #( .WIDTH(1) ) _53291_ ( .A(_maxi_write_idle), .B(1'h0), .S(_maxi_ram_w8_l2048_id11_1_write_start), .Y(_28392_) );
  \$mux  #( .WIDTH(1) ) _53292_ ( .A(_28392_), .B(1'h1), .S(axim_flag_1021), .Y(_28393_) );
  \$mux  #( .WIDTH(1) ) _53293_ ( .A(_28393_), .B(1'h0), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_28394_) );
  \$mux  #( .WIDTH(1) ) _53294_ ( .A(_28394_), .B(1'h0), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_28395_) );
  \$mux  #( .WIDTH(1) ) _53295_ ( .A(_28395_), .B(1'h1), .S(_RESETN_inv_2), .Y(_01793_) );
  \$mux  #( .WIDTH(32) ) _53296_ ( .A(_maxi_write_local_stride), .B(_maxi_ram_w8_l2048_id11_1_write_local_stride), .S(_maxi_ram_w8_l2048_id11_1_write_start), .Y(_28396_) );
  \$mux  #( .WIDTH(32) ) _53297_ ( .A(_28396_), .B(_maxi_ram_w8_l2048_id0_1_write_local_stride), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_28397_) );
  \$mux  #( .WIDTH(32) ) _53298_ ( .A(_28397_), .B(_maxi_ram_w8_l2048_id1_1_write_local_stride), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_28398_) );
  \$mux  #( .WIDTH(32) ) _53299_ ( .A(_28398_), .B(0), .S(_RESETN_inv_2), .Y(_01795_) );
  \$mux  #( .WIDTH(33) ) _53300_ ( .A(_maxi_write_size), .B(_maxi_ram_w8_l2048_id11_1_write_size), .S(_maxi_ram_w8_l2048_id11_1_write_start), .Y(_28399_) );
  \$mux  #( .WIDTH(33) ) _53301_ ( .A(_28399_), .B(_maxi_ram_w8_l2048_id0_1_write_size), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_28400_) );
  \$mux  #( .WIDTH(33) ) _53302_ ( .A(_28400_), .B(_maxi_ram_w8_l2048_id1_1_write_size), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_28401_) );
  \$mux  #( .WIDTH(33) ) _53303_ ( .A(_28401_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01798_) );
  \$mux  #( .WIDTH(32) ) _53304_ ( .A(_maxi_write_global_addr), .B(_maxi_ram_w8_l2048_id11_1_write_global_addr), .S(_maxi_ram_w8_l2048_id11_1_write_start), .Y(_28402_) );
  \$mux  #( .WIDTH(32) ) _53305_ ( .A(_28402_), .B(_maxi_ram_w8_l2048_id0_1_write_global_addr), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_28403_) );
  \$mux  #( .WIDTH(32) ) _53306_ ( .A(_28403_), .B(_maxi_ram_w8_l2048_id1_1_write_global_addr), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_28404_) );
  \$mux  #( .WIDTH(32) ) _53307_ ( .A(_28404_), .B(0), .S(_RESETN_inv_2), .Y(_01792_) );
  \$mux  #( .WIDTH(32) ) _53308_ ( .A(_maxi_write_local_addr), .B(_maxi_ram_w8_l2048_id11_1_write_local_addr), .S(_maxi_ram_w8_l2048_id11_1_write_start), .Y(_28405_) );
  \$mux  #( .WIDTH(32) ) _53309_ ( .A(_28405_), .B(_maxi_ram_w8_l2048_id0_1_write_local_addr), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_28406_) );
  \$mux  #( .WIDTH(32) ) _53310_ ( .A(_28406_), .B(_maxi_ram_w8_l2048_id1_1_write_local_addr), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_28407_) );
  \$mux  #( .WIDTH(32) ) _53311_ ( .A(_28407_), .B(0), .S(_RESETN_inv_2), .Y(_01794_) );
  \$mux  #( .WIDTH(8) ) _53312_ ( .A(_maxi_write_op_sel), .B(_maxi_ram_w8_l2048_id11_1_write_op_sel), .S(_maxi_ram_w8_l2048_id11_1_write_start), .Y(_28408_) );
  \$mux  #( .WIDTH(8) ) _53313_ ( .A(_28408_), .B(_maxi_ram_w8_l2048_id0_1_write_op_sel), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_28409_) );
  \$mux  #( .WIDTH(8) ) _53314_ ( .A(_28409_), .B(_maxi_ram_w8_l2048_id1_1_write_op_sel), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_28410_) );
  \$mux  #( .WIDTH(8) ) _53315_ ( .A(_28410_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01796_) );
  \$mux  #( .WIDTH(1) ) _53316_ ( .A(1'h0), .B(1'h1), .S(_maxi_ram_w8_l2048_id11_1_write_start), .Y(_28411_) );
  \$mux  #( .WIDTH(1) ) _53317_ ( .A(_28411_), .B(1'h1), .S(_maxi_ram_w8_l2048_id0_1_write_start), .Y(_28412_) );
  \$mux  #( .WIDTH(1) ) _53318_ ( .A(_28412_), .B(1'h1), .S(_maxi_ram_w8_l2048_id1_1_write_start), .Y(_28413_) );
  \$mux  #( .WIDTH(1) ) _53319_ ( .A(_28413_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01799_) );
  \$mux  #( .WIDTH(1) ) _53320_ ( .A(_maxi_read_idle), .B(1'h0), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_28414_) );
  \$mux  #( .WIDTH(1) ) _53321_ ( .A(_28414_), .B(1'h1), .S(axim_flag_21), .Y(_28415_) );
  \$mux  #( .WIDTH(1) ) _53322_ ( .A(_28415_), .B(1'h0), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_28416_) );
  \$mux  #( .WIDTH(1) ) _53323_ ( .A(_28416_), .B(1'h0), .S(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start), .Y(_28417_) );
  \$mux  #( .WIDTH(1) ) _53324_ ( .A(_28417_), .B(1'h0), .S(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start), .Y(_28418_) );
  \$mux  #( .WIDTH(1) ) _53325_ ( .A(_28418_), .B(1'h0), .S(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start), .Y(_28419_) );
  \$mux  #( .WIDTH(1) ) _53326_ ( .A(_28419_), .B(1'h0), .S(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start), .Y(_28420_) );
  \$mux  #( .WIDTH(1) ) _53327_ ( .A(_28420_), .B(1'h0), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_28421_) );
  \$mux  #( .WIDTH(1) ) _53328_ ( .A(_28421_), .B(1'h0), .S(_maxi_ram_w4_l8192_id0_1_read_start), .Y(_28422_) );
  \$mux  #( .WIDTH(1) ) _53329_ ( .A(_28422_), .B(1'h0), .S(_maxi_ram_w8_l2048_id3_1_read_start), .Y(_28423_) );
  \$mux  #( .WIDTH(1) ) _53330_ ( .A(_28423_), .B(1'h1), .S(_RESETN_inv_2), .Y(_01782_) );
  \$mux  #( .WIDTH(32) ) _53331_ ( .A(_maxi_read_local_stride), .B(_maxi_ram_w8_l2048_id1_1_read_local_stride), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_28424_) );
  \$mux  #( .WIDTH(32) ) _53332_ ( .A(_28424_), .B(_maxi_ram_w8_l2048_id0_1_read_local_stride), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_28425_) );
  \$mux  #( .WIDTH(32) ) _53333_ ( .A(_28425_), .B(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_stride), .S(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start), .Y(_28426_) );
  \$mux  #( .WIDTH(32) ) _53334_ ( .A(_28426_), .B(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_stride), .S(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start), .Y(_28427_) );
  \$mux  #( .WIDTH(32) ) _53335_ ( .A(_28427_), .B(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_stride), .S(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start), .Y(_28428_) );
  \$mux  #( .WIDTH(32) ) _53336_ ( .A(_28428_), .B(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_stride), .S(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start), .Y(_28429_) );
  \$mux  #( .WIDTH(32) ) _53337_ ( .A(_28429_), .B(_maxi_ram_w8_l2048_id2_1_read_local_stride), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_28430_) );
  \$mux  #( .WIDTH(32) ) _53338_ ( .A(_28430_), .B(_maxi_ram_w4_l8192_id0_1_read_local_stride), .S(_maxi_ram_w4_l8192_id0_1_read_start), .Y(_28431_) );
  \$mux  #( .WIDTH(32) ) _53339_ ( .A(_28431_), .B(_maxi_ram_w8_l2048_id3_1_read_local_stride), .S(_maxi_ram_w8_l2048_id3_1_read_start), .Y(_28432_) );
  \$mux  #( .WIDTH(32) ) _53340_ ( .A(_28432_), .B(0), .S(_RESETN_inv_2), .Y(_01784_) );
  \$mux  #( .WIDTH(33) ) _53341_ ( .A(_maxi_read_size), .B(_maxi_ram_w8_l2048_id1_1_read_size), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_28433_) );
  \$mux  #( .WIDTH(33) ) _53342_ ( .A(_28433_), .B(_maxi_ram_w8_l2048_id0_1_read_size), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_28434_) );
  \$mux  #( .WIDTH(33) ) _53343_ ( .A(_28434_), .B(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_size), .S(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start), .Y(_28435_) );
  \$mux  #( .WIDTH(33) ) _53344_ ( .A(_28435_), .B(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_size), .S(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start), .Y(_28436_) );
  \$mux  #( .WIDTH(33) ) _53345_ ( .A(_28436_), .B(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_size), .S(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start), .Y(_28437_) );
  \$mux  #( .WIDTH(33) ) _53346_ ( .A(_28437_), .B(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_size), .S(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start), .Y(_28438_) );
  \$mux  #( .WIDTH(33) ) _53347_ ( .A(_28438_), .B(_maxi_ram_w8_l2048_id2_1_read_size), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_28439_) );
  \$mux  #( .WIDTH(33) ) _53348_ ( .A(_28439_), .B(_maxi_ram_w4_l8192_id0_1_read_size), .S(_maxi_ram_w4_l8192_id0_1_read_start), .Y(_28440_) );
  \$mux  #( .WIDTH(33) ) _53349_ ( .A(_28440_), .B(_maxi_ram_w8_l2048_id3_1_read_size), .S(_maxi_ram_w8_l2048_id3_1_read_start), .Y(_28441_) );
  \$mux  #( .WIDTH(33) ) _53350_ ( .A(_28441_), .B(33'h000000000), .S(_RESETN_inv_2), .Y(_01787_) );
  \$mux  #( .WIDTH(32) ) _53351_ ( .A(_maxi_read_global_addr), .B(_maxi_ram_w8_l2048_id1_1_read_global_addr), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_28442_) );
  \$mux  #( .WIDTH(32) ) _53352_ ( .A(_28442_), .B(_maxi_ram_w8_l2048_id0_1_read_global_addr), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_28443_) );
  \$mux  #( .WIDTH(32) ) _53353_ ( .A(_28443_), .B(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_global_addr), .S(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start), .Y(_28444_) );
  \$mux  #( .WIDTH(32) ) _53354_ ( .A(_28444_), .B(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_global_addr), .S(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start), .Y(_28445_) );
  \$mux  #( .WIDTH(32) ) _53355_ ( .A(_28445_), .B(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_global_addr), .S(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start), .Y(_28446_) );
  \$mux  #( .WIDTH(32) ) _53356_ ( .A(_28446_), .B(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_global_addr), .S(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start), .Y(_28447_) );
  \$mux  #( .WIDTH(32) ) _53357_ ( .A(_28447_), .B(_maxi_ram_w8_l2048_id2_1_read_global_addr), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_28448_) );
  \$mux  #( .WIDTH(32) ) _53358_ ( .A(_28448_), .B(_maxi_ram_w4_l8192_id0_1_read_global_addr), .S(_maxi_ram_w4_l8192_id0_1_read_start), .Y(_28449_) );
  \$mux  #( .WIDTH(32) ) _53359_ ( .A(_28449_), .B(_maxi_ram_w8_l2048_id3_1_read_global_addr), .S(_maxi_ram_w8_l2048_id3_1_read_start), .Y(_28450_) );
  \$mux  #( .WIDTH(32) ) _53360_ ( .A(_28450_), .B(0), .S(_RESETN_inv_2), .Y(_01781_) );
  \$mux  #( .WIDTH(32) ) _53361_ ( .A(_maxi_read_local_addr), .B(_maxi_ram_w8_l2048_id1_1_read_local_addr), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_28451_) );
  \$mux  #( .WIDTH(32) ) _53362_ ( .A(_28451_), .B(_maxi_ram_w8_l2048_id0_1_read_local_addr), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_28452_) );
  \$mux  #( .WIDTH(32) ) _53363_ ( .A(_28452_), .B(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_addr), .S(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start), .Y(_28453_) );
  \$mux  #( .WIDTH(32) ) _53364_ ( .A(_28453_), .B(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_addr), .S(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start), .Y(_28454_) );
  \$mux  #( .WIDTH(32) ) _53365_ ( .A(_28454_), .B(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_addr), .S(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start), .Y(_28455_) );
  \$mux  #( .WIDTH(32) ) _53366_ ( .A(_28455_), .B(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_addr), .S(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start), .Y(_28456_) );
  \$mux  #( .WIDTH(32) ) _53367_ ( .A(_28456_), .B(_maxi_ram_w8_l2048_id2_1_read_local_addr), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_28457_) );
  \$mux  #( .WIDTH(32) ) _53368_ ( .A(_28457_), .B(_maxi_ram_w4_l8192_id0_1_read_local_addr), .S(_maxi_ram_w4_l8192_id0_1_read_start), .Y(_28458_) );
  \$mux  #( .WIDTH(32) ) _53369_ ( .A(_28458_), .B(_maxi_ram_w8_l2048_id3_1_read_local_addr), .S(_maxi_ram_w8_l2048_id3_1_read_start), .Y(_28459_) );
  \$mux  #( .WIDTH(32) ) _53370_ ( .A(_28459_), .B(0), .S(_RESETN_inv_2), .Y(_01783_) );
  \$mux  #( .WIDTH(8) ) _53371_ ( .A(_maxi_read_op_sel), .B(_maxi_ram_w8_l2048_id1_1_read_op_sel), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_28460_) );
  \$mux  #( .WIDTH(8) ) _53372_ ( .A(_28460_), .B(_maxi_ram_w8_l2048_id0_1_read_op_sel), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_28461_) );
  \$mux  #( .WIDTH(8) ) _53373_ ( .A(_28461_), .B(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_op_sel), .S(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start), .Y(_28462_) );
  \$mux  #( .WIDTH(8) ) _53374_ ( .A(_28462_), .B(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_op_sel), .S(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start), .Y(_28463_) );
  \$mux  #( .WIDTH(8) ) _53375_ ( .A(_28463_), .B(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_op_sel), .S(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start), .Y(_28464_) );
  \$mux  #( .WIDTH(8) ) _53376_ ( .A(_28464_), .B(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_op_sel), .S(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start), .Y(_28465_) );
  \$mux  #( .WIDTH(8) ) _53377_ ( .A(_28465_), .B(_maxi_ram_w8_l2048_id2_1_read_op_sel), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_28466_) );
  \$mux  #( .WIDTH(8) ) _53378_ ( .A(_28466_), .B(_maxi_ram_w4_l8192_id0_1_read_op_sel), .S(_maxi_ram_w4_l8192_id0_1_read_start), .Y(_28467_) );
  \$mux  #( .WIDTH(8) ) _53379_ ( .A(_28467_), .B(_maxi_ram_w8_l2048_id3_1_read_op_sel), .S(_maxi_ram_w8_l2048_id3_1_read_start), .Y(_28468_) );
  \$mux  #( .WIDTH(8) ) _53380_ ( .A(_28468_), .B(8'h00), .S(_RESETN_inv_2), .Y(_01785_) );
  \$mux  #( .WIDTH(1) ) _53381_ ( .A(1'h0), .B(1'h1), .S(_maxi_ram_w8_l2048_id1_1_read_start), .Y(_28469_) );
  \$mux  #( .WIDTH(1) ) _53382_ ( .A(_28469_), .B(1'h1), .S(_maxi_ram_w8_l2048_id0_1_read_start), .Y(_28470_) );
  \$mux  #( .WIDTH(1) ) _53383_ ( .A(_28470_), .B(1'h1), .S(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start), .Y(_28471_) );
  \$mux  #( .WIDTH(1) ) _53384_ ( .A(_28471_), .B(1'h1), .S(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start), .Y(_28472_) );
  \$mux  #( .WIDTH(1) ) _53385_ ( .A(_28472_), .B(1'h1), .S(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start), .Y(_28473_) );
  \$mux  #( .WIDTH(1) ) _53386_ ( .A(_28473_), .B(1'h1), .S(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start), .Y(_28474_) );
  \$mux  #( .WIDTH(1) ) _53387_ ( .A(_28474_), .B(1'h1), .S(_maxi_ram_w8_l2048_id2_1_read_start), .Y(_28475_) );
  \$mux  #( .WIDTH(1) ) _53388_ ( .A(_28475_), .B(1'h1), .S(_maxi_ram_w4_l8192_id0_1_read_start), .Y(_28476_) );
  \$mux  #( .WIDTH(1) ) _53389_ ( .A(_28476_), .B(1'h1), .S(_maxi_ram_w8_l2048_id3_1_read_start), .Y(_28477_) );
  \$mux  #( .WIDTH(1) ) _53390_ ( .A(_28477_), .B(1'h0), .S(_RESETN_inv_2), .Y(_01788_) );
  \$mux  #( .WIDTH(1) ) _53391_ ( .A(maxi_arvalid), .B(1'h0), .S(_saxi_cond_0_1), .Y(_28478_) );
  \$mux  #( .WIDTH(1) ) _53392_ ( .A(_28478_), .B(1'h1), .S(_06181_), .Y(_28479_) );
  \$mux  #( .WIDTH(1) ) _53393_ ( .A(_28479_), .B(maxi_arvalid), .S(_06182_), .Y(_28480_) );
  \$mux  #( .WIDTH(1) ) _53394_ ( .A(_28480_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03365_) );
  \$mux  #( .WIDTH(8) ) _53395_ ( .A(maxi_arlen), .B(_28532_[7:0]), .S(_06181_), .Y(_28481_) );
  \$mux  #( .WIDTH(8) ) _53396_ ( .A(_28481_), .B(8'h00), .S(_RESETN_inv_2), .Y(_03364_) );
  \$mux  #( .WIDTH(32) ) _53397_ ( .A(maxi_araddr), .B(_maxi_read_cur_global_addr), .S(_06181_), .Y(_28482_) );
  \$mux  #( .WIDTH(32) ) _53398_ ( .A(_28482_), .B(0), .S(_RESETN_inv_2), .Y(_03363_) );
  \$mux  #( .WIDTH(1) ) _53399_ ( .A(maxi_wvalid), .B(1'h0), .S(_saxi_cond_0_1), .Y(_28483_) );
  \$mux  #( .WIDTH(1) ) _53400_ ( .A(_28483_), .B(1'h1), .S(_06187_), .Y(_28484_) );
  \$mux  #( .WIDTH(1) ) _53401_ ( .A(_28484_), .B(1'h1), .S(_06190_), .Y(_28485_) );
  \$mux  #( .WIDTH(1) ) _53402_ ( .A(_28485_), .B(1'h1), .S(_06192_), .Y(_28486_) );
  \$mux  #( .WIDTH(1) ) _53403_ ( .A(_28486_), .B(maxi_wvalid), .S(_06189_), .Y(_28487_) );
  \$mux  #( .WIDTH(1) ) _53404_ ( .A(_28487_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03372_) );
  \$mux  #( .WIDTH(1) ) _53405_ ( .A(maxi_wlast), .B(1'h0), .S(_saxi_cond_0_1), .Y(_28488_) );
  \$mux  #( .WIDTH(1) ) _53406_ ( .A(_28488_), .B(1'h0), .S(_06187_), .Y(_28489_) );
  \$mux  #( .WIDTH(1) ) _53407_ ( .A(_28489_), .B(1'h1), .S(_06188_), .Y(_28490_) );
  \$mux  #( .WIDTH(1) ) _53408_ ( .A(_28490_), .B(1'h0), .S(_06190_), .Y(_28491_) );
  \$mux  #( .WIDTH(1) ) _53409_ ( .A(_28491_), .B(1'h1), .S(_06191_), .Y(_28492_) );
  \$mux  #( .WIDTH(1) ) _53410_ ( .A(_28492_), .B(1'h0), .S(_06192_), .Y(_28493_) );
  \$mux  #( .WIDTH(1) ) _53411_ ( .A(_28493_), .B(1'h1), .S(_06193_), .Y(_28494_) );
  \$mux  #( .WIDTH(1) ) _53412_ ( .A(_28494_), .B(maxi_wlast), .S(_06189_), .Y(_28495_) );
  \$mux  #( .WIDTH(1) ) _53413_ ( .A(_28495_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03370_) );
  \$mux  #( .WIDTH(4) ) _53414_ ( .A(maxi_wstrb), .B(4'hf), .S(_06187_), .Y(_28496_) );
  \$mux  #( .WIDTH(4) ) _53415_ ( .A(_28496_), .B(4'hf), .S(_06190_), .Y(_28497_) );
  \$mux  #( .WIDTH(4) ) _53416_ ( .A(_28497_), .B(4'hf), .S(_06192_), .Y(_28498_) );
  \$mux  #( .WIDTH(4) ) _53417_ ( .A(_28498_), .B(4'h0), .S(_RESETN_inv_2), .Y(_03371_) );
  \$mux  #( .WIDTH(32) ) _53418_ ( .A(maxi_wdata), .B(_dataflow_cat_data_98), .S(_06187_), .Y(_28499_) );
  \$mux  #( .WIDTH(32) ) _53419_ ( .A(_28499_), .B(_dataflow_cat_data_107), .S(_06190_), .Y(_28500_) );
  \$mux  #( .WIDTH(32) ) _53420_ ( .A(_28500_), .B(_dataflow_cat_data_167), .S(_06192_), .Y(_28501_) );
  \$mux  #( .WIDTH(32) ) _53421_ ( .A(_28501_), .B(0), .S(_RESETN_inv_2), .Y(_03369_) );
  \$mux  #( .WIDTH(1) ) _53422_ ( .A(maxi_awvalid), .B(1'h0), .S(_saxi_cond_0_1), .Y(_28502_) );
  \$mux  #( .WIDTH(1) ) _53423_ ( .A(_28502_), .B(1'h1), .S(_06184_), .Y(_28503_) );
  \$mux  #( .WIDTH(1) ) _53424_ ( .A(_28503_), .B(1'h0), .S(_06185_), .Y(_28504_) );
  \$mux  #( .WIDTH(1) ) _53425_ ( .A(_28504_), .B(maxi_awvalid), .S(_06186_), .Y(_28505_) );
  \$mux  #( .WIDTH(1) ) _53426_ ( .A(_28505_), .B(1'h0), .S(_RESETN_inv_2), .Y(_03368_) );
  \$mux  #( .WIDTH(8) ) _53427_ ( .A(maxi_awlen), .B(_28534_[7:0]), .S(_06184_), .Y(_28506_) );
  \$mux  #( .WIDTH(8) ) _53428_ ( .A(_28506_), .B(8'h00), .S(_RESETN_inv_2), .Y(_03367_) );
  \$mux  #( .WIDTH(32) ) _53429_ ( .A(maxi_awaddr), .B(_maxi_write_cur_global_addr), .S(_06184_), .Y(_28507_) );
  \$mux  #( .WIDTH(32) ) _53430_ ( .A(_28507_), .B(0), .S(_RESETN_inv_2), .Y(_03366_) );
  \$mux  #( .WIDTH(32) ) _53845_ ( .A(_stream_matmul_29_sink_21_sink_fsm_4), .B({ _13233_, _13232_, _13230_, _13229_, _13228_, _13227_, _13226_, _13225_, _13224_, _13223_, _13222_, _13221_, _13219_, _13218_, _13217_, _13216_, _13215_, _13214_, _13213_, _13212_, _13211_, _13210_, _13240_, _13239_, _13238_, _13237_, _13236_, _13235_, _13234_, _13231_, _13220_, _13209_ }), .S(_24030_), .Y(_24656_) );
  \$mux  #( .WIDTH(32) ) _53846_ ( .A(_stream_matmul_29_source_20_source_pat_fsm_3), .B({ _13297_, _13296_, _13294_, _13293_, _13292_, _13291_, _13290_, _13289_, _13288_, _13287_, _13286_, _13285_, _13283_, _13282_, _13281_, _13280_, _13279_, _13278_, _13277_, _13276_, _13275_, _13274_, _13304_, _13303_, _13302_, _13301_, _13300_, _13299_, _13298_, _13295_, _13284_, _13273_ }), .S(_24031_), .Y(_24657_) );
  \$mux  #( .WIDTH(32) ) _53847_ ( .A(_stream_matmul_29_source_19_source_pat_fsm_2), .B({ _13393_, _13392_, _13390_, _13389_, _13388_, _13387_, _13386_, _13385_, _13384_, _13383_, _13382_, _13381_, _13379_, _13378_, _13377_, _13376_, _13375_, _13374_, _13373_, _13372_, _13371_, _13370_, _13400_, _13399_, _13398_, _13397_, _13396_, _13395_, _13394_, _13391_, _13380_, _13369_ }), .S(_24032_), .Y(_24658_) );
  \$mux  #( .WIDTH(32) ) _53848_ ( .A(_stream_matmul_29_source_8_source_pat_fsm_1), .B({ _13489_, _13488_, _13486_, _13485_, _13484_, _13483_, _13482_, _13481_, _13480_, _13479_, _13478_, _13477_, _13475_, _13474_, _13473_, _13472_, _13471_, _13470_, _13469_, _13468_, _13467_, _13466_, _13496_, _13495_, _13494_, _13493_, _13492_, _13491_, _13490_, _13487_, _13476_, _13465_ }), .S(_24033_), .Y(_24659_) );
  \$mux  #( .WIDTH(32) ) _53849_ ( .A(_stream_matmul_29_source_6_source_pat_fsm_0), .B({ _13585_, _13584_, _13582_, _13581_, _13580_, _13579_, _13578_, _13577_, _13576_, _13575_, _13574_, _13573_, _13571_, _13570_, _13569_, _13568_, _13567_, _13566_, _13565_, _13564_, _13563_, _13562_, _13592_, _13591_, _13590_, _13589_, _13588_, _13587_, _13586_, _13583_, _13572_, _13561_ }), .S(_24034_), .Y(_24660_) );
  \$mux  #( .WIDTH(32) ) _53850_ ( .A(matmul_29_comp_fsm), .B({ _13681_, _13680_, _13678_, _13677_, _13676_, _13675_, _13674_, _13673_, _13672_, _13671_, _13670_, _13669_, _13667_, _13666_, _13665_, _13664_, _13663_, _13662_, _13661_, _13660_, _13659_, _13658_, _13688_, _13687_, _13686_, _13685_, _13684_, _13683_, _13682_, _13679_, _13668_, _13657_ }), .S(_24035_), .Y(_24668_) );
  \$mux  #( .WIDTH(32) ) _53851_ ( .A(matmul_29_stream_out_local_col), .B(0), .S(_24036_), .Y(_24669_) );
  \$mux  #( .WIDTH(32) ) _53852_ ( .A(matmul_29_stream_act_local_0), .B(0), .S(_24036_), .Y(_24670_) );
  \$mux  #( .WIDTH(1) ) _53853_ ( .A(matmul_29_col_select), .B(1'h0), .S(_24036_), .Y(_24671_) );
  \$mux  #( .WIDTH(32) ) _53854_ ( .A(matmul_29_col_count), .B(0), .S(_24036_), .Y(_24672_) );
  \$mux  #( .WIDTH(1) ) _53855_ ( .A(matmul_29_skip_write_out), .B(_13754_), .S(_05515_), .Y(_24696_) );
  \$mux  #( .WIDTH(1) ) _53856_ ( .A(matmul_29_skip_comp), .B(_13757_), .S(_05515_), .Y(_24697_) );
  \$mux  #( .WIDTH(1) ) _53857_ ( .A(matmul_29_skip_read_act), .B(_13755_), .S(_05515_), .Y(_24698_) );
  \$mux  #( .WIDTH(1) ) _53858_ ( .A(matmul_29_skip_read_filter), .B(_13759_), .S(_05515_), .Y(_24699_) );
  \$mux  #( .WIDTH(32) ) _53859_ ( .A(matmul_29_out_laddr_offset), .B({ _05644_, _05643_, _05640_, _05639_, _05642_, _05641_, _05638_, _05637_, _05636_, _05635_, _05634_, _05633_, _05632_, _05631_, _05630_, _05629_, _05628_, _05627_, _05626_, _05625_, _05624_, _05623_, _05622_, _05621_, _05620_, _05619_, _05618_, _05617_, _05616_, _05615_, _05614_, _05613_ }), .S(_24037_), .Y(_24700_) );
  \$mux  #( .WIDTH(32) ) _53860_ ( .A(matmul_29_out_page_dma_offset), .B({ _13880_, _13879_, _13877_, _13876_, _13875_, _13874_, _13873_, _13872_, _13871_, _13870_, _13869_, _13868_, _13866_, _13865_, _13864_, _13863_, _13862_, _13861_, _13860_, _13859_, _13858_, _13857_, _13887_, _13886_, _13885_, _13884_, _13883_, _13882_, _13881_, _13878_, _13867_, _13856_ }), .S(_05515_), .Y(_24701_) );
  \$mux  #( .WIDTH(32) ) _53861_ ( .A(matmul_29_out_page_comp_offset), .B({ _13944_, _13943_, _13941_, _13940_, _13939_, _13938_, _13937_, _13936_, _13935_, _13934_, _13933_, _13932_, _13930_, _13929_, _13928_, _13927_, _13926_, _13925_, _13924_, _13923_, _13922_, _13921_, _13951_, _13950_, _13949_, _13948_, _13947_, _13946_, _13945_, _13942_, _13931_, _13920_ }), .S(_05515_), .Y(_24702_) );
  \$mux  #( .WIDTH(1) ) _53862_ ( .A(matmul_29_out_page), .B(_13953_), .S(_05515_), .Y(_24703_) );
  \$mux  #( .WIDTH(32) ) _53863_ ( .A(matmul_29_filter_page_dma_offset), .B({ _14010_, _14009_, _14007_, _14006_, _14005_, _14004_, _14003_, _14002_, _14001_, _14000_, _13999_, _13998_, _13996_, _13995_, _13994_, _13993_, _13992_, _13991_, _13990_, _13989_, _13988_, _13987_, _14017_, _14016_, _14015_, _14014_, _14013_, _14012_, _14011_, _14008_, _13997_, _13986_ }), .S(_05515_), .Y(_24704_) );
  \$mux  #( .WIDTH(32) ) _53864_ ( .A(matmul_29_filter_page_comp_offset), .B({ _14074_, _14073_, _14071_, _14070_, _14069_, _14068_, _14067_, _14066_, _14065_, _14064_, _14063_, _14062_, _14060_, _14059_, _14058_, _14057_, _14056_, _14055_, _14054_, _14053_, _14052_, _14051_, _14081_, _14080_, _14079_, _14078_, _14077_, _14076_, _14075_, _14072_, _14061_, _14050_ }), .S(_05515_), .Y(_24705_) );
  \$mux  #( .WIDTH(32) ) _53865_ ( .A(matmul_29_act_page_dma_offset_0), .B(0), .S(_05515_), .Y(_24706_) );
  \$mux  #( .WIDTH(32) ) _53866_ ( .A(matmul_29_act_page_comp_offset_0), .B(0), .S(_05515_), .Y(_24707_) );
  \$mux  #( .WIDTH(32) ) _53867_ ( .A(matmul_29_prev_och_count), .B({ _14106_, _14105_, _14103_, _14102_, _14101_, _14100_, _14099_, _14098_, _14097_, _14096_, _14095_, _14094_, _14092_, _14091_, _14090_, _14089_, _14088_, _14087_, _14086_, _14085_, _14084_, _14083_, _14113_, _14112_, _14111_, _14110_, _14109_, _14108_, _14107_, _14104_, _14093_, _14082_ }), .S(_05515_), .Y(_24709_) );
  \$mux  #( .WIDTH(32) ) _53868_ ( .A(matmul_29_prev_bat_count), .B({ _14138_, _14137_, _14135_, _14134_, _14133_, _14132_, _14131_, _14130_, _14129_, _14128_, _14127_, _14126_, _14124_, _14123_, _14122_, _14121_, _14120_, _14119_, _14118_, _14117_, _14116_, _14115_, _14145_, _14144_, _14143_, _14142_, _14141_, _14140_, _14139_, _14136_, _14125_, _14114_ }), .S(_05515_), .Y(_24710_) );
  \$mux  #( .WIDTH(32) ) _53869_ ( .A(matmul_29_prev_row_count), .B({ _14170_, _14169_, _14167_, _14166_, _14165_, _14164_, _14163_, _14162_, _14161_, _14160_, _14159_, _14158_, _14156_, _14155_, _14154_, _14153_, _14152_, _14151_, _14150_, _14149_, _14148_, _14147_, _14177_, _14176_, _14175_, _14174_, _14173_, _14172_, _14171_, _14168_, _14157_, _14146_ }), .S(_05515_), .Y(_24711_) );
  \$mux  #( .WIDTH(32) ) _53870_ ( .A(matmul_29_out_ram_select), .B({ _05610_, _05612_, _05608_, _05611_, _05609_, _05606_, _05607_, _05603_, _05605_, _05604_, _05602_, _05596_, _05601_, _05600_, _05592_, _05599_, _05598_, _05597_, _05590_, _05595_, _05594_, _05593_, _05591_, _05589_, _05588_, _05587_, _05586_, _05581_, _05585_, _05584_, _05583_, _05582_ }), .S(_24037_), .Y(_24712_) );
  \$mux  #( .WIDTH(32) ) _53871_ ( .A(matmul_29_out_row_count), .B({ _14298_, _14297_, _14295_, _14294_, _14293_, _14292_, _14291_, _14290_, _14289_, _14288_, _14287_, _14286_, _14284_, _14283_, _14282_, _14281_, _14280_, _14279_, _14278_, _14277_, _14276_, _14275_, _14305_, _14304_, _14303_, _14302_, _14301_, _14300_, _14299_, _14296_, _14285_, _14274_ }), .S(_05515_), .Y(_24713_) );
  \$mux  #( .WIDTH(32) ) _53872_ ( .A(matmul_29_och_count), .B({ _14330_, _14329_, _14327_, _14326_, _14325_, _14324_, _14323_, _14322_, _14321_, _14320_, _14319_, _14318_, _14316_, _14315_, _14314_, _14313_, _14312_, _14311_, _14310_, _14309_, _14308_, _14307_, _14337_, _14336_, _14335_, _14334_, _14333_, _14332_, _14331_, _14328_, _14317_, _14306_ }), .S(_05515_), .Y(_24715_) );
  \$mux  #( .WIDTH(32) ) _53873_ ( .A(matmul_29_bat_count), .B(0), .S(_05515_), .Y(_24716_) );
  \$mux  #( .WIDTH(32) ) _53874_ ( .A(matmul_29_row_count), .B(0), .S(_05515_), .Y(_24717_) );
  \$mux  #( .WIDTH(32) ) _53875_ ( .A(matmul_29_sync_out_count), .B({ _14394_, _14393_, _14391_, _14390_, _14389_, _14388_, _14387_, _14386_, _14385_, _14384_, _14383_, _14382_, _14380_, _14379_, _14378_, _14377_, _14376_, _14375_, _14374_, _14373_, _14372_, _14371_, _14401_, _14400_, _14399_, _14398_, _14397_, _14396_, _14395_, _14392_, _14381_, _14370_ }), .S(_24038_), .Y(_24719_) );
  \$mux  #( .WIDTH(32) ) _53876_ ( .A(matmul_29_out_base_offset_och), .B({ _14458_, _14457_, _14455_, _14454_, _14453_, _14452_, _14451_, _14450_, _14449_, _14448_, _14447_, _14446_, _14444_, _14443_, _14442_, _14441_, _14440_, _14439_, _14438_, _14437_, _14436_, _14435_, _14465_, _14464_, _14463_, _14462_, _14461_, _14460_, _14459_, _14456_, _14445_, _14434_ }), .S(_05515_), .Y(_24721_) );
  \$mux  #( .WIDTH(32) ) _53877_ ( .A(matmul_29_out_base_offset_bat), .B({ _14522_, _14521_, _14519_, _14518_, _14517_, _14516_, _14515_, _14514_, _14513_, _14512_, _14511_, _14510_, _14508_, _14507_, _14506_, _14505_, _14504_, _14503_, _14502_, _14501_, _14500_, _14499_, _14529_, _14528_, _14527_, _14526_, _14525_, _14524_, _14523_, _14520_, _14509_, _14498_ }), .S(_05515_), .Y(_24722_) );
  \$mux  #( .WIDTH(32) ) _53878_ ( .A(matmul_29_out_base_offset_row), .B({ _14586_, _14585_, _14583_, _14582_, _14581_, _14580_, _14579_, _14578_, _14577_, _14576_, _14575_, _14574_, _14572_, _14571_, _14570_, _14569_, _14568_, _14567_, _14566_, _14565_, _14564_, _14563_, _14593_, _14592_, _14591_, _14590_, _14589_, _14588_, _14587_, _14584_, _14573_, _14562_ }), .S(_05515_), .Y(_24723_) );
  \$mux  #( .WIDTH(32) ) _53879_ ( .A(matmul_29_out_base_offset_col), .B({ _05580_, _05579_, _05578_, _05577_, _05576_, _05575_, _05574_, _05573_, _05572_, _05571_, _05570_, _05569_, _05568_, _05567_, _05566_, _05565_, _05564_, _05563_, _05562_, _05561_, _05560_, _05559_, _05558_, _05557_, _05556_, _05555_, _05554_, _05553_, _05552_, _05551_, _05550_, _05549_ }), .S(_24037_), .Y(_24724_) );
  \$mux  #( .WIDTH(32) ) _53880_ ( .A(matmul_29_filter_base_offset), .B({ _14682_, _14681_, _14679_, _14678_, _14677_, _14676_, _14675_, _14674_, _14673_, _14672_, _14671_, _14670_, _14668_, _14667_, _14666_, _14665_, _14664_, _14663_, _14662_, _14661_, _14660_, _14659_, _14689_, _14688_, _14687_, _14686_, _14685_, _14684_, _14683_, _14680_, _14669_, _14658_ }), .S(_05515_), .Y(_24726_) );
  \$mux  #( .WIDTH(32) ) _53881_ ( .A(matmul_29_act_base_offset_bat), .B(0), .S(_05515_), .Y(_24727_) );
  \$mux  #( .WIDTH(32) ) _53882_ ( .A(matmul_29_act_base_offset_row), .B(0), .S(_05515_), .Y(_24728_) );
  \$mux  #( .WIDTH(32) ) _53883_ ( .A(control_matmul_29), .B({ _14746_, _14745_, _14743_, _14742_, _14741_, _14740_, _14739_, _14738_, _14737_, _14736_, _14735_, _14734_, _14732_, _14731_, _14730_, _14729_, _14728_, _14727_, _14726_, _14725_, _14724_, _14723_, _14753_, _14752_, _14751_, _14750_, _14749_, _14748_, _14747_, _14744_, _14733_, _14722_ }), .S(_24039_), .Y(_24731_) );
  \$mux  #( .WIDTH(32) ) _53884_ ( .A(_stream_max_pool_serial_18_sink_3_sink_fsm_1), .B({ _15322_, _15321_, _15319_, _15318_, _15317_, _15316_, _15315_, _15314_, _15313_, _15312_, _15311_, _15310_, _15308_, _15307_, _15306_, _15305_, _15304_, _15303_, _15302_, _15301_, _15300_, _15299_, _15329_, _15328_, _15327_, _15326_, _15325_, _15324_, _15323_, _15320_, _15309_, _15298_ }), .S(_24040_), .Y(_24738_) );
  \$mux  #( .WIDTH(32) ) _53885_ ( .A(_stream_max_pool_serial_18_source_1_source_pat_fsm_0), .B({ _15386_, _15385_, _15383_, _15382_, _15381_, _15380_, _15379_, _15378_, _15377_, _15376_, _15375_, _15374_, _15372_, _15371_, _15370_, _15369_, _15368_, _15367_, _15366_, _15365_, _15364_, _15363_, _15393_, _15392_, _15391_, _15390_, _15389_, _15388_, _15387_, _15384_, _15373_, _15362_ }), .S(_24041_), .Y(_24739_) );
  \$mux  #( .WIDTH(32) ) _53886_ ( .A(max_pool_serial_18_comp_fsm), .B({ _15514_, _15513_, _15511_, _15510_, _15509_, _15508_, _15507_, _15506_, _15505_, _15504_, _15503_, _15502_, _15500_, _15499_, _15498_, _15497_, _15496_, _15495_, _15494_, _15493_, _15492_, _15491_, _15521_, _15520_, _15519_, _15518_, _15517_, _15516_, _15515_, _15512_, _15501_, _15490_ }), .S(_24042_), .Y(_24744_) );
  \$mux  #( .WIDTH(32) ) _53887_ ( .A(max_pool_serial_18_stream_out_local), .B({ _15642_, _15641_, _15639_, _15638_, _15637_, _15636_, _15635_, _15634_, _15633_, _15632_, _15631_, _15630_, _15628_, _15627_, _15626_, _15625_, _15624_, _15623_, _15622_, _15621_, _15620_, _15619_, _15649_, _15648_, _15647_, _15646_, _15645_, _15644_, _15643_, _15640_, _15629_, _15618_ }), .S(_24043_), .Y(_24747_) );
  \$mux  #( .WIDTH(32) ) _53888_ ( .A(max_pool_serial_18_stream_act_local), .B({ _15706_, _15705_, _15703_, _15702_, _15701_, _15700_, _15699_, _15698_, _15697_, _15696_, _15695_, _15694_, _15692_, _15691_, _15690_, _15689_, _15688_, _15687_, _15686_, _15685_, _15684_, _15683_, _15713_, _15712_, _15711_, _15710_, _15709_, _15708_, _15707_, _15704_, _15693_, _15682_ }), .S(_24043_), .Y(_24748_) );
  \$mux  #( .WIDTH(32) ) _53889_ ( .A(max_pool_serial_18_col_count), .B({ _15770_, _15769_, _15767_, _15766_, _15765_, _15764_, _15763_, _15762_, _15761_, _15760_, _15759_, _15758_, _15756_, _15755_, _15754_, _15753_, _15752_, _15751_, _15750_, _15749_, _15748_, _15747_, _15777_, _15776_, _15775_, _15774_, _15773_, _15772_, _15771_, _15768_, _15757_, _15746_ }), .S(_24043_), .Y(_24749_) );
  \$mux  #( .WIDTH(32) ) _53890_ ( .A(max_pool_serial_18_out_count), .B({ _15802_, _15801_, _15799_, _15798_, _15797_, _15796_, _15795_, _15794_, _15793_, _15792_, _15791_, _15790_, _15788_, _15787_, _15786_, _15785_, _15784_, _15783_, _15782_, _15781_, _15780_, _15779_, _15809_, _15808_, _15807_, _15806_, _15805_, _15804_, _15803_, _15800_, _15789_, _15778_ }), .S(_24044_), .Y(_24762_) );
  \$mux  #( .WIDTH(1) ) _53891_ ( .A(max_pool_serial_18_skip_write_out), .B(_15811_), .S(_24045_), .Y(_24763_) );
  \$mux  #( .WIDTH(1) ) _53892_ ( .A(max_pool_serial_18_skip_comp), .B(_15813_), .S(_24045_), .Y(_24764_) );
  \$mux  #( .WIDTH(1) ) _53893_ ( .A(max_pool_serial_18_skip_read_act), .B(_15815_), .S(_24045_), .Y(_24765_) );
  \$mux  #( .WIDTH(32) ) _53894_ ( .A(max_pool_serial_18_out_page_dma_offset), .B({ _15872_, _15871_, _15869_, _15868_, _15867_, _15866_, _15865_, _15864_, _15863_, _15862_, _15861_, _15860_, _15858_, _15857_, _15856_, _15855_, _15854_, _15853_, _15852_, _15851_, _15850_, _15849_, _15879_, _15878_, _15877_, _15876_, _15875_, _15874_, _15873_, _15870_, _15859_, _15848_ }), .S(_24045_), .Y(_24766_) );
  \$mux  #( .WIDTH(32) ) _53895_ ( .A(max_pool_serial_18_out_page_comp_offset), .B({ _15936_, _15935_, _15933_, _15932_, _15931_, _15930_, _15929_, _15928_, _15927_, _15926_, _15925_, _15924_, _15922_, _15921_, _15920_, _15919_, _15918_, _15917_, _15916_, _15915_, _15914_, _15913_, _15943_, _15942_, _15941_, _15940_, _15939_, _15938_, _15937_, _15934_, _15923_, _15912_ }), .S(_24045_), .Y(_24767_) );
  \$mux  #( .WIDTH(1) ) _53896_ ( .A(max_pool_serial_18_out_page), .B(_15945_), .S(_24045_), .Y(_24768_) );
  \$mux  #( .WIDTH(32) ) _53897_ ( .A(max_pool_serial_18_act_page_dma_offset), .B({ _16002_, _16001_, _15999_, _15998_, _15997_, _15996_, _15995_, _15994_, _15993_, _15992_, _15991_, _15990_, _15988_, _15987_, _15986_, _15985_, _15984_, _15983_, _15982_, _15981_, _15980_, _15979_, _16009_, _16008_, _16007_, _16006_, _16005_, _16004_, _16003_, _16000_, _15989_, _15978_ }), .S(_24045_), .Y(_24769_) );
  \$mux  #( .WIDTH(32) ) _53898_ ( .A(max_pool_serial_18_act_page_comp_offset), .B({ _16002_, _16001_, _15999_, _15998_, _15997_, _15996_, _15995_, _15994_, _15993_, _15992_, _15991_, _15990_, _15988_, _15987_, _15986_, _15985_, _15984_, _15983_, _15982_, _15981_, _15980_, _15979_, _16009_, _16008_, _16007_, _16006_, _16005_, _16004_, _16003_, _16000_, _15989_, _15978_ }), .S(_24045_), .Y(_24770_) );
  \$mux  #( .WIDTH(1) ) _53899_ ( .A(max_pool_serial_18_act_page), .B(_16011_), .S(_24045_), .Y(_24771_) );
  \$mux  #( .WIDTH(32) ) _53900_ ( .A(max_pool_serial_18_prev_bat_count), .B({ _16036_, _16035_, _16033_, _16032_, _16031_, _16030_, _16029_, _16028_, _16027_, _16026_, _16025_, _16024_, _16022_, _16021_, _16020_, _16019_, _16018_, _16017_, _16016_, _16015_, _16014_, _16013_, _16043_, _16042_, _16041_, _16040_, _16039_, _16038_, _16037_, _16034_, _16023_, _16012_ }), .S(_24045_), .Y(_24772_) );
  \$mux  #( .WIDTH(32) ) _53901_ ( .A(max_pool_serial_18_prev_row_count), .B({ _16068_, _16067_, _16065_, _16064_, _16063_, _16062_, _16061_, _16060_, _16059_, _16058_, _16057_, _16056_, _16054_, _16053_, _16052_, _16051_, _16050_, _16049_, _16048_, _16047_, _16046_, _16045_, _16075_, _16074_, _16073_, _16072_, _16071_, _16070_, _16069_, _16066_, _16055_, _16044_ }), .S(_24045_), .Y(_24773_) );
  \$mux  #( .WIDTH(32) ) _53902_ ( .A(max_pool_serial_18_bat_count), .B({ _16132_, _16131_, _16129_, _16128_, _16127_, _16126_, _16125_, _16124_, _16123_, _16122_, _16121_, _16120_, _16118_, _16117_, _16116_, _16115_, _16114_, _16113_, _16112_, _16111_, _16110_, _16109_, _16139_, _16138_, _16137_, _16136_, _16135_, _16134_, _16133_, _16130_, _16119_, _16108_ }), .S(_24045_), .Y(_24774_) );
  \$mux  #( .WIDTH(32) ) _53903_ ( .A(max_pool_serial_18_row_count), .B({ _16196_, _16195_, _16193_, _16192_, _16191_, _16190_, _16189_, _16188_, _16187_, _16186_, _16185_, _16184_, _16182_, _16181_, _16180_, _16179_, _16178_, _16177_, _16176_, _16175_, _16174_, _16173_, _16203_, _16202_, _16201_, _16200_, _16199_, _16198_, _16197_, _16194_, _16183_, _16172_ }), .S(_24045_), .Y(_24775_) );
  \$mux  #( .WIDTH(32) ) _53904_ ( .A(max_pool_serial_18_out_base_offset_bat), .B({ _16260_, _16259_, _16257_, _16256_, _16255_, _16254_, _16253_, _16252_, _16251_, _16250_, _16249_, _16248_, _16246_, _16245_, _16244_, _16243_, _16242_, _16241_, _16240_, _16239_, _16238_, _16237_, _16267_, _16266_, _16265_, _16264_, _16263_, _16262_, _16261_, _16258_, _16247_, _16236_ }), .S(_24045_), .Y(_24776_) );
  \$mux  #( .WIDTH(32) ) _53905_ ( .A(max_pool_serial_18_out_base_offset_row), .B({ _16324_, _16323_, _16321_, _16320_, _16319_, _16318_, _16317_, _16316_, _16315_, _16314_, _16313_, _16312_, _16310_, _16309_, _16308_, _16307_, _16306_, _16305_, _16304_, _16303_, _16302_, _16301_, _16331_, _16330_, _16329_, _16328_, _16327_, _16326_, _16325_, _16322_, _16311_, _16300_ }), .S(_24045_), .Y(_24778_) );
  \$mux  #( .WIDTH(32) ) _53906_ ( .A(max_pool_serial_18_act_base_offset_bat), .B({ _16388_, _16387_, _16385_, _16384_, _16383_, _16382_, _16381_, _16380_, _16379_, _16378_, _16377_, _16376_, _16374_, _16373_, _16372_, _16371_, _16370_, _16369_, _16368_, _16367_, _16366_, _16365_, _16395_, _16394_, _16393_, _16392_, _16391_, _16390_, _16389_, _16386_, _16375_, _16364_ }), .S(_24045_), .Y(_24779_) );
  \$mux  #( .WIDTH(32) ) _53907_ ( .A(max_pool_serial_18_act_base_offset_row), .B({ _16452_, _16451_, _16449_, _16448_, _16447_, _16446_, _16445_, _16444_, _16443_, _16442_, _16441_, _16440_, _16438_, _16437_, _16436_, _16435_, _16434_, _16433_, _16432_, _16431_, _16430_, _16429_, _16459_, _16458_, _16457_, _16456_, _16455_, _16454_, _16453_, _16450_, _16439_, _16428_ }), .S(_24045_), .Y(_24780_) );
  \$mux  #( .WIDTH(32) ) _53908_ ( .A(control_max_pool_serial_18), .B({ _16516_, _16515_, _16513_, _16512_, _16511_, _16510_, _16509_, _16508_, _16507_, _16506_, _16505_, _16504_, _16502_, _16501_, _16500_, _16499_, _16498_, _16497_, _16496_, _16495_, _16494_, _16493_, _16523_, _16522_, _16521_, _16520_, _16519_, _16518_, _16517_, _16514_, _16503_, _16492_ }), .S(_24046_), .Y(_24783_) );
  \$mux  #( .WIDTH(33) ) _53909_ ( .A(_maxi_write_rest_size), .B({ _16966_, _16965_, _16964_, _16962_, _16961_, _16960_, _16959_, _16958_, _16957_, _16956_, _16955_, _16954_, _16953_, _16951_, _16950_, _16949_, _16948_, _16947_, _16946_, _16945_, _16944_, _16943_, _16942_, _16973_, _16972_, _16971_, _16970_, _16969_, _16968_, _16967_, _16963_, _16952_, _16941_ }), .S(_05516_), .Y(_24794_) );
  \$mux  #( .WIDTH(32) ) _53910_ ( .A(_maxi_write_cur_global_addr), .B({ _17063_, _17062_, _17060_, _17059_, _17058_, _17057_, _17056_, _17055_, _17054_, _17053_, _17052_, _17051_, _17049_, _17048_, _17047_, _17046_, _17045_, _17044_, _17043_, _17042_, _17041_, _17040_, _17070_, _17069_, _17068_, _17067_, _17066_, _17065_, _17064_, _17061_, _17050_, _17039_ }), .S(_24047_), .Y(_24799_) );
  \$mux  #( .WIDTH(32) ) _53911_ ( .A(_maxi_write_fsm), .B({ _17127_, _17126_, _17124_, _17123_, _17122_, _17121_, _17120_, _17119_, _17118_, _17117_, _17116_, _17115_, _17113_, _17112_, _17111_, _17110_, _17109_, _17108_, _17107_, _17106_, _17105_, _17104_, _17134_, _17133_, _17132_, _17131_, _17130_, _17129_, _17128_, _17125_, _17114_, _17103_ }), .S(_24048_), .Y(_24800_) );
  \$mux  #( .WIDTH(32) ) _53912_ ( .A(_stream_conv2d_16_sink_37_sink_fsm_20), .B({ _17287_, _17286_, _17284_, _17283_, _17282_, _17281_, _17280_, _17279_, _17278_, _17277_, _17276_, _17275_, _17273_, _17272_, _17271_, _17270_, _17269_, _17268_, _17267_, _17266_, _17265_, _17264_, _17294_, _17293_, _17292_, _17291_, _17290_, _17289_, _17288_, _17285_, _17274_, _17263_ }), .S(_24049_), .Y(_24805_) );
  \$mux  #( .WIDTH(32) ) _53913_ ( .A(_stream_conv2d_16_source_36_source_pat_fsm_19), .B({ _17351_, _17350_, _17348_, _17347_, _17346_, _17345_, _17344_, _17343_, _17342_, _17341_, _17340_, _17339_, _17337_, _17336_, _17335_, _17334_, _17333_, _17332_, _17331_, _17330_, _17329_, _17328_, _17358_, _17357_, _17356_, _17355_, _17354_, _17353_, _17352_, _17349_, _17338_, _17327_ }), .S(_24050_), .Y(_24806_) );
  \$mux  #( .WIDTH(32) ) _53914_ ( .A(_stream_conv2d_16_source_35_source_pat_fsm_18), .B({ _17447_, _17446_, _17444_, _17443_, _17442_, _17441_, _17440_, _17439_, _17438_, _17437_, _17436_, _17435_, _17433_, _17432_, _17431_, _17430_, _17429_, _17428_, _17427_, _17426_, _17425_, _17424_, _17454_, _17453_, _17452_, _17451_, _17450_, _17449_, _17448_, _17445_, _17434_, _17423_ }), .S(_24051_), .Y(_24807_) );
  \$mux  #( .WIDTH(32) ) _53915_ ( .A(_stream_conv2d_16_source_34_source_pat_fsm_17), .B({ _17543_, _17542_, _17540_, _17539_, _17538_, _17537_, _17536_, _17535_, _17534_, _17533_, _17532_, _17531_, _17529_, _17528_, _17527_, _17526_, _17525_, _17524_, _17523_, _17522_, _17521_, _17520_, _17550_, _17549_, _17548_, _17547_, _17546_, _17545_, _17544_, _17541_, _17530_, _17519_ }), .S(_24052_), .Y(_24808_) );
  \$mux  #( .WIDTH(32) ) _53916_ ( .A(_stream_conv2d_16_source_33_source_pat_fsm_16), .B({ _17639_, _17638_, _17636_, _17635_, _17634_, _17633_, _17632_, _17631_, _17630_, _17629_, _17628_, _17627_, _17625_, _17624_, _17623_, _17622_, _17621_, _17620_, _17619_, _17618_, _17617_, _17616_, _17646_, _17645_, _17644_, _17643_, _17642_, _17641_, _17640_, _17637_, _17626_, _17615_ }), .S(_24053_), .Y(_24809_) );
  \$mux  #( .WIDTH(32) ) _53917_ ( .A(_stream_conv2d_16_source_32_source_pat_fsm_15), .B({ _17735_, _17734_, _17732_, _17731_, _17730_, _17729_, _17728_, _17727_, _17726_, _17725_, _17724_, _17723_, _17721_, _17720_, _17719_, _17718_, _17717_, _17716_, _17715_, _17714_, _17713_, _17712_, _17742_, _17741_, _17740_, _17739_, _17738_, _17737_, _17736_, _17733_, _17722_, _17711_ }), .S(_24054_), .Y(_24810_) );
  \$mux  #( .WIDTH(32) ) _53918_ ( .A(_stream_conv2d_16_source_31_source_pat_fsm_14), .B({ _17831_, _17830_, _17828_, _17827_, _17826_, _17825_, _17824_, _17823_, _17822_, _17821_, _17820_, _17819_, _17817_, _17816_, _17815_, _17814_, _17813_, _17812_, _17811_, _17810_, _17809_, _17808_, _17838_, _17837_, _17836_, _17835_, _17834_, _17833_, _17832_, _17829_, _17818_, _17807_ }), .S(_24055_), .Y(_24811_) );
  \$mux  #( .WIDTH(32) ) _53919_ ( .A(_stream_conv2d_16_source_30_source_pat_fsm_13), .B({ _17927_, _17926_, _17924_, _17923_, _17922_, _17921_, _17920_, _17919_, _17918_, _17917_, _17916_, _17915_, _17913_, _17912_, _17911_, _17910_, _17909_, _17908_, _17907_, _17906_, _17905_, _17904_, _17934_, _17933_, _17932_, _17931_, _17930_, _17929_, _17928_, _17925_, _17914_, _17903_ }), .S(_24056_), .Y(_24812_) );
  \$mux  #( .WIDTH(32) ) _53920_ ( .A(_stream_conv2d_16_source_29_source_pat_fsm_12), .B({ _18023_, _18022_, _18020_, _18019_, _18018_, _18017_, _18016_, _18015_, _18014_, _18013_, _18012_, _18011_, _18009_, _18008_, _18007_, _18006_, _18005_, _18004_, _18003_, _18002_, _18001_, _18000_, _18030_, _18029_, _18028_, _18027_, _18026_, _18025_, _18024_, _18021_, _18010_, _17999_ }), .S(_24057_), .Y(_24813_) );
  \$mux  #( .WIDTH(32) ) _53921_ ( .A(_stream_conv2d_16_source_28_source_pat_fsm_11), .B({ _18119_, _18118_, _18116_, _18115_, _18114_, _18113_, _18112_, _18111_, _18110_, _18109_, _18108_, _18107_, _18105_, _18104_, _18103_, _18102_, _18101_, _18100_, _18099_, _18098_, _18097_, _18096_, _18126_, _18125_, _18124_, _18123_, _18122_, _18121_, _18120_, _18117_, _18106_, _18095_ }), .S(_24058_), .Y(_24814_) );
  \$mux  #( .WIDTH(32) ) _53922_ ( .A(_stream_conv2d_16_source_27_source_pat_fsm_10), .B({ _18215_, _18214_, _18212_, _18211_, _18210_, _18209_, _18208_, _18207_, _18206_, _18205_, _18204_, _18203_, _18201_, _18200_, _18199_, _18198_, _18197_, _18196_, _18195_, _18194_, _18193_, _18192_, _18222_, _18221_, _18220_, _18219_, _18218_, _18217_, _18216_, _18213_, _18202_, _18191_ }), .S(_24059_), .Y(_24815_) );
  \$mux  #( .WIDTH(32) ) _53923_ ( .A(_stream_conv2d_16_source_26_source_pat_fsm_9), .B({ _18311_, _18310_, _18308_, _18307_, _18306_, _18305_, _18304_, _18303_, _18302_, _18301_, _18300_, _18299_, _18297_, _18296_, _18295_, _18294_, _18293_, _18292_, _18291_, _18290_, _18289_, _18288_, _18318_, _18317_, _18316_, _18315_, _18314_, _18313_, _18312_, _18309_, _18298_, _18287_ }), .S(_24060_), .Y(_24816_) );
  \$mux  #( .WIDTH(32) ) _53924_ ( .A(_stream_conv2d_16_source_25_source_pat_fsm_8), .B({ _18407_, _18406_, _18404_, _18403_, _18402_, _18401_, _18400_, _18399_, _18398_, _18397_, _18396_, _18395_, _18393_, _18392_, _18391_, _18390_, _18389_, _18388_, _18387_, _18386_, _18385_, _18384_, _18414_, _18413_, _18412_, _18411_, _18410_, _18409_, _18408_, _18405_, _18394_, _18383_ }), .S(_24061_), .Y(_24817_) );
  \$mux  #( .WIDTH(32) ) _53925_ ( .A(_stream_conv2d_16_source_24_source_pat_fsm_7), .B({ _18503_, _18502_, _18500_, _18499_, _18498_, _18497_, _18496_, _18495_, _18494_, _18493_, _18492_, _18491_, _18489_, _18488_, _18487_, _18486_, _18485_, _18484_, _18483_, _18482_, _18481_, _18480_, _18510_, _18509_, _18508_, _18507_, _18506_, _18505_, _18504_, _18501_, _18490_, _18479_ }), .S(_24062_), .Y(_24818_) );
  \$mux  #( .WIDTH(32) ) _53926_ ( .A(_stream_conv2d_16_source_23_source_pat_fsm_6), .B({ _18599_, _18598_, _18596_, _18595_, _18594_, _18593_, _18592_, _18591_, _18590_, _18589_, _18588_, _18587_, _18585_, _18584_, _18583_, _18582_, _18581_, _18580_, _18579_, _18578_, _18577_, _18576_, _18606_, _18605_, _18604_, _18603_, _18602_, _18601_, _18600_, _18597_, _18586_, _18575_ }), .S(_24063_), .Y(_24819_) );
  \$mux  #( .WIDTH(32) ) _53927_ ( .A(_stream_conv2d_16_source_22_source_pat_fsm_5), .B({ _18695_, _18694_, _18692_, _18691_, _18690_, _18689_, _18688_, _18687_, _18686_, _18685_, _18684_, _18683_, _18681_, _18680_, _18679_, _18678_, _18677_, _18676_, _18675_, _18674_, _18673_, _18672_, _18702_, _18701_, _18700_, _18699_, _18698_, _18697_, _18696_, _18693_, _18682_, _18671_ }), .S(_24064_), .Y(_24820_) );
  \$mux  #( .WIDTH(32) ) _53928_ ( .A(_stream_conv2d_16_source_21_source_pat_fsm_4), .B({ _18791_, _18790_, _18788_, _18787_, _18786_, _18785_, _18784_, _18783_, _18782_, _18781_, _18780_, _18779_, _18777_, _18776_, _18775_, _18774_, _18773_, _18772_, _18771_, _18770_, _18769_, _18768_, _18798_, _18797_, _18796_, _18795_, _18794_, _18793_, _18792_, _18789_, _18778_, _18767_ }), .S(_24065_), .Y(_24821_) );
  \$mux  #( .WIDTH(32) ) _53929_ ( .A(_stream_conv2d_16_source_20_source_pat_fsm_3), .B({ _18887_, _18886_, _18884_, _18883_, _18882_, _18881_, _18880_, _18879_, _18878_, _18877_, _18876_, _18875_, _18873_, _18872_, _18871_, _18870_, _18869_, _18868_, _18867_, _18866_, _18865_, _18864_, _18894_, _18893_, _18892_, _18891_, _18890_, _18889_, _18888_, _18885_, _18874_, _18863_ }), .S(_24066_), .Y(_24822_) );
  \$mux  #( .WIDTH(32) ) _53930_ ( .A(_stream_conv2d_16_source_19_source_pat_fsm_2), .B({ _18983_, _18982_, _18980_, _18979_, _18978_, _18977_, _18976_, _18975_, _18974_, _18973_, _18972_, _18971_, _18969_, _18968_, _18967_, _18966_, _18965_, _18964_, _18963_, _18962_, _18961_, _18960_, _18990_, _18989_, _18988_, _18987_, _18986_, _18985_, _18984_, _18981_, _18970_, _18959_ }), .S(_24067_), .Y(_24823_) );
  \$mux  #( .WIDTH(32) ) _53931_ ( .A(_stream_conv2d_16_source_8_source_pat_fsm_1), .B({ _19079_, _19078_, _19076_, _19075_, _19074_, _19073_, _19072_, _19071_, _19070_, _19069_, _19068_, _19067_, _19065_, _19064_, _19063_, _19062_, _19061_, _19060_, _19059_, _19058_, _19057_, _19056_, _19086_, _19085_, _19084_, _19083_, _19082_, _19081_, _19080_, _19077_, _19066_, _19055_ }), .S(_24068_), .Y(_24824_) );
  \$mux  #( .WIDTH(32) ) _53932_ ( .A(_stream_conv2d_16_source_6_source_pat_fsm_0), .B({ _19175_, _19174_, _19172_, _19171_, _19170_, _19169_, _19168_, _19167_, _19166_, _19165_, _19164_, _19163_, _19161_, _19160_, _19159_, _19158_, _19157_, _19156_, _19155_, _19154_, _19153_, _19152_, _19182_, _19181_, _19180_, _19179_, _19178_, _19177_, _19176_, _19173_, _19162_, _19151_ }), .S(_24069_), .Y(_24825_) );
  \$mux  #( .WIDTH(32) ) _53933_ ( .A(conv2d_16_comp_fsm), .B({ _19303_, _19302_, _19300_, _19299_, _19298_, _19297_, _19296_, _19295_, _19294_, _19293_, _19292_, _19291_, _19289_, _19288_, _19287_, _19286_, _19285_, _19284_, _19283_, _19282_, _19281_, _19280_, _19310_, _19309_, _19308_, _19307_, _19306_, _19305_, _19304_, _19301_, _19290_, _19279_ }), .S(_24070_), .Y(_24835_) );
  \$mux  #( .WIDTH(32) ) _53934_ ( .A(conv2d_16_stream_out_local_col), .B({ _19431_, _19430_, _19428_, _19427_, _19426_, _19425_, _19424_, _19423_, _19422_, _19421_, _19420_, _19419_, _19417_, _19416_, _19415_, _19414_, _19413_, _19412_, _19411_, _19410_, _19409_, _19408_, _19438_, _19437_, _19436_, _19435_, _19434_, _19433_, _19432_, _19429_, _19418_, _19407_ }), .S(_24071_), .Y(_24836_) );
  \$mux  #( .WIDTH(32) ) _53935_ ( .A(conv2d_16_stream_act_local_8), .B({ _19496_, _19495_, _19493_, _19492_, _19491_, _19490_, _19489_, _19488_, _19487_, _19486_, _19485_, _19484_, _19482_, _19481_, _19480_, _19479_, _19478_, _19477_, _19476_, _19475_, _19474_, _19473_, _19503_, _19502_, _19501_, _19500_, _19499_, _19498_, _19497_, _19494_, _19483_, _19472_ }), .S(_24071_), .Y(_24838_) );
  \$mux  #( .WIDTH(32) ) _53936_ ( .A(conv2d_16_stream_act_local_7), .B({ _19561_, _19560_, _19558_, _19557_, _19556_, _19555_, _19554_, _19553_, _19552_, _19551_, _19550_, _19549_, _19547_, _19546_, _19545_, _19544_, _19543_, _19542_, _19541_, _19540_, _19539_, _19538_, _19568_, _19567_, _19566_, _19565_, _19564_, _19563_, _19562_, _19559_, _19548_, _19537_ }), .S(_24071_), .Y(_24840_) );
  \$mux  #( .WIDTH(32) ) _53937_ ( .A(conv2d_16_stream_act_local_6), .B({ _19626_, _19625_, _19623_, _19622_, _19621_, _19620_, _19619_, _19618_, _19617_, _19616_, _19615_, _19614_, _19612_, _19611_, _19610_, _19609_, _19608_, _19607_, _19606_, _19605_, _19604_, _19603_, _19633_, _19632_, _19631_, _19630_, _19629_, _19628_, _19627_, _19624_, _19613_, _19602_ }), .S(_24071_), .Y(_24842_) );
  \$mux  #( .WIDTH(32) ) _53938_ ( .A(conv2d_16_stream_act_local_5), .B({ _19690_, _19689_, _19687_, _19686_, _19685_, _19684_, _19683_, _19682_, _19681_, _19680_, _19679_, _19678_, _19676_, _19675_, _19674_, _19673_, _19672_, _19671_, _19670_, _19669_, _19668_, _19667_, _19697_, _19696_, _19695_, _19694_, _19693_, _19692_, _19691_, _19688_, _19677_, _19666_ }), .S(_24071_), .Y(_24844_) );
  \$mux  #( .WIDTH(32) ) _53939_ ( .A(conv2d_16_stream_act_local_4), .B({ _19754_, _19753_, _19751_, _19750_, _19749_, _19748_, _19747_, _19746_, _19745_, _19744_, _19743_, _19742_, _19740_, _19739_, _19738_, _19737_, _19736_, _19735_, _19734_, _19733_, _19732_, _19731_, _19761_, _19760_, _19759_, _19758_, _19757_, _19756_, _19755_, _19752_, _19741_, _19730_ }), .S(_24071_), .Y(_24846_) );
  \$mux  #( .WIDTH(32) ) _53940_ ( .A(conv2d_16_stream_act_local_3), .B({ _19818_, _19817_, _19815_, _19814_, _19813_, _19812_, _19811_, _19810_, _19809_, _19808_, _19807_, _19806_, _19804_, _19803_, _19802_, _19801_, _19800_, _19799_, _19798_, _19797_, _19796_, _19795_, _19825_, _19824_, _19823_, _19822_, _19821_, _19820_, _19819_, _19816_, _19805_, _19794_ }), .S(_24071_), .Y(_24848_) );
  \$mux  #( .WIDTH(32) ) _53941_ ( .A(conv2d_16_stream_act_local_2), .B({ _19882_, _19881_, _19879_, _19878_, _19877_, _19876_, _19875_, _19874_, _19873_, _19872_, _19871_, _19870_, _19868_, _19867_, _19866_, _19865_, _19864_, _19863_, _19862_, _19861_, _19860_, _19859_, _19889_, _19888_, _19887_, _19886_, _19885_, _19884_, _19883_, _19880_, _19869_, _19858_ }), .S(_24071_), .Y(_24850_) );
  \$mux  #( .WIDTH(32) ) _53942_ ( .A(conv2d_16_stream_act_local_1), .B({ _19946_, _19945_, _19943_, _19942_, _19941_, _19940_, _19939_, _19938_, _19937_, _19936_, _19935_, _19934_, _19932_, _19931_, _19930_, _19929_, _19928_, _19927_, _19926_, _19925_, _19924_, _19923_, _19953_, _19952_, _19951_, _19950_, _19949_, _19948_, _19947_, _19944_, _19933_, _19922_ }), .S(_24071_), .Y(_24852_) );
  \$mux  #( .WIDTH(32) ) _53943_ ( .A(conv2d_16_stream_act_local_0), .B({ _20010_, _20009_, _20007_, _20006_, _20005_, _20004_, _20003_, _20002_, _20001_, _20000_, _19999_, _19998_, _19996_, _19995_, _19994_, _19993_, _19992_, _19991_, _19990_, _19989_, _19988_, _19987_, _20017_, _20016_, _20015_, _20014_, _20013_, _20012_, _20011_, _20008_, _19997_, _19986_ }), .S(_24071_), .Y(_24854_) );
  \$mux  #( .WIDTH(2) ) _53944_ ( .A(conv2d_16_col_select), .B({ _20021_, _20020_ }), .S(_24071_), .Y(_24856_) );
  \$mux  #( .WIDTH(32) ) _53945_ ( .A(conv2d_16_col_count), .B({ _20078_, _20077_, _20075_, _20074_, _20073_, _20072_, _20071_, _20070_, _20069_, _20068_, _20067_, _20066_, _20064_, _20063_, _20062_, _20061_, _20060_, _20059_, _20058_, _20057_, _20056_, _20055_, _20085_, _20084_, _20083_, _20082_, _20081_, _20080_, _20079_, _20076_, _20065_, _20054_ }), .S(_24071_), .Y(_24857_) );
  \$mux  #( .WIDTH(33) ) _53946_ ( .A(_maxi_read_rest_size), .B({ _20144_, _20143_, _20142_, _20140_, _20139_, _20138_, _20137_, _20136_, _20135_, _20134_, _20133_, _20132_, _20131_, _20129_, _20128_, _20127_, _20126_, _20125_, _20124_, _20123_, _20122_, _20121_, _20120_, _20151_, _20150_, _20149_, _20148_, _20147_, _20146_, _20145_, _20141_, _20130_, _20119_ }), .S(_05658_), .Y(_24934_) );
  \$mux  #( .WIDTH(32) ) _53947_ ( .A(_maxi_read_cur_global_addr), .B({ _20241_, _20240_, _20238_, _20237_, _20236_, _20235_, _20234_, _20233_, _20232_, _20231_, _20230_, _20229_, _20227_, _20226_, _20225_, _20224_, _20223_, _20222_, _20221_, _20220_, _20219_, _20218_, _20248_, _20247_, _20246_, _20245_, _20244_, _20243_, _20242_, _20239_, _20228_, _20217_ }), .S(_24072_), .Y(_24939_) );
  \$mux  #( .WIDTH(32) ) _53948_ ( .A(_maxi_read_fsm), .B({ _20305_, _20304_, _20302_, _20301_, _20300_, _20299_, _20298_, _20297_, _20296_, _20295_, _20294_, _20293_, _20291_, _20290_, _20289_, _20288_, _20287_, _20286_, _20285_, _20284_, _20283_, _20282_, _20312_, _20311_, _20310_, _20309_, _20308_, _20307_, _20306_, _20303_, _20292_, _20281_ }), .S(_24073_), .Y(_24940_) );
  \$mux  #( .WIDTH(1) ) _53949_ ( .A(conv2d_16_skip_write_out), .B(_20410_), .S(_05514_), .Y(_24994_) );
  \$mux  #( .WIDTH(1) ) _53950_ ( .A(conv2d_16_skip_comp), .B(_20412_), .S(_05514_), .Y(_24995_) );
  \$mux  #( .WIDTH(1) ) _53951_ ( .A(conv2d_16_skip_read_act), .B(_20414_), .S(_05514_), .Y(_24996_) );
  \$mux  #( .WIDTH(1) ) _53952_ ( .A(conv2d_16_skip_read_filter), .B(_20416_), .S(_05514_), .Y(_24997_) );
  \$mux  #( .WIDTH(32) ) _53953_ ( .A(conv2d_16_out_laddr_offset), .B({ _05659_, _05647_, _05648_, _05660_, _05661_, _05662_, _05649_, _05678_, _05663_, _05664_, _05665_, _05679_, _05650_, _05651_, _05666_, _05667_, _05652_, _05668_, _05653_, _05654_, _05669_, _05670_, _05671_, _05655_, _05656_, _05672_, _05673_, _05674_, _05657_, _05675_, _05676_, _05677_ }), .S(_24074_), .Y(_24998_) );
  \$mux  #( .WIDTH(32) ) _53954_ ( .A(conv2d_16_out_page_dma_offset), .B({ _20537_, _20536_, _20534_, _20533_, _20532_, _20531_, _20530_, _20529_, _20528_, _20527_, _20526_, _20525_, _20523_, _20522_, _20521_, _20520_, _20519_, _20518_, _20517_, _20516_, _20515_, _20514_, _20544_, _20543_, _20542_, _20541_, _20540_, _20539_, _20538_, _20535_, _20524_, _20513_ }), .S(_05514_), .Y(_24999_) );
  \$mux  #( .WIDTH(32) ) _53955_ ( .A(conv2d_16_out_page_comp_offset), .B({ _20601_, _20600_, _20598_, _20597_, _20596_, _20595_, _20594_, _20593_, _20592_, _20591_, _20590_, _20589_, _20587_, _20586_, _20585_, _20584_, _20583_, _20582_, _20581_, _20580_, _20579_, _20578_, _20608_, _20607_, _20606_, _20605_, _20604_, _20603_, _20602_, _20599_, _20588_, _20577_ }), .S(_05514_), .Y(_25000_) );
  \$mux  #( .WIDTH(1) ) _53956_ ( .A(conv2d_16_out_page), .B(_20610_), .S(_05514_), .Y(_25001_) );
  \$mux  #( .WIDTH(32) ) _53957_ ( .A(conv2d_16_filter_page_dma_offset), .B({ _20667_, _20666_, _20664_, _20663_, _20662_, _20661_, _20660_, _20659_, _20658_, _20657_, _20656_, _20655_, _20653_, _20652_, _20651_, _20650_, _20649_, _20648_, _20647_, _20646_, _20645_, _20644_, _20674_, _20673_, _20672_, _20671_, _20670_, _20669_, _20668_, _20665_, _20654_, _20643_ }), .S(_05514_), .Y(_25003_) );
  \$mux  #( .WIDTH(32) ) _53958_ ( .A(conv2d_16_filter_page_comp_offset), .B({ _20731_, _20730_, _20728_, _20727_, _20726_, _20725_, _20724_, _20723_, _20722_, _20721_, _20720_, _20719_, _20717_, _20716_, _20715_, _20714_, _20713_, _20712_, _20711_, _20710_, _20709_, _20708_, _20738_, _20737_, _20736_, _20735_, _20734_, _20733_, _20732_, _20729_, _20718_, _20707_ }), .S(_05514_), .Y(_25005_) );
  \$mux  #( .WIDTH(32) ) _53959_ ( .A(conv2d_16_act_page_dma_offset_2), .B({ _20795_, _20794_, _20792_, _20791_, _20790_, _20789_, _20788_, _20787_, _20786_, _20785_, _20784_, _20783_, _20781_, _20780_, _20779_, _20778_, _20777_, _20776_, _20775_, _20774_, _20773_, _20772_, _20802_, _20801_, _20800_, _20799_, _20798_, _20797_, _20796_, _20793_, _20782_, _20771_ }), .S(_05514_), .Y(_25008_) );
  \$mux  #( .WIDTH(32) ) _53960_ ( .A(conv2d_16_act_page_dma_offset_1), .B({ _20859_, _20858_, _20856_, _20855_, _20854_, _20853_, _20852_, _20851_, _20850_, _20849_, _20848_, _20847_, _20845_, _20844_, _20843_, _20842_, _20841_, _20840_, _20839_, _20838_, _20837_, _20836_, _20866_, _20865_, _20864_, _20863_, _20862_, _20861_, _20860_, _20857_, _20846_, _20835_ }), .S(_05514_), .Y(_25011_) );
  \$mux  #( .WIDTH(32) ) _53961_ ( .A(conv2d_16_act_page_dma_offset_0), .B({ _20923_, _20922_, _20920_, _20919_, _20918_, _20917_, _20916_, _20915_, _20914_, _20913_, _20912_, _20911_, _20909_, _20908_, _20907_, _20906_, _20905_, _20904_, _20903_, _20902_, _20901_, _20900_, _20930_, _20929_, _20928_, _20927_, _20926_, _20925_, _20924_, _20921_, _20910_, _20899_ }), .S(_05514_), .Y(_25014_) );
  \$mux  #( .WIDTH(32) ) _53962_ ( .A(conv2d_16_act_page_comp_offset_2), .B({ _20987_, _20986_, _20984_, _20983_, _20982_, _20981_, _20980_, _20979_, _20978_, _20977_, _20976_, _20975_, _20973_, _20972_, _20971_, _20970_, _20969_, _20968_, _20967_, _20966_, _20965_, _20964_, _20994_, _20993_, _20992_, _20991_, _20990_, _20989_, _20988_, _20985_, _20974_, _20963_ }), .S(_05514_), .Y(_25017_) );
  \$mux  #( .WIDTH(32) ) _53963_ ( .A(conv2d_16_act_page_comp_offset_1), .B({ _21051_, _21050_, _21048_, _21047_, _21046_, _21045_, _21044_, _21043_, _21042_, _21041_, _21040_, _21039_, _21037_, _21036_, _21035_, _21034_, _21033_, _21032_, _21031_, _21030_, _21029_, _21028_, _21058_, _21057_, _21056_, _21055_, _21054_, _21053_, _21052_, _21049_, _21038_, _21027_ }), .S(_05514_), .Y(_25020_) );
  \$mux  #( .WIDTH(32) ) _53964_ ( .A(conv2d_16_act_page_comp_offset_0), .B({ _21115_, _21114_, _21112_, _21111_, _21110_, _21109_, _21108_, _21107_, _21106_, _21105_, _21104_, _21103_, _21101_, _21100_, _21099_, _21098_, _21097_, _21096_, _21095_, _21094_, _21093_, _21092_, _21122_, _21121_, _21120_, _21119_, _21118_, _21117_, _21116_, _21113_, _21102_, _21091_ }), .S(_05514_), .Y(_25023_) );
  \$mux  #( .WIDTH(2) ) _53965_ ( .A(conv2d_16_prev_row_select), .B({ _21126_, _21125_ }), .S(_05514_), .Y(_25024_) );
  \$mux  #( .WIDTH(32) ) _53966_ ( .A(conv2d_16_prev_och_count), .B({ _21151_, _21150_, _21148_, _21147_, _21146_, _21145_, _21144_, _21143_, _21142_, _21141_, _21140_, _21139_, _21137_, _21136_, _21135_, _21134_, _21133_, _21132_, _21131_, _21130_, _21129_, _21128_, _21158_, _21157_, _21156_, _21155_, _21154_, _21153_, _21152_, _21149_, _21138_, _21127_ }), .S(_05514_), .Y(_25025_) );
  \$mux  #( .WIDTH(32) ) _53967_ ( .A(conv2d_16_prev_bat_count), .B({ _21183_, _21182_, _21180_, _21179_, _21178_, _21177_, _21176_, _21175_, _21174_, _21173_, _21172_, _21171_, _21169_, _21168_, _21167_, _21166_, _21165_, _21164_, _21163_, _21162_, _21161_, _21160_, _21190_, _21189_, _21188_, _21187_, _21186_, _21185_, _21184_, _21181_, _21170_, _21159_ }), .S(_05514_), .Y(_25026_) );
  \$mux  #( .WIDTH(32) ) _53968_ ( .A(conv2d_16_prev_row_count), .B({ _21215_, _21214_, _21212_, _21211_, _21210_, _21209_, _21208_, _21207_, _21206_, _21205_, _21204_, _21203_, _21201_, _21200_, _21199_, _21198_, _21197_, _21196_, _21195_, _21194_, _21193_, _21192_, _21222_, _21221_, _21220_, _21219_, _21218_, _21217_, _21216_, _21213_, _21202_, _21191_ }), .S(_05514_), .Y(_25027_) );
  \$mux  #( .WIDTH(32) ) _53969_ ( .A(conv2d_16_out_ram_select), .B({ _05517_, _05518_, _05519_, _05520_, _05521_, _05522_, _05523_, _05524_, _05525_, _05526_, _05527_, _05528_, _05529_, _05530_, _05531_, _05532_, _05533_, _05534_, _05535_, _05536_, _05537_, _05538_, _05539_, _05540_, _05541_, _05542_, _05543_, _05544_, _05545_, _05546_, _05547_, _05548_ }), .S(_24074_), .Y(_25028_) );
  \$mux  #( .WIDTH(32) ) _53970_ ( .A(conv2d_16_out_row_count), .B({ _21343_, _21342_, _21340_, _21339_, _21338_, _21337_, _21336_, _21335_, _21334_, _21333_, _21332_, _21331_, _21329_, _21328_, _21327_, _21326_, _21325_, _21324_, _21323_, _21322_, _21321_, _21320_, _21350_, _21349_, _21348_, _21347_, _21346_, _21345_, _21344_, _21341_, _21330_, _21319_ }), .S(_05514_), .Y(_25030_) );
  \$mux  #( .WIDTH(2) ) _53971_ ( .A(conv2d_16_row_select), .B({ _21354_, _21353_ }), .S(_05514_), .Y(_25032_) );
  \$mux  #( .WIDTH(32) ) _53972_ ( .A(conv2d_16_och_count), .B({ _21411_, _21410_, _21408_, _21407_, _21406_, _21405_, _21404_, _21403_, _21402_, _21401_, _21400_, _21399_, _21397_, _21396_, _21395_, _21394_, _21393_, _21392_, _21391_, _21390_, _21389_, _21388_, _21418_, _21417_, _21416_, _21415_, _21414_, _21413_, _21412_, _21409_, _21398_, _21387_ }), .S(_05514_), .Y(_25033_) );
  \$mux  #( .WIDTH(32) ) _53973_ ( .A(conv2d_16_bat_count), .B({ _21475_, _21474_, _21472_, _21471_, _21470_, _21469_, _21468_, _21467_, _21466_, _21465_, _21464_, _21463_, _21461_, _21460_, _21459_, _21458_, _21457_, _21456_, _21455_, _21454_, _21453_, _21452_, _21482_, _21481_, _21480_, _21479_, _21478_, _21477_, _21476_, _21473_, _21462_, _21451_ }), .S(_05514_), .Y(_25034_) );
  \$mux  #( .WIDTH(32) ) _53974_ ( .A(conv2d_16_row_count), .B({ _21539_, _21538_, _21536_, _21535_, _21534_, _21533_, _21532_, _21531_, _21530_, _21529_, _21528_, _21527_, _21525_, _21524_, _21523_, _21522_, _21521_, _21520_, _21519_, _21518_, _21517_, _21516_, _21546_, _21545_, _21544_, _21543_, _21542_, _21541_, _21540_, _21537_, _21526_, _21515_ }), .S(_05514_), .Y(_25035_) );
  \$mux  #( .WIDTH(32) ) _53975_ ( .A(conv2d_16_sync_out_count), .B({ _21571_, _21570_, _21568_, _21567_, _21566_, _21565_, _21564_, _21563_, _21562_, _21561_, _21560_, _21559_, _21557_, _21556_, _21555_, _21554_, _21553_, _21552_, _21551_, _21550_, _21549_, _21548_, _21578_, _21577_, _21576_, _21575_, _21574_, _21573_, _21572_, _21569_, _21558_, _21547_ }), .S(_24075_), .Y(_25037_) );
  \$mux  #( .WIDTH(1) ) _53976_ ( .A(conv2d_16_dma_flag_2), .B(_21580_), .S(_05514_), .Y(_25038_) );
  \$mux  #( .WIDTH(1) ) _53977_ ( .A(conv2d_16_dma_flag_1), .B(_21580_), .S(_05514_), .Y(_25039_) );
  \$mux  #( .WIDTH(32) ) _53978_ ( .A(conv2d_16_out_base_offset_och), .B({ _21637_, _21636_, _21634_, _21633_, _21632_, _21631_, _21630_, _21629_, _21628_, _21627_, _21626_, _21625_, _21623_, _21622_, _21621_, _21620_, _21619_, _21618_, _21617_, _21616_, _21615_, _21614_, _21644_, _21643_, _21642_, _21641_, _21640_, _21639_, _21638_, _21635_, _21624_, _21613_ }), .S(_05514_), .Y(_25041_) );
  \$mux  #( .WIDTH(32) ) _53979_ ( .A(conv2d_16_out_base_offset_bat), .B({ _21701_, _21700_, _21698_, _21697_, _21696_, _21695_, _21694_, _21693_, _21692_, _21691_, _21690_, _21689_, _21687_, _21686_, _21685_, _21684_, _21683_, _21682_, _21681_, _21680_, _21679_, _21678_, _21708_, _21707_, _21706_, _21705_, _21704_, _21703_, _21702_, _21699_, _21688_, _21677_ }), .S(_05514_), .Y(_25042_) );
  \$mux  #( .WIDTH(32) ) _53980_ ( .A(conv2d_16_out_base_offset_row), .B({ _21765_, _21764_, _21762_, _21761_, _21760_, _21759_, _21758_, _21757_, _21756_, _21755_, _21754_, _21753_, _21751_, _21750_, _21749_, _21748_, _21747_, _21746_, _21745_, _21744_, _21743_, _21742_, _21772_, _21771_, _21770_, _21769_, _21768_, _21767_, _21766_, _21763_, _21752_, _21741_ }), .S(_05514_), .Y(_25044_) );
  \$mux  #( .WIDTH(32) ) _53981_ ( .A(conv2d_16_out_base_offset_col), .B({ _21829_, _21828_, _21826_, _21825_, _21824_, _21823_, _21822_, _21821_, _21820_, _21819_, _21818_, _21817_, _21815_, _21814_, _21813_, _21812_, _21811_, _21810_, _21809_, _21808_, _21807_, _21806_, _21836_, _21835_, _21834_, _21833_, _21832_, _21831_, _21830_, _21827_, _21816_, _21805_ }), .S(_05514_), .Y(_25045_) );
  \$mux  #( .WIDTH(32) ) _53982_ ( .A(conv2d_16_filter_base_offset), .B({ _21893_, _21892_, _21890_, _21889_, _21888_, _21887_, _21886_, _21885_, _21884_, _21883_, _21882_, _21881_, _21879_, _21878_, _21877_, _21876_, _21875_, _21874_, _21873_, _21872_, _21871_, _21870_, _21900_, _21899_, _21898_, _21897_, _21896_, _21895_, _21894_, _21891_, _21880_, _21869_ }), .S(_05514_), .Y(_25047_) );
  \$mux  #( .WIDTH(32) ) _53983_ ( .A(conv2d_16_act_base_offset_bat), .B({ _21957_, _21956_, _21954_, _21953_, _21952_, _21951_, _21950_, _21949_, _21948_, _21947_, _21946_, _21945_, _21943_, _21942_, _21941_, _21940_, _21939_, _21938_, _21937_, _21936_, _21935_, _21934_, _21964_, _21963_, _21962_, _21961_, _21960_, _21959_, _21958_, _21955_, _21944_, _21933_ }), .S(_05514_), .Y(_25048_) );
  \$mux  #( .WIDTH(32) ) _53984_ ( .A(conv2d_16_act_base_offset_row), .B({ _22021_, _22020_, _22018_, _22017_, _22016_, _22015_, _22014_, _22013_, _22012_, _22011_, _22010_, _22009_, _22007_, _22006_, _22005_, _22004_, _22003_, _22002_, _22001_, _22000_, _21999_, _21998_, _22028_, _22027_, _22026_, _22025_, _22024_, _22023_, _22022_, _22019_, _22008_, _21997_ }), .S(_05514_), .Y(_25049_) );
  \$mux  #( .WIDTH(32) ) _53985_ ( .A(control_conv2d_16), .B({ _22085_, _22084_, _22082_, _22081_, _22080_, _22079_, _22078_, _22077_, _22076_, _22075_, _22074_, _22073_, _22071_, _22070_, _22069_, _22068_, _22067_, _22066_, _22065_, _22064_, _22063_, _22062_, _22092_, _22091_, _22090_, _22089_, _22088_, _22087_, _22086_, _22083_, _22072_, _22061_ }), .S(_24076_), .Y(_25052_) );
  \$mux  #( .WIDTH(32) ) _53986_ ( .A(matmul_29_arg_objaddr_3), .B({ _22821_, _22820_, _22818_, _22817_, _22816_, _22815_, _22814_, _22813_, _22812_, _22811_, _22810_, _22809_, _22807_, _22806_, _22805_, _22804_, _22803_, _22802_, _22801_, _22800_, _22799_, _22798_, _22828_, _22827_, _22826_, _22825_, _22824_, _22823_, _22822_, _22819_, _22808_, _22797_ }), .S(_24077_), .Y(_25059_) );
  \$mux  #( .WIDTH(32) ) _53987_ ( .A(matmul_29_arg_objaddr_2), .B({ _22853_, _22852_, _22850_, _22849_, _22848_, _22847_, _22846_, _22845_, _22844_, _22843_, _22842_, _22841_, _22839_, _22838_, _22837_, _22836_, _22835_, _22834_, _22833_, _22832_, _22831_, _22830_, _22860_, _22859_, _22858_, _22857_, _22856_, _22855_, _22854_, _22851_, _22840_, _22829_ }), .S(_24078_), .Y(_25060_) );
  \$mux  #( .WIDTH(32) ) _53988_ ( .A(matmul_29_arg_objaddr_1), .B({ _22885_, _22884_, _22882_, _22881_, _22880_, _22879_, _22878_, _22877_, _22876_, _22875_, _22874_, _22873_, _22871_, _22870_, _22869_, _22868_, _22867_, _22866_, _22865_, _22864_, _22863_, _22862_, _22892_, _22891_, _22890_, _22889_, _22888_, _22887_, _22886_, _22883_, _22872_, _22861_ }), .S(_24079_), .Y(_25061_) );
  \$mux  #( .WIDTH(32) ) _53989_ ( .A(matmul_29_arg_objaddr_0), .B({ _22917_, _22916_, _22914_, _22913_, _22912_, _22911_, _22910_, _22909_, _22908_, _22907_, _22906_, _22905_, _22903_, _22902_, _22901_, _22900_, _22899_, _22898_, _22897_, _22896_, _22895_, _22894_, _22924_, _22923_, _22922_, _22921_, _22920_, _22919_, _22918_, _22915_, _22904_, _22893_ }), .S(_24080_), .Y(_25062_) );
  \$mux  #( .WIDTH(32) ) _53990_ ( .A(matmul_29_objaddr), .B({ _22949_, _22948_, _22946_, _22945_, _22944_, _22943_, _22942_, _22941_, _22940_, _22939_, _22938_, _22937_, _22935_, _22934_, _22933_, _22932_, _22931_, _22930_, _22929_, _22928_, _22927_, _22926_, _22956_, _22955_, _22954_, _22953_, _22952_, _22951_, _22950_, _22947_, _22936_, _22925_ }), .S(_24081_), .Y(_25063_) );
  \$mux  #( .WIDTH(32) ) _53991_ ( .A(max_pool_serial_18_arg_objaddr_0), .B({ _22981_, _22980_, _22978_, _22977_, _22976_, _22975_, _22974_, _22973_, _22972_, _22971_, _22970_, _22969_, _22967_, _22966_, _22965_, _22964_, _22963_, _22962_, _22961_, _22960_, _22959_, _22958_, _22988_, _22987_, _22986_, _22985_, _22984_, _22983_, _22982_, _22979_, _22968_, _22957_ }), .S(_24082_), .Y(_25064_) );
  \$mux  #( .WIDTH(32) ) _53992_ ( .A(max_pool_serial_18_objaddr), .B({ _23013_, _23012_, _23010_, _23009_, _23008_, _23007_, _23006_, _23005_, _23004_, _23003_, _23002_, _23001_, _22999_, _22998_, _22997_, _22996_, _22995_, _22994_, _22993_, _22992_, _22991_, _22990_, _23020_, _23019_, _23018_, _23017_, _23016_, _23015_, _23014_, _23011_, _23000_, _22989_ }), .S(_24083_), .Y(_25065_) );
  \$mux  #( .WIDTH(32) ) _53993_ ( .A(conv2d_16_arg_objaddr_3), .B({ _23045_, _23044_, _23042_, _23041_, _23040_, _23039_, _23038_, _23037_, _23036_, _23035_, _23034_, _23033_, _23031_, _23030_, _23029_, _23028_, _23027_, _23026_, _23025_, _23024_, _23023_, _23022_, _23052_, _23051_, _23050_, _23049_, _23048_, _23047_, _23046_, _23043_, _23032_, _23021_ }), .S(_24084_), .Y(_25066_) );
  \$mux  #( .WIDTH(32) ) _53994_ ( .A(conv2d_16_arg_objaddr_2), .B({ _23077_, _23076_, _23074_, _23073_, _23072_, _23071_, _23070_, _23069_, _23068_, _23067_, _23066_, _23065_, _23063_, _23062_, _23061_, _23060_, _23059_, _23058_, _23057_, _23056_, _23055_, _23054_, _23084_, _23083_, _23082_, _23081_, _23080_, _23079_, _23078_, _23075_, _23064_, _23053_ }), .S(_24085_), .Y(_25067_) );
  \$mux  #( .WIDTH(32) ) _53995_ ( .A(conv2d_16_arg_objaddr_1), .B({ _23109_, _23108_, _23106_, _23105_, _23104_, _23103_, _23102_, _23101_, _23100_, _23099_, _23098_, _23097_, _23095_, _23094_, _23093_, _23092_, _23091_, _23090_, _23089_, _23088_, _23087_, _23086_, _23116_, _23115_, _23114_, _23113_, _23112_, _23111_, _23110_, _23107_, _23096_, _23085_ }), .S(_24086_), .Y(_25068_) );
  \$mux  #( .WIDTH(32) ) _53996_ ( .A(conv2d_16_arg_objaddr_0), .B({ _23141_, _23140_, _23138_, _23137_, _23136_, _23135_, _23134_, _23133_, _23132_, _23131_, _23130_, _23129_, _23127_, _23126_, _23125_, _23124_, _23123_, _23122_, _23121_, _23120_, _23119_, _23118_, _23148_, _23147_, _23146_, _23145_, _23144_, _23143_, _23142_, _23139_, _23128_, _23117_ }), .S(_24087_), .Y(_25069_) );
  \$mux  #( .WIDTH(32) ) _53997_ ( .A(conv2d_16_objaddr), .B({ _23173_, _23172_, _23170_, _23169_, _23168_, _23167_, _23166_, _23165_, _23164_, _23163_, _23162_, _23161_, _23159_, _23158_, _23157_, _23156_, _23155_, _23154_, _23153_, _23152_, _23151_, _23150_, _23180_, _23179_, _23178_, _23177_, _23176_, _23175_, _23174_, _23171_, _23160_, _23149_ }), .S(_24088_), .Y(_25070_) );
  \$mux  #( .WIDTH(32) ) _53998_ ( .A(main_fsm), .B({ _23205_, _23204_, _23202_, _23201_, _23200_, _23199_, _23198_, _23197_, _23196_, _23195_, _23194_, _23193_, _23191_, _23190_, _23189_, _23188_, _23187_, _23186_, _23185_, _23184_, _23183_, _23182_, _23212_, _23211_, _23210_, _23209_, _23208_, _23207_, _23206_, _23203_, _23192_, _23181_ }), .S(_24089_), .Y(_25071_) );
  \$mux  #( .WIDTH(2) ) _53999_ ( .A(matmul_29_control_param_index), .B({ _05680_, _05681_ }), .S(_24090_), .Y(_25072_) );
  \$mux  #( .WIDTH(2) ) _54000_ ( .A(max_pool_serial_18_control_param_index), .B({ _05682_, _05646_ }), .S(_24091_), .Y(_25073_) );
  \$mux  #( .WIDTH(2) ) _54001_ ( .A(conv2d_16_control_param_index), .B({ _05645_, _05683_ }), .S(_24092_), .Y(_25074_) );
  \$mux  #( .WIDTH(1) ) _54002_ ( .A(_stream_matmul_29_source_busy), .B(_23533_), .S(_24093_), .Y(_25075_) );
  \$mux  #( .WIDTH(32) ) _54003_ ( .A(_stream_matmul_29_fsm), .B({ _23559_, _23558_, _23556_, _23555_, _23554_, _23553_, _23552_, _23551_, _23550_, _23549_, _23548_, _23547_, _23545_, _23544_, _23543_, _23542_, _23541_, _23540_, _23539_, _23538_, _23537_, _23536_, _23566_, _23565_, _23564_, _23563_, _23562_, _23561_, _23560_, _23557_, _23546_, _23535_ }), .S(_24094_), .Y(_25080_) );
  \$mux  #( .WIDTH(1) ) _54004_ ( .A(_stream_max_pool_serial_18_source_busy), .B(_23631_), .S(_24095_), .Y(_25325_) );
  \$mux  #( .WIDTH(32) ) _54005_ ( .A(_stream_max_pool_serial_18_fsm), .B({ _23657_, _23656_, _23654_, _23653_, _23652_, _23651_, _23650_, _23649_, _23648_, _23647_, _23646_, _23645_, _23643_, _23642_, _23641_, _23640_, _23639_, _23638_, _23637_, _23636_, _23635_, _23634_, _23664_, _23663_, _23662_, _23661_, _23660_, _23659_, _23658_, _23655_, _23644_, _23633_ }), .S(_24096_), .Y(_25330_) );
  \$mux  #( .WIDTH(1) ) _54006_ ( .A(_stream_conv2d_16_source_busy), .B(_23729_), .S(_24097_), .Y(_25402_) );
  \$mux  #( .WIDTH(32) ) _54007_ ( .A(_stream_conv2d_16_fsm), .B({ _23755_, _23754_, _23752_, _23751_, _23750_, _23749_, _23748_, _23747_, _23746_, _23745_, _23744_, _23743_, _23741_, _23740_, _23739_, _23738_, _23737_, _23736_, _23735_, _23734_, _23733_, _23732_, _23762_, _23761_, _23760_, _23759_, _23758_, _23757_, _23756_, _23753_, _23742_, _23731_ }), .S(_24098_), .Y(_25407_) );
  \$mux  #( .WIDTH(32) ) _54008_ ( .A(_saxi_register_fsm), .B({ _23851_, _23850_, _23848_, _23847_, _23846_, _23845_, _23844_, _23843_, _23842_, _23841_, _23840_, _23839_, _23837_, _23836_, _23835_, _23834_, _23833_, _23832_, _23831_, _23830_, _23829_, _23828_, _23858_, _23857_, _23856_, _23855_, _23854_, _23853_, _23852_, _23849_, _23838_, _23827_ }), .S(_24099_), .Y(_28091_) );
  \$mux  #( .WIDTH(2) ) _54009_ ( .A({ 1'hx, _29054_ }), .B({ _29054_, 1'hx }), .S(_counter_data_782[31]), .Y(_28508_) );
  \$mux  #( .WIDTH(66) ) _54010_ ( .A({ _28949_[65:34], _28944_[65:32] }), .B({ _28944_[65:32], 32'h00000000 }), .S(_minus_data_5[5]), .Y(_28509_) );
  \$mux  #( .WIDTH(66) ) _54011_ ( .A({ _28948_[65:50], _28943_[65:16] }), .B({ _28943_[65:16], 16'h0000 }), .S(_minus_data_5[4]), .Y({ _28949_[65:34], _28944_[65:32] }) );
  \$mux  #( .WIDTH(66) ) _54012_ ( .A(_28947_), .B({ _28947_[57:0], 8'h00 }), .S(_minus_data_5[3]), .Y({ _28948_[65:50], _28943_[65:16] }) );
  \$mux  #( .WIDTH(66) ) _54013_ ( .A(_28946_), .B({ _28946_[61:0], 4'h0 }), .S(_minus_data_5[2]), .Y(_28947_) );
  \$mux  #( .WIDTH(66) ) _54014_ ( .A(_28945_), .B({ _28945_[63:0], 2'h0 }), .S(_minus_data_5[1]), .Y(_28946_) );
  \$mux  #( .WIDTH(66) ) _54015_ ( .A(66'h00000000000000001), .B(66'h00000000000000002), .S(_minus_data_5[0]), .Y(_28945_) );
  \$mux  #( .WIDTH(18) ) _54016_ ( .A(_28952_), .B({ _28952_[9:0], 8'h00 }), .S(_minus_data_59[3]), .Y(_28510_) );
  \$mux  #( .WIDTH(18) ) _54017_ ( .A(_28951_), .B({ _28951_[13:0], 4'h0 }), .S(_minus_data_59[2]), .Y(_28952_) );
  \$mux  #( .WIDTH(18) ) _54018_ ( .A(_28950_), .B({ _28950_[15:0], 2'h0 }), .S(_minus_data_59[1]), .Y(_28951_) );
  \$mux  #( .WIDTH(18) ) _54019_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_59[0]), .Y(_28950_) );
  \$mux  #( .WIDTH(18) ) _54020_ ( .A(_28955_), .B({ _28955_[9:0], 8'h00 }), .S(_minus_data_76[3]), .Y(_28511_) );
  \$mux  #( .WIDTH(18) ) _54021_ ( .A(_28954_), .B({ _28954_[13:0], 4'h0 }), .S(_minus_data_76[2]), .Y(_28955_) );
  \$mux  #( .WIDTH(18) ) _54022_ ( .A(_28953_), .B({ _28953_[15:0], 2'h0 }), .S(_minus_data_76[1]), .Y(_28954_) );
  \$mux  #( .WIDTH(18) ) _54023_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_76[0]), .Y(_28953_) );
  \$mux  #( .WIDTH(18) ) _54024_ ( .A(_28958_), .B({ _28958_[9:0], 8'h00 }), .S(_minus_data_93[3]), .Y(_28512_) );
  \$mux  #( .WIDTH(18) ) _54025_ ( .A(_28957_), .B({ _28957_[13:0], 4'h0 }), .S(_minus_data_93[2]), .Y(_28958_) );
  \$mux  #( .WIDTH(18) ) _54026_ ( .A(_28956_), .B({ _28956_[15:0], 2'h0 }), .S(_minus_data_93[1]), .Y(_28957_) );
  \$mux  #( .WIDTH(18) ) _54027_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_93[0]), .Y(_28956_) );
  \$mux  #( .WIDTH(18) ) _54028_ ( .A(_28961_), .B({ _28961_[9:0], 8'h00 }), .S(_minus_data_110[3]), .Y(_28513_) );
  \$mux  #( .WIDTH(18) ) _54029_ ( .A(_28960_), .B({ _28960_[13:0], 4'h0 }), .S(_minus_data_110[2]), .Y(_28961_) );
  \$mux  #( .WIDTH(18) ) _54030_ ( .A(_28959_), .B({ _28959_[15:0], 2'h0 }), .S(_minus_data_110[1]), .Y(_28960_) );
  \$mux  #( .WIDTH(18) ) _54031_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_110[0]), .Y(_28959_) );
  \$mux  #( .WIDTH(18) ) _54032_ ( .A(_28964_), .B({ _28964_[9:0], 8'h00 }), .S(_minus_data_127[3]), .Y(_28514_) );
  \$mux  #( .WIDTH(18) ) _54033_ ( .A(_28963_), .B({ _28963_[13:0], 4'h0 }), .S(_minus_data_127[2]), .Y(_28964_) );
  \$mux  #( .WIDTH(18) ) _54034_ ( .A(_28962_), .B({ _28962_[15:0], 2'h0 }), .S(_minus_data_127[1]), .Y(_28963_) );
  \$mux  #( .WIDTH(18) ) _54035_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_127[0]), .Y(_28962_) );
  \$mux  #( .WIDTH(18) ) _54036_ ( .A(_28967_), .B({ _28967_[9:0], 8'h00 }), .S(_minus_data_144[3]), .Y(_28515_) );
  \$mux  #( .WIDTH(18) ) _54037_ ( .A(_28966_), .B({ _28966_[13:0], 4'h0 }), .S(_minus_data_144[2]), .Y(_28967_) );
  \$mux  #( .WIDTH(18) ) _54038_ ( .A(_28965_), .B({ _28965_[15:0], 2'h0 }), .S(_minus_data_144[1]), .Y(_28966_) );
  \$mux  #( .WIDTH(18) ) _54039_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_144[0]), .Y(_28965_) );
  \$mux  #( .WIDTH(18) ) _54040_ ( .A(_28970_), .B({ _28970_[9:0], 8'h00 }), .S(_minus_data_161[3]), .Y(_28516_) );
  \$mux  #( .WIDTH(18) ) _54041_ ( .A(_28969_), .B({ _28969_[13:0], 4'h0 }), .S(_minus_data_161[2]), .Y(_28970_) );
  \$mux  #( .WIDTH(18) ) _54042_ ( .A(_28968_), .B({ _28968_[15:0], 2'h0 }), .S(_minus_data_161[1]), .Y(_28969_) );
  \$mux  #( .WIDTH(18) ) _54043_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_161[0]), .Y(_28968_) );
  \$mux  #( .WIDTH(18) ) _54044_ ( .A(_28973_), .B({ _28973_[9:0], 8'h00 }), .S(_minus_data_178[3]), .Y(_28517_) );
  \$mux  #( .WIDTH(18) ) _54045_ ( .A(_28972_), .B({ _28972_[13:0], 4'h0 }), .S(_minus_data_178[2]), .Y(_28973_) );
  \$mux  #( .WIDTH(18) ) _54046_ ( .A(_28971_), .B({ _28971_[15:0], 2'h0 }), .S(_minus_data_178[1]), .Y(_28972_) );
  \$mux  #( .WIDTH(18) ) _54047_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_178[0]), .Y(_28971_) );
  \$mux  #( .WIDTH(18) ) _54048_ ( .A(_28976_), .B({ _28976_[9:0], 8'h00 }), .S(_minus_data_195[3]), .Y(_28518_) );
  \$mux  #( .WIDTH(18) ) _54049_ ( .A(_28975_), .B({ _28975_[13:0], 4'h0 }), .S(_minus_data_195[2]), .Y(_28976_) );
  \$mux  #( .WIDTH(18) ) _54050_ ( .A(_28974_), .B({ _28974_[15:0], 2'h0 }), .S(_minus_data_195[1]), .Y(_28975_) );
  \$mux  #( .WIDTH(18) ) _54051_ ( .A(18'h00001), .B(18'h00002), .S(_minus_data_195[0]), .Y(_28974_) );
  \$mux  #( .WIDTH(32) ) _54052_ ( .A(_28979_), .B({ _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31], _28979_[31] }), .S(__delay_data_754[5]), .Y(_28521_) );
  \$mux  #( .WIDTH(32) ) _54053_ ( .A(_28977_), .B({ _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31], _28977_[31:16] }), .S(__delay_data_754[4]), .Y(_28979_) );
  \$mux  #( .WIDTH(32) ) _54054_ ( .A({ _28978_[31], _28978_[22:0], _28982_[7:0] }), .B({ _28978_[31], _28978_[31], _28978_[31], _28978_[31], _28978_[31], _28978_[31], _28978_[31], _28978_[31], _28978_[31], _28978_[22:0] }), .S(__delay_data_754[3]), .Y(_28977_) );
  \$mux  #( .WIDTH(32) ) _54055_ ( .A(_28981_), .B({ _28981_[31], _28981_[31], _28981_[31], _28981_[31], _28981_[31:4] }), .S(__delay_data_754[2]), .Y({ _28978_[31], _28978_[22:0], _28982_[7:0] }) );
  \$mux  #( .WIDTH(32) ) _54056_ ( .A(_28980_), .B({ _28980_[31], _28980_[31], _28980_[31:2] }), .S(__delay_data_754[1]), .Y(_28981_) );
  \$mux  #( .WIDTH(32) ) _54057_ ( .A(_plus_data_20), .B({ _plus_data_20[31], _plus_data_20[31:1] }), .S(__delay_data_754[0]), .Y(_28980_) );
  \$mux  #( .WIDTH(40) ) _54058_ ( .A(_28985_), .B({ _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39], _28985_[39:32] }), .S(__delay_data_767[5]), .Y(_28522_) );
  \$mux  #( .WIDTH(40) ) _54059_ ( .A(_28983_), .B({ _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39], _28983_[39:16] }), .S(__delay_data_767[4]), .Y(_28985_) );
  \$mux  #( .WIDTH(40) ) _54060_ ( .A({ _28984_[39], _28984_[30:0], _28988_[7:0] }), .B({ _28984_[39], _28984_[39], _28984_[39], _28984_[39], _28984_[39], _28984_[39], _28984_[39], _28984_[39], _28984_[39], _28984_[30:0] }), .S(__delay_data_767[3]), .Y(_28983_) );
  \$mux  #( .WIDTH(40) ) _54061_ ( .A(_28987_), .B({ _28987_[39], _28987_[39], _28987_[39], _28987_[39], _28987_[39:4] }), .S(__delay_data_767[2]), .Y({ _28984_[39], _28984_[30:0], _28988_[7:0] }) );
  \$mux  #( .WIDTH(40) ) _54062_ ( .A(_28986_), .B({ _28986_[39], _28986_[39], _28986_[39:2] }), .S(__delay_data_767[1]), .Y(_28987_) );
  \$mux  #( .WIDTH(40) ) _54063_ ( .A(_times_mul_odata_reg_41), .B({ _times_mul_odata_reg_41[39], _times_mul_odata_reg_41[39:1] }), .S(__delay_data_767[0]), .Y(_28986_) );
  \$mux  #( .WIDTH(12) ) _54064_ ( .A({ _28989_[11], _28989_[2:0], _28992_[7:0] }), .B({ _28989_[11], _28989_[11], _28989_[11], _28989_[11], _28989_[11], _28989_[11], _28989_[11], _28989_[11], _28989_[11], _28989_[2:0] }), .S(__delay_data_606[3]), .Y(_28523_) );
  \$mux  #( .WIDTH(12) ) _54065_ ( .A(_28991_), .B({ _28991_[11], _28991_[11], _28991_[11], _28991_[11], _28991_[11:4] }), .S(__delay_data_606[2]), .Y({ _28989_[11], _28989_[2:0], _28992_[7:0] }) );
  \$mux  #( .WIDTH(12) ) _54066_ ( .A(_28990_), .B({ _28990_[11], _28990_[11], _28990_[11:2] }), .S(__delay_data_606[1]), .Y(_28991_) );
  \$mux  #( .WIDTH(12) ) _54067_ ( .A(__muladd_madd_odata_reg_69), .B({ __muladd_madd_odata_reg_69[11], __muladd_madd_odata_reg_69[11:1] }), .S(__delay_data_606[0]), .Y(_28990_) );
  \$mux  #( .WIDTH(12) ) _54068_ ( .A({ _28993_[11], _28993_[2:0], _28996_[7:0] }), .B({ _28993_[11], _28993_[11], _28993_[11], _28993_[11], _28993_[11], _28993_[11], _28993_[11], _28993_[11], _28993_[11], _28993_[2:0] }), .S(__delay_data_623[3]), .Y(_28524_) );
  \$mux  #( .WIDTH(12) ) _54069_ ( .A(_28995_), .B({ _28995_[11], _28995_[11], _28995_[11], _28995_[11], _28995_[11:4] }), .S(__delay_data_623[2]), .Y({ _28993_[11], _28993_[2:0], _28996_[7:0] }) );
  \$mux  #( .WIDTH(12) ) _54070_ ( .A(_28994_), .B({ _28994_[11], _28994_[11], _28994_[11:2] }), .S(__delay_data_623[1]), .Y(_28995_) );
  \$mux  #( .WIDTH(12) ) _54071_ ( .A(__muladd_madd_odata_reg_86), .B({ __muladd_madd_odata_reg_86[11], __muladd_madd_odata_reg_86[11:1] }), .S(__delay_data_623[0]), .Y(_28994_) );
  \$mux  #( .WIDTH(12) ) _54072_ ( .A({ _28997_[11], _28997_[2:0], _29000_[7:0] }), .B({ _28997_[11], _28997_[11], _28997_[11], _28997_[11], _28997_[11], _28997_[11], _28997_[11], _28997_[11], _28997_[11], _28997_[2:0] }), .S(__delay_data_640[3]), .Y(_28525_) );
  \$mux  #( .WIDTH(12) ) _54073_ ( .A(_28999_), .B({ _28999_[11], _28999_[11], _28999_[11], _28999_[11], _28999_[11:4] }), .S(__delay_data_640[2]), .Y({ _28997_[11], _28997_[2:0], _29000_[7:0] }) );
  \$mux  #( .WIDTH(12) ) _54074_ ( .A(_28998_), .B({ _28998_[11], _28998_[11], _28998_[11:2] }), .S(__delay_data_640[1]), .Y(_28999_) );
  \$mux  #( .WIDTH(12) ) _54075_ ( .A(__muladd_madd_odata_reg_103), .B({ __muladd_madd_odata_reg_103[11], __muladd_madd_odata_reg_103[11:1] }), .S(__delay_data_640[0]), .Y(_28998_) );
  \$mux  #( .WIDTH(12) ) _54076_ ( .A({ _29001_[11], _29001_[2:0], _29004_[7:0] }), .B({ _29001_[11], _29001_[11], _29001_[11], _29001_[11], _29001_[11], _29001_[11], _29001_[11], _29001_[11], _29001_[11], _29001_[2:0] }), .S(__delay_data_657[3]), .Y(_28526_) );
  \$mux  #( .WIDTH(12) ) _54077_ ( .A(_29003_), .B({ _29003_[11], _29003_[11], _29003_[11], _29003_[11], _29003_[11:4] }), .S(__delay_data_657[2]), .Y({ _29001_[11], _29001_[2:0], _29004_[7:0] }) );
  \$mux  #( .WIDTH(12) ) _54078_ ( .A(_29002_), .B({ _29002_[11], _29002_[11], _29002_[11:2] }), .S(__delay_data_657[1]), .Y(_29003_) );
  \$mux  #( .WIDTH(12) ) _54079_ ( .A(__muladd_madd_odata_reg_120), .B({ __muladd_madd_odata_reg_120[11], __muladd_madd_odata_reg_120[11:1] }), .S(__delay_data_657[0]), .Y(_29002_) );
  \$mux  #( .WIDTH(12) ) _54080_ ( .A({ _29005_[11], _29005_[2:0], _29008_[7:0] }), .B({ _29005_[11], _29005_[11], _29005_[11], _29005_[11], _29005_[11], _29005_[11], _29005_[11], _29005_[11], _29005_[11], _29005_[2:0] }), .S(__delay_data_674[3]), .Y(_28527_) );
  \$mux  #( .WIDTH(12) ) _54081_ ( .A(_29007_), .B({ _29007_[11], _29007_[11], _29007_[11], _29007_[11], _29007_[11:4] }), .S(__delay_data_674[2]), .Y({ _29005_[11], _29005_[2:0], _29008_[7:0] }) );
  \$mux  #( .WIDTH(12) ) _54082_ ( .A(_29006_), .B({ _29006_[11], _29006_[11], _29006_[11:2] }), .S(__delay_data_674[1]), .Y(_29007_) );
  \$mux  #( .WIDTH(12) ) _54083_ ( .A(__muladd_madd_odata_reg_137), .B({ __muladd_madd_odata_reg_137[11], __muladd_madd_odata_reg_137[11:1] }), .S(__delay_data_674[0]), .Y(_29006_) );
  \$mux  #( .WIDTH(12) ) _54084_ ( .A({ _29009_[11], _29009_[2:0], _29012_[7:0] }), .B({ _29009_[11], _29009_[11], _29009_[11], _29009_[11], _29009_[11], _29009_[11], _29009_[11], _29009_[11], _29009_[11], _29009_[2:0] }), .S(__delay_data_691[3]), .Y(_28528_) );
  \$mux  #( .WIDTH(12) ) _54085_ ( .A(_29011_), .B({ _29011_[11], _29011_[11], _29011_[11], _29011_[11], _29011_[11:4] }), .S(__delay_data_691[2]), .Y({ _29009_[11], _29009_[2:0], _29012_[7:0] }) );
  \$mux  #( .WIDTH(12) ) _54086_ ( .A(_29010_), .B({ _29010_[11], _29010_[11], _29010_[11:2] }), .S(__delay_data_691[1]), .Y(_29011_) );
  \$mux  #( .WIDTH(12) ) _54087_ ( .A(__muladd_madd_odata_reg_154), .B({ __muladd_madd_odata_reg_154[11], __muladd_madd_odata_reg_154[11:1] }), .S(__delay_data_691[0]), .Y(_29010_) );
  \$mux  #( .WIDTH(12) ) _54088_ ( .A({ _29013_[11], _29013_[2:0], _29016_[7:0] }), .B({ _29013_[11], _29013_[11], _29013_[11], _29013_[11], _29013_[11], _29013_[11], _29013_[11], _29013_[11], _29013_[11], _29013_[2:0] }), .S(__delay_data_708[3]), .Y(_28529_) );
  \$mux  #( .WIDTH(12) ) _54089_ ( .A(_29015_), .B({ _29015_[11], _29015_[11], _29015_[11], _29015_[11], _29015_[11:4] }), .S(__delay_data_708[2]), .Y({ _29013_[11], _29013_[2:0], _29016_[7:0] }) );
  \$mux  #( .WIDTH(12) ) _54090_ ( .A(_29014_), .B({ _29014_[11], _29014_[11], _29014_[11:2] }), .S(__delay_data_708[1]), .Y(_29015_) );
  \$mux  #( .WIDTH(12) ) _54091_ ( .A(__muladd_madd_odata_reg_171), .B({ __muladd_madd_odata_reg_171[11], __muladd_madd_odata_reg_171[11:1] }), .S(__delay_data_708[0]), .Y(_29014_) );
  \$mux  #( .WIDTH(12) ) _54092_ ( .A({ _29017_[11], _29017_[2:0], _29020_[7:0] }), .B({ _29017_[11], _29017_[11], _29017_[11], _29017_[11], _29017_[11], _29017_[11], _29017_[11], _29017_[11], _29017_[11], _29017_[2:0] }), .S(__delay_data_725[3]), .Y(_28530_) );
  \$mux  #( .WIDTH(12) ) _54093_ ( .A(_29019_), .B({ _29019_[11], _29019_[11], _29019_[11], _29019_[11], _29019_[11:4] }), .S(__delay_data_725[2]), .Y({ _29017_[11], _29017_[2:0], _29020_[7:0] }) );
  \$mux  #( .WIDTH(12) ) _54094_ ( .A(_29018_), .B({ _29018_[11], _29018_[11], _29018_[11:2] }), .S(__delay_data_725[1]), .Y(_29019_) );
  \$mux  #( .WIDTH(12) ) _54095_ ( .A(__muladd_madd_odata_reg_188), .B({ __muladd_madd_odata_reg_188[11], __muladd_madd_odata_reg_188[11:1] }), .S(__delay_data_725[0]), .Y(_29018_) );
  \$mux  #( .WIDTH(12) ) _54096_ ( .A({ _29021_[11], _29021_[2:0], _29024_[7:0] }), .B({ _29021_[11], _29021_[11], _29021_[11], _29021_[11], _29021_[11], _29021_[11], _29021_[11], _29021_[11], _29021_[11], _29021_[2:0] }), .S(__delay_data_742[3]), .Y(_28531_) );
  \$mux  #( .WIDTH(12) ) _54097_ ( .A(_29023_), .B({ _29023_[11], _29023_[11], _29023_[11], _29023_[11], _29023_[11:4] }), .S(__delay_data_742[2]), .Y({ _29021_[11], _29021_[2:0], _29024_[7:0] }) );
  \$mux  #( .WIDTH(12) ) _54098_ ( .A(_29022_), .B({ _29022_[11], _29022_[11], _29022_[11:2] }), .S(__delay_data_742[1]), .Y(_29023_) );
  \$mux  #( .WIDTH(12) ) _54099_ ( .A(__muladd_madd_odata_reg_205), .B({ __muladd_madd_odata_reg_205[11], __muladd_madd_odata_reg_205[11:1] }), .S(__delay_data_742[0]), .Y(_29022_) );
  \$mux  #( .WIDTH(1) ) _54100_ ( .A(_29055_), .B(_29056_), .S(_counter_data_782[1]), .Y(_29025_) );
  \$mux  #( .WIDTH(1) ) _54101_ ( .A(_29025_), .B(1'hx), .S(_counter_data_782[2]), .Y(_29026_) );
  \$mux  #( .WIDTH(1) ) _54102_ ( .A(_29026_), .B(1'hx), .S(_counter_data_782[3]), .Y(_29027_) );
  \$mux  #( .WIDTH(1) ) _54103_ ( .A(_29027_), .B(1'hx), .S(_counter_data_782[4]), .Y(_29028_) );
  \$mux  #( .WIDTH(1) ) _54104_ ( .A(_29028_), .B(1'hx), .S(_counter_data_782[5]), .Y(_29029_) );
  \$mux  #( .WIDTH(1) ) _54105_ ( .A(_29029_), .B(1'hx), .S(_counter_data_782[6]), .Y(_29030_) );
  \$mux  #( .WIDTH(1) ) _54106_ ( .A(_29030_), .B(1'hx), .S(_counter_data_782[7]), .Y(_29031_) );
  \$mux  #( .WIDTH(1) ) _54107_ ( .A(_29031_), .B(1'hx), .S(_counter_data_782[8]), .Y(_29032_) );
  \$mux  #( .WIDTH(1) ) _54108_ ( .A(_29032_), .B(1'hx), .S(_counter_data_782[9]), .Y(_29033_) );
  \$mux  #( .WIDTH(1) ) _54109_ ( .A(_29033_), .B(1'hx), .S(_counter_data_782[10]), .Y(_29034_) );
  \$mux  #( .WIDTH(1) ) _54110_ ( .A(_29034_), .B(1'hx), .S(_counter_data_782[11]), .Y(_29035_) );
  \$mux  #( .WIDTH(1) ) _54111_ ( .A(_29035_), .B(1'hx), .S(_counter_data_782[12]), .Y(_29036_) );
  \$mux  #( .WIDTH(1) ) _54112_ ( .A(_29036_), .B(1'hx), .S(_counter_data_782[13]), .Y(_29037_) );
  \$mux  #( .WIDTH(1) ) _54113_ ( .A(_29037_), .B(1'hx), .S(_counter_data_782[14]), .Y(_29038_) );
  \$mux  #( .WIDTH(1) ) _54114_ ( .A(_29038_), .B(1'hx), .S(_counter_data_782[15]), .Y(_29039_) );
  \$mux  #( .WIDTH(1) ) _54115_ ( .A(_29039_), .B(1'hx), .S(_counter_data_782[16]), .Y(_29040_) );
  \$mux  #( .WIDTH(1) ) _54116_ ( .A(_29040_), .B(1'hx), .S(_counter_data_782[17]), .Y(_29041_) );
  \$mux  #( .WIDTH(1) ) _54117_ ( .A(_29041_), .B(1'hx), .S(_counter_data_782[18]), .Y(_29042_) );
  \$mux  #( .WIDTH(1) ) _54118_ ( .A(_29042_), .B(1'hx), .S(_counter_data_782[19]), .Y(_29043_) );
  \$mux  #( .WIDTH(1) ) _54119_ ( .A(_29043_), .B(1'hx), .S(_counter_data_782[20]), .Y(_29044_) );
  \$mux  #( .WIDTH(1) ) _54120_ ( .A(_29044_), .B(1'hx), .S(_counter_data_782[21]), .Y(_29045_) );
  \$mux  #( .WIDTH(1) ) _54121_ ( .A(_29045_), .B(1'hx), .S(_counter_data_782[22]), .Y(_29046_) );
  \$mux  #( .WIDTH(1) ) _54122_ ( .A(_29046_), .B(1'hx), .S(_counter_data_782[23]), .Y(_29047_) );
  \$mux  #( .WIDTH(1) ) _54123_ ( .A(_29047_), .B(1'hx), .S(_counter_data_782[24]), .Y(_29048_) );
  \$mux  #( .WIDTH(1) ) _54124_ ( .A(_29048_), .B(1'hx), .S(_counter_data_782[25]), .Y(_29049_) );
  \$mux  #( .WIDTH(1) ) _54125_ ( .A(_29049_), .B(1'hx), .S(_counter_data_782[26]), .Y(_29050_) );
  \$mux  #( .WIDTH(1) ) _54126_ ( .A(_29050_), .B(1'hx), .S(_counter_data_782[27]), .Y(_29051_) );
  \$mux  #( .WIDTH(1) ) _54127_ ( .A(_29051_), .B(1'hx), .S(_counter_data_782[28]), .Y(_29052_) );
  \$mux  #( .WIDTH(1) ) _54128_ ( .A(_29052_), .B(1'hx), .S(_counter_data_782[29]), .Y(_29053_) );
  \$mux  #( .WIDTH(1) ) _54129_ ( .A(_29053_), .B(1'hx), .S(_counter_data_782[30]), .Y(_29054_) );
  \$mux  #( .WIDTH(1) ) _54130_ ( .A(__delay_data_1411[0]), .B(__delay_data_1411[1]), .S(_counter_data_782[0]), .Y(_29055_) );
  \$mux  #( .WIDTH(1) ) _54131_ ( .A(__delay_data_1411[2]), .B(__delay_data_1411[3]), .S(_counter_data_782[0]), .Y(_29056_) );
  \$mux  #( .WIDTH(8) ) _54200_ ( .A(__tmp_977_1), .B(ram_w8_l2048_id11_0_1_rdata), .S(__tmp_976_1), .Y(_tmp_977) );
  \$mux  #( .WIDTH(8) ) _54201_ ( .A(__tmp_989_1), .B(ram_w8_l2048_id11_1_1_rdata), .S(__tmp_988_1), .Y(_tmp_989) );
  \$mux  #( .WIDTH(8) ) _54202_ ( .A(__tmp_1001_1), .B(ram_w8_l2048_id11_2_1_rdata), .S(__tmp_1000_1), .Y(_tmp_1001) );
  \$mux  #( .WIDTH(8) ) _54203_ ( .A(__tmp_1013_1), .B(ram_w8_l2048_id11_3_1_rdata), .S(__tmp_1012_1), .Y(_tmp_1013) );
  \$mux  #( .WIDTH(32) ) _54204_ ( .A(_29057_), .B(_29058_), .S(_05845_), .Y(_29059_) );
  \$mux  #( .WIDTH(32) ) _54205_ ( .A(1), .B(_29059_), .S(_05713_), .Y({ _29060_[31:1], conv2d_16_mux_next_dma_flag_0 }) );
  \$mux  #( .WIDTH(32) ) _54206_ ( .A(_29057_), .B(0), .S(_05846_), .Y(_29058_) );
  \$mux  #( .WIDTH(32) ) _54207_ ( .A(1), .B(_29058_), .S(_05845_), .Y(_29061_) );
  \$mux  #( .WIDTH(32) ) _54208_ ( .A(_29057_), .B(_29061_), .S(_05713_), .Y({ _29062_[31:1], conv2d_16_mux_next_dma_flag_1 }) );
  \$mux  #( .WIDTH(32) ) _54209_ ( .A(0), .B(1), .S(conv2d_16_update_filter), .Y(_29057_) );
  \$mux  #( .WIDTH(32) ) _54210_ ( .A(1), .B(0), .S(_05846_), .Y(_29063_) );
  \$mux  #( .WIDTH(32) ) _54211_ ( .A(_29057_), .B(_29063_), .S(_05845_), .Y(_29064_) );
  \$mux  #( .WIDTH(32) ) _54212_ ( .A(_29057_), .B(_29064_), .S(_05713_), .Y({ _29065_[31:1], conv2d_16_mux_next_dma_flag_2 }) );
  \$mux  #( .WIDTH(32) ) _54213_ ( .A({ 24'h000000, ram_w8_l2048_id1_3_0_rdata }), .B(0), .S(_05849_), .Y(_29066_) );
  \$mux  #( .WIDTH(32) ) _54214_ ( .A({ 24'h000000, ram_w8_l2048_id1_2_0_rdata }), .B(_29066_), .S(_05848_), .Y(_29067_) );
  \$mux  #( .WIDTH(32) ) _54215_ ( .A({ 24'h000000, ram_w8_l2048_id1_1_0_rdata }), .B(_29067_), .S(_05847_), .Y(_29068_) );
  \$mux  #( .WIDTH(32) ) _54216_ ( .A({ 24'h000000, ram_w8_l2048_id1_0_0_rdata }), .B(_29068_), .S(_05714_), .Y({ _29069_[31:8], _tmp_1032 }) );
  \$mux  #( .WIDTH(32) ) _54217_ ( .A({ _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032[7], _tmp_1032 }), .B(0), .S(_05892_), .Y({ _29070_[31:8], _stream_max_pool_serial_18_source_1_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54218_ ( .A(0), .B(1), .S(_set_flag_1038), .Y({ _29071_[31:1], _stream_max_pool_serial_18_start_flag }) );
  \$mux  #( .WIDTH(8) ) _54219_ ( .A(__tmp_1078_1), .B(ram_w8_l2048_id0_0_1_rdata), .S(__tmp_1077_1), .Y(_tmp_1078) );
  \$mux  #( .WIDTH(8) ) _54220_ ( .A(__tmp_1090_1), .B(ram_w8_l2048_id0_1_1_rdata), .S(__tmp_1089_1), .Y(_tmp_1090) );
  \$mux  #( .WIDTH(8) ) _54221_ ( .A(__tmp_1102_1), .B(ram_w8_l2048_id0_2_1_rdata), .S(__tmp_1101_1), .Y(_tmp_1102) );
  \$mux  #( .WIDTH(8) ) _54222_ ( .A(__tmp_1114_1), .B(ram_w8_l2048_id0_3_1_rdata), .S(__tmp_1113_1), .Y(_tmp_1114) );
  \$mux  #( .WIDTH(32) ) _54223_ ( .A(_24202_), .B(0), .S(matmul_29_row_select), .Y(matmul_29_mux_act_gaddr_0) );
  \$mux  #( .WIDTH(1) ) _54224_ ( .A(matmul_29_dma_pad_mask_0), .B(1'h0), .S(matmul_29_row_select), .Y(matmul_29_mux_dma_pad_mask_0) );
  \$mux  #( .WIDTH(1) ) _54225_ ( .A(matmul_29_dma_flag_0), .B(1'h0), .S(matmul_29_prev_row_select), .Y(matmul_29_mux_dma_flag_0) );
  \$mux  #( .WIDTH(32) ) _54226_ ( .A({ 24'h000000, ram_w8_l2048_id2_3_0_rdata }), .B(0), .S(_05852_), .Y(_29072_) );
  \$mux  #( .WIDTH(32) ) _54227_ ( .A({ 24'h000000, ram_w8_l2048_id2_2_0_rdata }), .B(_29072_), .S(_05851_), .Y(_29073_) );
  \$mux  #( .WIDTH(32) ) _54228_ ( .A({ 24'h000000, ram_w8_l2048_id2_1_0_rdata }), .B(_29073_), .S(_05850_), .Y(_29074_) );
  \$mux  #( .WIDTH(32) ) _54229_ ( .A({ 24'h000000, ram_w8_l2048_id2_0_0_rdata }), .B(_29074_), .S(_05715_), .Y({ _29075_[31:8], _tmp_1175 }) );
  \$mux  #( .WIDTH(32) ) _54230_ ( .A({ _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175[7], _tmp_1175 }), .B(0), .S(_05894_), .Y({ _29076_[31:8], _stream_matmul_29_source_6_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54231_ ( .A({ 24'h000000, ram_w8_l2048_id0_3_0_rdata }), .B(0), .S(_05855_), .Y(_29077_) );
  \$mux  #( .WIDTH(32) ) _54232_ ( .A({ 24'h000000, ram_w8_l2048_id0_2_0_rdata }), .B(_29077_), .S(_05854_), .Y(_29078_) );
  \$mux  #( .WIDTH(32) ) _54233_ ( .A({ 24'h000000, ram_w8_l2048_id0_1_0_rdata }), .B(_29078_), .S(_05853_), .Y(_29079_) );
  \$mux  #( .WIDTH(32) ) _54234_ ( .A({ 24'h000000, ram_w8_l2048_id0_0_0_rdata }), .B(_29079_), .S(_05716_), .Y({ _29080_[31:8], _tmp_1186 }) );
  \$mux  #( .WIDTH(32) ) _54235_ ( .A({ _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186[7], _tmp_1186 }), .B(0), .S(_05890_), .Y({ _29081_[31:8], _stream_matmul_29_source_8_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54236_ ( .A({ 24'h000000, ram_w8_l2048_id3_3_0_rdata }), .B(0), .S(_05858_), .Y(_29082_) );
  \$mux  #( .WIDTH(32) ) _54237_ ( .A({ 24'h000000, ram_w8_l2048_id3_2_0_rdata }), .B(_29082_), .S(_05857_), .Y(_29083_) );
  \$mux  #( .WIDTH(32) ) _54238_ ( .A({ 24'h000000, ram_w8_l2048_id3_1_0_rdata }), .B(_29083_), .S(_05856_), .Y(_29084_) );
  \$mux  #( .WIDTH(32) ) _54239_ ( .A({ 24'h000000, ram_w8_l2048_id3_0_0_rdata }), .B(_29084_), .S(_05717_), .Y({ _29085_[31:8], _tmp_1206 }) );
  \$mux  #( .WIDTH(32) ) _54240_ ( .A({ _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206[7], _tmp_1206 }), .B(0), .S(_05896_), .Y({ _29086_[31:8], _stream_matmul_29_source_19_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54241_ ( .A({ 28'h0000000, ram_w4_l8192_id0_7_0_rdata }), .B(0), .S(_05865_), .Y(_29087_) );
  \$mux  #( .WIDTH(32) ) _54242_ ( .A({ 28'h0000000, ram_w4_l8192_id0_6_0_rdata }), .B(_29087_), .S(_05864_), .Y(_29088_) );
  \$mux  #( .WIDTH(32) ) _54243_ ( .A({ 28'h0000000, ram_w4_l8192_id0_5_0_rdata }), .B(_29088_), .S(_05863_), .Y(_29089_) );
  \$mux  #( .WIDTH(32) ) _54244_ ( .A({ 28'h0000000, ram_w4_l8192_id0_4_0_rdata }), .B(_29089_), .S(_05862_), .Y(_29090_) );
  \$mux  #( .WIDTH(32) ) _54245_ ( .A({ 28'h0000000, ram_w4_l8192_id0_3_0_rdata }), .B(_29090_), .S(_05861_), .Y(_29091_) );
  \$mux  #( .WIDTH(32) ) _54246_ ( .A({ 28'h0000000, ram_w4_l8192_id0_2_0_rdata }), .B(_29091_), .S(_05860_), .Y(_29092_) );
  \$mux  #( .WIDTH(32) ) _54247_ ( .A({ 28'h0000000, ram_w4_l8192_id0_1_0_rdata }), .B(_29092_), .S(_05859_), .Y(_29093_) );
  \$mux  #( .WIDTH(32) ) _54248_ ( .A({ 28'h0000000, ram_w4_l8192_id0_0_0_rdata }), .B(_29093_), .S(_05718_), .Y({ _29094_[31:4], _tmp_1220 }) );
  \$mux  #( .WIDTH(32) ) _54249_ ( .A({ _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220[3], _tmp_1220 }), .B(0), .S(_05880_), .Y({ _29095_[31:4], _stream_matmul_29_source_20_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54250_ ( .A(0), .B(1), .S(_06177_), .Y({ _29096_[31:1], _stream_matmul_29_start_flag }) );
  \$mux  #( .WIDTH(8) ) _54251_ ( .A(__tmp_1315_1), .B(ram_w8_l2048_id1_0_1_rdata), .S(__tmp_1314_1), .Y(_tmp_1315) );
  \$mux  #( .WIDTH(8) ) _54252_ ( .A(__tmp_1327_1), .B(ram_w8_l2048_id1_1_1_rdata), .S(__tmp_1326_1), .Y(_tmp_1327) );
  \$mux  #( .WIDTH(8) ) _54253_ ( .A(__tmp_1339_1), .B(ram_w8_l2048_id1_2_1_rdata), .S(__tmp_1338_1), .Y(_tmp_1339) );
  \$mux  #( .WIDTH(8) ) _54254_ ( .A(__tmp_1351_1), .B(ram_w8_l2048_id1_3_1_rdata), .S(__tmp_1350_1), .Y(_tmp_1351) );
  \$mux  #( .WIDTH(32) ) _54255_ ( .A(0), .B(1), .S(_06180_), .Y(_29097_) );
  \$mux  #( .WIDTH(32) ) _54256_ ( .A(_29097_), .B(1), .S(_06179_), .Y(_29098_) );
  \$mux  #( .WIDTH(32) ) _54257_ ( .A(_29098_), .B(1), .S(_06178_), .Y({ _29099_[31:1], _maxi_write_data_done }) );
  \$mux  #( .WIDTH(32) ) _54258_ ( .A(1), .B(0), .S(_24020_), .Y(_29100_) );
  \$mux  #( .WIDTH(32) ) _54259_ ( .A(1), .B(0), .S(_24021_), .Y(_29101_) );
  \$mux  #( .WIDTH(32) ) _54260_ ( .A(1), .B(0), .S(_24022_), .Y(_29102_) );
  \$mux  #( .WIDTH(32) ) _54261_ ( .A(1), .B(0), .S(_24023_), .Y(_29103_) );
  \$mux  #( .WIDTH(32) ) _54262_ ( .A(1), .B(0), .S(_24024_), .Y(_29104_) );
  \$mux  #( .WIDTH(32) ) _54263_ ( .A(1), .B(0), .S(_24025_), .Y(_29105_) );
  \$mux  #( .WIDTH(32) ) _54264_ ( .A(1), .B(0), .S(_24026_), .Y(_29106_) );
  \$mux  #( .WIDTH(32) ) _54265_ ( .A(1), .B(0), .S(_24027_), .Y(_29107_) );
  \$mux  #( .WIDTH(32) ) _54266_ ( .A(_saxi_register_13), .B(32'hxxxxxxxx), .S(_05878_), .Y(_29108_) );
  \$mux  #( .WIDTH(32) ) _54267_ ( .A(_saxi_register_12), .B(_29108_), .S(_05877_), .Y(_29109_) );
  \$mux  #( .WIDTH(32) ) _54268_ ( .A(_saxi_register_11), .B(_29109_), .S(_05876_), .Y(_29110_) );
  \$mux  #( .WIDTH(32) ) _54269_ ( .A(_saxi_register_10), .B(_29110_), .S(_05875_), .Y(_29111_) );
  \$mux  #( .WIDTH(32) ) _54270_ ( .A(_saxi_register_9), .B(_29111_), .S(_05874_), .Y(_29112_) );
  \$mux  #( .WIDTH(32) ) _54271_ ( .A(_saxi_register_8), .B(_29112_), .S(_05873_), .Y(_29113_) );
  \$mux  #( .WIDTH(32) ) _54272_ ( .A(_saxi_register_7), .B(_29113_), .S(_05872_), .Y(_29114_) );
  \$mux  #( .WIDTH(32) ) _54273_ ( .A(_saxi_register_6), .B(_29114_), .S(_05871_), .Y(_29115_) );
  \$mux  #( .WIDTH(32) ) _54274_ ( .A(_saxi_register_5), .B(_29115_), .S(_05870_), .Y(_29116_) );
  \$mux  #( .WIDTH(32) ) _54275_ ( .A(_saxi_register_4), .B(_29116_), .S(_05869_), .Y(_29117_) );
  \$mux  #( .WIDTH(32) ) _54276_ ( .A(_saxi_register_3), .B(_29117_), .S(_05868_), .Y(_29118_) );
  \$mux  #( .WIDTH(32) ) _54277_ ( .A(_saxi_register_2), .B(_29118_), .S(_05867_), .Y(_29119_) );
  \$mux  #( .WIDTH(32) ) _54278_ ( .A(_saxi_register_1), .B(_29119_), .S(_05866_), .Y(_29120_) );
  \$mux  #( .WIDTH(32) ) _54279_ ( .A(_saxi_register_0), .B(_29120_), .S(_05719_), .Y(_tmp_6) );
  \$mux  #( .WIDTH(32) ) _54280_ ( .A({ 31'h00000000, _saxi_flag_13 }), .B(32'hxxxxxxxx), .S(_05878_), .Y(_29121_) );
  \$mux  #( .WIDTH(32) ) _54281_ ( .A({ 31'h00000000, _saxi_flag_12 }), .B(_29121_), .S(_05877_), .Y(_29122_) );
  \$mux  #( .WIDTH(32) ) _54282_ ( .A({ 31'h00000000, _saxi_flag_11 }), .B(_29122_), .S(_05876_), .Y(_29123_) );
  \$mux  #( .WIDTH(32) ) _54283_ ( .A({ 31'h00000000, _saxi_flag_10 }), .B(_29123_), .S(_05875_), .Y(_29124_) );
  \$mux  #( .WIDTH(32) ) _54284_ ( .A({ 31'h00000000, _saxi_flag_9 }), .B(_29124_), .S(_05874_), .Y(_29125_) );
  \$mux  #( .WIDTH(32) ) _54285_ ( .A({ 31'h00000000, _saxi_flag_8 }), .B(_29125_), .S(_05873_), .Y(_29126_) );
  \$mux  #( .WIDTH(32) ) _54286_ ( .A({ 31'h00000000, _saxi_flag_7 }), .B(_29126_), .S(_05872_), .Y(_29127_) );
  \$mux  #( .WIDTH(32) ) _54287_ ( .A({ 31'h00000000, _saxi_flag_6 }), .B(_29127_), .S(_05871_), .Y(_29128_) );
  \$mux  #( .WIDTH(32) ) _54288_ ( .A({ 31'h00000000, _saxi_flag_5 }), .B(_29128_), .S(_05870_), .Y(_29129_) );
  \$mux  #( .WIDTH(32) ) _54289_ ( .A({ 31'h00000000, _saxi_flag_4 }), .B(_29129_), .S(_05869_), .Y(_29130_) );
  \$mux  #( .WIDTH(32) ) _54290_ ( .A({ 31'h00000000, _saxi_flag_3 }), .B(_29130_), .S(_05868_), .Y(_29131_) );
  \$mux  #( .WIDTH(32) ) _54291_ ( .A({ 31'h00000000, _saxi_flag_2 }), .B(_29131_), .S(_05867_), .Y(_29132_) );
  \$mux  #( .WIDTH(32) ) _54292_ ( .A({ 31'h00000000, _saxi_flag_1 }), .B(_29132_), .S(_05866_), .Y(_29133_) );
  \$mux  #( .WIDTH(32) ) _54293_ ( .A({ 31'h00000000, _saxi_flag_0 }), .B(_29133_), .S(_05719_), .Y({ _29134_[31:1], _tmp_7 }) );
  \$mux  #( .WIDTH(32) ) _54294_ ( .A(_saxi_resetval_13), .B(32'hxxxxxxxx), .S(_05878_), .Y(_29135_) );
  \$mux  #( .WIDTH(32) ) _54295_ ( .A(_saxi_resetval_12), .B(_29135_), .S(_05877_), .Y(_29136_) );
  \$mux  #( .WIDTH(32) ) _54296_ ( .A(_saxi_resetval_11), .B(_29136_), .S(_05876_), .Y(_29137_) );
  \$mux  #( .WIDTH(32) ) _54297_ ( .A(_saxi_resetval_10), .B(_29137_), .S(_05875_), .Y(_29138_) );
  \$mux  #( .WIDTH(32) ) _54298_ ( .A(_saxi_resetval_9), .B(_29138_), .S(_05874_), .Y(_29139_) );
  \$mux  #( .WIDTH(32) ) _54299_ ( .A(_saxi_resetval_8), .B(_29139_), .S(_05873_), .Y(_29140_) );
  \$mux  #( .WIDTH(32) ) _54300_ ( .A(_saxi_resetval_7), .B(_29140_), .S(_05872_), .Y(_29141_) );
  \$mux  #( .WIDTH(32) ) _54301_ ( .A(_saxi_resetval_6), .B(_29141_), .S(_05871_), .Y(_29142_) );
  \$mux  #( .WIDTH(32) ) _54302_ ( .A(_saxi_resetval_5), .B(_29142_), .S(_05870_), .Y(_29143_) );
  \$mux  #( .WIDTH(32) ) _54303_ ( .A(_saxi_resetval_4), .B(_29143_), .S(_05869_), .Y(_29144_) );
  \$mux  #( .WIDTH(32) ) _54304_ ( .A(_saxi_resetval_3), .B(_29144_), .S(_05868_), .Y(_29145_) );
  \$mux  #( .WIDTH(32) ) _54305_ ( .A(_saxi_resetval_2), .B(_29145_), .S(_05867_), .Y(_29146_) );
  \$mux  #( .WIDTH(32) ) _54306_ ( .A(_saxi_resetval_1), .B(_29146_), .S(_05866_), .Y(_29147_) );
  \$mux  #( .WIDTH(32) ) _54307_ ( .A(_saxi_resetval_0), .B(_29147_), .S(_05719_), .Y(_tmp_8) );
  \$mux  #( .WIDTH(33) ) _54308_ ( .A(_24291_), .B(33'h000000000), .S(_06147_), .Y(_29148_) );
  \$mux  #( .WIDTH(33) ) _54309_ ( .A(_24292_), .B(33'h000000000), .S(_06148_), .Y(_29149_) );
  \$mux  #( .WIDTH(66) ) _54310_ ( .A(66'h00000000000000000), .B(_sll_data_7), .S(__delay_data_748), .Y(_29150_) );
  \$mux  #( .WIDTH(40) ) _54311_ ( .A(__delay_data_768), .B(40'h000000007f), .S(_greaterthan_data_43), .Y(_29151_) );
  \$mux  #( .WIDTH(40) ) _54312_ ( .A(__delay_data_768), .B(40'hffffffff81), .S(_lessthan_data_47), .Y(_29152_) );
  \$mux  #( .WIDTH(40) ) _54313_ ( .A(_cond_data_49), .B(_cond_data_45), .S(__delay_data_769), .Y(_29153_) );
  \$mux  #( .WIDTH(18) ) _54314_ ( .A(18'h00000), .B(_sll_data_61), .S(__delay_data_593), .Y(_29154_) );
  \$mux  #( .WIDTH(18) ) _54315_ ( .A(18'h00000), .B(_sll_data_78), .S(__delay_data_610), .Y(_29155_) );
  \$mux  #( .WIDTH(18) ) _54316_ ( .A(18'h00000), .B(_sll_data_95), .S(__delay_data_627), .Y(_29156_) );
  \$mux  #( .WIDTH(18) ) _54317_ ( .A(18'h00000), .B(_sll_data_112), .S(__delay_data_644), .Y(_29157_) );
  \$mux  #( .WIDTH(18) ) _54318_ ( .A(18'h00000), .B(_sll_data_129), .S(__delay_data_661), .Y(_29158_) );
  \$mux  #( .WIDTH(18) ) _54319_ ( .A(18'h00000), .B(_sll_data_146), .S(__delay_data_678), .Y(_29159_) );
  \$mux  #( .WIDTH(18) ) _54320_ ( .A(18'h00000), .B(_sll_data_163), .S(__delay_data_695), .Y(_29160_) );
  \$mux  #( .WIDTH(18) ) _54321_ ( .A(18'h00000), .B(_sll_data_180), .S(__delay_data_712), .Y(_29161_) );
  \$mux  #( .WIDTH(18) ) _54322_ ( .A(18'h00000), .B(_sll_data_197), .S(__delay_data_729), .Y(_29162_) );
  \$mux  #( .WIDTH(8) ) _54323_ ( .A(_reducemax_data_211), .B(__variable_wdata_207), .S(_06884_), .Y(_29163_) );
  \$mux  #( .WIDTH(32) ) _54324_ ( .A(_24302_), .B(0), .S(_06150_), .Y(_29164_) );
  \$mux  #( .WIDTH(9) ) _54325_ ( .A({ __variable_wdata_207[7], __variable_wdata_207 }), .B(9'h180), .S(_24029_), .Y(_29165_) );
  \$mux  #( .WIDTH(32) ) _54326_ ( .A(_24303_), .B(0), .S(_06151_), .Y(_29166_) );
  \$mux  #( .WIDTH(8) ) _54327_ ( .A(8'h00), .B(__delay_data_898), .S(_eq_data_357), .Y(_29167_) );
  \$mux  #( .WIDTH(8) ) _54328_ ( .A(8'h00), .B(__delay_data_904), .S(_eq_data_357), .Y(_29168_) );
  \$mux  #( .WIDTH(8) ) _54329_ ( .A(8'h00), .B(__delay_data_900), .S(_eq_data_357), .Y(_29169_) );
  \$mux  #( .WIDTH(8) ) _54330_ ( .A(8'h00), .B(__delay_data_907), .S(_eq_data_357), .Y(_29170_) );
  \$mux  #( .WIDTH(8) ) _54331_ ( .A(8'h00), .B(__delay_data_913), .S(_eq_data_357), .Y(_29171_) );
  \$mux  #( .WIDTH(8) ) _54332_ ( .A(8'h00), .B(__delay_data_909), .S(_eq_data_357), .Y(_29172_) );
  \$mux  #( .WIDTH(8) ) _54333_ ( .A(8'h00), .B(__delay_data_916), .S(_eq_data_357), .Y(_29173_) );
  \$mux  #( .WIDTH(8) ) _54334_ ( .A(8'h00), .B(__delay_data_922), .S(_eq_data_357), .Y(_29174_) );
  \$mux  #( .WIDTH(8) ) _54335_ ( .A(8'h00), .B(__delay_data_918), .S(_eq_data_357), .Y(_29175_) );
  \$mux  #( .WIDTH(8) ) _54336_ ( .A(_cond_data_279), .B(__delay_data_901), .S(__delay_data_1021), .Y(_29176_) );
  \$mux  #( .WIDTH(8) ) _54337_ ( .A(_cond_data_289), .B(__delay_data_963), .S(__delay_data_1021), .Y(_29177_) );
  \$mux  #( .WIDTH(8) ) _54338_ ( .A(_cond_data_299), .B(__delay_data_905), .S(__delay_data_1021), .Y(_29178_) );
  \$mux  #( .WIDTH(8) ) _54339_ ( .A(_cond_data_309), .B(__delay_data_910), .S(__delay_data_1021), .Y(_29179_) );
  \$mux  #( .WIDTH(8) ) _54340_ ( .A(_cond_data_319), .B(__delay_data_968), .S(__delay_data_1021), .Y(_29180_) );
  \$mux  #( .WIDTH(8) ) _54341_ ( .A(_cond_data_329), .B(__delay_data_914), .S(__delay_data_1021), .Y(_29181_) );
  \$mux  #( .WIDTH(8) ) _54342_ ( .A(_cond_data_339), .B(__delay_data_919), .S(__delay_data_1021), .Y(_29182_) );
  \$mux  #( .WIDTH(8) ) _54343_ ( .A(_cond_data_349), .B(__delay_data_973), .S(__delay_data_1021), .Y(_29183_) );
  \$mux  #( .WIDTH(8) ) _54344_ ( .A(_cond_data_359), .B(__delay_data_923), .S(__delay_data_1021), .Y(_29184_) );
  \$mux  #( .WIDTH(8) ) _54345_ ( .A(_cond_data_283), .B(__delay_data_906), .S(__delay_data_1023), .Y(_29185_) );
  \$mux  #( .WIDTH(8) ) _54346_ ( .A(_cond_data_293), .B(__delay_data_966), .S(__delay_data_1023), .Y(_29186_) );
  \$mux  #( .WIDTH(8) ) _54347_ ( .A(_cond_data_303), .B(__delay_data_1016), .S(__delay_data_1023), .Y(_29187_) );
  \$mux  #( .WIDTH(8) ) _54348_ ( .A(_cond_data_313), .B(__delay_data_915), .S(__delay_data_1023), .Y(_29188_) );
  \$mux  #( .WIDTH(8) ) _54349_ ( .A(_cond_data_323), .B(__delay_data_971), .S(__delay_data_1023), .Y(_29189_) );
  \$mux  #( .WIDTH(8) ) _54350_ ( .A(_cond_data_333), .B(__delay_data_1020), .S(__delay_data_1023), .Y(_29190_) );
  \$mux  #( .WIDTH(8) ) _54351_ ( .A(_cond_data_343), .B(__delay_data_924), .S(__delay_data_1023), .Y(_29191_) );
  \$mux  #( .WIDTH(8) ) _54352_ ( .A(_cond_data_353), .B(__delay_data_976), .S(__delay_data_1023), .Y(_29192_) );
  \$mux  #( .WIDTH(8) ) _54353_ ( .A(_cond_data_363), .B(__delay_data_1024), .S(__delay_data_1023), .Y(_29193_) );
  \$mux  #( .WIDTH(8) ) _54354_ ( .A(8'h00), .B(_cond_data_346), .S(__delay_data_1236), .Y(_29194_) );
  \$mux  #( .WIDTH(8) ) _54355_ ( .A(8'h00), .B(_cond_data_286), .S(__delay_data_1236), .Y(_29195_) );
  \$mux  #( .WIDTH(8) ) _54356_ ( .A(8'h00), .B(_cond_data_316), .S(__delay_data_1236), .Y(_29196_) );
  \$mux  #( .WIDTH(8) ) _54357_ ( .A(8'h00), .B(_cond_data_356), .S(__delay_data_1236), .Y(_29197_) );
  \$mux  #( .WIDTH(8) ) _54358_ ( .A(8'h00), .B(_cond_data_296), .S(__delay_data_1236), .Y(_29198_) );
  \$mux  #( .WIDTH(8) ) _54359_ ( .A(8'h00), .B(_cond_data_326), .S(__delay_data_1236), .Y(_29199_) );
  \$mux  #( .WIDTH(8) ) _54360_ ( .A(8'h00), .B(_cond_data_366), .S(__delay_data_1236), .Y(_29200_) );
  \$mux  #( .WIDTH(8) ) _54361_ ( .A(8'h00), .B(_cond_data_306), .S(__delay_data_1236), .Y(_29201_) );
  \$mux  #( .WIDTH(8) ) _54362_ ( .A(8'h00), .B(_cond_data_336), .S(__delay_data_1236), .Y(_29202_) );
  \$mux  #( .WIDTH(8) ) _54363_ ( .A(_cond_data_369), .B(__delay_data_932), .S(__delay_data_1240), .Y(_29203_) );
  \$mux  #( .WIDTH(8) ) _54364_ ( .A(_cond_data_379), .B(__delay_data_1068), .S(__delay_data_1240), .Y(_29204_) );
  \$mux  #( .WIDTH(8) ) _54365_ ( .A(_cond_data_389), .B(__delay_data_938), .S(__delay_data_1240), .Y(_29205_) );
  \$mux  #( .WIDTH(8) ) _54366_ ( .A(_cond_data_399), .B(__delay_data_984), .S(__delay_data_1240), .Y(_29206_) );
  \$mux  #( .WIDTH(8) ) _54367_ ( .A(_cond_data_409), .B(__delay_data_1103), .S(__delay_data_1240), .Y(_29207_) );
  \$mux  #( .WIDTH(8) ) _54368_ ( .A(_cond_data_419), .B(__delay_data_990), .S(__delay_data_1240), .Y(_29208_) );
  \$mux  #( .WIDTH(8) ) _54369_ ( .A(_cond_data_429), .B(__delay_data_1032), .S(__delay_data_1240), .Y(_29209_) );
  \$mux  #( .WIDTH(8) ) _54370_ ( .A(_cond_data_439), .B(__delay_data_1138), .S(__delay_data_1240), .Y(_29210_) );
  \$mux  #( .WIDTH(8) ) _54371_ ( .A(_cond_data_449), .B(__delay_data_1038), .S(__delay_data_1240), .Y(_29211_) );
  \$mux  #( .WIDTH(8) ) _54372_ ( .A(_cond_data_373), .B(__delay_data_939), .S(__delay_data_1245), .Y(_29212_) );
  \$mux  #( .WIDTH(8) ) _54373_ ( .A(_cond_data_383), .B(__delay_data_1074), .S(__delay_data_1245), .Y(_29213_) );
  \$mux  #( .WIDTH(8) ) _54374_ ( .A(_cond_data_393), .B(__delay_data_1178), .S(__delay_data_1245), .Y(_29214_) );
  \$mux  #( .WIDTH(8) ) _54375_ ( .A(_cond_data_403), .B(__delay_data_991), .S(__delay_data_1245), .Y(_29215_) );
  \$mux  #( .WIDTH(8) ) _54376_ ( .A(_cond_data_413), .B(__delay_data_1109), .S(__delay_data_1245), .Y(_29216_) );
  \$mux  #( .WIDTH(8) ) _54377_ ( .A(_cond_data_423), .B(__delay_data_1212), .S(__delay_data_1245), .Y(_29217_) );
  \$mux  #( .WIDTH(8) ) _54378_ ( .A(_cond_data_433), .B(__delay_data_1039), .S(__delay_data_1245), .Y(_29218_) );
  \$mux  #( .WIDTH(8) ) _54379_ ( .A(_cond_data_443), .B(__delay_data_1144), .S(__delay_data_1245), .Y(_29219_) );
  \$mux  #( .WIDTH(8) ) _54380_ ( .A(_cond_data_453), .B(__delay_data_1246), .S(__delay_data_1245), .Y(_29220_) );
  \$mux  #( .WIDTH(8) ) _54381_ ( .A(_cond_data_376), .B(8'h00), .S(__delay_data_946), .Y(_29221_) );
  \$mux  #( .WIDTH(8) ) _54382_ ( .A(_cond_data_406), .B(8'h00), .S(__delay_data_998), .Y(_29222_) );
  \$mux  #( .WIDTH(8) ) _54383_ ( .A(_cond_data_436), .B(8'h00), .S(__delay_data_1046), .Y(_29223_) );
  \$mux  #( .WIDTH(8) ) _54384_ ( .A(_cond_data_386), .B(8'h00), .S(__delay_data_1081), .Y(_29224_) );
  \$mux  #( .WIDTH(8) ) _54385_ ( .A(_cond_data_416), .B(8'h00), .S(__delay_data_1116), .Y(_29225_) );
  \$mux  #( .WIDTH(8) ) _54386_ ( .A(_cond_data_446), .B(8'h00), .S(__delay_data_1151), .Y(_29226_) );
  \$mux  #( .WIDTH(8) ) _54387_ ( .A(_cond_data_396), .B(8'h00), .S(__delay_data_1185), .Y(_29227_) );
  \$mux  #( .WIDTH(8) ) _54388_ ( .A(_cond_data_426), .B(8'h00), .S(__delay_data_1219), .Y(_29228_) );
  \$mux  #( .WIDTH(8) ) _54389_ ( .A(_cond_data_456), .B(8'h00), .S(__delay_data_1253), .Y(_29229_) );
  \$mux  #( .WIDTH(32) ) _54390_ ( .A(0), .B(conv2d_16_och_count_buf), .S(_05904_), .Y(_29231_) );
  \$mux  #( .WIDTH(32) ) _54391_ ( .A(0), .B(1), .S(_05904_), .Y(_29232_) );
  \$mux  #( .WIDTH(32) ) _54392_ ( .A(10), .B(11), .S(_05744_), .Y(_29237_) );
  \$mux  #( .WIDTH(32) ) _54393_ ( .A(12), .B(_29237_), .S(_05689_), .Y({ _29238_[31:4], cparam_conv2d_16_cshamt_out_value }) );
  \$mux  #( .WIDTH(32) ) _54394_ ( .A(15), .B(7), .S(_05744_), .Y(_29239_) );
  \$mux  #( .WIDTH(32) ) _54395_ ( .A(31), .B(_29239_), .S(_05689_), .Y({ _29240_[31:5], cparam_conv2d_16_max_col_count }) );
  \$mux  #( .WIDTH(32) ) _54396_ ( .A(64), .B(128), .S(_05744_), .Y(_29241_) );
  \$mux  #( .WIDTH(32) ) _54397_ ( .A(32), .B(_29241_), .S(_05689_), .Y({ _29242_[31:8], cparam_conv2d_16_och_count_step }) );
  \$mux  #( .WIDTH(32) ) _54398_ ( .A(-128), .B(-256), .S(_05689_), .Y(cparam_conv2d_16_act_offset_values_0) );
  \$mux  #( .WIDTH(32) ) _54399_ ( .A(128), .B(256), .S(_05689_), .Y(cparam_conv2d_16_act_offset_values_2) );
  \$mux  #( .WIDTH(32) ) _54400_ ( .A(44), .B(96), .S(_05689_), .Y({ _29245_[31:7], cparam_conv2d_16_act_read_step }) );
  \$mux  #( .WIDTH(32) ) _54401_ ( .A(2304), .B(9216), .S(_05744_), .Y(_29246_) );
  \$mux  #( .WIDTH(32) ) _54402_ ( .A(576), .B(_29246_), .S(_05689_), .Y({ _29247_[31:14], cparam_conv2d_16_filter_base_step }) );
  \$mux  #( .WIDTH(32) ) _54403_ ( .A(4608), .B(18432), .S(_05744_), .Y(_29248_) );
  \$mux  #( .WIDTH(32) ) _54404_ ( .A(1152), .B(_29248_), .S(_05689_), .Y({ _29249_[31:15], cparam_conv2d_16_filter_read_size }) );
  \$mux  #( .WIDTH(32) ) _54405_ ( .A(512), .B(2048), .S(_05744_), .Y(_29251_) );
  \$mux  #( .WIDTH(32) ) _54406_ ( .A(128), .B(_29251_), .S(_05689_), .Y({ _29252_[31:12], cparam_conv2d_16_filter_read_step }) );
  \$mux  #( .WIDTH(32) ) _54407_ ( .A(3), .B(_29243_), .S(_05689_), .Y({ _29253_[31:6], cparam_conv2d_16_stream_reduce_size }) );
  \$mux  #( .WIDTH(32) ) _54408_ ( .A(8), .B(_29243_), .S(_05689_), .Y({ _29250_[31:6], cparam_conv2d_16_filter_read_block }) );
  \$mux  #( .WIDTH(32) ) _54409_ ( .A(16), .B(32), .S(_05744_), .Y(_29243_) );
  \$mux  #( .WIDTH(32) ) _54410_ ( .A(4), .B(_29243_), .S(_05689_), .Y({ _29244_[31:6], cparam_conv2d_16_inc_act_laddr_large }) );
  \$mux  #( .WIDTH(32) ) _54411_ ( .A(32), .B(64), .S(_05744_), .Y(_29235_) );
  \$mux  #( .WIDTH(32) ) _54412_ ( .A(16), .B(_29235_), .S(_05689_), .Y({ _29236_[31:7], cparam_conv2d_16_bias_num }) );
  \$mux  #( .WIDTH(32) ) _54413_ ( .A(-16), .B(-32), .S(_05744_), .Y(_29254_) );
  \$mux  #( .WIDTH(32) ) _54414_ ( .A(-4), .B(_29254_), .S(_05689_), .Y({ _29255_[31:7], cparam_conv2d_16_stream_act_local_large_offset }) );
  \$mux  #( .WIDTH(32) ) _54415_ ( .A(16), .B(8), .S(_05744_), .Y(_29233_) );
  \$mux  #( .WIDTH(32) ) _54416_ ( .A(32), .B(_29233_), .S(_05689_), .Y({ _29234_[31:6], cparam_conv2d_16_act_num_row }) );
  \$mux  #( .WIDTH(32) ) _54417_ ( .A(16), .B(8), .S(_05745_), .Y(_29256_) );
  \$mux  #( .WIDTH(32) ) _54418_ ( .A(32), .B(_29256_), .S(_05690_), .Y({ _29257_[31:6], cparam_max_pool_serial_18_act_num_col }) );
  \$mux  #( .WIDTH(32) ) _54419_ ( .A(13), .B(5), .S(_05745_), .Y(_29258_) );
  \$mux  #( .WIDTH(32) ) _54420_ ( .A(29), .B(_29258_), .S(_05690_), .Y({ _29259_[31:5], cparam_max_pool_serial_18_max_col_count }) );
  \$mux  #( .WIDTH(32) ) _54421_ ( .A(64), .B(128), .S(_05745_), .Y(_29262_) );
  \$mux  #( .WIDTH(32) ) _54422_ ( .A(32), .B(_29262_), .S(_05690_), .Y({ _29263_[31:8], cparam_max_pool_serial_18_inc_act_laddr }) );
  \$mux  #( .WIDTH(32) ) _54423_ ( .A(32), .B(64), .S(_05745_), .Y(_29260_) );
  \$mux  #( .WIDTH(32) ) _54424_ ( .A(16), .B(_29260_), .S(_05690_), .Y({ _29261_[31:7], cparam_max_pool_serial_18_inc_out_laddr }) );
  \$mux  #( .WIDTH(32) ) _54425_ ( .A(10), .B(13), .S(_05746_), .Y(_29266_) );
  \$mux  #( .WIDTH(32) ) _54426_ ( .A(12), .B(_29266_), .S(_05691_), .Y({ _29267_[31:4], cparam_matmul_29_cshamt_out_value }) );
  \$mux  #( .WIDTH(32) ) _54427_ ( .A(112), .B(0), .S(_05746_), .Y(_29270_) );
  \$mux  #( .WIDTH(32) ) _54428_ ( .A(252), .B(_29270_), .S(_05691_), .Y({ _29271_[31:8], cparam_matmul_29_max_och_count }) );
  \$mux  #( .WIDTH(32) ) _54429_ ( .A(16), .B(32), .S(_05746_), .Y(_29272_) );
  \$mux  #( .WIDTH(32) ) _54430_ ( .A(4), .B(_29272_), .S(_05691_), .Y({ _29273_[31:6], cparam_matmul_29_och_count_step }) );
  \$mux  #( .WIDTH(32) ) _54431_ ( .A(2048), .B(640), .S(_05746_), .Y(_29276_) );
  \$mux  #( .WIDTH(32) ) _54432_ ( .A(2048), .B(_29276_), .S(_05691_), .Y({ _29277_[31:12], cparam_matmul_29_filter_base_step }) );
  \$mux  #( .WIDTH(32) ) _54433_ ( .A(_24399_), .B(_28870_), .S(_06152_), .Y(_29280_) );
  \$mux  #( .WIDTH(32) ) _54434_ ( .A(4096), .B(1280), .S(_05746_), .Y(_29278_) );
  \$mux  #( .WIDTH(32) ) _54435_ ( .A(4096), .B(_29278_), .S(_05691_), .Y({ _29279_[31:13], cparam_matmul_29_filter_read_size }) );
  \$mux  #( .WIDTH(9) ) _54436_ ( .A({ __delay_data_1413[7], __delay_data_1413 }), .B(9'h180), .S(_pointer_data_784), .Y(_29281_) );
  \$mux  #( .WIDTH(32) ) _54437_ ( .A(128), .B(12), .S(_05746_), .Y(_29282_) );
  \$mux  #( .WIDTH(32) ) _54438_ ( .A(256), .B(_29282_), .S(_05691_), .Y({ _29283_[31:9], cparam_matmul_29_out_bat_step }) );
  \$mux  #( .WIDTH(32) ) _54439_ ( .A(16), .B(10), .S(_05746_), .Y(_29284_) );
  \$mux  #( .WIDTH(32) ) _54440_ ( .A(4), .B(_29284_), .S(_05691_), .Y({ _29285_[31:5], cparam_matmul_29_out_och_step }) );
  \$mux  #( .WIDTH(32) ) _54441_ ( .A(0), .B(1), .S(_05746_), .Y(_29268_) );
  \$mux  #( .WIDTH(32) ) _54442_ ( .A(0), .B(_29268_), .S(_05691_), .Y({ _29269_[31:1], cparam_matmul_29_keep_filter }) );
  \$mux  #( .WIDTH(32) ) _54443_ ( .A(16), .B(12), .S(_05746_), .Y(_29286_) );
  \$mux  #( .WIDTH(32) ) _54444_ ( .A(4), .B(_29286_), .S(_05691_), .Y({ _29287_[31:5], cparam_matmul_29_out_write_size }) );
  \$mux  #( .WIDTH(32) ) _54445_ ( .A(256), .B(128), .S(_05746_), .Y(_29274_) );
  \$mux  #( .WIDTH(32) ) _54446_ ( .A(1024), .B(_29274_), .S(_05691_), .Y({ _29275_[31:11], cparam_matmul_29_act_bat_step }) );
  \$mux  #( .WIDTH(32) ) _54447_ ( .A(128), .B(10), .S(_05746_), .Y(_29264_) );
  \$mux  #( .WIDTH(32) ) _54448_ ( .A(256), .B(_29264_), .S(_05691_), .Y({ _29265_[31:9], cparam_matmul_29_bias_num }) );
  \$mux  #( .WIDTH(8) ) _54449_ ( .A(8'h00), .B(__delay_data_1417), .S(_eq_data_851), .Y(_29288_) );
  \$mux  #( .WIDTH(8) ) _54450_ ( .A(8'h00), .B(_cond_data_853), .S(__delay_data_1418), .Y(_29289_) );
  \$mux  #( .WIDTH(8) ) _54451_ ( .A(_cond_data_857), .B(8'h00), .S(__delay_data_1421), .Y(_29290_) );
  \$mux  #( .WIDTH(8) ) _54452_ ( .A(8'h00), .B(__delay_data_1528), .S(_greaterthan_data_888), .Y(_29230_) );
  \$mux  #( .WIDTH(8) ) _54453_ ( .A(__delay_data_1564), .B(_cond_data_890), .S(__delay_data_1563), .Y(_29291_) );
  \$mux  #( .WIDTH(8) ) _54454_ ( .A(_cond_data_893), .B(__delay_data_1601), .S(__delay_data_1600), .Y(_29292_) );
  \$mux  #( .WIDTH(32) ) _54455_ ( .A(0), .B(matmul_29_och_count_buf), .S(_05905_), .Y(_29293_) );
  \$mux  #( .WIDTH(32) ) _54456_ ( .A(0), .B(1), .S(_05905_), .Y(_29294_) );
  \$mux  #( .WIDTH(32) ) _54457_ ( .A(1), .B(0), .S(_05723_), .Y({ _24124_, _24123_, _24121_, _24120_, _24119_, _24118_, _24117_, _24116_, _24115_, _24114_, _24113_, _24112_, _24110_, _24109_, _24108_, _24107_, _24106_, _24105_, _24104_, _24103_, _24102_, _24101_, _24131_, _24130_, _24129_, _24128_, _24127_, _24126_, _24125_, _24122_, _24111_, _24100_ }) );
  \$mux  #( .WIDTH(32) ) _54458_ ( .A(1), .B(0), .S(_05906_), .Y(_29295_) );
  \$mux  #( .WIDTH(32) ) _54459_ ( .A(0), .B(_29295_), .S(_05723_), .Y({ _24156_, _24155_, _24153_, _24152_, _24151_, _24150_, _24149_, _24148_, _24147_, _24146_, _24145_, _24144_, _24142_, _24141_, _24140_, _24139_, _24138_, _24137_, _24136_, _24135_, _24134_, _24133_, _24163_, _24162_, _24161_, _24160_, _24159_, _24158_, _24157_, _24154_, _24143_, _24132_ }) );
  \$mux  #( .WIDTH(32) ) _54460_ ( .A(1), .B(0), .S(_05907_), .Y(_29296_) );
  \$mux  #( .WIDTH(32) ) _54461_ ( .A(0), .B(_29296_), .S(_05906_), .Y(_29297_) );
  \$mux  #( .WIDTH(32) ) _54462_ ( .A(0), .B(_29297_), .S(_05723_), .Y({ _24188_, _24187_, _24185_, _24184_, _24183_, _24182_, _24181_, _24180_, _24179_, _24178_, _24177_, _24176_, _24174_, _24173_, _24172_, _24171_, _24170_, _24169_, _24168_, _24167_, _24166_, _24165_, _24195_, _24194_, _24193_, _24192_, _24191_, _24190_, _24189_, _24186_, _24175_, _24164_ }) );
  \$mux  #( .WIDTH(32) ) _54463_ ( .A(_24558_), .B(0), .S(_05846_), .Y(_29298_) );
  \$mux  #( .WIDTH(32) ) _54464_ ( .A(_24557_), .B(_29298_), .S(_05845_), .Y(_29299_) );
  \$mux  #( .WIDTH(32) ) _54465_ ( .A(_24555_), .B(_29299_), .S(_05713_), .Y(conv2d_16_mux_act_gaddr_0) );
  \$mux  #( .WIDTH(32) ) _54466_ ( .A(_24557_), .B(0), .S(_05846_), .Y(_29300_) );
  \$mux  #( .WIDTH(32) ) _54467_ ( .A(_24555_), .B(_29300_), .S(_05845_), .Y(_29301_) );
  \$mux  #( .WIDTH(32) ) _54468_ ( .A(_24558_), .B(_29301_), .S(_05713_), .Y(conv2d_16_mux_act_gaddr_1) );
  \$mux  #( .WIDTH(32) ) _54469_ ( .A(_24555_), .B(0), .S(_05846_), .Y(_29302_) );
  \$mux  #( .WIDTH(32) ) _54470_ ( .A(_24558_), .B(_29302_), .S(_05845_), .Y(_29303_) );
  \$mux  #( .WIDTH(32) ) _54471_ ( .A(_24557_), .B(_29303_), .S(_05713_), .Y(conv2d_16_mux_act_gaddr_2) );
  \$mux  #( .WIDTH(1) ) _54472_ ( .A(conv2d_16_dma_pad_mask_1), .B(1'h0), .S(_05846_), .Y(_29304_) );
  \$mux  #( .WIDTH(1) ) _54473_ ( .A(conv2d_16_dma_pad_mask_2), .B(_29304_), .S(_05845_), .Y(_29305_) );
  \$mux  #( .WIDTH(1) ) _54474_ ( .A(conv2d_16_dma_pad_mask_0), .B(_29305_), .S(_05713_), .Y(conv2d_16_mux_dma_pad_mask_0) );
  \$mux  #( .WIDTH(1) ) _54475_ ( .A(conv2d_16_dma_pad_mask_2), .B(1'h0), .S(_05846_), .Y(_29306_) );
  \$mux  #( .WIDTH(1) ) _54476_ ( .A(conv2d_16_dma_pad_mask_0), .B(_29306_), .S(_05845_), .Y(_29307_) );
  \$mux  #( .WIDTH(1) ) _54477_ ( .A(conv2d_16_dma_pad_mask_1), .B(_29307_), .S(_05713_), .Y(conv2d_16_mux_dma_pad_mask_1) );
  \$mux  #( .WIDTH(1) ) _54478_ ( .A(conv2d_16_dma_pad_mask_0), .B(1'h0), .S(_05846_), .Y(_29308_) );
  \$mux  #( .WIDTH(1) ) _54479_ ( .A(conv2d_16_dma_pad_mask_1), .B(_29308_), .S(_05845_), .Y(_29309_) );
  \$mux  #( .WIDTH(1) ) _54480_ ( .A(conv2d_16_dma_pad_mask_2), .B(_29309_), .S(_05713_), .Y(conv2d_16_mux_dma_pad_mask_2) );
  \$mux  #( .WIDTH(1) ) _54481_ ( .A(conv2d_16_dma_flag_1), .B(1'h0), .S(_05748_), .Y(_29310_) );
  \$mux  #( .WIDTH(1) ) _54482_ ( .A(conv2d_16_dma_flag_2), .B(_29310_), .S(_05747_), .Y(_29311_) );
  \$mux  #( .WIDTH(1) ) _54483_ ( .A(conv2d_16_dma_flag_0), .B(_29311_), .S(_05692_), .Y(conv2d_16_mux_dma_flag_0) );
  \$mux  #( .WIDTH(1) ) _54484_ ( .A(conv2d_16_dma_flag_2), .B(1'h0), .S(_05748_), .Y(_29312_) );
  \$mux  #( .WIDTH(1) ) _54485_ ( .A(conv2d_16_dma_flag_0), .B(_29312_), .S(_05747_), .Y(_29313_) );
  \$mux  #( .WIDTH(1) ) _54486_ ( .A(conv2d_16_dma_flag_1), .B(_29313_), .S(_05692_), .Y(conv2d_16_mux_dma_flag_1) );
  \$mux  #( .WIDTH(1) ) _54487_ ( .A(conv2d_16_dma_flag_0), .B(1'h0), .S(_05748_), .Y(_29314_) );
  \$mux  #( .WIDTH(1) ) _54488_ ( .A(conv2d_16_dma_flag_1), .B(_29314_), .S(_05747_), .Y(_29315_) );
  \$mux  #( .WIDTH(1) ) _54489_ ( .A(conv2d_16_dma_flag_2), .B(_29315_), .S(_05692_), .Y(conv2d_16_mux_dma_flag_2) );
  \$mux  #( .WIDTH(32) ) _54490_ ( .A({ 24'h000000, ram_w8_l2048_id1_3_0_rdata }), .B(0), .S(_05751_), .Y(_29316_) );
  \$mux  #( .WIDTH(32) ) _54491_ ( .A({ 24'h000000, ram_w8_l2048_id1_2_0_rdata }), .B(_29316_), .S(_05750_), .Y(_29317_) );
  \$mux  #( .WIDTH(32) ) _54492_ ( .A({ 24'h000000, ram_w8_l2048_id1_1_0_rdata }), .B(_29317_), .S(_05749_), .Y(_29318_) );
  \$mux  #( .WIDTH(32) ) _54493_ ( .A({ 24'h000000, ram_w8_l2048_id1_0_0_rdata }), .B(_29318_), .S(_05693_), .Y({ _29319_[31:8], _tmp_469 }) );
  \$mux  #( .WIDTH(32) ) _54494_ ( .A({ _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469[7], _tmp_469 }), .B(0), .S(_05891_), .Y({ _29320_[31:8], _stream_conv2d_16_source_6_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54495_ ( .A({ 24'h000000, ram_w8_l2048_id0_3_0_rdata }), .B(0), .S(_05754_), .Y(_29321_) );
  \$mux  #( .WIDTH(32) ) _54496_ ( .A({ 24'h000000, ram_w8_l2048_id0_2_0_rdata }), .B(_29321_), .S(_05753_), .Y(_29322_) );
  \$mux  #( .WIDTH(32) ) _54497_ ( .A({ 24'h000000, ram_w8_l2048_id0_1_0_rdata }), .B(_29322_), .S(_05752_), .Y(_29323_) );
  \$mux  #( .WIDTH(32) ) _54498_ ( .A({ 24'h000000, ram_w8_l2048_id0_0_0_rdata }), .B(_29323_), .S(_05694_), .Y({ _29324_[31:8], _tmp_480 }) );
  \$mux  #( .WIDTH(32) ) _54499_ ( .A({ _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480[7], _tmp_480 }), .B(0), .S(_05889_), .Y({ _29325_[31:8], _stream_conv2d_16_source_8_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54500_ ( .A({ 24'h000000, ram_w8_l2048_id2_3_0_rdata }), .B(0), .S(_05757_), .Y(_29326_) );
  \$mux  #( .WIDTH(32) ) _54501_ ( .A({ 24'h000000, ram_w8_l2048_id2_2_0_rdata }), .B(_29326_), .S(_05756_), .Y(_29327_) );
  \$mux  #( .WIDTH(32) ) _54502_ ( .A({ 24'h000000, ram_w8_l2048_id2_1_0_rdata }), .B(_29327_), .S(_05755_), .Y(_29328_) );
  \$mux  #( .WIDTH(32) ) _54503_ ( .A({ 24'h000000, ram_w8_l2048_id2_0_0_rdata }), .B(_29328_), .S(_05695_), .Y({ _29329_[31:8], _tmp_500 }) );
  \$mux  #( .WIDTH(32) ) _54504_ ( .A({ _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500[7], _tmp_500 }), .B(0), .S(_05893_), .Y({ _29330_[31:8], _stream_conv2d_16_source_19_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54505_ ( .A({ 24'h000000, ram_w8_l2048_id3_3_0_rdata }), .B(0), .S(_05760_), .Y(_29331_) );
  \$mux  #( .WIDTH(32) ) _54506_ ( .A({ 24'h000000, ram_w8_l2048_id3_2_0_rdata }), .B(_29331_), .S(_05759_), .Y(_29332_) );
  \$mux  #( .WIDTH(32) ) _54507_ ( .A({ 24'h000000, ram_w8_l2048_id3_1_0_rdata }), .B(_29332_), .S(_05758_), .Y(_29333_) );
  \$mux  #( .WIDTH(32) ) _54508_ ( .A({ 24'h000000, ram_w8_l2048_id3_0_0_rdata }), .B(_29333_), .S(_05696_), .Y({ _29334_[31:8], _tmp_510 }) );
  \$mux  #( .WIDTH(32) ) _54509_ ( .A({ _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510[7], _tmp_510 }), .B(0), .S(_05895_), .Y({ _29335_[31:8], _stream_conv2d_16_source_20_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54510_ ( .A({ 24'h000000, ram_w8_l2048_id4_3_0_rdata }), .B(0), .S(_05763_), .Y(_29336_) );
  \$mux  #( .WIDTH(32) ) _54511_ ( .A({ 24'h000000, ram_w8_l2048_id4_2_0_rdata }), .B(_29336_), .S(_05762_), .Y(_29337_) );
  \$mux  #( .WIDTH(32) ) _54512_ ( .A({ 24'h000000, ram_w8_l2048_id4_1_0_rdata }), .B(_29337_), .S(_05761_), .Y(_29338_) );
  \$mux  #( .WIDTH(32) ) _54513_ ( .A({ 24'h000000, ram_w8_l2048_id4_0_0_rdata }), .B(_29338_), .S(_05697_), .Y({ _29339_[31:8], _tmp_520 }) );
  \$mux  #( .WIDTH(32) ) _54514_ ( .A({ _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520[7], _tmp_520 }), .B(0), .S(_05897_), .Y({ _29340_[31:8], _stream_conv2d_16_source_21_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54515_ ( .A({ 24'h000000, ram_w8_l2048_id5_3_0_rdata }), .B(0), .S(_05766_), .Y(_29341_) );
  \$mux  #( .WIDTH(32) ) _54516_ ( .A({ 24'h000000, ram_w8_l2048_id5_2_0_rdata }), .B(_29341_), .S(_05765_), .Y(_29342_) );
  \$mux  #( .WIDTH(32) ) _54517_ ( .A({ 24'h000000, ram_w8_l2048_id5_1_0_rdata }), .B(_29342_), .S(_05764_), .Y(_29343_) );
  \$mux  #( .WIDTH(32) ) _54518_ ( .A({ 24'h000000, ram_w8_l2048_id5_0_0_rdata }), .B(_29343_), .S(_05698_), .Y({ _29344_[31:8], _tmp_530 }) );
  \$mux  #( .WIDTH(32) ) _54519_ ( .A({ _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530[7], _tmp_530 }), .B(0), .S(_05898_), .Y({ _29345_[31:8], _stream_conv2d_16_source_22_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54520_ ( .A({ 24'h000000, ram_w8_l2048_id6_3_0_rdata }), .B(0), .S(_05769_), .Y(_29346_) );
  \$mux  #( .WIDTH(32) ) _54521_ ( .A({ 24'h000000, ram_w8_l2048_id6_2_0_rdata }), .B(_29346_), .S(_05768_), .Y(_29347_) );
  \$mux  #( .WIDTH(32) ) _54522_ ( .A({ 24'h000000, ram_w8_l2048_id6_1_0_rdata }), .B(_29347_), .S(_05767_), .Y(_29348_) );
  \$mux  #( .WIDTH(32) ) _54523_ ( .A({ 24'h000000, ram_w8_l2048_id6_0_0_rdata }), .B(_29348_), .S(_05699_), .Y({ _29349_[31:8], _tmp_540 }) );
  \$mux  #( .WIDTH(32) ) _54524_ ( .A({ _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540[7], _tmp_540 }), .B(0), .S(_05899_), .Y({ _29350_[31:8], _stream_conv2d_16_source_23_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54525_ ( .A({ 24'h000000, ram_w8_l2048_id7_3_0_rdata }), .B(0), .S(_05772_), .Y(_29351_) );
  \$mux  #( .WIDTH(32) ) _54526_ ( .A({ 24'h000000, ram_w8_l2048_id7_2_0_rdata }), .B(_29351_), .S(_05771_), .Y(_29352_) );
  \$mux  #( .WIDTH(32) ) _54527_ ( .A({ 24'h000000, ram_w8_l2048_id7_1_0_rdata }), .B(_29352_), .S(_05770_), .Y(_29353_) );
  \$mux  #( .WIDTH(32) ) _54528_ ( .A({ 24'h000000, ram_w8_l2048_id7_0_0_rdata }), .B(_29353_), .S(_05700_), .Y({ _29354_[31:8], _tmp_550 }) );
  \$mux  #( .WIDTH(32) ) _54529_ ( .A({ _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550[7], _tmp_550 }), .B(0), .S(_05900_), .Y({ _29355_[31:8], _stream_conv2d_16_source_24_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54530_ ( .A({ 24'h000000, ram_w8_l2048_id8_3_0_rdata }), .B(0), .S(_05775_), .Y(_29356_) );
  \$mux  #( .WIDTH(32) ) _54531_ ( .A({ 24'h000000, ram_w8_l2048_id8_2_0_rdata }), .B(_29356_), .S(_05774_), .Y(_29357_) );
  \$mux  #( .WIDTH(32) ) _54532_ ( .A({ 24'h000000, ram_w8_l2048_id8_1_0_rdata }), .B(_29357_), .S(_05773_), .Y(_29358_) );
  \$mux  #( .WIDTH(32) ) _54533_ ( .A({ 24'h000000, ram_w8_l2048_id8_0_0_rdata }), .B(_29358_), .S(_05701_), .Y({ _29359_[31:8], _tmp_560 }) );
  \$mux  #( .WIDTH(32) ) _54534_ ( .A({ _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560[7], _tmp_560 }), .B(0), .S(_05901_), .Y({ _29360_[31:8], _stream_conv2d_16_source_25_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54535_ ( .A({ 24'h000000, ram_w8_l2048_id9_3_0_rdata }), .B(0), .S(_05778_), .Y(_29361_) );
  \$mux  #( .WIDTH(32) ) _54536_ ( .A({ 24'h000000, ram_w8_l2048_id9_2_0_rdata }), .B(_29361_), .S(_05777_), .Y(_29362_) );
  \$mux  #( .WIDTH(32) ) _54537_ ( .A({ 24'h000000, ram_w8_l2048_id9_1_0_rdata }), .B(_29362_), .S(_05776_), .Y(_29363_) );
  \$mux  #( .WIDTH(32) ) _54538_ ( .A({ 24'h000000, ram_w8_l2048_id9_0_0_rdata }), .B(_29363_), .S(_05702_), .Y({ _29364_[31:8], _tmp_570 }) );
  \$mux  #( .WIDTH(32) ) _54539_ ( .A({ _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570[7], _tmp_570 }), .B(0), .S(_05902_), .Y({ _29365_[31:8], _stream_conv2d_16_source_26_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54540_ ( .A({ 24'h000000, ram_w8_l2048_id10_3_0_rdata }), .B(0), .S(_05781_), .Y(_29366_) );
  \$mux  #( .WIDTH(32) ) _54541_ ( .A({ 24'h000000, ram_w8_l2048_id10_2_0_rdata }), .B(_29366_), .S(_05780_), .Y(_29367_) );
  \$mux  #( .WIDTH(32) ) _54542_ ( .A({ 24'h000000, ram_w8_l2048_id10_1_0_rdata }), .B(_29367_), .S(_05779_), .Y(_29368_) );
  \$mux  #( .WIDTH(32) ) _54543_ ( .A({ 24'h000000, ram_w8_l2048_id10_0_0_rdata }), .B(_29368_), .S(_05703_), .Y({ _29369_[31:8], _tmp_580 }) );
  \$mux  #( .WIDTH(32) ) _54544_ ( .A({ _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580[7], _tmp_580 }), .B(0), .S(_05903_), .Y({ _29370_[31:8], _stream_conv2d_16_source_27_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54545_ ( .A({ 28'h0000000, ram_w4_l8192_id0_7_0_rdata }), .B(0), .S(_05788_), .Y(_29371_) );
  \$mux  #( .WIDTH(32) ) _54546_ ( .A({ 28'h0000000, ram_w4_l8192_id0_6_0_rdata }), .B(_29371_), .S(_05787_), .Y(_29372_) );
  \$mux  #( .WIDTH(32) ) _54547_ ( .A({ 28'h0000000, ram_w4_l8192_id0_5_0_rdata }), .B(_29372_), .S(_05786_), .Y(_29373_) );
  \$mux  #( .WIDTH(32) ) _54548_ ( .A({ 28'h0000000, ram_w4_l8192_id0_4_0_rdata }), .B(_29373_), .S(_05785_), .Y(_29374_) );
  \$mux  #( .WIDTH(32) ) _54549_ ( .A({ 28'h0000000, ram_w4_l8192_id0_3_0_rdata }), .B(_29374_), .S(_05784_), .Y(_29375_) );
  \$mux  #( .WIDTH(32) ) _54550_ ( .A({ 28'h0000000, ram_w4_l8192_id0_2_0_rdata }), .B(_29375_), .S(_05783_), .Y(_29376_) );
  \$mux  #( .WIDTH(32) ) _54551_ ( .A({ 28'h0000000, ram_w4_l8192_id0_1_0_rdata }), .B(_29376_), .S(_05782_), .Y(_29377_) );
  \$mux  #( .WIDTH(32) ) _54552_ ( .A({ 28'h0000000, ram_w4_l8192_id0_0_0_rdata }), .B(_29377_), .S(_05704_), .Y({ _29378_[31:4], _tmp_594 }) );
  \$mux  #( .WIDTH(32) ) _54553_ ( .A({ _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594[3], _tmp_594 }), .B(0), .S(_05879_), .Y({ _29379_[31:4], _stream_conv2d_16_source_28_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54554_ ( .A({ 28'h0000000, ram_w4_l8192_id1_7_0_rdata }), .B(0), .S(_05795_), .Y(_29380_) );
  \$mux  #( .WIDTH(32) ) _54555_ ( .A({ 28'h0000000, ram_w4_l8192_id1_6_0_rdata }), .B(_29380_), .S(_05794_), .Y(_29381_) );
  \$mux  #( .WIDTH(32) ) _54556_ ( .A({ 28'h0000000, ram_w4_l8192_id1_5_0_rdata }), .B(_29381_), .S(_05793_), .Y(_29382_) );
  \$mux  #( .WIDTH(32) ) _54557_ ( .A({ 28'h0000000, ram_w4_l8192_id1_4_0_rdata }), .B(_29382_), .S(_05792_), .Y(_29383_) );
  \$mux  #( .WIDTH(32) ) _54558_ ( .A({ 28'h0000000, ram_w4_l8192_id1_3_0_rdata }), .B(_29383_), .S(_05791_), .Y(_29384_) );
  \$mux  #( .WIDTH(32) ) _54559_ ( .A({ 28'h0000000, ram_w4_l8192_id1_2_0_rdata }), .B(_29384_), .S(_05790_), .Y(_29385_) );
  \$mux  #( .WIDTH(32) ) _54560_ ( .A({ 28'h0000000, ram_w4_l8192_id1_1_0_rdata }), .B(_29385_), .S(_05789_), .Y(_29386_) );
  \$mux  #( .WIDTH(32) ) _54561_ ( .A({ 28'h0000000, ram_w4_l8192_id1_0_0_rdata }), .B(_29386_), .S(_05705_), .Y({ _29387_[31:4], _tmp_608 }) );
  \$mux  #( .WIDTH(32) ) _54562_ ( .A({ _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608[3], _tmp_608 }), .B(0), .S(_05881_), .Y({ _29388_[31:4], _stream_conv2d_16_source_29_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54563_ ( .A({ 28'h0000000, ram_w4_l8192_id2_7_0_rdata }), .B(0), .S(_05802_), .Y(_29389_) );
  \$mux  #( .WIDTH(32) ) _54564_ ( .A({ 28'h0000000, ram_w4_l8192_id2_6_0_rdata }), .B(_29389_), .S(_05801_), .Y(_29390_) );
  \$mux  #( .WIDTH(32) ) _54565_ ( .A({ 28'h0000000, ram_w4_l8192_id2_5_0_rdata }), .B(_29390_), .S(_05800_), .Y(_29391_) );
  \$mux  #( .WIDTH(32) ) _54566_ ( .A({ 28'h0000000, ram_w4_l8192_id2_4_0_rdata }), .B(_29391_), .S(_05799_), .Y(_29392_) );
  \$mux  #( .WIDTH(32) ) _54567_ ( .A({ 28'h0000000, ram_w4_l8192_id2_3_0_rdata }), .B(_29392_), .S(_05798_), .Y(_29393_) );
  \$mux  #( .WIDTH(32) ) _54568_ ( .A({ 28'h0000000, ram_w4_l8192_id2_2_0_rdata }), .B(_29393_), .S(_05797_), .Y(_29394_) );
  \$mux  #( .WIDTH(32) ) _54569_ ( .A({ 28'h0000000, ram_w4_l8192_id2_1_0_rdata }), .B(_29394_), .S(_05796_), .Y(_29395_) );
  \$mux  #( .WIDTH(32) ) _54570_ ( .A({ 28'h0000000, ram_w4_l8192_id2_0_0_rdata }), .B(_29395_), .S(_05706_), .Y({ _29396_[31:4], _tmp_622 }) );
  \$mux  #( .WIDTH(32) ) _54571_ ( .A({ _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622[3], _tmp_622 }), .B(0), .S(_05882_), .Y({ _29397_[31:4], _stream_conv2d_16_source_30_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54572_ ( .A({ 28'h0000000, ram_w4_l8192_id3_7_0_rdata }), .B(0), .S(_05809_), .Y(_29398_) );
  \$mux  #( .WIDTH(32) ) _54573_ ( .A({ 28'h0000000, ram_w4_l8192_id3_6_0_rdata }), .B(_29398_), .S(_05808_), .Y(_29399_) );
  \$mux  #( .WIDTH(32) ) _54574_ ( .A({ 28'h0000000, ram_w4_l8192_id3_5_0_rdata }), .B(_29399_), .S(_05807_), .Y(_29400_) );
  \$mux  #( .WIDTH(32) ) _54575_ ( .A({ 28'h0000000, ram_w4_l8192_id3_4_0_rdata }), .B(_29400_), .S(_05806_), .Y(_29401_) );
  \$mux  #( .WIDTH(32) ) _54576_ ( .A({ 28'h0000000, ram_w4_l8192_id3_3_0_rdata }), .B(_29401_), .S(_05805_), .Y(_29402_) );
  \$mux  #( .WIDTH(32) ) _54577_ ( .A({ 28'h0000000, ram_w4_l8192_id3_2_0_rdata }), .B(_29402_), .S(_05804_), .Y(_29403_) );
  \$mux  #( .WIDTH(32) ) _54578_ ( .A({ 28'h0000000, ram_w4_l8192_id3_1_0_rdata }), .B(_29403_), .S(_05803_), .Y(_29404_) );
  \$mux  #( .WIDTH(32) ) _54579_ ( .A({ 28'h0000000, ram_w4_l8192_id3_0_0_rdata }), .B(_29404_), .S(_05707_), .Y({ _29405_[31:4], _tmp_636 }) );
  \$mux  #( .WIDTH(32) ) _54580_ ( .A({ _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636[3], _tmp_636 }), .B(0), .S(_05883_), .Y({ _29406_[31:4], _stream_conv2d_16_source_31_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54581_ ( .A({ 28'h0000000, ram_w4_l8192_id4_7_0_rdata }), .B(0), .S(_05816_), .Y(_29407_) );
  \$mux  #( .WIDTH(32) ) _54582_ ( .A({ 28'h0000000, ram_w4_l8192_id4_6_0_rdata }), .B(_29407_), .S(_05815_), .Y(_29408_) );
  \$mux  #( .WIDTH(32) ) _54583_ ( .A({ 28'h0000000, ram_w4_l8192_id4_5_0_rdata }), .B(_29408_), .S(_05814_), .Y(_29409_) );
  \$mux  #( .WIDTH(32) ) _54584_ ( .A({ 28'h0000000, ram_w4_l8192_id4_4_0_rdata }), .B(_29409_), .S(_05813_), .Y(_29410_) );
  \$mux  #( .WIDTH(32) ) _54585_ ( .A({ 28'h0000000, ram_w4_l8192_id4_3_0_rdata }), .B(_29410_), .S(_05812_), .Y(_29411_) );
  \$mux  #( .WIDTH(32) ) _54586_ ( .A({ 28'h0000000, ram_w4_l8192_id4_2_0_rdata }), .B(_29411_), .S(_05811_), .Y(_29412_) );
  \$mux  #( .WIDTH(32) ) _54587_ ( .A({ 28'h0000000, ram_w4_l8192_id4_1_0_rdata }), .B(_29412_), .S(_05810_), .Y(_29413_) );
  \$mux  #( .WIDTH(32) ) _54588_ ( .A({ 28'h0000000, ram_w4_l8192_id4_0_0_rdata }), .B(_29413_), .S(_05708_), .Y({ _29414_[31:4], _tmp_650 }) );
  \$mux  #( .WIDTH(32) ) _54589_ ( .A({ _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650[3], _tmp_650 }), .B(0), .S(_05884_), .Y({ _29415_[31:4], _stream_conv2d_16_source_32_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54590_ ( .A({ 28'h0000000, ram_w4_l8192_id5_7_0_rdata }), .B(0), .S(_05823_), .Y(_29416_) );
  \$mux  #( .WIDTH(32) ) _54591_ ( .A({ 28'h0000000, ram_w4_l8192_id5_6_0_rdata }), .B(_29416_), .S(_05822_), .Y(_29417_) );
  \$mux  #( .WIDTH(32) ) _54592_ ( .A({ 28'h0000000, ram_w4_l8192_id5_5_0_rdata }), .B(_29417_), .S(_05821_), .Y(_29418_) );
  \$mux  #( .WIDTH(32) ) _54593_ ( .A({ 28'h0000000, ram_w4_l8192_id5_4_0_rdata }), .B(_29418_), .S(_05820_), .Y(_29419_) );
  \$mux  #( .WIDTH(32) ) _54594_ ( .A({ 28'h0000000, ram_w4_l8192_id5_3_0_rdata }), .B(_29419_), .S(_05819_), .Y(_29420_) );
  \$mux  #( .WIDTH(32) ) _54595_ ( .A({ 28'h0000000, ram_w4_l8192_id5_2_0_rdata }), .B(_29420_), .S(_05818_), .Y(_29421_) );
  \$mux  #( .WIDTH(32) ) _54596_ ( .A({ 28'h0000000, ram_w4_l8192_id5_1_0_rdata }), .B(_29421_), .S(_05817_), .Y(_29422_) );
  \$mux  #( .WIDTH(32) ) _54597_ ( .A({ 28'h0000000, ram_w4_l8192_id5_0_0_rdata }), .B(_29422_), .S(_05709_), .Y({ _29423_[31:4], _tmp_664 }) );
  \$mux  #( .WIDTH(32) ) _54598_ ( .A({ _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664[3], _tmp_664 }), .B(0), .S(_05885_), .Y({ _29424_[31:4], _stream_conv2d_16_source_33_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54599_ ( .A({ 28'h0000000, ram_w4_l8192_id6_7_0_rdata }), .B(0), .S(_05830_), .Y(_29425_) );
  \$mux  #( .WIDTH(32) ) _54600_ ( .A({ 28'h0000000, ram_w4_l8192_id6_6_0_rdata }), .B(_29425_), .S(_05829_), .Y(_29426_) );
  \$mux  #( .WIDTH(32) ) _54601_ ( .A({ 28'h0000000, ram_w4_l8192_id6_5_0_rdata }), .B(_29426_), .S(_05828_), .Y(_29427_) );
  \$mux  #( .WIDTH(32) ) _54602_ ( .A({ 28'h0000000, ram_w4_l8192_id6_4_0_rdata }), .B(_29427_), .S(_05827_), .Y(_29428_) );
  \$mux  #( .WIDTH(32) ) _54603_ ( .A({ 28'h0000000, ram_w4_l8192_id6_3_0_rdata }), .B(_29428_), .S(_05826_), .Y(_29429_) );
  \$mux  #( .WIDTH(32) ) _54604_ ( .A({ 28'h0000000, ram_w4_l8192_id6_2_0_rdata }), .B(_29429_), .S(_05825_), .Y(_29430_) );
  \$mux  #( .WIDTH(32) ) _54605_ ( .A({ 28'h0000000, ram_w4_l8192_id6_1_0_rdata }), .B(_29430_), .S(_05824_), .Y(_29431_) );
  \$mux  #( .WIDTH(32) ) _54606_ ( .A({ 28'h0000000, ram_w4_l8192_id6_0_0_rdata }), .B(_29431_), .S(_05710_), .Y({ _29432_[31:4], _tmp_678 }) );
  \$mux  #( .WIDTH(32) ) _54607_ ( .A({ _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678[3], _tmp_678 }), .B(0), .S(_05886_), .Y({ _29433_[31:4], _stream_conv2d_16_source_34_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54608_ ( .A({ 28'h0000000, ram_w4_l8192_id7_7_0_rdata }), .B(0), .S(_05837_), .Y(_29434_) );
  \$mux  #( .WIDTH(32) ) _54609_ ( .A({ 28'h0000000, ram_w4_l8192_id7_6_0_rdata }), .B(_29434_), .S(_05836_), .Y(_29435_) );
  \$mux  #( .WIDTH(32) ) _54610_ ( .A({ 28'h0000000, ram_w4_l8192_id7_5_0_rdata }), .B(_29435_), .S(_05835_), .Y(_29436_) );
  \$mux  #( .WIDTH(32) ) _54611_ ( .A({ 28'h0000000, ram_w4_l8192_id7_4_0_rdata }), .B(_29436_), .S(_05834_), .Y(_29437_) );
  \$mux  #( .WIDTH(32) ) _54612_ ( .A({ 28'h0000000, ram_w4_l8192_id7_3_0_rdata }), .B(_29437_), .S(_05833_), .Y(_29438_) );
  \$mux  #( .WIDTH(32) ) _54613_ ( .A({ 28'h0000000, ram_w4_l8192_id7_2_0_rdata }), .B(_29438_), .S(_05832_), .Y(_29439_) );
  \$mux  #( .WIDTH(32) ) _54614_ ( .A({ 28'h0000000, ram_w4_l8192_id7_1_0_rdata }), .B(_29439_), .S(_05831_), .Y(_29440_) );
  \$mux  #( .WIDTH(32) ) _54615_ ( .A({ 28'h0000000, ram_w4_l8192_id7_0_0_rdata }), .B(_29440_), .S(_05711_), .Y({ _29441_[31:4], _tmp_692 }) );
  \$mux  #( .WIDTH(32) ) _54616_ ( .A({ _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692[3], _tmp_692 }), .B(0), .S(_05887_), .Y({ _29442_[31:4], _stream_conv2d_16_source_35_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54617_ ( .A({ 28'h0000000, ram_w4_l8192_id8_7_0_rdata }), .B(0), .S(_05844_), .Y(_29443_) );
  \$mux  #( .WIDTH(32) ) _54618_ ( .A({ 28'h0000000, ram_w4_l8192_id8_6_0_rdata }), .B(_29443_), .S(_05843_), .Y(_29444_) );
  \$mux  #( .WIDTH(32) ) _54619_ ( .A({ 28'h0000000, ram_w4_l8192_id8_5_0_rdata }), .B(_29444_), .S(_05842_), .Y(_29445_) );
  \$mux  #( .WIDTH(32) ) _54620_ ( .A({ 28'h0000000, ram_w4_l8192_id8_4_0_rdata }), .B(_29445_), .S(_05841_), .Y(_29446_) );
  \$mux  #( .WIDTH(32) ) _54621_ ( .A({ 28'h0000000, ram_w4_l8192_id8_3_0_rdata }), .B(_29446_), .S(_05840_), .Y(_29447_) );
  \$mux  #( .WIDTH(32) ) _54622_ ( .A({ 28'h0000000, ram_w4_l8192_id8_2_0_rdata }), .B(_29447_), .S(_05839_), .Y(_29448_) );
  \$mux  #( .WIDTH(32) ) _54623_ ( .A({ 28'h0000000, ram_w4_l8192_id8_1_0_rdata }), .B(_29448_), .S(_05838_), .Y(_29449_) );
  \$mux  #( .WIDTH(32) ) _54624_ ( .A({ 28'h0000000, ram_w4_l8192_id8_0_0_rdata }), .B(_29449_), .S(_05712_), .Y({ _29450_[31:4], _tmp_706 }) );
  \$mux  #( .WIDTH(32) ) _54625_ ( .A({ _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706[3], _tmp_706 }), .B(0), .S(_05888_), .Y({ _29451_[31:4], _stream_conv2d_16_source_36_source_ram_rdata }) );
  \$mux  #( .WIDTH(32) ) _54626_ ( .A(0), .B(1), .S(_06874_), .Y({ _29452_[31:1], _stream_conv2d_16_start_flag }) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41747_ ( .CLK(CLK), .D(_02715_), .Q(_stream_matmul_29_sink_21_sink_fsm_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41748_ ( .CLK(CLK), .D(_02744_), .Q(_stream_matmul_29_source_20_source_pat_fsm_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41749_ ( .CLK(CLK), .D(_02735_), .Q(_stream_matmul_29_source_19_source_pat_fsm_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41750_ ( .CLK(CLK), .D(_02762_), .Q(_stream_matmul_29_source_8_source_pat_fsm_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41751_ ( .CLK(CLK), .D(_02753_), .Q(_stream_matmul_29_source_6_source_pat_fsm_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41752_ ( .CLK(CLK), .D(_03300_), .Q(matmul_29_next_stream_num_ops) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41753_ ( .CLK(CLK), .D(_03331_), .Q(matmul_29_sync_comp_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41754_ ( .CLK(CLK), .D(_03290_), .Q(matmul_29_col_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) matmul_29_col_select_reg  ( .CLK(CLK), .D(_03291_), .Q(matmul_29_col_select) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41756_ ( .CLK(CLK), .D(_03328_), .Q(matmul_29_stream_act_local_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41757_ ( .CLK(CLK), .D(_03329_), .Q(matmul_29_stream_out_local_col) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41758_ ( .CLK(CLK), .D(_03292_), .Q(matmul_29_comp_fsm) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41759_ ( .CLK(CLK), .D(_03297_), .Q(matmul_29_filter_page_comp_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41760_ ( .CLK(CLK), .D(_03283_), .Q(matmul_29_act_page_comp_offset_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41761_ ( .CLK(CLK), .D(_03312_), .Q(matmul_29_out_page_comp_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41762_ ( .CLK(CLK), .D(_03321_), .Q(matmul_29_row_count_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) matmul_29_row_select_buf_reg  ( .CLK(CLK), .D(_03323_), .Q(matmul_29_row_select_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41764_ ( .CLK(CLK), .D(_03303_), .Q(matmul_29_och_count_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) matmul_29_stream_pad_masks_reg  ( .CLK(CLK), .D(_03330_), .Q(matmul_29_stream_pad_masks) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41766_ ( .CLK(CLK), .D(_03208_), .Q(control_matmul_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41767_ ( .CLK(CLK), .D(_03281_), .Q(matmul_29_act_base_offset_row) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41768_ ( .CLK(CLK), .D(_03280_), .Q(matmul_29_act_base_offset_bat) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41769_ ( .CLK(CLK), .D(_03295_), .Q(matmul_29_filter_base_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41770_ ( .CLK(CLK), .D(_03308_), .Q(matmul_29_out_base_offset_val) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41771_ ( .CLK(CLK), .D(_03305_), .Q(matmul_29_out_base_offset_col) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41772_ ( .CLK(CLK), .D(_03307_), .Q(matmul_29_out_base_offset_row) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41773_ ( .CLK(CLK), .D(_03304_), .Q(matmul_29_out_base_offset_bat) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41774_ ( .CLK(CLK), .D(_03306_), .Q(matmul_29_out_base_offset_och) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) matmul_29_dma_flag_0_reg  ( .CLK(CLK), .D(_03294_), .Q(matmul_29_dma_flag_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41776_ ( .CLK(CLK), .D(_03332_), .Q(matmul_29_sync_out_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41777_ ( .CLK(CLK), .D(_03299_), .Q(matmul_29_next_out_write_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41778_ ( .CLK(CLK), .D(_03320_), .Q(matmul_29_row_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41779_ ( .CLK(CLK), .D(_03289_), .Q(matmul_29_bat_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41780_ ( .CLK(CLK), .D(_03302_), .Q(matmul_29_och_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) matmul_29_row_select_reg  ( .CLK(CLK), .D(_03322_), .Q(matmul_29_row_select) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41782_ ( .CLK(CLK), .D(_03315_), .Q(matmul_29_out_row_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41783_ ( .CLK(CLK), .D(_03314_), .Q(matmul_29_out_ram_select) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41784_ ( .CLK(CLK), .D(_03318_), .Q(matmul_29_prev_row_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41785_ ( .CLK(CLK), .D(_03316_), .Q(matmul_29_prev_bat_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41786_ ( .CLK(CLK), .D(_03317_), .Q(matmul_29_prev_och_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) matmul_29_prev_row_select_reg  ( .CLK(CLK), .D(_03319_), .Q(matmul_29_prev_row_select) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41788_ ( .CLK(CLK), .D(_03282_), .Q(matmul_29_act_page_comp_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41789_ ( .CLK(CLK), .D(_03284_), .Q(matmul_29_act_page_dma_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41790_ ( .CLK(CLK), .D(_03296_), .Q(matmul_29_filter_page_comp_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41791_ ( .CLK(CLK), .D(_03298_), .Q(matmul_29_filter_page_dma_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) matmul_29_out_page_reg  ( .CLK(CLK), .D(_03310_), .Q(matmul_29_out_page) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41793_ ( .CLK(CLK), .D(_03311_), .Q(matmul_29_out_page_comp_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41794_ ( .CLK(CLK), .D(_03313_), .Q(matmul_29_out_page_dma_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41795_ ( .CLK(CLK), .D(_03309_), .Q(matmul_29_out_laddr_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) matmul_29_skip_read_filter_reg  ( .CLK(CLK), .D(_03326_), .Q(matmul_29_skip_read_filter) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) matmul_29_skip_read_act_reg  ( .CLK(CLK), .D(_03325_), .Q(matmul_29_skip_read_act) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) matmul_29_skip_comp_reg  ( .CLK(CLK), .D(_03324_), .Q(matmul_29_skip_comp) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) matmul_29_skip_write_out_reg  ( .CLK(CLK), .D(_03327_), .Q(matmul_29_skip_write_out) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_1121_reg  ( .CLK(CLK), .D(_03194_), .Q(axim_flag_1121) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41801_ ( .CLK(CLK), .D(_01584_), .Q(_d1_control_matmul_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_matmul_29_cond_3_0_1_reg  ( .CLK(CLK), .D(_01574_), .Q(_control_matmul_29_cond_3_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_1132_reg  ( .CLK(CLK), .D(_03195_), .Q(axim_flag_1132) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_matmul_29_cond_8_1_1_reg  ( .CLK(CLK), .D(_01575_), .Q(_control_matmul_29_cond_8_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_1133_reg  ( .CLK(CLK), .D(_03196_), .Q(axim_flag_1133) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_matmul_29_cond_14_2_1_reg  ( .CLK(CLK), .D(_01571_), .Q(_control_matmul_29_cond_14_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_1152_reg  ( .CLK(CLK), .D(_03197_), .Q(axim_flag_1152) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_matmul_29_cond_22_3_1_reg  ( .CLK(CLK), .D(_01572_), .Q(_control_matmul_29_cond_22_3_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_1308_reg  ( .CLK(CLK), .D(_03198_), .Q(axim_flag_1308) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_matmul_29_cond_32_4_1_reg  ( .CLK(CLK), .D(_01573_), .Q(_control_matmul_29_cond_32_4_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41811_ ( .CLK(CLK), .D(_02776_), .Q(_stream_max_pool_serial_18_sink_3_sink_fsm_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41812_ ( .CLK(CLK), .D(_02790_), .Q(_stream_max_pool_serial_18_source_1_source_pat_fsm_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41813_ ( .CLK(CLK), .D(_03341_), .Q(max_pool_serial_18_col_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41814_ ( .CLK(CLK), .D(_03360_), .Q(max_pool_serial_18_stream_act_local) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41815_ ( .CLK(CLK), .D(_03361_), .Q(max_pool_serial_18_stream_out_local) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41816_ ( .CLK(CLK), .D(_03342_), .Q(max_pool_serial_18_comp_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41817_ ( .CLK(CLK), .D(_03343_), .Q(max_pool_serial_18_comp_fsm) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41818_ ( .CLK(CLK), .D(_03337_), .Q(max_pool_serial_18_act_page_comp_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41819_ ( .CLK(CLK), .D(_03351_), .Q(max_pool_serial_18_out_page_comp_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41820_ ( .CLK(CLK), .D(_03356_), .Q(max_pool_serial_18_row_count_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _41821_ ( .CLK(CLK), .D(_03362_), .Q(max_pool_serial_18_stream_pad_masks) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41822_ ( .CLK(CLK), .D(_03209_), .Q(control_max_pool_serial_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41823_ ( .CLK(CLK), .D(_03334_), .Q(max_pool_serial_18_act_base_offset_row) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41824_ ( .CLK(CLK), .D(_03333_), .Q(max_pool_serial_18_act_base_offset_bat) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41825_ ( .CLK(CLK), .D(_03347_), .Q(max_pool_serial_18_out_base_offset_row) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41826_ ( .CLK(CLK), .D(_03346_), .Q(max_pool_serial_18_out_base_offset_bat) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41827_ ( .CLK(CLK), .D(_03355_), .Q(max_pool_serial_18_row_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41828_ ( .CLK(CLK), .D(_03340_), .Q(max_pool_serial_18_bat_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41829_ ( .CLK(CLK), .D(_03354_), .Q(max_pool_serial_18_prev_row_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41830_ ( .CLK(CLK), .D(_03353_), .Q(max_pool_serial_18_prev_bat_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) max_pool_serial_18_act_page_reg  ( .CLK(CLK), .D(_03335_), .Q(max_pool_serial_18_act_page) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41832_ ( .CLK(CLK), .D(_03336_), .Q(max_pool_serial_18_act_page_comp_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41833_ ( .CLK(CLK), .D(_03338_), .Q(max_pool_serial_18_act_page_dma_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) max_pool_serial_18_out_page_reg  ( .CLK(CLK), .D(_03349_), .Q(max_pool_serial_18_out_page) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41835_ ( .CLK(CLK), .D(_03350_), .Q(max_pool_serial_18_out_page_comp_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41836_ ( .CLK(CLK), .D(_03352_), .Q(max_pool_serial_18_out_page_dma_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) max_pool_serial_18_skip_read_act_reg  ( .CLK(CLK), .D(_03358_), .Q(max_pool_serial_18_skip_read_act) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) max_pool_serial_18_skip_comp_reg  ( .CLK(CLK), .D(_03357_), .Q(max_pool_serial_18_skip_comp) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) max_pool_serial_18_skip_write_out_reg  ( .CLK(CLK), .D(_03359_), .Q(max_pool_serial_18_skip_write_out) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41840_ ( .CLK(CLK), .D(_03348_), .Q(max_pool_serial_18_out_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_1022_reg  ( .CLK(CLK), .D(_03191_), .Q(axim_flag_1022) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41842_ ( .CLK(CLK), .D(_01585_), .Q(_d1_control_max_pool_serial_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_max_pool_serial_18_cond_5_0_1_reg  ( .CLK(CLK), .D(_01578_), .Q(_control_max_pool_serial_18_cond_5_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_1023_reg  ( .CLK(CLK), .D(_03192_), .Q(axim_flag_1023) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_max_pool_serial_18_cond_11_1_1_reg  ( .CLK(CLK), .D(_01576_), .Q(_control_max_pool_serial_18_cond_11_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_1071_reg  ( .CLK(CLK), .D(_03193_), .Q(axim_flag_1071) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_max_pool_serial_18_cond_19_2_1_reg  ( .CLK(CLK), .D(_01577_), .Q(_control_max_pool_serial_18_cond_19_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41848_ ( .CLK(CLK), .D(_01791_), .Q(_maxi_write_fsm) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41849_ ( .CLK(CLK), .D(_01789_), .Q(_maxi_write_cur_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _41850_ ( .CLK(CLK), .D(_01790_), .Q(_maxi_write_cur_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _41851_ ( .CLK(CLK), .D(_01797_), .Q(_maxi_write_rest_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_1021_reg  ( .CLK(CLK), .D(_03190_), .Q(axim_flag_1021) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41853_ ( .CLK(CLK), .D(_01582_), .Q(_d1__maxi_write_fsm) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __maxi_write_fsm_cond_4_0_1_reg  ( .CLK(CLK), .D(_00691_), .Q(__maxi_write_fsm_cond_4_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41855_ ( .CLK(CLK), .D(_02505_), .Q(_stream_conv2d_16_sink_37_sink_fsm_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41856_ ( .CLK(CLK), .D(_02678_), .Q(_stream_conv2d_16_source_36_source_pat_fsm_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41857_ ( .CLK(CLK), .D(_01286_), .Q(__tmp_697_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41858_ ( .CLK(CLK), .D(_01287_), .Q(__tmp_697_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41859_ ( .CLK(CLK), .D(_02669_), .Q(_stream_conv2d_16_source_35_source_pat_fsm_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41860_ ( .CLK(CLK), .D(_01283_), .Q(__tmp_683_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41861_ ( .CLK(CLK), .D(_01284_), .Q(__tmp_683_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41862_ ( .CLK(CLK), .D(_02660_), .Q(_stream_conv2d_16_source_34_source_pat_fsm_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41863_ ( .CLK(CLK), .D(_01280_), .Q(__tmp_669_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41864_ ( .CLK(CLK), .D(_01281_), .Q(__tmp_669_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41865_ ( .CLK(CLK), .D(_02651_), .Q(_stream_conv2d_16_source_33_source_pat_fsm_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41866_ ( .CLK(CLK), .D(_01277_), .Q(__tmp_655_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41867_ ( .CLK(CLK), .D(_01278_), .Q(__tmp_655_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41868_ ( .CLK(CLK), .D(_02642_), .Q(_stream_conv2d_16_source_32_source_pat_fsm_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41869_ ( .CLK(CLK), .D(_01274_), .Q(__tmp_641_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41870_ ( .CLK(CLK), .D(_01275_), .Q(__tmp_641_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41871_ ( .CLK(CLK), .D(_02633_), .Q(_stream_conv2d_16_source_31_source_pat_fsm_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41872_ ( .CLK(CLK), .D(_01271_), .Q(__tmp_627_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41873_ ( .CLK(CLK), .D(_01272_), .Q(__tmp_627_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41874_ ( .CLK(CLK), .D(_02624_), .Q(_stream_conv2d_16_source_30_source_pat_fsm_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41875_ ( .CLK(CLK), .D(_01268_), .Q(__tmp_613_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41876_ ( .CLK(CLK), .D(_01269_), .Q(__tmp_613_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41877_ ( .CLK(CLK), .D(_02615_), .Q(_stream_conv2d_16_source_29_source_pat_fsm_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41878_ ( .CLK(CLK), .D(_01265_), .Q(__tmp_599_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41879_ ( .CLK(CLK), .D(_01266_), .Q(__tmp_599_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41880_ ( .CLK(CLK), .D(_02606_), .Q(_stream_conv2d_16_source_28_source_pat_fsm_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41881_ ( .CLK(CLK), .D(_01262_), .Q(__tmp_585_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41882_ ( .CLK(CLK), .D(_01263_), .Q(__tmp_585_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41883_ ( .CLK(CLK), .D(_01148_), .Q(__tmp_1211_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _41884_ ( .CLK(CLK), .D(_01149_), .Q(__tmp_1211_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41885_ ( .CLK(CLK), .D(_02597_), .Q(_stream_conv2d_16_source_27_source_pat_fsm_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41886_ ( .CLK(CLK), .D(_01259_), .Q(__tmp_575_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41887_ ( .CLK(CLK), .D(_01260_), .Q(__tmp_575_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41888_ ( .CLK(CLK), .D(_02588_), .Q(_stream_conv2d_16_source_26_source_pat_fsm_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41889_ ( .CLK(CLK), .D(_01256_), .Q(__tmp_565_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41890_ ( .CLK(CLK), .D(_01257_), .Q(__tmp_565_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41891_ ( .CLK(CLK), .D(_02579_), .Q(_stream_conv2d_16_source_25_source_pat_fsm_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41892_ ( .CLK(CLK), .D(_01253_), .Q(__tmp_555_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41893_ ( .CLK(CLK), .D(_01254_), .Q(__tmp_555_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41894_ ( .CLK(CLK), .D(_02570_), .Q(_stream_conv2d_16_source_24_source_pat_fsm_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41895_ ( .CLK(CLK), .D(_01250_), .Q(__tmp_545_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41896_ ( .CLK(CLK), .D(_01251_), .Q(__tmp_545_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41897_ ( .CLK(CLK), .D(_02561_), .Q(_stream_conv2d_16_source_23_source_pat_fsm_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41898_ ( .CLK(CLK), .D(_01247_), .Q(__tmp_535_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41899_ ( .CLK(CLK), .D(_01248_), .Q(__tmp_535_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41900_ ( .CLK(CLK), .D(_02552_), .Q(_stream_conv2d_16_source_22_source_pat_fsm_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41901_ ( .CLK(CLK), .D(_01244_), .Q(__tmp_525_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41902_ ( .CLK(CLK), .D(_01245_), .Q(__tmp_525_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41903_ ( .CLK(CLK), .D(_02543_), .Q(_stream_conv2d_16_source_21_source_pat_fsm_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41904_ ( .CLK(CLK), .D(_01241_), .Q(__tmp_515_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41905_ ( .CLK(CLK), .D(_01242_), .Q(__tmp_515_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41906_ ( .CLK(CLK), .D(_02534_), .Q(_stream_conv2d_16_source_20_source_pat_fsm_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41907_ ( .CLK(CLK), .D(_01238_), .Q(__tmp_505_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41908_ ( .CLK(CLK), .D(_01239_), .Q(__tmp_505_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41909_ ( .CLK(CLK), .D(_01145_), .Q(__tmp_1201_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41910_ ( .CLK(CLK), .D(_01146_), .Q(__tmp_1201_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41911_ ( .CLK(CLK), .D(_02525_), .Q(_stream_conv2d_16_source_19_source_pat_fsm_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41912_ ( .CLK(CLK), .D(_01235_), .Q(__tmp_495_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41913_ ( .CLK(CLK), .D(_01236_), .Q(__tmp_495_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41914_ ( .CLK(CLK), .D(_01139_), .Q(__tmp_1170_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41915_ ( .CLK(CLK), .D(_01140_), .Q(__tmp_1170_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41916_ ( .CLK(CLK), .D(_02696_), .Q(_stream_conv2d_16_source_8_source_pat_fsm_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41917_ ( .CLK(CLK), .D(_01232_), .Q(__tmp_475_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41918_ ( .CLK(CLK), .D(_01233_), .Q(__tmp_475_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41919_ ( .CLK(CLK), .D(_01142_), .Q(__tmp_1181_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41920_ ( .CLK(CLK), .D(_01143_), .Q(__tmp_1181_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41921_ ( .CLK(CLK), .D(_02687_), .Q(_stream_conv2d_16_source_6_source_pat_fsm_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41922_ ( .CLK(CLK), .D(_01229_), .Q(__tmp_464_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41923_ ( .CLK(CLK), .D(_01230_), .Q(__tmp_464_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41924_ ( .CLK(CLK), .D(_01109_), .Q(__tmp_1027_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41925_ ( .CLK(CLK), .D(_01110_), .Q(__tmp_1027_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41926_ ( .CLK(CLK), .D(_03238_), .Q(conv2d_16_next_stream_num_ops) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41927_ ( .CLK(CLK), .D(_03277_), .Q(conv2d_16_sync_comp_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41928_ ( .CLK(CLK), .D(_03226_), .Q(conv2d_16_col_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41929_ ( .CLK(CLK), .D(_03227_), .Q(conv2d_16_col_select) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41930_ ( .CLK(CLK), .D(_03266_), .Q(conv2d_16_stream_act_local_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41931_ ( .CLK(CLK), .D(_03267_), .Q(conv2d_16_stream_act_local_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41932_ ( .CLK(CLK), .D(_03268_), .Q(conv2d_16_stream_act_local_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41933_ ( .CLK(CLK), .D(_03269_), .Q(conv2d_16_stream_act_local_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41934_ ( .CLK(CLK), .D(_03270_), .Q(conv2d_16_stream_act_local_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41935_ ( .CLK(CLK), .D(_03271_), .Q(conv2d_16_stream_act_local_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41936_ ( .CLK(CLK), .D(_03272_), .Q(conv2d_16_stream_act_local_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41937_ ( .CLK(CLK), .D(_03273_), .Q(conv2d_16_stream_act_local_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41938_ ( .CLK(CLK), .D(_03274_), .Q(conv2d_16_stream_act_local_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41939_ ( .CLK(CLK), .D(_03275_), .Q(conv2d_16_stream_out_local_col) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41940_ ( .CLK(CLK), .D(_03228_), .Q(conv2d_16_comp_fsm) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41941_ ( .CLK(CLK), .D(_03235_), .Q(conv2d_16_filter_page_comp_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41942_ ( .CLK(CLK), .D(_03215_), .Q(conv2d_16_act_page_comp_offset_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41943_ ( .CLK(CLK), .D(_03216_), .Q(conv2d_16_act_page_comp_offset_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41944_ ( .CLK(CLK), .D(_03217_), .Q(conv2d_16_act_page_comp_offset_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41945_ ( .CLK(CLK), .D(_03250_), .Q(conv2d_16_out_page_comp_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41946_ ( .CLK(CLK), .D(_03259_), .Q(conv2d_16_row_count_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _41947_ ( .CLK(CLK), .D(_03261_), .Q(conv2d_16_row_select_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41948_ ( .CLK(CLK), .D(_03241_), .Q(conv2d_16_och_count_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _41949_ ( .CLK(CLK), .D(_03276_), .Q(conv2d_16_stream_pad_masks) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _41950_ ( .CLK(CLK), .D(_03872_), .Q(req_block_size_400) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _41951_ ( .CLK(CLK), .D(_03871_), .Q(req_block_size_343) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _41952_ ( .CLK(CLK), .D(_03869_), .Q(req_block_size_286) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _41953_ ( .CLK(CLK), .D(_03870_), .Q(req_block_size_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41954_ ( .CLK(CLK), .D(_01780_), .Q(_maxi_read_fsm) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41955_ ( .CLK(CLK), .D(_01778_), .Q(_maxi_read_cur_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _41956_ ( .CLK(CLK), .D(_01779_), .Q(_maxi_read_cur_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _41957_ ( .CLK(CLK), .D(_01786_), .Q(_maxi_read_rest_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41958_ ( .CLK(CLK), .D(_03172_), .Q(_wdata_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _wvalid_11_reg  ( .CLK(CLK), .D(_03184_), .Q(_wvalid_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41960_ ( .CLK(CLK), .D(_01581_), .Q(_d1__maxi_read_fsm) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __maxi_read_fsm_cond_3_0_1_reg  ( .CLK(CLK), .D(_00681_), .Q(__maxi_read_fsm_cond_3_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_21_reg  ( .CLK(CLK), .D(_03199_), .Q(axim_flag_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __maxi_read_fsm_cond_4_1_1_reg  ( .CLK(CLK), .D(_00690_), .Q(__maxi_read_fsm_cond_4_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41964_ ( .CLK(CLK), .D(_03176_), .Q(_wdata_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _wvalid_24_reg  ( .CLK(CLK), .D(_03185_), .Q(_wvalid_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __maxi_read_fsm_cond_3_2_1_reg  ( .CLK(CLK), .D(_00682_), .Q(__maxi_read_fsm_cond_3_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41967_ ( .CLK(CLK), .D(_03179_), .Q(_wdata_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _wvalid_37_reg  ( .CLK(CLK), .D(_03188_), .Q(_wvalid_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __maxi_read_fsm_cond_3_3_1_reg  ( .CLK(CLK), .D(_00683_), .Q(__maxi_read_fsm_cond_3_3_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41970_ ( .CLK(CLK), .D(_03177_), .Q(_wdata_289) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _wvalid_290_reg  ( .CLK(CLK), .D(_03186_), .Q(_wvalid_290) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __maxi_read_fsm_cond_3_4_1_reg  ( .CLK(CLK), .D(_00684_), .Q(__maxi_read_fsm_cond_3_4_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41973_ ( .CLK(CLK), .D(_03178_), .Q(_wdata_346) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _wvalid_347_reg  ( .CLK(CLK), .D(_03187_), .Q(_wvalid_347) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __maxi_read_fsm_cond_3_5_1_reg  ( .CLK(CLK), .D(_00685_), .Q(__maxi_read_fsm_cond_3_5_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41976_ ( .CLK(CLK), .D(_03180_), .Q(_wdata_403) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _wvalid_404_reg  ( .CLK(CLK), .D(_03189_), .Q(_wvalid_404) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __maxi_read_fsm_cond_3_6_1_reg  ( .CLK(CLK), .D(_00686_), .Q(__maxi_read_fsm_cond_3_6_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41979_ ( .CLK(CLK), .D(_03173_), .Q(_wdata_1122) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _wvalid_1123_reg  ( .CLK(CLK), .D(_03181_), .Q(_wvalid_1123) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __maxi_read_fsm_cond_3_7_1_reg  ( .CLK(CLK), .D(_00687_), .Q(__maxi_read_fsm_cond_3_7_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41982_ ( .CLK(CLK), .D(_03174_), .Q(_wdata_1134) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _wvalid_1135_reg  ( .CLK(CLK), .D(_03182_), .Q(_wvalid_1135) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __maxi_read_fsm_cond_3_8_1_reg  ( .CLK(CLK), .D(_00688_), .Q(__maxi_read_fsm_cond_3_8_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41985_ ( .CLK(CLK), .D(_03175_), .Q(_wdata_1153) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _wvalid_1154_reg  ( .CLK(CLK), .D(_03183_), .Q(_wvalid_1154) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __maxi_read_fsm_cond_3_9_1_reg  ( .CLK(CLK), .D(_00689_), .Q(__maxi_read_fsm_cond_3_9_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41988_ ( .CLK(CLK), .D(_03207_), .Q(control_conv2d_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41989_ ( .CLK(CLK), .D(_03211_), .Q(conv2d_16_act_base_offset_row) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41990_ ( .CLK(CLK), .D(_03210_), .Q(conv2d_16_act_base_offset_bat) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41991_ ( .CLK(CLK), .D(_03233_), .Q(conv2d_16_filter_base_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41992_ ( .CLK(CLK), .D(_03246_), .Q(conv2d_16_out_base_offset_val) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41993_ ( .CLK(CLK), .D(_03243_), .Q(conv2d_16_out_base_offset_col) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41994_ ( .CLK(CLK), .D(_03245_), .Q(conv2d_16_out_base_offset_row) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41995_ ( .CLK(CLK), .D(_03242_), .Q(conv2d_16_out_base_offset_bat) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _41996_ ( .CLK(CLK), .D(_03244_), .Q(conv2d_16_out_base_offset_och) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) conv2d_16_dma_flag_0_reg  ( .CLK(CLK), .D(_03230_), .Q(conv2d_16_dma_flag_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) conv2d_16_dma_flag_1_reg  ( .CLK(CLK), .D(_03231_), .Q(conv2d_16_dma_flag_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) conv2d_16_dma_flag_2_reg  ( .CLK(CLK), .D(_03232_), .Q(conv2d_16_dma_flag_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42000_ ( .CLK(CLK), .D(_03278_), .Q(conv2d_16_sync_out_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42001_ ( .CLK(CLK), .D(_03237_), .Q(conv2d_16_next_out_write_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42002_ ( .CLK(CLK), .D(_03258_), .Q(conv2d_16_row_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42003_ ( .CLK(CLK), .D(_03225_), .Q(conv2d_16_bat_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42004_ ( .CLK(CLK), .D(_03240_), .Q(conv2d_16_och_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _42005_ ( .CLK(CLK), .D(_03260_), .Q(conv2d_16_row_select) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42006_ ( .CLK(CLK), .D(_03253_), .Q(conv2d_16_out_row_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42007_ ( .CLK(CLK), .D(_03252_), .Q(conv2d_16_out_ram_select) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42008_ ( .CLK(CLK), .D(_03256_), .Q(conv2d_16_prev_row_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42009_ ( .CLK(CLK), .D(_03254_), .Q(conv2d_16_prev_bat_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42010_ ( .CLK(CLK), .D(_03255_), .Q(conv2d_16_prev_och_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _42011_ ( .CLK(CLK), .D(_03257_), .Q(conv2d_16_prev_row_select) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42012_ ( .CLK(CLK), .D(_03212_), .Q(conv2d_16_act_page_comp_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42013_ ( .CLK(CLK), .D(_03213_), .Q(conv2d_16_act_page_comp_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42014_ ( .CLK(CLK), .D(_03214_), .Q(conv2d_16_act_page_comp_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42015_ ( .CLK(CLK), .D(_03218_), .Q(conv2d_16_act_page_dma_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42016_ ( .CLK(CLK), .D(_03219_), .Q(conv2d_16_act_page_dma_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42017_ ( .CLK(CLK), .D(_03220_), .Q(conv2d_16_act_page_dma_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42018_ ( .CLK(CLK), .D(_03234_), .Q(conv2d_16_filter_page_comp_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42019_ ( .CLK(CLK), .D(_03236_), .Q(conv2d_16_filter_page_dma_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) conv2d_16_out_page_reg  ( .CLK(CLK), .D(_03248_), .Q(conv2d_16_out_page) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42021_ ( .CLK(CLK), .D(_03249_), .Q(conv2d_16_out_page_comp_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42022_ ( .CLK(CLK), .D(_03251_), .Q(conv2d_16_out_page_dma_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42023_ ( .CLK(CLK), .D(_03247_), .Q(conv2d_16_out_laddr_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) conv2d_16_skip_read_filter_reg  ( .CLK(CLK), .D(_03264_), .Q(conv2d_16_skip_read_filter) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) conv2d_16_skip_read_act_reg  ( .CLK(CLK), .D(_03263_), .Q(conv2d_16_skip_read_act) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) conv2d_16_skip_comp_reg  ( .CLK(CLK), .D(_03262_), .Q(conv2d_16_skip_comp) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) conv2d_16_skip_write_out_reg  ( .CLK(CLK), .D(_03265_), .Q(conv2d_16_skip_write_out) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_9_reg  ( .CLK(CLK), .D(_03206_), .Q(axim_flag_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42029_ ( .CLK(CLK), .D(_01583_), .Q(_d1_control_conv2d_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_conv2d_16_cond_3_0_1_reg  ( .CLK(CLK), .D(_01568_), .Q(_control_conv2d_16_cond_3_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_22_reg  ( .CLK(CLK), .D(_03200_), .Q(axim_flag_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_conv2d_16_cond_8_1_1_reg  ( .CLK(CLK), .D(_01570_), .Q(_control_conv2d_16_cond_8_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) set_req_34_reg  ( .CLK(CLK), .D(_03878_), .Q(set_req_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_conv2d_16_cond_14_2_1_reg  ( .CLK(CLK), .D(_01560_), .Q(_control_conv2d_16_cond_14_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_35_reg  ( .CLK(CLK), .D(_03203_), .Q(axim_flag_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_conv2d_16_cond_15_3_1_reg  ( .CLK(CLK), .D(_01561_), .Q(_control_conv2d_16_cond_15_3_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) set_req_287_reg  ( .CLK(CLK), .D(_03876_), .Q(set_req_287) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_conv2d_16_cond_23_4_1_reg  ( .CLK(CLK), .D(_01562_), .Q(_control_conv2d_16_cond_23_4_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_288_reg  ( .CLK(CLK), .D(_03201_), .Q(axim_flag_288) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_conv2d_16_cond_24_5_1_reg  ( .CLK(CLK), .D(_01563_), .Q(_control_conv2d_16_cond_24_5_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) set_req_344_reg  ( .CLK(CLK), .D(_03877_), .Q(set_req_344) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_conv2d_16_cond_30_6_1_reg  ( .CLK(CLK), .D(_01564_), .Q(_control_conv2d_16_cond_30_6_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_345_reg  ( .CLK(CLK), .D(_03202_), .Q(axim_flag_345) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_conv2d_16_cond_31_7_1_reg  ( .CLK(CLK), .D(_01565_), .Q(_control_conv2d_16_cond_31_7_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) set_req_401_reg  ( .CLK(CLK), .D(_03879_), .Q(set_req_401) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_conv2d_16_cond_37_8_1_reg  ( .CLK(CLK), .D(_01566_), .Q(_control_conv2d_16_cond_37_8_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_402_reg  ( .CLK(CLK), .D(_03204_), .Q(axim_flag_402) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_conv2d_16_cond_38_9_1_reg  ( .CLK(CLK), .D(_01567_), .Q(_control_conv2d_16_cond_38_9_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) axim_flag_970_reg  ( .CLK(CLK), .D(_03205_), .Q(axim_flag_970) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _control_conv2d_16_cond_48_10_1_reg  ( .CLK(CLK), .D(_01569_), .Q(_control_conv2d_16_cond_48_10_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _42051_ ( .CLK(CLK), .D(_03229_), .Q(conv2d_16_control_param_index) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _42052_ ( .CLK(CLK), .D(_03344_), .Q(max_pool_serial_18_control_param_index) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _42053_ ( .CLK(CLK), .D(_03293_), .Q(matmul_29_control_param_index) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42054_ ( .CLK(CLK), .D(_03279_), .Q(main_fsm) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42055_ ( .CLK(CLK), .D(_03239_), .Q(conv2d_16_objaddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42056_ ( .CLK(CLK), .D(_03221_), .Q(conv2d_16_arg_objaddr_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42057_ ( .CLK(CLK), .D(_03222_), .Q(conv2d_16_arg_objaddr_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42058_ ( .CLK(CLK), .D(_03223_), .Q(conv2d_16_arg_objaddr_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42059_ ( .CLK(CLK), .D(_03224_), .Q(conv2d_16_arg_objaddr_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42060_ ( .CLK(CLK), .D(_03345_), .Q(max_pool_serial_18_objaddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42061_ ( .CLK(CLK), .D(_03339_), .Q(max_pool_serial_18_arg_objaddr_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42062_ ( .CLK(CLK), .D(_03301_), .Q(matmul_29_objaddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42063_ ( .CLK(CLK), .D(_03285_), .Q(matmul_29_arg_objaddr_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42064_ ( .CLK(CLK), .D(_03286_), .Q(matmul_29_arg_objaddr_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42065_ ( .CLK(CLK), .D(_03287_), .Q(matmul_29_arg_objaddr_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42066_ ( .CLK(CLK), .D(_03288_), .Q(matmul_29_arg_objaddr_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42067_ ( .CLK(CLK), .D(_02713_), .Q(_stream_matmul_29_fsm) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_start_reg  ( .CLK(CLK), .D(_02768_), .Q(_stream_matmul_29_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_end_flag_reg  ( .CLK(CLK), .D(_02712_), .Q(_stream_matmul_29_end_flag) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_term_sink_reg  ( .CLK(CLK), .D(_02769_), .Q(_stream_matmul_29_term_sink) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_busy_reg  ( .CLK(CLK), .D(_02767_), .Q(_stream_matmul_29_source_busy) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42072_ ( .CLK(CLK), .D(_02704_), .Q(_stream_matmul_29_constant_0_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_constant_1_next_constant_data_reg  ( .CLK(CLK), .D(_02709_), .Q(_stream_matmul_29_constant_1_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_constant_2_next_constant_data_reg  ( .CLK(CLK), .D(_02710_), .Q(_stream_matmul_29_constant_2_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_constant_3_next_constant_data_reg  ( .CLK(CLK), .D(_02711_), .Q(_stream_matmul_29_constant_3_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_6_idle_reg  ( .CLK(CLK), .D(_02749_), .Q(_stream_matmul_29_source_6_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42077_ ( .CLK(CLK), .D(_02750_), .Q(_stream_matmul_29_source_6_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42078_ ( .CLK(CLK), .D(_02751_), .Q(_stream_matmul_29_source_6_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42079_ ( .CLK(CLK), .D(_02752_), .Q(_stream_matmul_29_source_6_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42080_ ( .CLK(CLK), .D(_02757_), .Q(_stream_matmul_29_source_6_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42081_ ( .CLK(CLK), .D(_02754_), .Q(_stream_matmul_29_source_6_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_6_source_ram_renable_reg  ( .CLK(CLK), .D(_02755_), .Q(_stream_matmul_29_source_6_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_6_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02756_), .Q(_stream_matmul_29_source_6_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_8_idle_reg  ( .CLK(CLK), .D(_02758_), .Q(_stream_matmul_29_source_8_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42085_ ( .CLK(CLK), .D(_02759_), .Q(_stream_matmul_29_source_8_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42086_ ( .CLK(CLK), .D(_02760_), .Q(_stream_matmul_29_source_8_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42087_ ( .CLK(CLK), .D(_02761_), .Q(_stream_matmul_29_source_8_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42088_ ( .CLK(CLK), .D(_02766_), .Q(_stream_matmul_29_source_8_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42089_ ( .CLK(CLK), .D(_02763_), .Q(_stream_matmul_29_source_8_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_8_source_ram_renable_reg  ( .CLK(CLK), .D(_02764_), .Q(_stream_matmul_29_source_8_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_8_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02765_), .Q(_stream_matmul_29_source_8_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_10_idle_reg  ( .CLK(CLK), .D(_02725_), .Q(_stream_matmul_29_source_10_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42093_ ( .CLK(CLK), .D(_02726_), .Q(_stream_matmul_29_source_10_source_empty_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_12_idle_reg  ( .CLK(CLK), .D(_02727_), .Q(_stream_matmul_29_source_12_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42095_ ( .CLK(CLK), .D(_02728_), .Q(_stream_matmul_29_source_12_source_empty_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_14_idle_reg  ( .CLK(CLK), .D(_02729_), .Q(_stream_matmul_29_source_14_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42097_ ( .CLK(CLK), .D(_02730_), .Q(_stream_matmul_29_source_14_source_empty_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_constant_15_next_constant_data_reg  ( .CLK(CLK), .D(_02705_), .Q(_stream_matmul_29_constant_15_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_constant_16_next_constant_data_reg  ( .CLK(CLK), .D(_02706_), .Q(_stream_matmul_29_constant_16_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _42100_ ( .CLK(CLK), .D(_02707_), .Q(_stream_matmul_29_constant_17_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _42101_ ( .CLK(CLK), .D(_02708_), .Q(_stream_matmul_29_constant_18_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_19_idle_reg  ( .CLK(CLK), .D(_02731_), .Q(_stream_matmul_29_source_19_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42103_ ( .CLK(CLK), .D(_02732_), .Q(_stream_matmul_29_source_19_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42104_ ( .CLK(CLK), .D(_02733_), .Q(_stream_matmul_29_source_19_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42105_ ( .CLK(CLK), .D(_02734_), .Q(_stream_matmul_29_source_19_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42106_ ( .CLK(CLK), .D(_02739_), .Q(_stream_matmul_29_source_19_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42107_ ( .CLK(CLK), .D(_02736_), .Q(_stream_matmul_29_source_19_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_19_source_ram_renable_reg  ( .CLK(CLK), .D(_02737_), .Q(_stream_matmul_29_source_19_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_19_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02738_), .Q(_stream_matmul_29_source_19_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_20_idle_reg  ( .CLK(CLK), .D(_02740_), .Q(_stream_matmul_29_source_20_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42111_ ( .CLK(CLK), .D(_02741_), .Q(_stream_matmul_29_source_20_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42112_ ( .CLK(CLK), .D(_02742_), .Q(_stream_matmul_29_source_20_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42113_ ( .CLK(CLK), .D(_02743_), .Q(_stream_matmul_29_source_20_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42114_ ( .CLK(CLK), .D(_02748_), .Q(_stream_matmul_29_source_20_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42115_ ( .CLK(CLK), .D(_02745_), .Q(_stream_matmul_29_source_20_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_20_source_ram_renable_reg  ( .CLK(CLK), .D(_02746_), .Q(_stream_matmul_29_source_20_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_source_20_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02747_), .Q(_stream_matmul_29_source_20_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42118_ ( .CLK(CLK), .D(_02716_), .Q(_stream_matmul_29_sink_21_sink_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42119_ ( .CLK(CLK), .D(_02717_), .Q(_stream_matmul_29_sink_21_sink_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42120_ ( .CLK(CLK), .D(_02719_), .Q(_stream_matmul_29_sink_21_sink_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42121_ ( .CLK(CLK), .D(_02720_), .Q(_stream_matmul_29_sink_21_sink_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42122_ ( .CLK(CLK), .D(_02714_), .Q(_stream_matmul_29_sink_21_sink_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42123_ ( .CLK(CLK), .D(_02721_), .Q(_stream_matmul_29_sink_21_sink_stride_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42124_ ( .CLK(CLK), .D(_02718_), .Q(_stream_matmul_29_sink_21_sink_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42125_ ( .CLK(CLK), .D(_02722_), .Q(_stream_matmul_29_sink_21_sink_waddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_matmul_29_sink_21_sink_wenable_reg  ( .CLK(CLK), .D(_02724_), .Q(_stream_matmul_29_sink_21_sink_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42127_ ( .CLK(CLK), .D(_02723_), .Q(_stream_matmul_29_sink_21_sink_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42128_ ( .CLK(CLK), .D(_01549_), .Q(_cond_data_817) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42129_ ( .CLK(CLK), .D(_01550_), .Q(_cond_data_824) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42130_ ( .CLK(CLK), .D(_01551_), .Q(_cond_data_831) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42131_ ( .CLK(CLK), .D(_01552_), .Q(_cond_data_838) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42132_ ( .CLK(CLK), .D(_01553_), .Q(_cond_data_845) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _eq_data_851_reg  ( .CLK(CLK), .D(_01686_), .Q(_eq_data_851) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _eq_data_855_reg  ( .CLK(CLK), .D(_01687_), .Q(_eq_data_855) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _eq_data_891_reg  ( .CLK(CLK), .D(_01688_), .Q(_eq_data_891) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _eq_data_894_reg  ( .CLK(CLK), .D(_01689_), .Q(_eq_data_894) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42137_ ( .CLK(CLK), .D(_00298_), .Q(__delay_data_1417) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1419_reg  ( .CLK(CLK), .D(_00300_), .Q(__delay_data_1419) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1422_reg  ( .CLK(CLK), .D(_00303_), .Q(__delay_data_1422) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _42140_ ( .CLK(CLK), .D(_00304_), .Q(__delay_data_1423) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1429_reg  ( .CLK(CLK), .D(_00310_), .Q(__delay_data_1429) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42142_ ( .CLK(CLK), .D(_00325_), .Q(__delay_data_1444) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _42143_ ( .CLK(CLK), .D(_00363_), .Q(__delay_data_1482) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42144_ ( .CLK(CLK), .D(_01555_), .Q(_cond_data_853) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42145_ ( .CLK(CLK), .D(_01815_), .Q(_plus_data_875) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42146_ ( .CLK(CLK), .D(_01816_), .Q(_plus_data_880) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42147_ ( .CLK(CLK), .D(_01818_), .Q(_plus_data_885) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1418_reg  ( .CLK(CLK), .D(_00299_), .Q(__delay_data_1418) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1420_reg  ( .CLK(CLK), .D(_00301_), .Q(__delay_data_1420) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _42150_ ( .CLK(CLK), .D(_00305_), .Q(__delay_data_1424) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42151_ ( .CLK(CLK), .D(_00326_), .Q(__delay_data_1445) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42152_ ( .CLK(CLK), .D(_00341_), .Q(__delay_data_1460) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42153_ ( .CLK(CLK), .D(_00364_), .Q(__delay_data_1483) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1529_reg  ( .CLK(CLK), .D(_00409_), .Q(__delay_data_1529) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1565_reg  ( .CLK(CLK), .D(_00445_), .Q(__delay_data_1565) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42156_ ( .CLK(CLK), .D(_01556_), .Q(_cond_data_857) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1421_reg  ( .CLK(CLK), .D(_00302_), .Q(__delay_data_1421) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _42158_ ( .CLK(CLK), .D(_00306_), .Q(__delay_data_1425) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42159_ ( .CLK(CLK), .D(_00308_), .Q(__delay_data_1427) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42160_ ( .CLK(CLK), .D(_00311_), .Q(__delay_data_1430) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42161_ ( .CLK(CLK), .D(_00327_), .Q(__delay_data_1446) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42162_ ( .CLK(CLK), .D(_00342_), .Q(__delay_data_1461) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42163_ ( .CLK(CLK), .D(_00365_), .Q(__delay_data_1484) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42164_ ( .CLK(CLK), .D(_00387_), .Q(__delay_data_1506) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1530_reg  ( .CLK(CLK), .D(_00410_), .Q(__delay_data_1530) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1566_reg  ( .CLK(CLK), .D(_00446_), .Q(__delay_data_1566) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42167_ ( .CLK(CLK), .D(_01557_), .Q(_cond_data_873) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _42168_ ( .CLK(CLK), .D(_00307_), .Q(__delay_data_1426) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42169_ ( .CLK(CLK), .D(_00309_), .Q(__delay_data_1428) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42170_ ( .CLK(CLK), .D(_00312_), .Q(__delay_data_1431) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42171_ ( .CLK(CLK), .D(_00328_), .Q(__delay_data_1447) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42172_ ( .CLK(CLK), .D(_00343_), .Q(__delay_data_1462) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42173_ ( .CLK(CLK), .D(_00366_), .Q(__delay_data_1485) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42174_ ( .CLK(CLK), .D(_00388_), .Q(__delay_data_1507) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1531_reg  ( .CLK(CLK), .D(_00411_), .Q(__delay_data_1531) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1567_reg  ( .CLK(CLK), .D(_00447_), .Q(__delay_data_1567) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42177_ ( .CLK(CLK), .D(_00313_), .Q(__delay_data_1432) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42178_ ( .CLK(CLK), .D(_00329_), .Q(__delay_data_1448) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42179_ ( .CLK(CLK), .D(_00344_), .Q(__delay_data_1463) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42180_ ( .CLK(CLK), .D(_00367_), .Q(__delay_data_1486) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42181_ ( .CLK(CLK), .D(_00389_), .Q(__delay_data_1508) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1532_reg  ( .CLK(CLK), .D(_00412_), .Q(__delay_data_1532) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1568_reg  ( .CLK(CLK), .D(_00448_), .Q(__delay_data_1568) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42184_ ( .CLK(CLK), .D(_00314_), .Q(__delay_data_1433) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42185_ ( .CLK(CLK), .D(_00330_), .Q(__delay_data_1449) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42186_ ( .CLK(CLK), .D(_00345_), .Q(__delay_data_1464) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42187_ ( .CLK(CLK), .D(_00368_), .Q(__delay_data_1487) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42188_ ( .CLK(CLK), .D(_00390_), .Q(__delay_data_1509) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1533_reg  ( .CLK(CLK), .D(_00413_), .Q(__delay_data_1533) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1569_reg  ( .CLK(CLK), .D(_00449_), .Q(__delay_data_1569) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42191_ ( .CLK(CLK), .D(_00315_), .Q(__delay_data_1434) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42192_ ( .CLK(CLK), .D(_00331_), .Q(__delay_data_1450) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42193_ ( .CLK(CLK), .D(_00346_), .Q(__delay_data_1465) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42194_ ( .CLK(CLK), .D(_00369_), .Q(__delay_data_1488) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42195_ ( .CLK(CLK), .D(_00391_), .Q(__delay_data_1510) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1534_reg  ( .CLK(CLK), .D(_00414_), .Q(__delay_data_1534) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1570_reg  ( .CLK(CLK), .D(_00450_), .Q(__delay_data_1570) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42198_ ( .CLK(CLK), .D(_00316_), .Q(__delay_data_1435) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42199_ ( .CLK(CLK), .D(_00332_), .Q(__delay_data_1451) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42200_ ( .CLK(CLK), .D(_00347_), .Q(__delay_data_1466) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42201_ ( .CLK(CLK), .D(_00370_), .Q(__delay_data_1489) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42202_ ( .CLK(CLK), .D(_00392_), .Q(__delay_data_1511) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1535_reg  ( .CLK(CLK), .D(_00415_), .Q(__delay_data_1535) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1571_reg  ( .CLK(CLK), .D(_00451_), .Q(__delay_data_1571) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42205_ ( .CLK(CLK), .D(_00317_), .Q(__delay_data_1436) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42206_ ( .CLK(CLK), .D(_00333_), .Q(__delay_data_1452) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42207_ ( .CLK(CLK), .D(_00348_), .Q(__delay_data_1467) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42208_ ( .CLK(CLK), .D(_00371_), .Q(__delay_data_1490) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42209_ ( .CLK(CLK), .D(_00393_), .Q(__delay_data_1512) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1536_reg  ( .CLK(CLK), .D(_00416_), .Q(__delay_data_1536) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1572_reg  ( .CLK(CLK), .D(_00452_), .Q(__delay_data_1572) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42212_ ( .CLK(CLK), .D(_00318_), .Q(__delay_data_1437) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42213_ ( .CLK(CLK), .D(_00334_), .Q(__delay_data_1453) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42214_ ( .CLK(CLK), .D(_00349_), .Q(__delay_data_1468) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42215_ ( .CLK(CLK), .D(_00372_), .Q(__delay_data_1491) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42216_ ( .CLK(CLK), .D(_00394_), .Q(__delay_data_1513) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1537_reg  ( .CLK(CLK), .D(_00417_), .Q(__delay_data_1537) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1573_reg  ( .CLK(CLK), .D(_00453_), .Q(__delay_data_1573) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42219_ ( .CLK(CLK), .D(_00319_), .Q(__delay_data_1438) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42220_ ( .CLK(CLK), .D(_00335_), .Q(__delay_data_1454) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42221_ ( .CLK(CLK), .D(_00350_), .Q(__delay_data_1469) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42222_ ( .CLK(CLK), .D(_00373_), .Q(__delay_data_1492) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42223_ ( .CLK(CLK), .D(_00395_), .Q(__delay_data_1514) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1538_reg  ( .CLK(CLK), .D(_00418_), .Q(__delay_data_1538) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1574_reg  ( .CLK(CLK), .D(_00454_), .Q(__delay_data_1574) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42226_ ( .CLK(CLK), .D(_00320_), .Q(__delay_data_1439) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42227_ ( .CLK(CLK), .D(_00336_), .Q(__delay_data_1455) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42228_ ( .CLK(CLK), .D(_00351_), .Q(__delay_data_1470) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42229_ ( .CLK(CLK), .D(_00374_), .Q(__delay_data_1493) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42230_ ( .CLK(CLK), .D(_00396_), .Q(__delay_data_1515) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1539_reg  ( .CLK(CLK), .D(_00419_), .Q(__delay_data_1539) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1575_reg  ( .CLK(CLK), .D(_00455_), .Q(__delay_data_1575) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42233_ ( .CLK(CLK), .D(_00321_), .Q(__delay_data_1440) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42234_ ( .CLK(CLK), .D(_00337_), .Q(__delay_data_1456) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42235_ ( .CLK(CLK), .D(_00352_), .Q(__delay_data_1471) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42236_ ( .CLK(CLK), .D(_00375_), .Q(__delay_data_1494) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42237_ ( .CLK(CLK), .D(_00397_), .Q(__delay_data_1516) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1540_reg  ( .CLK(CLK), .D(_00420_), .Q(__delay_data_1540) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1576_reg  ( .CLK(CLK), .D(_00456_), .Q(__delay_data_1576) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _42240_ ( .CLK(CLK), .D(_01089_), .Q(__substreamoutput_data_876) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42241_ ( .CLK(CLK), .D(_00322_), .Q(__delay_data_1441) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42242_ ( .CLK(CLK), .D(_00338_), .Q(__delay_data_1457) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42243_ ( .CLK(CLK), .D(_00353_), .Q(__delay_data_1472) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42244_ ( .CLK(CLK), .D(_00376_), .Q(__delay_data_1495) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42245_ ( .CLK(CLK), .D(_00398_), .Q(__delay_data_1517) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1541_reg  ( .CLK(CLK), .D(_00421_), .Q(__delay_data_1541) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1577_reg  ( .CLK(CLK), .D(_00457_), .Q(__delay_data_1577) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42248_ ( .CLK(CLK), .D(_00323_), .Q(__delay_data_1442) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42249_ ( .CLK(CLK), .D(_00339_), .Q(__delay_data_1458) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42250_ ( .CLK(CLK), .D(_00354_), .Q(__delay_data_1473) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42251_ ( .CLK(CLK), .D(_00377_), .Q(__delay_data_1496) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42252_ ( .CLK(CLK), .D(_00399_), .Q(__delay_data_1518) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1542_reg  ( .CLK(CLK), .D(_00422_), .Q(__delay_data_1542) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1578_reg  ( .CLK(CLK), .D(_00458_), .Q(__delay_data_1578) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42255_ ( .CLK(CLK), .D(_01104_), .Q(__substreamoutput_data_878) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42256_ ( .CLK(CLK), .D(_00324_), .Q(__delay_data_1443) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42257_ ( .CLK(CLK), .D(_00340_), .Q(__delay_data_1459) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42258_ ( .CLK(CLK), .D(_00355_), .Q(__delay_data_1474) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42259_ ( .CLK(CLK), .D(_00378_), .Q(__delay_data_1497) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42260_ ( .CLK(CLK), .D(_00400_), .Q(__delay_data_1519) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1543_reg  ( .CLK(CLK), .D(_00423_), .Q(__delay_data_1543) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1579_reg  ( .CLK(CLK), .D(_00459_), .Q(__delay_data_1579) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42263_ ( .CLK(CLK), .D(_00356_), .Q(__delay_data_1475) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42264_ ( .CLK(CLK), .D(_00379_), .Q(__delay_data_1498) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42265_ ( .CLK(CLK), .D(_00401_), .Q(__delay_data_1520) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1544_reg  ( .CLK(CLK), .D(_00424_), .Q(__delay_data_1544) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1580_reg  ( .CLK(CLK), .D(_00460_), .Q(__delay_data_1580) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42268_ ( .CLK(CLK), .D(_00357_), .Q(__delay_data_1476) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42269_ ( .CLK(CLK), .D(_00380_), .Q(__delay_data_1499) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42270_ ( .CLK(CLK), .D(_00402_), .Q(__delay_data_1521) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1545_reg  ( .CLK(CLK), .D(_00425_), .Q(__delay_data_1545) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1581_reg  ( .CLK(CLK), .D(_00461_), .Q(__delay_data_1581) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42273_ ( .CLK(CLK), .D(_00358_), .Q(__delay_data_1477) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42274_ ( .CLK(CLK), .D(_00381_), .Q(__delay_data_1500) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42275_ ( .CLK(CLK), .D(_00403_), .Q(__delay_data_1522) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1546_reg  ( .CLK(CLK), .D(_00426_), .Q(__delay_data_1546) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1582_reg  ( .CLK(CLK), .D(_00462_), .Q(__delay_data_1582) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42278_ ( .CLK(CLK), .D(_00359_), .Q(__delay_data_1478) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42279_ ( .CLK(CLK), .D(_00382_), .Q(__delay_data_1501) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42280_ ( .CLK(CLK), .D(_00404_), .Q(__delay_data_1523) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1547_reg  ( .CLK(CLK), .D(_00427_), .Q(__delay_data_1547) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1583_reg  ( .CLK(CLK), .D(_00463_), .Q(__delay_data_1583) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42283_ ( .CLK(CLK), .D(_00360_), .Q(__delay_data_1479) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42284_ ( .CLK(CLK), .D(_00383_), .Q(__delay_data_1502) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42285_ ( .CLK(CLK), .D(_00405_), .Q(__delay_data_1524) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1548_reg  ( .CLK(CLK), .D(_00428_), .Q(__delay_data_1548) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1584_reg  ( .CLK(CLK), .D(_00464_), .Q(__delay_data_1584) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42288_ ( .CLK(CLK), .D(_00361_), .Q(__delay_data_1480) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42289_ ( .CLK(CLK), .D(_00384_), .Q(__delay_data_1503) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42290_ ( .CLK(CLK), .D(_00406_), .Q(__delay_data_1525) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1549_reg  ( .CLK(CLK), .D(_00429_), .Q(__delay_data_1549) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1585_reg  ( .CLK(CLK), .D(_00465_), .Q(__delay_data_1585) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42293_ ( .CLK(CLK), .D(_01099_), .Q(__substreamoutput_data_881) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __substreamoutput_data_882_reg  ( .CLK(CLK), .D(_01100_), .Q(__substreamoutput_data_882) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42295_ ( .CLK(CLK), .D(_00362_), .Q(__delay_data_1481) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42296_ ( .CLK(CLK), .D(_00385_), .Q(__delay_data_1504) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42297_ ( .CLK(CLK), .D(_00407_), .Q(__delay_data_1526) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1550_reg  ( .CLK(CLK), .D(_00430_), .Q(__delay_data_1550) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1586_reg  ( .CLK(CLK), .D(_00466_), .Q(__delay_data_1586) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42300_ ( .CLK(CLK), .D(_01817_), .Q(_plus_data_883) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42301_ ( .CLK(CLK), .D(_00386_), .Q(__delay_data_1505) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42302_ ( .CLK(CLK), .D(_00408_), .Q(__delay_data_1527) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1551_reg  ( .CLK(CLK), .D(_00431_), .Q(__delay_data_1551) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1587_reg  ( .CLK(CLK), .D(_00467_), .Q(__delay_data_1587) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1602_reg  ( .CLK(CLK), .D(_00279_), .Q(__delay_data_1602) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1552_reg  ( .CLK(CLK), .D(_00432_), .Q(__delay_data_1552) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1588_reg  ( .CLK(CLK), .D(_00468_), .Q(__delay_data_1588) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1603_reg  ( .CLK(CLK), .D(_00280_), .Q(__delay_data_1603) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1553_reg  ( .CLK(CLK), .D(_00433_), .Q(__delay_data_1553) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1589_reg  ( .CLK(CLK), .D(_00469_), .Q(__delay_data_1589) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1604_reg  ( .CLK(CLK), .D(_00281_), .Q(__delay_data_1604) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1554_reg  ( .CLK(CLK), .D(_00434_), .Q(__delay_data_1554) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1590_reg  ( .CLK(CLK), .D(_00470_), .Q(__delay_data_1590) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1605_reg  ( .CLK(CLK), .D(_00282_), .Q(__delay_data_1605) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1555_reg  ( .CLK(CLK), .D(_00435_), .Q(__delay_data_1555) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1591_reg  ( .CLK(CLK), .D(_00471_), .Q(__delay_data_1591) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1606_reg  ( .CLK(CLK), .D(_00283_), .Q(__delay_data_1606) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1556_reg  ( .CLK(CLK), .D(_00436_), .Q(__delay_data_1556) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1592_reg  ( .CLK(CLK), .D(_00472_), .Q(__delay_data_1592) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1607_reg  ( .CLK(CLK), .D(_00284_), .Q(__delay_data_1607) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1557_reg  ( .CLK(CLK), .D(_00437_), .Q(__delay_data_1557) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1593_reg  ( .CLK(CLK), .D(_00473_), .Q(__delay_data_1593) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1608_reg  ( .CLK(CLK), .D(_00285_), .Q(__delay_data_1608) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1558_reg  ( .CLK(CLK), .D(_00438_), .Q(__delay_data_1558) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1594_reg  ( .CLK(CLK), .D(_00474_), .Q(__delay_data_1594) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1609_reg  ( .CLK(CLK), .D(_00286_), .Q(__delay_data_1609) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1559_reg  ( .CLK(CLK), .D(_00439_), .Q(__delay_data_1559) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1595_reg  ( .CLK(CLK), .D(_00475_), .Q(__delay_data_1595) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1610_reg  ( .CLK(CLK), .D(_00287_), .Q(__delay_data_1610) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1560_reg  ( .CLK(CLK), .D(_00440_), .Q(__delay_data_1560) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1596_reg  ( .CLK(CLK), .D(_00476_), .Q(__delay_data_1596) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1611_reg  ( .CLK(CLK), .D(_00288_), .Q(__delay_data_1611) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42333_ ( .CLK(CLK), .D(_01101_), .Q(__substreamoutput_data_886) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1561_reg  ( .CLK(CLK), .D(_00441_), .Q(__delay_data_1561) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1597_reg  ( .CLK(CLK), .D(_00477_), .Q(__delay_data_1597) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1612_reg  ( .CLK(CLK), .D(_00289_), .Q(__delay_data_1612) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greaterthan_data_888_reg  ( .CLK(CLK), .D(_01701_), .Q(_greaterthan_data_888) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42338_ ( .CLK(CLK), .D(_00278_), .Q(__delay_data_1528) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1562_reg  ( .CLK(CLK), .D(_00442_), .Q(__delay_data_1562) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1598_reg  ( .CLK(CLK), .D(_00478_), .Q(__delay_data_1598) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1613_reg  ( .CLK(CLK), .D(_00290_), .Q(__delay_data_1613) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42342_ ( .CLK(CLK), .D(_01547_), .Q(_cond_data_890) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1563_reg  ( .CLK(CLK), .D(_00443_), .Q(__delay_data_1563) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42344_ ( .CLK(CLK), .D(_00444_), .Q(__delay_data_1564) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1599_reg  ( .CLK(CLK), .D(_00479_), .Q(__delay_data_1599) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1614_reg  ( .CLK(CLK), .D(_00291_), .Q(__delay_data_1614) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42347_ ( .CLK(CLK), .D(_01558_), .Q(_cond_data_893) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1600_reg  ( .CLK(CLK), .D(_00480_), .Q(__delay_data_1600) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42349_ ( .CLK(CLK), .D(_00481_), .Q(__delay_data_1601) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1615_reg  ( .CLK(CLK), .D(_00482_), .Q(__delay_data_1615) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42351_ ( .CLK(CLK), .D(_01559_), .Q(_cond_data_896) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1616_reg  ( .CLK(CLK), .D(_00483_), .Q(__delay_data_1616) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _42353_ ( .CLK(CLK), .D(_01448_), .Q(__variable_wdata_796) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __variable_wdata_797_reg  ( .CLK(CLK), .D(_01449_), .Q(__variable_wdata_797) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __variable_wdata_798_reg  ( .CLK(CLK), .D(_01450_), .Q(__variable_wdata_798) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __variable_wdata_799_reg  ( .CLK(CLK), .D(_01451_), .Q(__variable_wdata_799) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42357_ ( .CLK(CLK), .D(_02416_), .Q(_source_stream_matmul_29_source_6_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42358_ ( .CLK(CLK), .D(_02417_), .Q(_source_stream_matmul_29_source_6_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42359_ ( .CLK(CLK), .D(_02418_), .Q(_source_stream_matmul_29_source_6_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42360_ ( .CLK(CLK), .D(_02419_), .Q(_source_stream_matmul_29_source_6_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42361_ ( .CLK(CLK), .D(_02420_), .Q(_source_stream_matmul_29_source_6_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42362_ ( .CLK(CLK), .D(_02421_), .Q(_source_stream_matmul_29_source_6_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42363_ ( .CLK(CLK), .D(_02422_), .Q(_source_stream_matmul_29_source_6_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42364_ ( .CLK(CLK), .D(_02423_), .Q(_source_stream_matmul_29_source_6_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42365_ ( .CLK(CLK), .D(_02428_), .Q(_source_stream_matmul_29_source_6_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42366_ ( .CLK(CLK), .D(_02429_), .Q(_source_stream_matmul_29_source_6_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42367_ ( .CLK(CLK), .D(_02430_), .Q(_source_stream_matmul_29_source_6_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42368_ ( .CLK(CLK), .D(_02431_), .Q(_source_stream_matmul_29_source_6_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42369_ ( .CLK(CLK), .D(_02412_), .Q(_source_stream_matmul_29_source_6_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42370_ ( .CLK(CLK), .D(_02413_), .Q(_source_stream_matmul_29_source_6_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42371_ ( .CLK(CLK), .D(_02414_), .Q(_source_stream_matmul_29_source_6_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42372_ ( .CLK(CLK), .D(_02415_), .Q(_source_stream_matmul_29_source_6_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42373_ ( .CLK(CLK), .D(_02424_), .Q(_source_stream_matmul_29_source_6_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42374_ ( .CLK(CLK), .D(_02425_), .Q(_source_stream_matmul_29_source_6_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42375_ ( .CLK(CLK), .D(_02426_), .Q(_source_stream_matmul_29_source_6_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42376_ ( .CLK(CLK), .D(_02427_), .Q(_source_stream_matmul_29_source_6_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42377_ ( .CLK(CLK), .D(_02432_), .Q(_source_stream_matmul_29_source_6_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42378_ ( .CLK(CLK), .D(_02433_), .Q(_source_stream_matmul_29_source_6_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42379_ ( .CLK(CLK), .D(_02434_), .Q(_source_stream_matmul_29_source_6_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42380_ ( .CLK(CLK), .D(_02435_), .Q(_source_stream_matmul_29_source_6_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42381_ ( .CLK(CLK), .D(_01452_), .Q(__variable_wdata_812) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42382_ ( .CLK(CLK), .D(_02440_), .Q(_source_stream_matmul_29_source_8_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42383_ ( .CLK(CLK), .D(_02441_), .Q(_source_stream_matmul_29_source_8_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42384_ ( .CLK(CLK), .D(_02442_), .Q(_source_stream_matmul_29_source_8_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42385_ ( .CLK(CLK), .D(_02443_), .Q(_source_stream_matmul_29_source_8_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42386_ ( .CLK(CLK), .D(_02444_), .Q(_source_stream_matmul_29_source_8_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42387_ ( .CLK(CLK), .D(_02445_), .Q(_source_stream_matmul_29_source_8_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42388_ ( .CLK(CLK), .D(_02446_), .Q(_source_stream_matmul_29_source_8_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42389_ ( .CLK(CLK), .D(_02447_), .Q(_source_stream_matmul_29_source_8_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42390_ ( .CLK(CLK), .D(_02452_), .Q(_source_stream_matmul_29_source_8_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42391_ ( .CLK(CLK), .D(_02453_), .Q(_source_stream_matmul_29_source_8_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42392_ ( .CLK(CLK), .D(_02454_), .Q(_source_stream_matmul_29_source_8_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42393_ ( .CLK(CLK), .D(_02455_), .Q(_source_stream_matmul_29_source_8_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42394_ ( .CLK(CLK), .D(_02436_), .Q(_source_stream_matmul_29_source_8_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42395_ ( .CLK(CLK), .D(_02437_), .Q(_source_stream_matmul_29_source_8_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42396_ ( .CLK(CLK), .D(_02438_), .Q(_source_stream_matmul_29_source_8_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42397_ ( .CLK(CLK), .D(_02439_), .Q(_source_stream_matmul_29_source_8_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42398_ ( .CLK(CLK), .D(_02448_), .Q(_source_stream_matmul_29_source_8_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42399_ ( .CLK(CLK), .D(_02449_), .Q(_source_stream_matmul_29_source_8_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42400_ ( .CLK(CLK), .D(_02450_), .Q(_source_stream_matmul_29_source_8_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42401_ ( .CLK(CLK), .D(_02451_), .Q(_source_stream_matmul_29_source_8_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42402_ ( .CLK(CLK), .D(_02456_), .Q(_source_stream_matmul_29_source_8_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42403_ ( .CLK(CLK), .D(_02457_), .Q(_source_stream_matmul_29_source_8_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42404_ ( .CLK(CLK), .D(_02458_), .Q(_source_stream_matmul_29_source_8_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42405_ ( .CLK(CLK), .D(_02459_), .Q(_source_stream_matmul_29_source_8_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42406_ ( .CLK(CLK), .D(_01453_), .Q(__variable_wdata_819) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42407_ ( .CLK(CLK), .D(_01454_), .Q(__variable_wdata_826) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42408_ ( .CLK(CLK), .D(_01455_), .Q(__variable_wdata_833) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42409_ ( .CLK(CLK), .D(_01456_), .Q(__variable_wdata_840) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __variable_wdata_846_reg  ( .CLK(CLK), .D(_01457_), .Q(__variable_wdata_846) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __variable_wdata_847_reg  ( .CLK(CLK), .D(_01458_), .Q(__variable_wdata_847) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _42412_ ( .CLK(CLK), .D(_01459_), .Q(__variable_wdata_848) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _42413_ ( .CLK(CLK), .D(_01460_), .Q(__variable_wdata_849) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42414_ ( .CLK(CLK), .D(_02368_), .Q(_source_stream_matmul_29_source_19_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42415_ ( .CLK(CLK), .D(_02369_), .Q(_source_stream_matmul_29_source_19_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42416_ ( .CLK(CLK), .D(_02370_), .Q(_source_stream_matmul_29_source_19_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42417_ ( .CLK(CLK), .D(_02371_), .Q(_source_stream_matmul_29_source_19_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42418_ ( .CLK(CLK), .D(_02372_), .Q(_source_stream_matmul_29_source_19_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42419_ ( .CLK(CLK), .D(_02373_), .Q(_source_stream_matmul_29_source_19_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42420_ ( .CLK(CLK), .D(_02374_), .Q(_source_stream_matmul_29_source_19_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42421_ ( .CLK(CLK), .D(_02375_), .Q(_source_stream_matmul_29_source_19_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42422_ ( .CLK(CLK), .D(_02380_), .Q(_source_stream_matmul_29_source_19_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42423_ ( .CLK(CLK), .D(_02381_), .Q(_source_stream_matmul_29_source_19_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42424_ ( .CLK(CLK), .D(_02382_), .Q(_source_stream_matmul_29_source_19_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42425_ ( .CLK(CLK), .D(_02383_), .Q(_source_stream_matmul_29_source_19_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42426_ ( .CLK(CLK), .D(_02364_), .Q(_source_stream_matmul_29_source_19_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42427_ ( .CLK(CLK), .D(_02365_), .Q(_source_stream_matmul_29_source_19_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42428_ ( .CLK(CLK), .D(_02366_), .Q(_source_stream_matmul_29_source_19_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42429_ ( .CLK(CLK), .D(_02367_), .Q(_source_stream_matmul_29_source_19_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42430_ ( .CLK(CLK), .D(_02376_), .Q(_source_stream_matmul_29_source_19_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42431_ ( .CLK(CLK), .D(_02377_), .Q(_source_stream_matmul_29_source_19_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42432_ ( .CLK(CLK), .D(_02378_), .Q(_source_stream_matmul_29_source_19_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42433_ ( .CLK(CLK), .D(_02379_), .Q(_source_stream_matmul_29_source_19_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42434_ ( .CLK(CLK), .D(_02384_), .Q(_source_stream_matmul_29_source_19_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42435_ ( .CLK(CLK), .D(_02385_), .Q(_source_stream_matmul_29_source_19_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42436_ ( .CLK(CLK), .D(_02386_), .Q(_source_stream_matmul_29_source_19_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42437_ ( .CLK(CLK), .D(_02387_), .Q(_source_stream_matmul_29_source_19_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42438_ ( .CLK(CLK), .D(_01461_), .Q(__variable_wdata_850) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42439_ ( .CLK(CLK), .D(_02392_), .Q(_source_stream_matmul_29_source_20_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42440_ ( .CLK(CLK), .D(_02393_), .Q(_source_stream_matmul_29_source_20_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42441_ ( .CLK(CLK), .D(_02394_), .Q(_source_stream_matmul_29_source_20_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42442_ ( .CLK(CLK), .D(_02395_), .Q(_source_stream_matmul_29_source_20_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42443_ ( .CLK(CLK), .D(_02396_), .Q(_source_stream_matmul_29_source_20_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42444_ ( .CLK(CLK), .D(_02397_), .Q(_source_stream_matmul_29_source_20_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42445_ ( .CLK(CLK), .D(_02398_), .Q(_source_stream_matmul_29_source_20_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42446_ ( .CLK(CLK), .D(_02399_), .Q(_source_stream_matmul_29_source_20_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42447_ ( .CLK(CLK), .D(_02404_), .Q(_source_stream_matmul_29_source_20_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42448_ ( .CLK(CLK), .D(_02405_), .Q(_source_stream_matmul_29_source_20_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42449_ ( .CLK(CLK), .D(_02406_), .Q(_source_stream_matmul_29_source_20_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42450_ ( .CLK(CLK), .D(_02407_), .Q(_source_stream_matmul_29_source_20_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42451_ ( .CLK(CLK), .D(_02388_), .Q(_source_stream_matmul_29_source_20_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42452_ ( .CLK(CLK), .D(_02389_), .Q(_source_stream_matmul_29_source_20_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42453_ ( .CLK(CLK), .D(_02390_), .Q(_source_stream_matmul_29_source_20_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42454_ ( .CLK(CLK), .D(_02391_), .Q(_source_stream_matmul_29_source_20_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42455_ ( .CLK(CLK), .D(_02400_), .Q(_source_stream_matmul_29_source_20_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42456_ ( .CLK(CLK), .D(_02401_), .Q(_source_stream_matmul_29_source_20_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42457_ ( .CLK(CLK), .D(_02402_), .Q(_source_stream_matmul_29_source_20_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42458_ ( .CLK(CLK), .D(_02403_), .Q(_source_stream_matmul_29_source_20_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42459_ ( .CLK(CLK), .D(_02408_), .Q(_source_stream_matmul_29_source_20_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42460_ ( .CLK(CLK), .D(_02409_), .Q(_source_stream_matmul_29_source_20_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42461_ ( .CLK(CLK), .D(_02410_), .Q(_source_stream_matmul_29_source_20_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42462_ ( .CLK(CLK), .D(_02411_), .Q(_source_stream_matmul_29_source_20_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1223_1_reg  ( .CLK(CLK), .D(_01150_), .Q(__tmp_1223_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _42464_ ( .CLK(CLK), .D(_01462_), .Q(__variable_wdata_864) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _set_flag_1224_reg  ( .CLK(CLK), .D(_01872_), .Q(_set_flag_1224) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42466_ ( .CLK(CLK), .D(_00947_), .Q(__stream_matmul_29_sink_21_sink_offset_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42467_ ( .CLK(CLK), .D(_00958_), .Q(__stream_matmul_29_sink_21_sink_offset_0_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42468_ ( .CLK(CLK), .D(_00969_), .Q(__stream_matmul_29_sink_21_sink_offset_0_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42469_ ( .CLK(CLK), .D(_00972_), .Q(__stream_matmul_29_sink_21_sink_offset_0_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42470_ ( .CLK(CLK), .D(_00973_), .Q(__stream_matmul_29_sink_21_sink_offset_0_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42471_ ( .CLK(CLK), .D(_00974_), .Q(__stream_matmul_29_sink_21_sink_offset_0_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42472_ ( .CLK(CLK), .D(_00975_), .Q(__stream_matmul_29_sink_21_sink_offset_0_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42473_ ( .CLK(CLK), .D(_00976_), .Q(__stream_matmul_29_sink_21_sink_offset_0_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42474_ ( .CLK(CLK), .D(_00977_), .Q(__stream_matmul_29_sink_21_sink_offset_0_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42475_ ( .CLK(CLK), .D(_00937_), .Q(__stream_matmul_29_sink_21_sink_offset_0_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42476_ ( .CLK(CLK), .D(_00938_), .Q(__stream_matmul_29_sink_21_sink_offset_0_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42477_ ( .CLK(CLK), .D(_00939_), .Q(__stream_matmul_29_sink_21_sink_offset_0_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42478_ ( .CLK(CLK), .D(_00940_), .Q(__stream_matmul_29_sink_21_sink_offset_0_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42479_ ( .CLK(CLK), .D(_00941_), .Q(__stream_matmul_29_sink_21_sink_offset_0_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42480_ ( .CLK(CLK), .D(_00942_), .Q(__stream_matmul_29_sink_21_sink_offset_0_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42481_ ( .CLK(CLK), .D(_00943_), .Q(__stream_matmul_29_sink_21_sink_offset_0_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42482_ ( .CLK(CLK), .D(_00944_), .Q(__stream_matmul_29_sink_21_sink_offset_0_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42483_ ( .CLK(CLK), .D(_00945_), .Q(__stream_matmul_29_sink_21_sink_offset_0_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42484_ ( .CLK(CLK), .D(_00946_), .Q(__stream_matmul_29_sink_21_sink_offset_0_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42485_ ( .CLK(CLK), .D(_00948_), .Q(__stream_matmul_29_sink_21_sink_offset_0_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42486_ ( .CLK(CLK), .D(_00949_), .Q(__stream_matmul_29_sink_21_sink_offset_0_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42487_ ( .CLK(CLK), .D(_00950_), .Q(__stream_matmul_29_sink_21_sink_offset_0_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42488_ ( .CLK(CLK), .D(_00951_), .Q(__stream_matmul_29_sink_21_sink_offset_0_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42489_ ( .CLK(CLK), .D(_00952_), .Q(__stream_matmul_29_sink_21_sink_offset_0_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42490_ ( .CLK(CLK), .D(_00953_), .Q(__stream_matmul_29_sink_21_sink_offset_0_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42491_ ( .CLK(CLK), .D(_00954_), .Q(__stream_matmul_29_sink_21_sink_offset_0_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42492_ ( .CLK(CLK), .D(_00955_), .Q(__stream_matmul_29_sink_21_sink_offset_0_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42493_ ( .CLK(CLK), .D(_00956_), .Q(__stream_matmul_29_sink_21_sink_offset_0_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42494_ ( .CLK(CLK), .D(_00957_), .Q(__stream_matmul_29_sink_21_sink_offset_0_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42495_ ( .CLK(CLK), .D(_00959_), .Q(__stream_matmul_29_sink_21_sink_offset_0_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42496_ ( .CLK(CLK), .D(_00960_), .Q(__stream_matmul_29_sink_21_sink_offset_0_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42497_ ( .CLK(CLK), .D(_00961_), .Q(__stream_matmul_29_sink_21_sink_offset_0_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42498_ ( .CLK(CLK), .D(_00962_), .Q(__stream_matmul_29_sink_21_sink_offset_0_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42499_ ( .CLK(CLK), .D(_00963_), .Q(__stream_matmul_29_sink_21_sink_offset_0_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42500_ ( .CLK(CLK), .D(_00964_), .Q(__stream_matmul_29_sink_21_sink_offset_0_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42501_ ( .CLK(CLK), .D(_00965_), .Q(__stream_matmul_29_sink_21_sink_offset_0_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42502_ ( .CLK(CLK), .D(_00966_), .Q(__stream_matmul_29_sink_21_sink_offset_0_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42503_ ( .CLK(CLK), .D(_00967_), .Q(__stream_matmul_29_sink_21_sink_offset_0_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42504_ ( .CLK(CLK), .D(_00968_), .Q(__stream_matmul_29_sink_21_sink_offset_0_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42505_ ( .CLK(CLK), .D(_00970_), .Q(__stream_matmul_29_sink_21_sink_offset_0_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42506_ ( .CLK(CLK), .D(_00971_), .Q(__stream_matmul_29_sink_21_sink_offset_0_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42507_ ( .CLK(CLK), .D(_00988_), .Q(__stream_matmul_29_sink_21_sink_size_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42508_ ( .CLK(CLK), .D(_00999_), .Q(__stream_matmul_29_sink_21_sink_size_1_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42509_ ( .CLK(CLK), .D(_01010_), .Q(__stream_matmul_29_sink_21_sink_size_1_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42510_ ( .CLK(CLK), .D(_01013_), .Q(__stream_matmul_29_sink_21_sink_size_1_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42511_ ( .CLK(CLK), .D(_01014_), .Q(__stream_matmul_29_sink_21_sink_size_1_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42512_ ( .CLK(CLK), .D(_01015_), .Q(__stream_matmul_29_sink_21_sink_size_1_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42513_ ( .CLK(CLK), .D(_01016_), .Q(__stream_matmul_29_sink_21_sink_size_1_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42514_ ( .CLK(CLK), .D(_01017_), .Q(__stream_matmul_29_sink_21_sink_size_1_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42515_ ( .CLK(CLK), .D(_01018_), .Q(__stream_matmul_29_sink_21_sink_size_1_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42516_ ( .CLK(CLK), .D(_00978_), .Q(__stream_matmul_29_sink_21_sink_size_1_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42517_ ( .CLK(CLK), .D(_00979_), .Q(__stream_matmul_29_sink_21_sink_size_1_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42518_ ( .CLK(CLK), .D(_00980_), .Q(__stream_matmul_29_sink_21_sink_size_1_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42519_ ( .CLK(CLK), .D(_00981_), .Q(__stream_matmul_29_sink_21_sink_size_1_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42520_ ( .CLK(CLK), .D(_00982_), .Q(__stream_matmul_29_sink_21_sink_size_1_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42521_ ( .CLK(CLK), .D(_00983_), .Q(__stream_matmul_29_sink_21_sink_size_1_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42522_ ( .CLK(CLK), .D(_00984_), .Q(__stream_matmul_29_sink_21_sink_size_1_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42523_ ( .CLK(CLK), .D(_00985_), .Q(__stream_matmul_29_sink_21_sink_size_1_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42524_ ( .CLK(CLK), .D(_00986_), .Q(__stream_matmul_29_sink_21_sink_size_1_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42525_ ( .CLK(CLK), .D(_00987_), .Q(__stream_matmul_29_sink_21_sink_size_1_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42526_ ( .CLK(CLK), .D(_00989_), .Q(__stream_matmul_29_sink_21_sink_size_1_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42527_ ( .CLK(CLK), .D(_00990_), .Q(__stream_matmul_29_sink_21_sink_size_1_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42528_ ( .CLK(CLK), .D(_00991_), .Q(__stream_matmul_29_sink_21_sink_size_1_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42529_ ( .CLK(CLK), .D(_00992_), .Q(__stream_matmul_29_sink_21_sink_size_1_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42530_ ( .CLK(CLK), .D(_00993_), .Q(__stream_matmul_29_sink_21_sink_size_1_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42531_ ( .CLK(CLK), .D(_00994_), .Q(__stream_matmul_29_sink_21_sink_size_1_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42532_ ( .CLK(CLK), .D(_00995_), .Q(__stream_matmul_29_sink_21_sink_size_1_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42533_ ( .CLK(CLK), .D(_00996_), .Q(__stream_matmul_29_sink_21_sink_size_1_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42534_ ( .CLK(CLK), .D(_00997_), .Q(__stream_matmul_29_sink_21_sink_size_1_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42535_ ( .CLK(CLK), .D(_00998_), .Q(__stream_matmul_29_sink_21_sink_size_1_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42536_ ( .CLK(CLK), .D(_01000_), .Q(__stream_matmul_29_sink_21_sink_size_1_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42537_ ( .CLK(CLK), .D(_01001_), .Q(__stream_matmul_29_sink_21_sink_size_1_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42538_ ( .CLK(CLK), .D(_01002_), .Q(__stream_matmul_29_sink_21_sink_size_1_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42539_ ( .CLK(CLK), .D(_01003_), .Q(__stream_matmul_29_sink_21_sink_size_1_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42540_ ( .CLK(CLK), .D(_01004_), .Q(__stream_matmul_29_sink_21_sink_size_1_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42541_ ( .CLK(CLK), .D(_01005_), .Q(__stream_matmul_29_sink_21_sink_size_1_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42542_ ( .CLK(CLK), .D(_01006_), .Q(__stream_matmul_29_sink_21_sink_size_1_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42543_ ( .CLK(CLK), .D(_01007_), .Q(__stream_matmul_29_sink_21_sink_size_1_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42544_ ( .CLK(CLK), .D(_01008_), .Q(__stream_matmul_29_sink_21_sink_size_1_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42545_ ( .CLK(CLK), .D(_01009_), .Q(__stream_matmul_29_sink_21_sink_size_1_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42546_ ( .CLK(CLK), .D(_01011_), .Q(__stream_matmul_29_sink_21_sink_size_1_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42547_ ( .CLK(CLK), .D(_01012_), .Q(__stream_matmul_29_sink_21_sink_size_1_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_1_reg  ( .CLK(CLK), .D(_00725_), .Q(__set_flag_1224_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_2_reg  ( .CLK(CLK), .D(_00736_), .Q(__set_flag_1224_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_3_reg  ( .CLK(CLK), .D(_00747_), .Q(__set_flag_1224_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_4_reg  ( .CLK(CLK), .D(_00750_), .Q(__set_flag_1224_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_5_reg  ( .CLK(CLK), .D(_00751_), .Q(__set_flag_1224_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_6_reg  ( .CLK(CLK), .D(_00752_), .Q(__set_flag_1224_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_7_reg  ( .CLK(CLK), .D(_00753_), .Q(__set_flag_1224_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_8_reg  ( .CLK(CLK), .D(_00754_), .Q(__set_flag_1224_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_9_reg  ( .CLK(CLK), .D(_00755_), .Q(__set_flag_1224_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_10_reg  ( .CLK(CLK), .D(_00715_), .Q(__set_flag_1224_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_11_reg  ( .CLK(CLK), .D(_00716_), .Q(__set_flag_1224_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_12_reg  ( .CLK(CLK), .D(_00717_), .Q(__set_flag_1224_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_13_reg  ( .CLK(CLK), .D(_00718_), .Q(__set_flag_1224_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_14_reg  ( .CLK(CLK), .D(_00719_), .Q(__set_flag_1224_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_15_reg  ( .CLK(CLK), .D(_00720_), .Q(__set_flag_1224_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_16_reg  ( .CLK(CLK), .D(_00721_), .Q(__set_flag_1224_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_17_reg  ( .CLK(CLK), .D(_00722_), .Q(__set_flag_1224_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_18_reg  ( .CLK(CLK), .D(_00723_), .Q(__set_flag_1224_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_19_reg  ( .CLK(CLK), .D(_00724_), .Q(__set_flag_1224_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_20_reg  ( .CLK(CLK), .D(_00726_), .Q(__set_flag_1224_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_21_reg  ( .CLK(CLK), .D(_00727_), .Q(__set_flag_1224_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_22_reg  ( .CLK(CLK), .D(_00728_), .Q(__set_flag_1224_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_23_reg  ( .CLK(CLK), .D(_00729_), .Q(__set_flag_1224_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_24_reg  ( .CLK(CLK), .D(_00730_), .Q(__set_flag_1224_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_25_reg  ( .CLK(CLK), .D(_00731_), .Q(__set_flag_1224_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_26_reg  ( .CLK(CLK), .D(_00732_), .Q(__set_flag_1224_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_27_reg  ( .CLK(CLK), .D(_00733_), .Q(__set_flag_1224_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_28_reg  ( .CLK(CLK), .D(_00734_), .Q(__set_flag_1224_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_29_reg  ( .CLK(CLK), .D(_00735_), .Q(__set_flag_1224_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_30_reg  ( .CLK(CLK), .D(_00737_), .Q(__set_flag_1224_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_31_reg  ( .CLK(CLK), .D(_00738_), .Q(__set_flag_1224_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_32_reg  ( .CLK(CLK), .D(_00739_), .Q(__set_flag_1224_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_33_reg  ( .CLK(CLK), .D(_00740_), .Q(__set_flag_1224_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_34_reg  ( .CLK(CLK), .D(_00741_), .Q(__set_flag_1224_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_35_reg  ( .CLK(CLK), .D(_00742_), .Q(__set_flag_1224_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_36_reg  ( .CLK(CLK), .D(_00743_), .Q(__set_flag_1224_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_37_reg  ( .CLK(CLK), .D(_00744_), .Q(__set_flag_1224_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_38_reg  ( .CLK(CLK), .D(_00745_), .Q(__set_flag_1224_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_39_reg  ( .CLK(CLK), .D(_00746_), .Q(__set_flag_1224_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_40_reg  ( .CLK(CLK), .D(_00748_), .Q(__set_flag_1224_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1224_41_reg  ( .CLK(CLK), .D(_00749_), .Q(__set_flag_1224_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_1_reg  ( .CLK(CLK), .D(_01029_), .Q(__stream_matmul_29_start_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_2_reg  ( .CLK(CLK), .D(_01040_), .Q(__stream_matmul_29_start_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_3_reg  ( .CLK(CLK), .D(_01051_), .Q(__stream_matmul_29_start_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_4_reg  ( .CLK(CLK), .D(_01055_), .Q(__stream_matmul_29_start_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_5_reg  ( .CLK(CLK), .D(_01056_), .Q(__stream_matmul_29_start_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_6_reg  ( .CLK(CLK), .D(_01057_), .Q(__stream_matmul_29_start_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_7_reg  ( .CLK(CLK), .D(_01058_), .Q(__stream_matmul_29_start_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_8_reg  ( .CLK(CLK), .D(_01059_), .Q(__stream_matmul_29_start_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_9_reg  ( .CLK(CLK), .D(_01060_), .Q(__stream_matmul_29_start_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_10_reg  ( .CLK(CLK), .D(_01019_), .Q(__stream_matmul_29_start_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_11_reg  ( .CLK(CLK), .D(_01020_), .Q(__stream_matmul_29_start_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_12_reg  ( .CLK(CLK), .D(_01021_), .Q(__stream_matmul_29_start_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_13_reg  ( .CLK(CLK), .D(_01022_), .Q(__stream_matmul_29_start_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_14_reg  ( .CLK(CLK), .D(_01023_), .Q(__stream_matmul_29_start_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_15_reg  ( .CLK(CLK), .D(_01024_), .Q(__stream_matmul_29_start_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_16_reg  ( .CLK(CLK), .D(_01025_), .Q(__stream_matmul_29_start_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_17_reg  ( .CLK(CLK), .D(_01026_), .Q(__stream_matmul_29_start_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_18_reg  ( .CLK(CLK), .D(_01027_), .Q(__stream_matmul_29_start_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_19_reg  ( .CLK(CLK), .D(_01028_), .Q(__stream_matmul_29_start_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_20_reg  ( .CLK(CLK), .D(_01030_), .Q(__stream_matmul_29_start_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_21_reg  ( .CLK(CLK), .D(_01031_), .Q(__stream_matmul_29_start_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_22_reg  ( .CLK(CLK), .D(_01032_), .Q(__stream_matmul_29_start_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_23_reg  ( .CLK(CLK), .D(_01033_), .Q(__stream_matmul_29_start_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_24_reg  ( .CLK(CLK), .D(_01034_), .Q(__stream_matmul_29_start_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_25_reg  ( .CLK(CLK), .D(_01035_), .Q(__stream_matmul_29_start_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_26_reg  ( .CLK(CLK), .D(_01036_), .Q(__stream_matmul_29_start_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_27_reg  ( .CLK(CLK), .D(_01037_), .Q(__stream_matmul_29_start_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_28_reg  ( .CLK(CLK), .D(_01038_), .Q(__stream_matmul_29_start_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_29_reg  ( .CLK(CLK), .D(_01039_), .Q(__stream_matmul_29_start_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_30_reg  ( .CLK(CLK), .D(_01041_), .Q(__stream_matmul_29_start_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_31_reg  ( .CLK(CLK), .D(_01042_), .Q(__stream_matmul_29_start_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_32_reg  ( .CLK(CLK), .D(_01043_), .Q(__stream_matmul_29_start_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_33_reg  ( .CLK(CLK), .D(_01044_), .Q(__stream_matmul_29_start_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_34_reg  ( .CLK(CLK), .D(_01045_), .Q(__stream_matmul_29_start_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_35_reg  ( .CLK(CLK), .D(_01046_), .Q(__stream_matmul_29_start_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_36_reg  ( .CLK(CLK), .D(_01047_), .Q(__stream_matmul_29_start_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_37_reg  ( .CLK(CLK), .D(_01048_), .Q(__stream_matmul_29_start_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_38_reg  ( .CLK(CLK), .D(_01049_), .Q(__stream_matmul_29_start_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_39_reg  ( .CLK(CLK), .D(_01050_), .Q(__stream_matmul_29_start_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_40_reg  ( .CLK(CLK), .D(_01052_), .Q(__stream_matmul_29_start_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_41_reg  ( .CLK(CLK), .D(_01053_), .Q(__stream_matmul_29_start_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_matmul_29_start_42_reg  ( .CLK(CLK), .D(_01054_), .Q(__stream_matmul_29_start_42) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_1_reg  ( .CLK(CLK), .D(_01151_), .Q(__tmp_1249_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_2_reg  ( .CLK(CLK), .D(_01152_), .Q(__tmp_1249_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_3_reg  ( .CLK(CLK), .D(_01153_), .Q(__tmp_1249_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_4_reg  ( .CLK(CLK), .D(_01154_), .Q(__tmp_1249_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_5_reg  ( .CLK(CLK), .D(_01155_), .Q(__tmp_1249_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_6_reg  ( .CLK(CLK), .D(_01156_), .Q(__tmp_1249_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_7_reg  ( .CLK(CLK), .D(_01157_), .Q(__tmp_1249_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_8_reg  ( .CLK(CLK), .D(_01158_), .Q(__tmp_1249_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_9_reg  ( .CLK(CLK), .D(_01168_), .Q(__tmp_1249_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_10_reg  ( .CLK(CLK), .D(_01159_), .Q(__tmp_1249_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_11_reg  ( .CLK(CLK), .D(_01160_), .Q(__tmp_1249_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_12_reg  ( .CLK(CLK), .D(_01161_), .Q(__tmp_1249_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_13_reg  ( .CLK(CLK), .D(_01162_), .Q(__tmp_1249_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_14_reg  ( .CLK(CLK), .D(_01163_), .Q(__tmp_1249_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_15_reg  ( .CLK(CLK), .D(_01164_), .Q(__tmp_1249_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_16_reg  ( .CLK(CLK), .D(_01165_), .Q(__tmp_1249_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_17_reg  ( .CLK(CLK), .D(_01166_), .Q(__tmp_1249_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_18_reg  ( .CLK(CLK), .D(_01167_), .Q(__tmp_1249_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_19_reg  ( .CLK(CLK), .D(_01169_), .Q(__tmp_1249_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_20_reg  ( .CLK(CLK), .D(_01170_), .Q(__tmp_1249_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_21_reg  ( .CLK(CLK), .D(_01171_), .Q(__tmp_1249_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_22_reg  ( .CLK(CLK), .D(_01172_), .Q(__tmp_1249_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_23_reg  ( .CLK(CLK), .D(_01173_), .Q(__tmp_1249_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_24_reg  ( .CLK(CLK), .D(_01174_), .Q(__tmp_1249_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_25_reg  ( .CLK(CLK), .D(_01175_), .Q(__tmp_1249_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_26_reg  ( .CLK(CLK), .D(_01176_), .Q(__tmp_1249_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_27_reg  ( .CLK(CLK), .D(_01177_), .Q(__tmp_1249_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1249_28_reg  ( .CLK(CLK), .D(_01178_), .Q(__tmp_1249_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1291_20_reg  ( .CLK(CLK), .D(_01198_), .Q(__tmp_1291_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1291_21_reg  ( .CLK(CLK), .D(_01199_), .Q(__tmp_1291_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1291_22_reg  ( .CLK(CLK), .D(_01200_), .Q(__tmp_1291_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1291_23_reg  ( .CLK(CLK), .D(_01201_), .Q(__tmp_1291_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1291_24_reg  ( .CLK(CLK), .D(_01202_), .Q(__tmp_1291_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1291_25_reg  ( .CLK(CLK), .D(_01203_), .Q(__tmp_1291_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_1_reg  ( .CLK(CLK), .D(_01179_), .Q(__tmp_1299_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_2_reg  ( .CLK(CLK), .D(_01180_), .Q(__tmp_1299_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_3_reg  ( .CLK(CLK), .D(_01181_), .Q(__tmp_1299_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_4_reg  ( .CLK(CLK), .D(_01182_), .Q(__tmp_1299_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_5_reg  ( .CLK(CLK), .D(_01183_), .Q(__tmp_1299_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_6_reg  ( .CLK(CLK), .D(_01187_), .Q(__tmp_1299_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_7_reg  ( .CLK(CLK), .D(_01188_), .Q(__tmp_1299_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_8_reg  ( .CLK(CLK), .D(_01189_), .Q(__tmp_1299_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_9_reg  ( .CLK(CLK), .D(_01190_), .Q(__tmp_1299_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_10_reg  ( .CLK(CLK), .D(_01184_), .Q(__tmp_1299_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_11_reg  ( .CLK(CLK), .D(_01185_), .Q(__tmp_1299_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_12_reg  ( .CLK(CLK), .D(_01186_), .Q(__tmp_1299_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_13_reg  ( .CLK(CLK), .D(_01191_), .Q(__tmp_1299_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_14_reg  ( .CLK(CLK), .D(_01192_), .Q(__tmp_1299_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_15_reg  ( .CLK(CLK), .D(_01193_), .Q(__tmp_1299_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_16_reg  ( .CLK(CLK), .D(_01194_), .Q(__tmp_1299_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_17_reg  ( .CLK(CLK), .D(_01195_), .Q(__tmp_1299_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_18_reg  ( .CLK(CLK), .D(_01196_), .Q(__tmp_1299_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1299_19_reg  ( .CLK(CLK), .D(_01197_), .Q(__tmp_1299_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1305_39_reg  ( .CLK(CLK), .D(_01217_), .Q(__tmp_1305_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1305_40_reg  ( .CLK(CLK), .D(_01218_), .Q(__tmp_1305_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1305_41_reg  ( .CLK(CLK), .D(_01219_), .Q(__tmp_1305_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1305_42_reg  ( .CLK(CLK), .D(_01220_), .Q(__tmp_1305_42) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_26_reg  ( .CLK(CLK), .D(_01204_), .Q(__tmp_1307_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_27_reg  ( .CLK(CLK), .D(_01205_), .Q(__tmp_1307_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_28_reg  ( .CLK(CLK), .D(_01206_), .Q(__tmp_1307_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_29_reg  ( .CLK(CLK), .D(_01207_), .Q(__tmp_1307_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_30_reg  ( .CLK(CLK), .D(_01208_), .Q(__tmp_1307_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_31_reg  ( .CLK(CLK), .D(_01209_), .Q(__tmp_1307_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_32_reg  ( .CLK(CLK), .D(_01210_), .Q(__tmp_1307_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_33_reg  ( .CLK(CLK), .D(_01211_), .Q(__tmp_1307_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_34_reg  ( .CLK(CLK), .D(_01212_), .Q(__tmp_1307_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_35_reg  ( .CLK(CLK), .D(_01213_), .Q(__tmp_1307_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_36_reg  ( .CLK(CLK), .D(_01214_), .Q(__tmp_1307_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_37_reg  ( .CLK(CLK), .D(_01215_), .Q(__tmp_1307_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1307_38_reg  ( .CLK(CLK), .D(_01216_), .Q(__tmp_1307_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42701_ ( .CLK(CLK), .D(_02773_), .Q(_stream_max_pool_serial_18_fsm) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_max_pool_serial_18_start_reg  ( .CLK(CLK), .D(_02796_), .Q(_stream_max_pool_serial_18_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_max_pool_serial_18_end_flag_reg  ( .CLK(CLK), .D(_02772_), .Q(_stream_max_pool_serial_18_end_flag) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_max_pool_serial_18_term_sink_reg  ( .CLK(CLK), .D(_02797_), .Q(_stream_max_pool_serial_18_term_sink) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_max_pool_serial_18_source_busy_reg  ( .CLK(CLK), .D(_02795_), .Q(_stream_max_pool_serial_18_source_busy) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_max_pool_serial_18_reduce_reset_reg  ( .CLK(CLK), .D(_02774_), .Q(_stream_max_pool_serial_18_reduce_reset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42707_ ( .CLK(CLK), .D(_02770_), .Q(_stream_max_pool_serial_18_constant_0_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_max_pool_serial_18_source_1_idle_reg  ( .CLK(CLK), .D(_02786_), .Q(_stream_max_pool_serial_18_source_1_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42709_ ( .CLK(CLK), .D(_02787_), .Q(_stream_max_pool_serial_18_source_1_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42710_ ( .CLK(CLK), .D(_02788_), .Q(_stream_max_pool_serial_18_source_1_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42711_ ( .CLK(CLK), .D(_02789_), .Q(_stream_max_pool_serial_18_source_1_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42712_ ( .CLK(CLK), .D(_02794_), .Q(_stream_max_pool_serial_18_source_1_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42713_ ( .CLK(CLK), .D(_02791_), .Q(_stream_max_pool_serial_18_source_1_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_max_pool_serial_18_source_1_source_ram_renable_reg  ( .CLK(CLK), .D(_02792_), .Q(_stream_max_pool_serial_18_source_1_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_max_pool_serial_18_source_1_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02793_), .Q(_stream_max_pool_serial_18_source_1_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _42716_ ( .CLK(CLK), .D(_02771_), .Q(_stream_max_pool_serial_18_constant_2_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42717_ ( .CLK(CLK), .D(_02777_), .Q(_stream_max_pool_serial_18_sink_3_sink_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42718_ ( .CLK(CLK), .D(_02778_), .Q(_stream_max_pool_serial_18_sink_3_sink_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42719_ ( .CLK(CLK), .D(_02780_), .Q(_stream_max_pool_serial_18_sink_3_sink_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42720_ ( .CLK(CLK), .D(_02781_), .Q(_stream_max_pool_serial_18_sink_3_sink_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42721_ ( .CLK(CLK), .D(_02775_), .Q(_stream_max_pool_serial_18_sink_3_sink_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42722_ ( .CLK(CLK), .D(_02782_), .Q(_stream_max_pool_serial_18_sink_3_sink_stride_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42723_ ( .CLK(CLK), .D(_02779_), .Q(_stream_max_pool_serial_18_sink_3_sink_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42724_ ( .CLK(CLK), .D(_02783_), .Q(_stream_max_pool_serial_18_sink_3_sink_waddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_max_pool_serial_18_sink_3_sink_wenable_reg  ( .CLK(CLK), .D(_02785_), .Q(_stream_max_pool_serial_18_sink_3_sink_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42726_ ( .CLK(CLK), .D(_02784_), .Q(_stream_max_pool_serial_18_sink_3_sink_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42727_ ( .CLK(CLK), .D(_01580_), .Q(_counter_data_782) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42728_ ( .CLK(CLK), .D(_01579_), .Q(_counter_count_782) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _42729_ ( .CLK(CLK), .D(_00292_), .Q(__delay_data_1411) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42730_ ( .CLK(CLK), .D(_00293_), .Q(__delay_data_1412) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42731_ ( .CLK(CLK), .D(_00295_), .Q(__delay_data_1414) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _pointer_data_784_reg  ( .CLK(CLK), .D(_01819_), .Q(_pointer_data_784) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42733_ ( .CLK(CLK), .D(_00294_), .Q(__delay_data_1413) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42734_ ( .CLK(CLK), .D(_00296_), .Q(__delay_data_1415) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _42735_ ( .CLK(CLK), .D(_01548_), .Q(_cond_data_791) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42736_ ( .CLK(CLK), .D(_00297_), .Q(__delay_data_1416) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42737_ ( .CLK(CLK), .D(_01102_), .Q(__substreamoutput_data_793) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __substreamoutput_data_794_reg  ( .CLK(CLK), .D(_01103_), .Q(__substreamoutput_data_794) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42739_ ( .CLK(CLK), .D(_01445_), .Q(__variable_wdata_777) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _42740_ ( .CLK(CLK), .D(_01447_), .Q(__variable_wdata_779) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42741_ ( .CLK(CLK), .D(_02464_), .Q(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42742_ ( .CLK(CLK), .D(_02465_), .Q(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42743_ ( .CLK(CLK), .D(_02466_), .Q(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42744_ ( .CLK(CLK), .D(_02467_), .Q(_source_stream_max_pool_serial_18_source_1_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42745_ ( .CLK(CLK), .D(_02468_), .Q(_source_stream_max_pool_serial_18_source_1_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42746_ ( .CLK(CLK), .D(_02469_), .Q(_source_stream_max_pool_serial_18_source_1_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42747_ ( .CLK(CLK), .D(_02470_), .Q(_source_stream_max_pool_serial_18_source_1_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42748_ ( .CLK(CLK), .D(_02471_), .Q(_source_stream_max_pool_serial_18_source_1_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42749_ ( .CLK(CLK), .D(_02476_), .Q(_source_stream_max_pool_serial_18_source_1_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42750_ ( .CLK(CLK), .D(_02477_), .Q(_source_stream_max_pool_serial_18_source_1_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42751_ ( .CLK(CLK), .D(_02478_), .Q(_source_stream_max_pool_serial_18_source_1_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42752_ ( .CLK(CLK), .D(_02479_), .Q(_source_stream_max_pool_serial_18_source_1_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42753_ ( .CLK(CLK), .D(_02460_), .Q(_source_stream_max_pool_serial_18_source_1_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42754_ ( .CLK(CLK), .D(_02461_), .Q(_source_stream_max_pool_serial_18_source_1_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42755_ ( .CLK(CLK), .D(_02462_), .Q(_source_stream_max_pool_serial_18_source_1_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42756_ ( .CLK(CLK), .D(_02463_), .Q(_source_stream_max_pool_serial_18_source_1_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42757_ ( .CLK(CLK), .D(_02472_), .Q(_source_stream_max_pool_serial_18_source_1_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42758_ ( .CLK(CLK), .D(_02473_), .Q(_source_stream_max_pool_serial_18_source_1_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42759_ ( .CLK(CLK), .D(_02474_), .Q(_source_stream_max_pool_serial_18_source_1_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42760_ ( .CLK(CLK), .D(_02475_), .Q(_source_stream_max_pool_serial_18_source_1_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42761_ ( .CLK(CLK), .D(_02480_), .Q(_source_stream_max_pool_serial_18_source_1_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42762_ ( .CLK(CLK), .D(_02481_), .Q(_source_stream_max_pool_serial_18_source_1_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42763_ ( .CLK(CLK), .D(_02482_), .Q(_source_stream_max_pool_serial_18_source_1_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42764_ ( .CLK(CLK), .D(_02483_), .Q(_source_stream_max_pool_serial_18_source_1_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42765_ ( .CLK(CLK), .D(_01446_), .Q(__variable_wdata_778) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _set_flag_1036_reg  ( .CLK(CLK), .D(_01870_), .Q(_set_flag_1036) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42767_ ( .CLK(CLK), .D(_01061_), .Q(__stream_max_pool_serial_18_sink_3_sink_offset_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42768_ ( .CLK(CLK), .D(_01062_), .Q(__stream_max_pool_serial_18_sink_3_sink_offset_0_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42769_ ( .CLK(CLK), .D(_01063_), .Q(__stream_max_pool_serial_18_sink_3_sink_offset_0_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42770_ ( .CLK(CLK), .D(_01064_), .Q(__stream_max_pool_serial_18_sink_3_sink_offset_0_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42771_ ( .CLK(CLK), .D(_01065_), .Q(__stream_max_pool_serial_18_sink_3_sink_offset_0_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42772_ ( .CLK(CLK), .D(_01066_), .Q(__stream_max_pool_serial_18_sink_3_sink_offset_0_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42773_ ( .CLK(CLK), .D(_01067_), .Q(__stream_max_pool_serial_18_sink_3_sink_offset_0_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42774_ ( .CLK(CLK), .D(_01068_), .Q(__stream_max_pool_serial_18_sink_3_sink_offset_0_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42775_ ( .CLK(CLK), .D(_01069_), .Q(__stream_max_pool_serial_18_sink_3_sink_offset_0_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42776_ ( .CLK(CLK), .D(_01070_), .Q(__stream_max_pool_serial_18_sink_3_sink_size_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42777_ ( .CLK(CLK), .D(_01071_), .Q(__stream_max_pool_serial_18_sink_3_sink_size_1_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42778_ ( .CLK(CLK), .D(_01072_), .Q(__stream_max_pool_serial_18_sink_3_sink_size_1_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42779_ ( .CLK(CLK), .D(_01073_), .Q(__stream_max_pool_serial_18_sink_3_sink_size_1_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42780_ ( .CLK(CLK), .D(_01074_), .Q(__stream_max_pool_serial_18_sink_3_sink_size_1_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42781_ ( .CLK(CLK), .D(_01075_), .Q(__stream_max_pool_serial_18_sink_3_sink_size_1_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42782_ ( .CLK(CLK), .D(_01076_), .Q(__stream_max_pool_serial_18_sink_3_sink_size_1_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42783_ ( .CLK(CLK), .D(_01077_), .Q(__stream_max_pool_serial_18_sink_3_sink_size_1_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42784_ ( .CLK(CLK), .D(_01078_), .Q(__stream_max_pool_serial_18_sink_3_sink_size_1_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1036_1_reg  ( .CLK(CLK), .D(_00706_), .Q(__set_flag_1036_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1036_2_reg  ( .CLK(CLK), .D(_00707_), .Q(__set_flag_1036_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1036_3_reg  ( .CLK(CLK), .D(_00708_), .Q(__set_flag_1036_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1036_4_reg  ( .CLK(CLK), .D(_00709_), .Q(__set_flag_1036_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1036_5_reg  ( .CLK(CLK), .D(_00710_), .Q(__set_flag_1036_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1036_6_reg  ( .CLK(CLK), .D(_00711_), .Q(__set_flag_1036_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1036_7_reg  ( .CLK(CLK), .D(_00712_), .Q(__set_flag_1036_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1036_8_reg  ( .CLK(CLK), .D(_00713_), .Q(__set_flag_1036_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_1036_9_reg  ( .CLK(CLK), .D(_00714_), .Q(__set_flag_1036_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_max_pool_serial_18_start_1_reg  ( .CLK(CLK), .D(_01080_), .Q(__stream_max_pool_serial_18_start_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_max_pool_serial_18_start_2_reg  ( .CLK(CLK), .D(_01081_), .Q(__stream_max_pool_serial_18_start_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_max_pool_serial_18_start_3_reg  ( .CLK(CLK), .D(_01082_), .Q(__stream_max_pool_serial_18_start_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_max_pool_serial_18_start_4_reg  ( .CLK(CLK), .D(_01083_), .Q(__stream_max_pool_serial_18_start_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_max_pool_serial_18_start_5_reg  ( .CLK(CLK), .D(_01084_), .Q(__stream_max_pool_serial_18_start_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_max_pool_serial_18_start_6_reg  ( .CLK(CLK), .D(_01085_), .Q(__stream_max_pool_serial_18_start_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_max_pool_serial_18_start_7_reg  ( .CLK(CLK), .D(_01086_), .Q(__stream_max_pool_serial_18_start_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_max_pool_serial_18_start_8_reg  ( .CLK(CLK), .D(_01087_), .Q(__stream_max_pool_serial_18_start_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_max_pool_serial_18_start_9_reg  ( .CLK(CLK), .D(_01088_), .Q(__stream_max_pool_serial_18_start_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_max_pool_serial_18_start_10_reg  ( .CLK(CLK), .D(_01079_), .Q(__stream_max_pool_serial_18_start_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _set_flag_1038_reg  ( .CLK(CLK), .D(_01871_), .Q(_set_flag_1038) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1042_8_reg  ( .CLK(CLK), .D(_01119_), .Q(__tmp_1042_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1042_9_reg  ( .CLK(CLK), .D(_01120_), .Q(__tmp_1042_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1046_1_reg  ( .CLK(CLK), .D(_01112_), .Q(__tmp_1046_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1046_2_reg  ( .CLK(CLK), .D(_01113_), .Q(__tmp_1046_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1046_3_reg  ( .CLK(CLK), .D(_01114_), .Q(__tmp_1046_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1046_4_reg  ( .CLK(CLK), .D(_01115_), .Q(__tmp_1046_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1046_5_reg  ( .CLK(CLK), .D(_01116_), .Q(__tmp_1046_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1046_6_reg  ( .CLK(CLK), .D(_01117_), .Q(__tmp_1046_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1046_7_reg  ( .CLK(CLK), .D(_01118_), .Q(__tmp_1046_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1068_7_reg  ( .CLK(CLK), .D(_01128_), .Q(__tmp_1068_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1068_8_reg  ( .CLK(CLK), .D(_01129_), .Q(__tmp_1068_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1068_9_reg  ( .CLK(CLK), .D(_01130_), .Q(__tmp_1068_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1068_10_reg  ( .CLK(CLK), .D(_01126_), .Q(__tmp_1068_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1070_6_reg  ( .CLK(CLK), .D(_01127_), .Q(__tmp_1070_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42819_ ( .CLK(CLK), .D(_02503_), .Q(_stream_conv2d_16_fsm) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_start_reg  ( .CLK(CLK), .D(_02702_), .Q(_stream_conv2d_16_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_end_flag_reg  ( .CLK(CLK), .D(_02502_), .Q(_stream_conv2d_16_end_flag) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_term_sink_reg  ( .CLK(CLK), .D(_02703_), .Q(_stream_conv2d_16_term_sink) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_busy_reg  ( .CLK(CLK), .D(_02701_), .Q(_stream_conv2d_16_source_busy) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _42824_ ( .CLK(CLK), .D(_02495_), .Q(_stream_conv2d_16_constant_0_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _42825_ ( .CLK(CLK), .D(_02499_), .Q(_stream_conv2d_16_constant_1_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _42826_ ( .CLK(CLK), .D(_02500_), .Q(_stream_conv2d_16_constant_2_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _42827_ ( .CLK(CLK), .D(_02501_), .Q(_stream_conv2d_16_constant_3_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_6_idle_reg  ( .CLK(CLK), .D(_02683_), .Q(_stream_conv2d_16_source_6_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42829_ ( .CLK(CLK), .D(_02684_), .Q(_stream_conv2d_16_source_6_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42830_ ( .CLK(CLK), .D(_02685_), .Q(_stream_conv2d_16_source_6_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42831_ ( .CLK(CLK), .D(_02686_), .Q(_stream_conv2d_16_source_6_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42832_ ( .CLK(CLK), .D(_02691_), .Q(_stream_conv2d_16_source_6_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42833_ ( .CLK(CLK), .D(_02688_), .Q(_stream_conv2d_16_source_6_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_6_source_ram_renable_reg  ( .CLK(CLK), .D(_02689_), .Q(_stream_conv2d_16_source_6_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_6_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02690_), .Q(_stream_conv2d_16_source_6_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_8_idle_reg  ( .CLK(CLK), .D(_02692_), .Q(_stream_conv2d_16_source_8_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42837_ ( .CLK(CLK), .D(_02693_), .Q(_stream_conv2d_16_source_8_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42838_ ( .CLK(CLK), .D(_02694_), .Q(_stream_conv2d_16_source_8_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42839_ ( .CLK(CLK), .D(_02695_), .Q(_stream_conv2d_16_source_8_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42840_ ( .CLK(CLK), .D(_02700_), .Q(_stream_conv2d_16_source_8_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42841_ ( .CLK(CLK), .D(_02697_), .Q(_stream_conv2d_16_source_8_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_8_source_ram_renable_reg  ( .CLK(CLK), .D(_02698_), .Q(_stream_conv2d_16_source_8_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_8_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02699_), .Q(_stream_conv2d_16_source_8_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_10_idle_reg  ( .CLK(CLK), .D(_02515_), .Q(_stream_conv2d_16_source_10_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42845_ ( .CLK(CLK), .D(_02516_), .Q(_stream_conv2d_16_source_10_source_empty_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_12_idle_reg  ( .CLK(CLK), .D(_02517_), .Q(_stream_conv2d_16_source_12_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42847_ ( .CLK(CLK), .D(_02518_), .Q(_stream_conv2d_16_source_12_source_empty_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_14_idle_reg  ( .CLK(CLK), .D(_02519_), .Q(_stream_conv2d_16_source_14_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42849_ ( .CLK(CLK), .D(_02520_), .Q(_stream_conv2d_16_source_14_source_empty_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_constant_15_next_constant_data_reg  ( .CLK(CLK), .D(_02496_), .Q(_stream_conv2d_16_constant_15_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_constant_16_next_constant_data_reg  ( .CLK(CLK), .D(_02497_), .Q(_stream_conv2d_16_constant_16_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _42852_ ( .CLK(CLK), .D(_02498_), .Q(_stream_conv2d_16_constant_17_next_constant_data) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_19_idle_reg  ( .CLK(CLK), .D(_02521_), .Q(_stream_conv2d_16_source_19_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42854_ ( .CLK(CLK), .D(_02522_), .Q(_stream_conv2d_16_source_19_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42855_ ( .CLK(CLK), .D(_02523_), .Q(_stream_conv2d_16_source_19_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42856_ ( .CLK(CLK), .D(_02524_), .Q(_stream_conv2d_16_source_19_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42857_ ( .CLK(CLK), .D(_02529_), .Q(_stream_conv2d_16_source_19_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42858_ ( .CLK(CLK), .D(_02526_), .Q(_stream_conv2d_16_source_19_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_19_source_ram_renable_reg  ( .CLK(CLK), .D(_02527_), .Q(_stream_conv2d_16_source_19_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_19_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02528_), .Q(_stream_conv2d_16_source_19_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_20_idle_reg  ( .CLK(CLK), .D(_02530_), .Q(_stream_conv2d_16_source_20_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42862_ ( .CLK(CLK), .D(_02531_), .Q(_stream_conv2d_16_source_20_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42863_ ( .CLK(CLK), .D(_02532_), .Q(_stream_conv2d_16_source_20_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42864_ ( .CLK(CLK), .D(_02533_), .Q(_stream_conv2d_16_source_20_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42865_ ( .CLK(CLK), .D(_02538_), .Q(_stream_conv2d_16_source_20_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42866_ ( .CLK(CLK), .D(_02535_), .Q(_stream_conv2d_16_source_20_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_20_source_ram_renable_reg  ( .CLK(CLK), .D(_02536_), .Q(_stream_conv2d_16_source_20_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_20_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02537_), .Q(_stream_conv2d_16_source_20_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_21_idle_reg  ( .CLK(CLK), .D(_02539_), .Q(_stream_conv2d_16_source_21_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42870_ ( .CLK(CLK), .D(_02540_), .Q(_stream_conv2d_16_source_21_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42871_ ( .CLK(CLK), .D(_02541_), .Q(_stream_conv2d_16_source_21_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42872_ ( .CLK(CLK), .D(_02542_), .Q(_stream_conv2d_16_source_21_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42873_ ( .CLK(CLK), .D(_02547_), .Q(_stream_conv2d_16_source_21_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42874_ ( .CLK(CLK), .D(_02544_), .Q(_stream_conv2d_16_source_21_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_21_source_ram_renable_reg  ( .CLK(CLK), .D(_02545_), .Q(_stream_conv2d_16_source_21_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_21_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02546_), .Q(_stream_conv2d_16_source_21_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_22_idle_reg  ( .CLK(CLK), .D(_02548_), .Q(_stream_conv2d_16_source_22_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42878_ ( .CLK(CLK), .D(_02549_), .Q(_stream_conv2d_16_source_22_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42879_ ( .CLK(CLK), .D(_02550_), .Q(_stream_conv2d_16_source_22_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42880_ ( .CLK(CLK), .D(_02551_), .Q(_stream_conv2d_16_source_22_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42881_ ( .CLK(CLK), .D(_02556_), .Q(_stream_conv2d_16_source_22_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42882_ ( .CLK(CLK), .D(_02553_), .Q(_stream_conv2d_16_source_22_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_22_source_ram_renable_reg  ( .CLK(CLK), .D(_02554_), .Q(_stream_conv2d_16_source_22_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_22_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02555_), .Q(_stream_conv2d_16_source_22_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_23_idle_reg  ( .CLK(CLK), .D(_02557_), .Q(_stream_conv2d_16_source_23_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42886_ ( .CLK(CLK), .D(_02558_), .Q(_stream_conv2d_16_source_23_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42887_ ( .CLK(CLK), .D(_02559_), .Q(_stream_conv2d_16_source_23_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42888_ ( .CLK(CLK), .D(_02560_), .Q(_stream_conv2d_16_source_23_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42889_ ( .CLK(CLK), .D(_02565_), .Q(_stream_conv2d_16_source_23_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42890_ ( .CLK(CLK), .D(_02562_), .Q(_stream_conv2d_16_source_23_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_23_source_ram_renable_reg  ( .CLK(CLK), .D(_02563_), .Q(_stream_conv2d_16_source_23_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_23_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02564_), .Q(_stream_conv2d_16_source_23_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_24_idle_reg  ( .CLK(CLK), .D(_02566_), .Q(_stream_conv2d_16_source_24_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42894_ ( .CLK(CLK), .D(_02567_), .Q(_stream_conv2d_16_source_24_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42895_ ( .CLK(CLK), .D(_02568_), .Q(_stream_conv2d_16_source_24_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42896_ ( .CLK(CLK), .D(_02569_), .Q(_stream_conv2d_16_source_24_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42897_ ( .CLK(CLK), .D(_02574_), .Q(_stream_conv2d_16_source_24_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42898_ ( .CLK(CLK), .D(_02571_), .Q(_stream_conv2d_16_source_24_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_24_source_ram_renable_reg  ( .CLK(CLK), .D(_02572_), .Q(_stream_conv2d_16_source_24_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_24_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02573_), .Q(_stream_conv2d_16_source_24_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_25_idle_reg  ( .CLK(CLK), .D(_02575_), .Q(_stream_conv2d_16_source_25_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42902_ ( .CLK(CLK), .D(_02576_), .Q(_stream_conv2d_16_source_25_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42903_ ( .CLK(CLK), .D(_02577_), .Q(_stream_conv2d_16_source_25_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42904_ ( .CLK(CLK), .D(_02578_), .Q(_stream_conv2d_16_source_25_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42905_ ( .CLK(CLK), .D(_02583_), .Q(_stream_conv2d_16_source_25_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42906_ ( .CLK(CLK), .D(_02580_), .Q(_stream_conv2d_16_source_25_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_25_source_ram_renable_reg  ( .CLK(CLK), .D(_02581_), .Q(_stream_conv2d_16_source_25_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_25_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02582_), .Q(_stream_conv2d_16_source_25_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_26_idle_reg  ( .CLK(CLK), .D(_02584_), .Q(_stream_conv2d_16_source_26_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42910_ ( .CLK(CLK), .D(_02585_), .Q(_stream_conv2d_16_source_26_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42911_ ( .CLK(CLK), .D(_02586_), .Q(_stream_conv2d_16_source_26_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42912_ ( .CLK(CLK), .D(_02587_), .Q(_stream_conv2d_16_source_26_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42913_ ( .CLK(CLK), .D(_02592_), .Q(_stream_conv2d_16_source_26_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42914_ ( .CLK(CLK), .D(_02589_), .Q(_stream_conv2d_16_source_26_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_26_source_ram_renable_reg  ( .CLK(CLK), .D(_02590_), .Q(_stream_conv2d_16_source_26_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_26_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02591_), .Q(_stream_conv2d_16_source_26_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_27_idle_reg  ( .CLK(CLK), .D(_02593_), .Q(_stream_conv2d_16_source_27_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42918_ ( .CLK(CLK), .D(_02594_), .Q(_stream_conv2d_16_source_27_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42919_ ( .CLK(CLK), .D(_02595_), .Q(_stream_conv2d_16_source_27_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42920_ ( .CLK(CLK), .D(_02596_), .Q(_stream_conv2d_16_source_27_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42921_ ( .CLK(CLK), .D(_02601_), .Q(_stream_conv2d_16_source_27_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42922_ ( .CLK(CLK), .D(_02598_), .Q(_stream_conv2d_16_source_27_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_27_source_ram_renable_reg  ( .CLK(CLK), .D(_02599_), .Q(_stream_conv2d_16_source_27_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_27_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02600_), .Q(_stream_conv2d_16_source_27_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_28_idle_reg  ( .CLK(CLK), .D(_02602_), .Q(_stream_conv2d_16_source_28_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42926_ ( .CLK(CLK), .D(_02603_), .Q(_stream_conv2d_16_source_28_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42927_ ( .CLK(CLK), .D(_02604_), .Q(_stream_conv2d_16_source_28_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42928_ ( .CLK(CLK), .D(_02605_), .Q(_stream_conv2d_16_source_28_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42929_ ( .CLK(CLK), .D(_02610_), .Q(_stream_conv2d_16_source_28_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42930_ ( .CLK(CLK), .D(_02607_), .Q(_stream_conv2d_16_source_28_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_28_source_ram_renable_reg  ( .CLK(CLK), .D(_02608_), .Q(_stream_conv2d_16_source_28_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_28_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02609_), .Q(_stream_conv2d_16_source_28_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_29_idle_reg  ( .CLK(CLK), .D(_02611_), .Q(_stream_conv2d_16_source_29_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42934_ ( .CLK(CLK), .D(_02612_), .Q(_stream_conv2d_16_source_29_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42935_ ( .CLK(CLK), .D(_02613_), .Q(_stream_conv2d_16_source_29_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42936_ ( .CLK(CLK), .D(_02614_), .Q(_stream_conv2d_16_source_29_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42937_ ( .CLK(CLK), .D(_02619_), .Q(_stream_conv2d_16_source_29_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42938_ ( .CLK(CLK), .D(_02616_), .Q(_stream_conv2d_16_source_29_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_29_source_ram_renable_reg  ( .CLK(CLK), .D(_02617_), .Q(_stream_conv2d_16_source_29_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_29_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02618_), .Q(_stream_conv2d_16_source_29_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_30_idle_reg  ( .CLK(CLK), .D(_02620_), .Q(_stream_conv2d_16_source_30_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42942_ ( .CLK(CLK), .D(_02621_), .Q(_stream_conv2d_16_source_30_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42943_ ( .CLK(CLK), .D(_02622_), .Q(_stream_conv2d_16_source_30_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42944_ ( .CLK(CLK), .D(_02623_), .Q(_stream_conv2d_16_source_30_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42945_ ( .CLK(CLK), .D(_02628_), .Q(_stream_conv2d_16_source_30_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42946_ ( .CLK(CLK), .D(_02625_), .Q(_stream_conv2d_16_source_30_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_30_source_ram_renable_reg  ( .CLK(CLK), .D(_02626_), .Q(_stream_conv2d_16_source_30_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_30_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02627_), .Q(_stream_conv2d_16_source_30_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_31_idle_reg  ( .CLK(CLK), .D(_02629_), .Q(_stream_conv2d_16_source_31_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42950_ ( .CLK(CLK), .D(_02630_), .Q(_stream_conv2d_16_source_31_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42951_ ( .CLK(CLK), .D(_02631_), .Q(_stream_conv2d_16_source_31_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42952_ ( .CLK(CLK), .D(_02632_), .Q(_stream_conv2d_16_source_31_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42953_ ( .CLK(CLK), .D(_02637_), .Q(_stream_conv2d_16_source_31_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42954_ ( .CLK(CLK), .D(_02634_), .Q(_stream_conv2d_16_source_31_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_31_source_ram_renable_reg  ( .CLK(CLK), .D(_02635_), .Q(_stream_conv2d_16_source_31_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_31_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02636_), .Q(_stream_conv2d_16_source_31_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_32_idle_reg  ( .CLK(CLK), .D(_02638_), .Q(_stream_conv2d_16_source_32_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42958_ ( .CLK(CLK), .D(_02639_), .Q(_stream_conv2d_16_source_32_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42959_ ( .CLK(CLK), .D(_02640_), .Q(_stream_conv2d_16_source_32_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42960_ ( .CLK(CLK), .D(_02641_), .Q(_stream_conv2d_16_source_32_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42961_ ( .CLK(CLK), .D(_02646_), .Q(_stream_conv2d_16_source_32_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42962_ ( .CLK(CLK), .D(_02643_), .Q(_stream_conv2d_16_source_32_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_32_source_ram_renable_reg  ( .CLK(CLK), .D(_02644_), .Q(_stream_conv2d_16_source_32_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_32_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02645_), .Q(_stream_conv2d_16_source_32_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_33_idle_reg  ( .CLK(CLK), .D(_02647_), .Q(_stream_conv2d_16_source_33_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42966_ ( .CLK(CLK), .D(_02648_), .Q(_stream_conv2d_16_source_33_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42967_ ( .CLK(CLK), .D(_02649_), .Q(_stream_conv2d_16_source_33_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42968_ ( .CLK(CLK), .D(_02650_), .Q(_stream_conv2d_16_source_33_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42969_ ( .CLK(CLK), .D(_02655_), .Q(_stream_conv2d_16_source_33_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42970_ ( .CLK(CLK), .D(_02652_), .Q(_stream_conv2d_16_source_33_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_33_source_ram_renable_reg  ( .CLK(CLK), .D(_02653_), .Q(_stream_conv2d_16_source_33_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_33_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02654_), .Q(_stream_conv2d_16_source_33_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_34_idle_reg  ( .CLK(CLK), .D(_02656_), .Q(_stream_conv2d_16_source_34_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42974_ ( .CLK(CLK), .D(_02657_), .Q(_stream_conv2d_16_source_34_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42975_ ( .CLK(CLK), .D(_02658_), .Q(_stream_conv2d_16_source_34_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42976_ ( .CLK(CLK), .D(_02659_), .Q(_stream_conv2d_16_source_34_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42977_ ( .CLK(CLK), .D(_02664_), .Q(_stream_conv2d_16_source_34_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42978_ ( .CLK(CLK), .D(_02661_), .Q(_stream_conv2d_16_source_34_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_34_source_ram_renable_reg  ( .CLK(CLK), .D(_02662_), .Q(_stream_conv2d_16_source_34_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_34_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02663_), .Q(_stream_conv2d_16_source_34_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_35_idle_reg  ( .CLK(CLK), .D(_02665_), .Q(_stream_conv2d_16_source_35_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42982_ ( .CLK(CLK), .D(_02666_), .Q(_stream_conv2d_16_source_35_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42983_ ( .CLK(CLK), .D(_02667_), .Q(_stream_conv2d_16_source_35_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42984_ ( .CLK(CLK), .D(_02668_), .Q(_stream_conv2d_16_source_35_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42985_ ( .CLK(CLK), .D(_02673_), .Q(_stream_conv2d_16_source_35_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42986_ ( .CLK(CLK), .D(_02670_), .Q(_stream_conv2d_16_source_35_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_35_source_ram_renable_reg  ( .CLK(CLK), .D(_02671_), .Q(_stream_conv2d_16_source_35_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_35_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02672_), .Q(_stream_conv2d_16_source_35_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_36_idle_reg  ( .CLK(CLK), .D(_02674_), .Q(_stream_conv2d_16_source_36_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42990_ ( .CLK(CLK), .D(_02675_), .Q(_stream_conv2d_16_source_36_source_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42991_ ( .CLK(CLK), .D(_02676_), .Q(_stream_conv2d_16_source_36_source_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42992_ ( .CLK(CLK), .D(_02677_), .Q(_stream_conv2d_16_source_36_source_offset_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _42993_ ( .CLK(CLK), .D(_02682_), .Q(_stream_conv2d_16_source_36_source_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42994_ ( .CLK(CLK), .D(_02679_), .Q(_stream_conv2d_16_source_36_source_ram_raddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_36_source_ram_renable_reg  ( .CLK(CLK), .D(_02680_), .Q(_stream_conv2d_16_source_36_source_ram_renable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_source_36_source_ram_rvalid_reg  ( .CLK(CLK), .D(_02681_), .Q(_stream_conv2d_16_source_36_source_ram_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(3) ) _42997_ ( .CLK(CLK), .D(_02506_), .Q(_stream_conv2d_16_sink_37_sink_mode) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _42998_ ( .CLK(CLK), .D(_02507_), .Q(_stream_conv2d_16_sink_37_sink_offset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _42999_ ( .CLK(CLK), .D(_02509_), .Q(_stream_conv2d_16_sink_37_sink_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43000_ ( .CLK(CLK), .D(_02510_), .Q(_stream_conv2d_16_sink_37_sink_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43001_ ( .CLK(CLK), .D(_02504_), .Q(_stream_conv2d_16_sink_37_sink_count) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43002_ ( .CLK(CLK), .D(_02511_), .Q(_stream_conv2d_16_sink_37_sink_stride_buf) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43003_ ( .CLK(CLK), .D(_02508_), .Q(_stream_conv2d_16_sink_37_sink_ram_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43004_ ( .CLK(CLK), .D(_02512_), .Q(_stream_conv2d_16_sink_37_sink_waddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _stream_conv2d_16_sink_37_sink_wenable_reg  ( .CLK(CLK), .D(_02514_), .Q(_stream_conv2d_16_sink_37_sink_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43006_ ( .CLK(CLK), .D(_02513_), .Q(_stream_conv2d_16_sink_37_sink_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43007_ ( .CLK(CLK), .D(_01475_), .Q(_cond_data_235) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43008_ ( .CLK(CLK), .D(_01476_), .Q(_cond_data_242) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43009_ ( .CLK(CLK), .D(_01477_), .Q(_cond_data_249) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43010_ ( .CLK(CLK), .D(_01478_), .Q(_cond_data_256) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43011_ ( .CLK(CLK), .D(_01479_), .Q(_cond_data_263) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _eq_data_357_reg  ( .CLK(CLK), .D(_01680_), .Q(_eq_data_357) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _eq_data_361_reg  ( .CLK(CLK), .D(_01681_), .Q(_eq_data_361) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _eq_data_364_reg  ( .CLK(CLK), .D(_01682_), .Q(_eq_data_364) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _eq_data_447_reg  ( .CLK(CLK), .D(_01683_), .Q(_eq_data_447) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _eq_data_451_reg  ( .CLK(CLK), .D(_01684_), .Q(_eq_data_451) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _eq_data_454_reg  ( .CLK(CLK), .D(_01685_), .Q(_eq_data_454) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43018_ ( .CLK(CLK), .D(_00627_), .Q(__delay_data_898) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43019_ ( .CLK(CLK), .D(_00628_), .Q(__delay_data_900) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43020_ ( .CLK(CLK), .D(_00630_), .Q(__delay_data_904) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43021_ ( .CLK(CLK), .D(_00633_), .Q(__delay_data_907) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43022_ ( .CLK(CLK), .D(_00634_), .Q(__delay_data_909) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43023_ ( .CLK(CLK), .D(_00636_), .Q(__delay_data_913) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43024_ ( .CLK(CLK), .D(_00639_), .Q(__delay_data_916) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43025_ ( .CLK(CLK), .D(_00640_), .Q(__delay_data_918) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43026_ ( .CLK(CLK), .D(_00642_), .Q(__delay_data_922) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_940_reg  ( .CLK(CLK), .D(_00648_), .Q(__delay_data_940) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_947_reg  ( .CLK(CLK), .D(_00655_), .Q(__delay_data_947) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43029_ ( .CLK(CLK), .D(_00656_), .Q(__delay_data_948) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_992_reg  ( .CLK(CLK), .D(_00673_), .Q(__delay_data_992) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43031_ ( .CLK(CLK), .D(_00680_), .Q(__delay_data_999) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1040_reg  ( .CLK(CLK), .D(_00035_), .Q(__delay_data_1040) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43033_ ( .CLK(CLK), .D(_00042_), .Q(__delay_data_1047) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1075_reg  ( .CLK(CLK), .D(_00052_), .Q(__delay_data_1075) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43035_ ( .CLK(CLK), .D(_00059_), .Q(__delay_data_1082) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1110_reg  ( .CLK(CLK), .D(_00069_), .Q(__delay_data_1110) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43037_ ( .CLK(CLK), .D(_00076_), .Q(__delay_data_1117) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1145_reg  ( .CLK(CLK), .D(_00086_), .Q(__delay_data_1145) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43039_ ( .CLK(CLK), .D(_00093_), .Q(__delay_data_1152) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1179_reg  ( .CLK(CLK), .D(_00102_), .Q(__delay_data_1179) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43041_ ( .CLK(CLK), .D(_00109_), .Q(__delay_data_1186) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1213_reg  ( .CLK(CLK), .D(_00118_), .Q(__delay_data_1213) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43043_ ( .CLK(CLK), .D(_00125_), .Q(__delay_data_1220) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1247_reg  ( .CLK(CLK), .D(_00134_), .Q(__delay_data_1247) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43045_ ( .CLK(CLK), .D(_00141_), .Q(__delay_data_1254) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1268_reg  ( .CLK(CLK), .D(_00149_), .Q(__delay_data_1268) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43047_ ( .CLK(CLK), .D(_00170_), .Q(__delay_data_1289) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43048_ ( .CLK(CLK), .D(_00220_), .Q(__delay_data_1339) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43049_ ( .CLK(CLK), .D(_01480_), .Q(_cond_data_279) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43050_ ( .CLK(CLK), .D(_01483_), .Q(_cond_data_289) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43051_ ( .CLK(CLK), .D(_01486_), .Q(_cond_data_299) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43052_ ( .CLK(CLK), .D(_01489_), .Q(_cond_data_309) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43053_ ( .CLK(CLK), .D(_01492_), .Q(_cond_data_319) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43054_ ( .CLK(CLK), .D(_01495_), .Q(_cond_data_329) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43055_ ( .CLK(CLK), .D(_01498_), .Q(_cond_data_339) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43056_ ( .CLK(CLK), .D(_01501_), .Q(_cond_data_349) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43057_ ( .CLK(CLK), .D(_01504_), .Q(_cond_data_359) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43058_ ( .CLK(CLK), .D(_01811_), .Q(_plus_data_743) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43059_ ( .CLK(CLK), .D(_01812_), .Q(_plus_data_759) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43060_ ( .CLK(CLK), .D(_01814_), .Q(_plus_data_770) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43061_ ( .CLK(CLK), .D(_00629_), .Q(__delay_data_901) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43062_ ( .CLK(CLK), .D(_00631_), .Q(__delay_data_905) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43063_ ( .CLK(CLK), .D(_00635_), .Q(__delay_data_910) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43064_ ( .CLK(CLK), .D(_00637_), .Q(__delay_data_914) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43065_ ( .CLK(CLK), .D(_00641_), .Q(__delay_data_919) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43066_ ( .CLK(CLK), .D(_00643_), .Q(__delay_data_923) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_941_reg  ( .CLK(CLK), .D(_00649_), .Q(__delay_data_941) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43068_ ( .CLK(CLK), .D(_00657_), .Q(__delay_data_949) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43069_ ( .CLK(CLK), .D(_00664_), .Q(__delay_data_963) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43070_ ( .CLK(CLK), .D(_00666_), .Q(__delay_data_968) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43071_ ( .CLK(CLK), .D(_00668_), .Q(__delay_data_973) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_993_reg  ( .CLK(CLK), .D(_00674_), .Q(__delay_data_993) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43073_ ( .CLK(CLK), .D(_00001_), .Q(__delay_data_1000) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1021_reg  ( .CLK(CLK), .D(_00014_), .Q(__delay_data_1021) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1022_reg  ( .CLK(CLK), .D(_00015_), .Q(__delay_data_1022) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1041_reg  ( .CLK(CLK), .D(_00036_), .Q(__delay_data_1041) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43077_ ( .CLK(CLK), .D(_00043_), .Q(__delay_data_1048) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1076_reg  ( .CLK(CLK), .D(_00053_), .Q(__delay_data_1076) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43079_ ( .CLK(CLK), .D(_00060_), .Q(__delay_data_1083) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1111_reg  ( .CLK(CLK), .D(_00070_), .Q(__delay_data_1111) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43081_ ( .CLK(CLK), .D(_00077_), .Q(__delay_data_1118) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1146_reg  ( .CLK(CLK), .D(_00087_), .Q(__delay_data_1146) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43083_ ( .CLK(CLK), .D(_00094_), .Q(__delay_data_1153) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1180_reg  ( .CLK(CLK), .D(_00103_), .Q(__delay_data_1180) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43085_ ( .CLK(CLK), .D(_00110_), .Q(__delay_data_1187) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1214_reg  ( .CLK(CLK), .D(_00119_), .Q(__delay_data_1214) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43087_ ( .CLK(CLK), .D(_00126_), .Q(__delay_data_1221) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1234_reg  ( .CLK(CLK), .D(_00020_), .Q(__delay_data_1234) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1237_reg  ( .CLK(CLK), .D(_00023_), .Q(__delay_data_1237) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1241_reg  ( .CLK(CLK), .D(_00028_), .Q(__delay_data_1241) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1248_reg  ( .CLK(CLK), .D(_00135_), .Q(__delay_data_1248) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43092_ ( .CLK(CLK), .D(_00142_), .Q(__delay_data_1255) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43093_ ( .CLK(CLK), .D(_00171_), .Q(__delay_data_1290) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43094_ ( .CLK(CLK), .D(_00192_), .Q(__delay_data_1311) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43095_ ( .CLK(CLK), .D(_00221_), .Q(__delay_data_1340) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43096_ ( .CLK(CLK), .D(_01481_), .Q(_cond_data_283) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43097_ ( .CLK(CLK), .D(_01484_), .Q(_cond_data_293) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43098_ ( .CLK(CLK), .D(_01487_), .Q(_cond_data_303) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43099_ ( .CLK(CLK), .D(_01490_), .Q(_cond_data_313) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43100_ ( .CLK(CLK), .D(_01493_), .Q(_cond_data_323) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43101_ ( .CLK(CLK), .D(_01496_), .Q(_cond_data_333) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43102_ ( .CLK(CLK), .D(_01499_), .Q(_cond_data_343) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43103_ ( .CLK(CLK), .D(_01502_), .Q(_cond_data_353) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43104_ ( .CLK(CLK), .D(_01505_), .Q(_cond_data_363) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43105_ ( .CLK(CLK), .D(_00632_), .Q(__delay_data_906) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43106_ ( .CLK(CLK), .D(_00638_), .Q(__delay_data_915) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43107_ ( .CLK(CLK), .D(_00644_), .Q(__delay_data_924) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_942_reg  ( .CLK(CLK), .D(_00650_), .Q(__delay_data_942) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43109_ ( .CLK(CLK), .D(_00658_), .Q(__delay_data_950) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43110_ ( .CLK(CLK), .D(_00665_), .Q(__delay_data_966) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43111_ ( .CLK(CLK), .D(_00667_), .Q(__delay_data_971) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43112_ ( .CLK(CLK), .D(_00669_), .Q(__delay_data_976) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_994_reg  ( .CLK(CLK), .D(_00675_), .Q(__delay_data_994) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43114_ ( .CLK(CLK), .D(_00002_), .Q(__delay_data_1001) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43115_ ( .CLK(CLK), .D(_00017_), .Q(__delay_data_1016) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43116_ ( .CLK(CLK), .D(_00018_), .Q(__delay_data_1020) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1023_reg  ( .CLK(CLK), .D(_00016_), .Q(__delay_data_1023) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43118_ ( .CLK(CLK), .D(_00019_), .Q(__delay_data_1024) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1042_reg  ( .CLK(CLK), .D(_00037_), .Q(__delay_data_1042) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43120_ ( .CLK(CLK), .D(_00044_), .Q(__delay_data_1049) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1077_reg  ( .CLK(CLK), .D(_00054_), .Q(__delay_data_1077) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43122_ ( .CLK(CLK), .D(_00061_), .Q(__delay_data_1084) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1112_reg  ( .CLK(CLK), .D(_00071_), .Q(__delay_data_1112) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43124_ ( .CLK(CLK), .D(_00078_), .Q(__delay_data_1119) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1147_reg  ( .CLK(CLK), .D(_00088_), .Q(__delay_data_1147) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43126_ ( .CLK(CLK), .D(_00095_), .Q(__delay_data_1154) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1181_reg  ( .CLK(CLK), .D(_00104_), .Q(__delay_data_1181) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43128_ ( .CLK(CLK), .D(_00111_), .Q(__delay_data_1188) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1215_reg  ( .CLK(CLK), .D(_00120_), .Q(__delay_data_1215) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43130_ ( .CLK(CLK), .D(_00127_), .Q(__delay_data_1222) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1235_reg  ( .CLK(CLK), .D(_00021_), .Q(__delay_data_1235) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1238_reg  ( .CLK(CLK), .D(_00024_), .Q(__delay_data_1238) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1242_reg  ( .CLK(CLK), .D(_00029_), .Q(__delay_data_1242) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1249_reg  ( .CLK(CLK), .D(_00136_), .Q(__delay_data_1249) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43135_ ( .CLK(CLK), .D(_00143_), .Q(__delay_data_1256) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43136_ ( .CLK(CLK), .D(_00008_), .Q(__delay_data_1262) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43137_ ( .CLK(CLK), .D(_00150_), .Q(__delay_data_1269) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43138_ ( .CLK(CLK), .D(_00172_), .Q(__delay_data_1291) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43139_ ( .CLK(CLK), .D(_00193_), .Q(__delay_data_1312) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43140_ ( .CLK(CLK), .D(_00222_), .Q(__delay_data_1341) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43141_ ( .CLK(CLK), .D(_00250_), .Q(__delay_data_1369) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43142_ ( .CLK(CLK), .D(_01482_), .Q(_cond_data_286) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43143_ ( .CLK(CLK), .D(_01485_), .Q(_cond_data_296) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43144_ ( .CLK(CLK), .D(_01488_), .Q(_cond_data_306) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43145_ ( .CLK(CLK), .D(_01491_), .Q(_cond_data_316) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43146_ ( .CLK(CLK), .D(_01494_), .Q(_cond_data_326) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43147_ ( .CLK(CLK), .D(_01497_), .Q(_cond_data_336) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43148_ ( .CLK(CLK), .D(_01500_), .Q(_cond_data_346) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43149_ ( .CLK(CLK), .D(_01503_), .Q(_cond_data_356) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43150_ ( .CLK(CLK), .D(_01506_), .Q(_cond_data_366) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_943_reg  ( .CLK(CLK), .D(_00651_), .Q(__delay_data_943) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43152_ ( .CLK(CLK), .D(_00659_), .Q(__delay_data_951) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_995_reg  ( .CLK(CLK), .D(_00676_), .Q(__delay_data_995) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43154_ ( .CLK(CLK), .D(_00003_), .Q(__delay_data_1002) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1043_reg  ( .CLK(CLK), .D(_00038_), .Q(__delay_data_1043) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43156_ ( .CLK(CLK), .D(_00045_), .Q(__delay_data_1050) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1078_reg  ( .CLK(CLK), .D(_00055_), .Q(__delay_data_1078) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43158_ ( .CLK(CLK), .D(_00062_), .Q(__delay_data_1085) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1113_reg  ( .CLK(CLK), .D(_00072_), .Q(__delay_data_1113) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43160_ ( .CLK(CLK), .D(_00079_), .Q(__delay_data_1120) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1148_reg  ( .CLK(CLK), .D(_00089_), .Q(__delay_data_1148) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43162_ ( .CLK(CLK), .D(_00096_), .Q(__delay_data_1155) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1182_reg  ( .CLK(CLK), .D(_00105_), .Q(__delay_data_1182) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43164_ ( .CLK(CLK), .D(_00112_), .Q(__delay_data_1189) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1216_reg  ( .CLK(CLK), .D(_00121_), .Q(__delay_data_1216) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43166_ ( .CLK(CLK), .D(_00128_), .Q(__delay_data_1223) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1236_reg  ( .CLK(CLK), .D(_00022_), .Q(__delay_data_1236) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1239_reg  ( .CLK(CLK), .D(_00025_), .Q(__delay_data_1239) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1243_reg  ( .CLK(CLK), .D(_00030_), .Q(__delay_data_1243) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1250_reg  ( .CLK(CLK), .D(_00137_), .Q(__delay_data_1250) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43171_ ( .CLK(CLK), .D(_00144_), .Q(__delay_data_1257) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43172_ ( .CLK(CLK), .D(_00009_), .Q(__delay_data_1263) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43173_ ( .CLK(CLK), .D(_00151_), .Q(__delay_data_1270) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43174_ ( .CLK(CLK), .D(_00173_), .Q(__delay_data_1292) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43175_ ( .CLK(CLK), .D(_00194_), .Q(__delay_data_1313) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43176_ ( .CLK(CLK), .D(_00223_), .Q(__delay_data_1342) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43177_ ( .CLK(CLK), .D(_00251_), .Q(__delay_data_1370) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43178_ ( .CLK(CLK), .D(_01507_), .Q(_cond_data_369) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43179_ ( .CLK(CLK), .D(_01510_), .Q(_cond_data_379) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43180_ ( .CLK(CLK), .D(_01513_), .Q(_cond_data_389) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43181_ ( .CLK(CLK), .D(_01516_), .Q(_cond_data_399) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43182_ ( .CLK(CLK), .D(_01519_), .Q(_cond_data_409) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43183_ ( .CLK(CLK), .D(_01522_), .Q(_cond_data_419) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43184_ ( .CLK(CLK), .D(_01525_), .Q(_cond_data_429) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43185_ ( .CLK(CLK), .D(_01528_), .Q(_cond_data_439) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43186_ ( .CLK(CLK), .D(_01531_), .Q(_cond_data_449) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43187_ ( .CLK(CLK), .D(_00645_), .Q(__delay_data_932) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43188_ ( .CLK(CLK), .D(_00646_), .Q(__delay_data_938) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_944_reg  ( .CLK(CLK), .D(_00652_), .Q(__delay_data_944) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43190_ ( .CLK(CLK), .D(_00660_), .Q(__delay_data_952) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43191_ ( .CLK(CLK), .D(_00670_), .Q(__delay_data_984) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43192_ ( .CLK(CLK), .D(_00671_), .Q(__delay_data_990) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_996_reg  ( .CLK(CLK), .D(_00677_), .Q(__delay_data_996) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43194_ ( .CLK(CLK), .D(_00004_), .Q(__delay_data_1003) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43195_ ( .CLK(CLK), .D(_00027_), .Q(__delay_data_1032) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43196_ ( .CLK(CLK), .D(_00033_), .Q(__delay_data_1038) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1044_reg  ( .CLK(CLK), .D(_00039_), .Q(__delay_data_1044) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43198_ ( .CLK(CLK), .D(_00046_), .Q(__delay_data_1051) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43199_ ( .CLK(CLK), .D(_00050_), .Q(__delay_data_1068) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1079_reg  ( .CLK(CLK), .D(_00056_), .Q(__delay_data_1079) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43201_ ( .CLK(CLK), .D(_00063_), .Q(__delay_data_1086) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43202_ ( .CLK(CLK), .D(_00067_), .Q(__delay_data_1103) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1114_reg  ( .CLK(CLK), .D(_00073_), .Q(__delay_data_1114) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43204_ ( .CLK(CLK), .D(_00080_), .Q(__delay_data_1121) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43205_ ( .CLK(CLK), .D(_00084_), .Q(__delay_data_1138) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1149_reg  ( .CLK(CLK), .D(_00090_), .Q(__delay_data_1149) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43207_ ( .CLK(CLK), .D(_00097_), .Q(__delay_data_1156) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1183_reg  ( .CLK(CLK), .D(_00106_), .Q(__delay_data_1183) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43209_ ( .CLK(CLK), .D(_00113_), .Q(__delay_data_1190) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1217_reg  ( .CLK(CLK), .D(_00122_), .Q(__delay_data_1217) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43211_ ( .CLK(CLK), .D(_00129_), .Q(__delay_data_1224) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1240_reg  ( .CLK(CLK), .D(_00026_), .Q(__delay_data_1240) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1244_reg  ( .CLK(CLK), .D(_00031_), .Q(__delay_data_1244) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1251_reg  ( .CLK(CLK), .D(_00138_), .Q(__delay_data_1251) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43215_ ( .CLK(CLK), .D(_00145_), .Q(__delay_data_1258) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43216_ ( .CLK(CLK), .D(_00010_), .Q(__delay_data_1264) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43217_ ( .CLK(CLK), .D(_00152_), .Q(__delay_data_1271) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43218_ ( .CLK(CLK), .D(_00174_), .Q(__delay_data_1293) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43219_ ( .CLK(CLK), .D(_00195_), .Q(__delay_data_1314) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43220_ ( .CLK(CLK), .D(_00224_), .Q(__delay_data_1343) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43221_ ( .CLK(CLK), .D(_00252_), .Q(__delay_data_1371) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43222_ ( .CLK(CLK), .D(_01508_), .Q(_cond_data_373) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43223_ ( .CLK(CLK), .D(_01511_), .Q(_cond_data_383) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43224_ ( .CLK(CLK), .D(_01514_), .Q(_cond_data_393) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43225_ ( .CLK(CLK), .D(_01517_), .Q(_cond_data_403) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43226_ ( .CLK(CLK), .D(_01520_), .Q(_cond_data_413) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43227_ ( .CLK(CLK), .D(_01523_), .Q(_cond_data_423) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43228_ ( .CLK(CLK), .D(_01526_), .Q(_cond_data_433) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43229_ ( .CLK(CLK), .D(_01529_), .Q(_cond_data_443) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43230_ ( .CLK(CLK), .D(_01532_), .Q(_cond_data_453) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43231_ ( .CLK(CLK), .D(_00647_), .Q(__delay_data_939) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_945_reg  ( .CLK(CLK), .D(_00653_), .Q(__delay_data_945) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43233_ ( .CLK(CLK), .D(_00661_), .Q(__delay_data_953) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43234_ ( .CLK(CLK), .D(_00672_), .Q(__delay_data_991) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_997_reg  ( .CLK(CLK), .D(_00678_), .Q(__delay_data_997) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43236_ ( .CLK(CLK), .D(_00005_), .Q(__delay_data_1004) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43237_ ( .CLK(CLK), .D(_00034_), .Q(__delay_data_1039) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1045_reg  ( .CLK(CLK), .D(_00040_), .Q(__delay_data_1045) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43239_ ( .CLK(CLK), .D(_00047_), .Q(__delay_data_1052) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43240_ ( .CLK(CLK), .D(_00051_), .Q(__delay_data_1074) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1080_reg  ( .CLK(CLK), .D(_00057_), .Q(__delay_data_1080) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43242_ ( .CLK(CLK), .D(_00064_), .Q(__delay_data_1087) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43243_ ( .CLK(CLK), .D(_00068_), .Q(__delay_data_1109) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1115_reg  ( .CLK(CLK), .D(_00074_), .Q(__delay_data_1115) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43245_ ( .CLK(CLK), .D(_00081_), .Q(__delay_data_1122) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43246_ ( .CLK(CLK), .D(_00085_), .Q(__delay_data_1144) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1150_reg  ( .CLK(CLK), .D(_00091_), .Q(__delay_data_1150) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43248_ ( .CLK(CLK), .D(_00098_), .Q(__delay_data_1157) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43249_ ( .CLK(CLK), .D(_00101_), .Q(__delay_data_1178) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1184_reg  ( .CLK(CLK), .D(_00107_), .Q(__delay_data_1184) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43251_ ( .CLK(CLK), .D(_00114_), .Q(__delay_data_1191) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43252_ ( .CLK(CLK), .D(_00117_), .Q(__delay_data_1212) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1218_reg  ( .CLK(CLK), .D(_00123_), .Q(__delay_data_1218) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43254_ ( .CLK(CLK), .D(_00130_), .Q(__delay_data_1225) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1245_reg  ( .CLK(CLK), .D(_00032_), .Q(__delay_data_1245) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43256_ ( .CLK(CLK), .D(_00133_), .Q(__delay_data_1246) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1252_reg  ( .CLK(CLK), .D(_00139_), .Q(__delay_data_1252) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43258_ ( .CLK(CLK), .D(_00146_), .Q(__delay_data_1259) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43259_ ( .CLK(CLK), .D(_00011_), .Q(__delay_data_1265) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43260_ ( .CLK(CLK), .D(_00153_), .Q(__delay_data_1272) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43261_ ( .CLK(CLK), .D(_00175_), .Q(__delay_data_1294) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43262_ ( .CLK(CLK), .D(_00196_), .Q(__delay_data_1315) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43263_ ( .CLK(CLK), .D(_00225_), .Q(__delay_data_1344) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43264_ ( .CLK(CLK), .D(_00253_), .Q(__delay_data_1372) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43265_ ( .CLK(CLK), .D(_01509_), .Q(_cond_data_376) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43266_ ( .CLK(CLK), .D(_01512_), .Q(_cond_data_386) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43267_ ( .CLK(CLK), .D(_01515_), .Q(_cond_data_396) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43268_ ( .CLK(CLK), .D(_01518_), .Q(_cond_data_406) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43269_ ( .CLK(CLK), .D(_01521_), .Q(_cond_data_416) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43270_ ( .CLK(CLK), .D(_01524_), .Q(_cond_data_426) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43271_ ( .CLK(CLK), .D(_01527_), .Q(_cond_data_436) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43272_ ( .CLK(CLK), .D(_01530_), .Q(_cond_data_446) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43273_ ( .CLK(CLK), .D(_01533_), .Q(_cond_data_456) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_946_reg  ( .CLK(CLK), .D(_00654_), .Q(__delay_data_946) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43275_ ( .CLK(CLK), .D(_00662_), .Q(__delay_data_954) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_998_reg  ( .CLK(CLK), .D(_00679_), .Q(__delay_data_998) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43277_ ( .CLK(CLK), .D(_00006_), .Q(__delay_data_1005) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1046_reg  ( .CLK(CLK), .D(_00041_), .Q(__delay_data_1046) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43279_ ( .CLK(CLK), .D(_00048_), .Q(__delay_data_1053) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1081_reg  ( .CLK(CLK), .D(_00058_), .Q(__delay_data_1081) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43281_ ( .CLK(CLK), .D(_00065_), .Q(__delay_data_1088) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1116_reg  ( .CLK(CLK), .D(_00075_), .Q(__delay_data_1116) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43283_ ( .CLK(CLK), .D(_00082_), .Q(__delay_data_1123) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1151_reg  ( .CLK(CLK), .D(_00092_), .Q(__delay_data_1151) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43285_ ( .CLK(CLK), .D(_00099_), .Q(__delay_data_1158) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1185_reg  ( .CLK(CLK), .D(_00108_), .Q(__delay_data_1185) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43287_ ( .CLK(CLK), .D(_00115_), .Q(__delay_data_1192) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1219_reg  ( .CLK(CLK), .D(_00124_), .Q(__delay_data_1219) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43289_ ( .CLK(CLK), .D(_00131_), .Q(__delay_data_1226) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_1253_reg  ( .CLK(CLK), .D(_00140_), .Q(__delay_data_1253) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43291_ ( .CLK(CLK), .D(_00147_), .Q(__delay_data_1260) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43292_ ( .CLK(CLK), .D(_00012_), .Q(__delay_data_1266) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43293_ ( .CLK(CLK), .D(_00154_), .Q(__delay_data_1273) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43294_ ( .CLK(CLK), .D(_00176_), .Q(__delay_data_1295) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43295_ ( .CLK(CLK), .D(_00197_), .Q(__delay_data_1316) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43296_ ( .CLK(CLK), .D(_00226_), .Q(__delay_data_1345) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43297_ ( .CLK(CLK), .D(_00254_), .Q(__delay_data_1373) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43298_ ( .CLK(CLK), .D(_01537_), .Q(_cond_data_575) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43299_ ( .CLK(CLK), .D(_01538_), .Q(_cond_data_577) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43300_ ( .CLK(CLK), .D(_01539_), .Q(_cond_data_579) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43301_ ( .CLK(CLK), .D(_01540_), .Q(_cond_data_581) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43302_ ( .CLK(CLK), .D(_01541_), .Q(_cond_data_583) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43303_ ( .CLK(CLK), .D(_01542_), .Q(_cond_data_585) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43304_ ( .CLK(CLK), .D(_01543_), .Q(_cond_data_587) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43305_ ( .CLK(CLK), .D(_01544_), .Q(_cond_data_589) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43306_ ( .CLK(CLK), .D(_01545_), .Q(_cond_data_591) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43307_ ( .CLK(CLK), .D(_00663_), .Q(__delay_data_955) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43308_ ( .CLK(CLK), .D(_00007_), .Q(__delay_data_1006) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43309_ ( .CLK(CLK), .D(_00049_), .Q(__delay_data_1054) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43310_ ( .CLK(CLK), .D(_00066_), .Q(__delay_data_1089) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43311_ ( .CLK(CLK), .D(_00083_), .Q(__delay_data_1124) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43312_ ( .CLK(CLK), .D(_00100_), .Q(__delay_data_1159) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43313_ ( .CLK(CLK), .D(_00116_), .Q(__delay_data_1193) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43314_ ( .CLK(CLK), .D(_00132_), .Q(__delay_data_1227) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43315_ ( .CLK(CLK), .D(_00148_), .Q(__delay_data_1261) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43316_ ( .CLK(CLK), .D(_00013_), .Q(__delay_data_1267) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43317_ ( .CLK(CLK), .D(_00155_), .Q(__delay_data_1274) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43318_ ( .CLK(CLK), .D(_00177_), .Q(__delay_data_1296) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43319_ ( .CLK(CLK), .D(_00198_), .Q(__delay_data_1317) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43320_ ( .CLK(CLK), .D(_00227_), .Q(__delay_data_1346) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43321_ ( .CLK(CLK), .D(_00255_), .Q(__delay_data_1374) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43322_ ( .CLK(CLK), .D(_00156_), .Q(__delay_data_1275) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43323_ ( .CLK(CLK), .D(_00178_), .Q(__delay_data_1297) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43324_ ( .CLK(CLK), .D(_00199_), .Q(__delay_data_1318) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43325_ ( .CLK(CLK), .D(_00228_), .Q(__delay_data_1347) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43326_ ( .CLK(CLK), .D(_00256_), .Q(__delay_data_1375) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43327_ ( .CLK(CLK), .D(_00157_), .Q(__delay_data_1276) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43328_ ( .CLK(CLK), .D(_00179_), .Q(__delay_data_1298) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43329_ ( .CLK(CLK), .D(_00200_), .Q(__delay_data_1319) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43330_ ( .CLK(CLK), .D(_00229_), .Q(__delay_data_1348) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43331_ ( .CLK(CLK), .D(_00257_), .Q(__delay_data_1376) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43332_ ( .CLK(CLK), .D(_00158_), .Q(__delay_data_1277) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43333_ ( .CLK(CLK), .D(_00180_), .Q(__delay_data_1299) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43334_ ( .CLK(CLK), .D(_00201_), .Q(__delay_data_1320) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43335_ ( .CLK(CLK), .D(_00230_), .Q(__delay_data_1349) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43336_ ( .CLK(CLK), .D(_00258_), .Q(__delay_data_1377) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43337_ ( .CLK(CLK), .D(_00159_), .Q(__delay_data_1278) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43338_ ( .CLK(CLK), .D(_00181_), .Q(__delay_data_1300) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43339_ ( .CLK(CLK), .D(_00202_), .Q(__delay_data_1321) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43340_ ( .CLK(CLK), .D(_00231_), .Q(__delay_data_1350) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43341_ ( .CLK(CLK), .D(_00259_), .Q(__delay_data_1378) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43342_ ( .CLK(CLK), .D(_00160_), .Q(__delay_data_1279) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43343_ ( .CLK(CLK), .D(_00182_), .Q(__delay_data_1301) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43344_ ( .CLK(CLK), .D(_00203_), .Q(__delay_data_1322) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43345_ ( .CLK(CLK), .D(_00232_), .Q(__delay_data_1351) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43346_ ( .CLK(CLK), .D(_00260_), .Q(__delay_data_1379) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43347_ ( .CLK(CLK), .D(_00161_), .Q(__delay_data_1280) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43348_ ( .CLK(CLK), .D(_00183_), .Q(__delay_data_1302) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43349_ ( .CLK(CLK), .D(_00204_), .Q(__delay_data_1323) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43350_ ( .CLK(CLK), .D(_00233_), .Q(__delay_data_1352) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43351_ ( .CLK(CLK), .D(_00261_), .Q(__delay_data_1380) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43352_ ( .CLK(CLK), .D(_00162_), .Q(__delay_data_1281) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43353_ ( .CLK(CLK), .D(_00184_), .Q(__delay_data_1303) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43354_ ( .CLK(CLK), .D(_00205_), .Q(__delay_data_1324) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43355_ ( .CLK(CLK), .D(_00234_), .Q(__delay_data_1353) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43356_ ( .CLK(CLK), .D(_00262_), .Q(__delay_data_1381) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43357_ ( .CLK(CLK), .D(_00163_), .Q(__delay_data_1282) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43358_ ( .CLK(CLK), .D(_00185_), .Q(__delay_data_1304) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43359_ ( .CLK(CLK), .D(_00206_), .Q(__delay_data_1325) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43360_ ( .CLK(CLK), .D(_00235_), .Q(__delay_data_1354) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43361_ ( .CLK(CLK), .D(_00263_), .Q(__delay_data_1382) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43362_ ( .CLK(CLK), .D(_00164_), .Q(__delay_data_1283) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43363_ ( .CLK(CLK), .D(_00186_), .Q(__delay_data_1305) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43364_ ( .CLK(CLK), .D(_00207_), .Q(__delay_data_1326) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43365_ ( .CLK(CLK), .D(_00236_), .Q(__delay_data_1355) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43366_ ( .CLK(CLK), .D(_00264_), .Q(__delay_data_1383) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _43367_ ( .CLK(CLK), .D(_01090_), .Q(__substreamoutput_data_625) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _43368_ ( .CLK(CLK), .D(_01091_), .Q(__substreamoutput_data_642) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _43369_ ( .CLK(CLK), .D(_01092_), .Q(__substreamoutput_data_659) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _43370_ ( .CLK(CLK), .D(_01093_), .Q(__substreamoutput_data_676) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _43371_ ( .CLK(CLK), .D(_01094_), .Q(__substreamoutput_data_693) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _43372_ ( .CLK(CLK), .D(_01095_), .Q(__substreamoutput_data_710) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _43373_ ( .CLK(CLK), .D(_01096_), .Q(__substreamoutput_data_727) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _43374_ ( .CLK(CLK), .D(_01097_), .Q(__substreamoutput_data_744) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43375_ ( .CLK(CLK), .D(_00165_), .Q(__delay_data_1284) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43376_ ( .CLK(CLK), .D(_00187_), .Q(__delay_data_1306) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43377_ ( .CLK(CLK), .D(_00208_), .Q(__delay_data_1327) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43378_ ( .CLK(CLK), .D(_00237_), .Q(__delay_data_1356) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43379_ ( .CLK(CLK), .D(_00265_), .Q(__delay_data_1384) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43380_ ( .CLK(CLK), .D(_00166_), .Q(__delay_data_1285) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43381_ ( .CLK(CLK), .D(_00188_), .Q(__delay_data_1307) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43382_ ( .CLK(CLK), .D(_00209_), .Q(__delay_data_1328) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43383_ ( .CLK(CLK), .D(_00238_), .Q(__delay_data_1357) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43384_ ( .CLK(CLK), .D(_00266_), .Q(__delay_data_1385) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43385_ ( .CLK(CLK), .D(_00167_), .Q(__delay_data_1286) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43386_ ( .CLK(CLK), .D(_00189_), .Q(__delay_data_1308) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43387_ ( .CLK(CLK), .D(_00210_), .Q(__delay_data_1329) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43388_ ( .CLK(CLK), .D(_00239_), .Q(__delay_data_1358) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43389_ ( .CLK(CLK), .D(_00267_), .Q(__delay_data_1386) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43390_ ( .CLK(CLK), .D(_00168_), .Q(__delay_data_1287) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43391_ ( .CLK(CLK), .D(_00190_), .Q(__delay_data_1309) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43392_ ( .CLK(CLK), .D(_00211_), .Q(__delay_data_1330) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43393_ ( .CLK(CLK), .D(_00240_), .Q(__delay_data_1359) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43394_ ( .CLK(CLK), .D(_00268_), .Q(__delay_data_1387) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43395_ ( .CLK(CLK), .D(_01098_), .Q(__substreamoutput_data_746) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43396_ ( .CLK(CLK), .D(_00169_), .Q(__delay_data_1288) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43397_ ( .CLK(CLK), .D(_00191_), .Q(__delay_data_1310) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43398_ ( .CLK(CLK), .D(_00212_), .Q(__delay_data_1331) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43399_ ( .CLK(CLK), .D(_00241_), .Q(__delay_data_1360) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43400_ ( .CLK(CLK), .D(_00269_), .Q(__delay_data_1388) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43401_ ( .CLK(CLK), .D(_00213_), .Q(__delay_data_1332) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43402_ ( .CLK(CLK), .D(_00242_), .Q(__delay_data_1361) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43403_ ( .CLK(CLK), .D(_00270_), .Q(__delay_data_1389) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43404_ ( .CLK(CLK), .D(_00214_), .Q(__delay_data_1333) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43405_ ( .CLK(CLK), .D(_00243_), .Q(__delay_data_1362) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43406_ ( .CLK(CLK), .D(_00271_), .Q(__delay_data_1390) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43407_ ( .CLK(CLK), .D(_00215_), .Q(__delay_data_1334) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43408_ ( .CLK(CLK), .D(_00244_), .Q(__delay_data_1363) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43409_ ( .CLK(CLK), .D(_00272_), .Q(__delay_data_1391) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43410_ ( .CLK(CLK), .D(_00216_), .Q(__delay_data_1335) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43411_ ( .CLK(CLK), .D(_00245_), .Q(__delay_data_1364) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43412_ ( .CLK(CLK), .D(_00273_), .Q(__delay_data_1392) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43413_ ( .CLK(CLK), .D(_00217_), .Q(__delay_data_1336) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43414_ ( .CLK(CLK), .D(_00246_), .Q(__delay_data_1365) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43415_ ( .CLK(CLK), .D(_00274_), .Q(__delay_data_1393) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43416_ ( .CLK(CLK), .D(_00218_), .Q(__delay_data_1337) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43417_ ( .CLK(CLK), .D(_00247_), .Q(__delay_data_1366) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43418_ ( .CLK(CLK), .D(_00275_), .Q(__delay_data_1394) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43419_ ( .CLK(CLK), .D(_00219_), .Q(__delay_data_1338) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43420_ ( .CLK(CLK), .D(_00248_), .Q(__delay_data_1367) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43421_ ( .CLK(CLK), .D(_00276_), .Q(__delay_data_1395) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43422_ ( .CLK(CLK), .D(_01813_), .Q(_plus_data_762) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43423_ ( .CLK(CLK), .D(_00249_), .Q(__delay_data_1368) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43424_ ( .CLK(CLK), .D(_00277_), .Q(__delay_data_1396) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _43425_ ( .CLK(CLK), .D(_01395_), .Q(__variable_wdata_214) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _43426_ ( .CLK(CLK), .D(_01396_), .Q(__variable_wdata_215) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _43427_ ( .CLK(CLK), .D(_01397_), .Q(__variable_wdata_216) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _43428_ ( .CLK(CLK), .D(_01398_), .Q(__variable_wdata_217) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43429_ ( .CLK(CLK), .D(_02320_), .Q(_source_stream_conv2d_16_source_6_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43430_ ( .CLK(CLK), .D(_02321_), .Q(_source_stream_conv2d_16_source_6_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43431_ ( .CLK(CLK), .D(_02322_), .Q(_source_stream_conv2d_16_source_6_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43432_ ( .CLK(CLK), .D(_02323_), .Q(_source_stream_conv2d_16_source_6_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43433_ ( .CLK(CLK), .D(_02324_), .Q(_source_stream_conv2d_16_source_6_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43434_ ( .CLK(CLK), .D(_02325_), .Q(_source_stream_conv2d_16_source_6_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43435_ ( .CLK(CLK), .D(_02326_), .Q(_source_stream_conv2d_16_source_6_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43436_ ( .CLK(CLK), .D(_02327_), .Q(_source_stream_conv2d_16_source_6_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43437_ ( .CLK(CLK), .D(_02332_), .Q(_source_stream_conv2d_16_source_6_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43438_ ( .CLK(CLK), .D(_02333_), .Q(_source_stream_conv2d_16_source_6_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43439_ ( .CLK(CLK), .D(_02334_), .Q(_source_stream_conv2d_16_source_6_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43440_ ( .CLK(CLK), .D(_02335_), .Q(_source_stream_conv2d_16_source_6_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43441_ ( .CLK(CLK), .D(_02316_), .Q(_source_stream_conv2d_16_source_6_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43442_ ( .CLK(CLK), .D(_02317_), .Q(_source_stream_conv2d_16_source_6_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43443_ ( .CLK(CLK), .D(_02318_), .Q(_source_stream_conv2d_16_source_6_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43444_ ( .CLK(CLK), .D(_02319_), .Q(_source_stream_conv2d_16_source_6_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43445_ ( .CLK(CLK), .D(_02328_), .Q(_source_stream_conv2d_16_source_6_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43446_ ( .CLK(CLK), .D(_02329_), .Q(_source_stream_conv2d_16_source_6_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43447_ ( .CLK(CLK), .D(_02330_), .Q(_source_stream_conv2d_16_source_6_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43448_ ( .CLK(CLK), .D(_02331_), .Q(_source_stream_conv2d_16_source_6_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43449_ ( .CLK(CLK), .D(_02336_), .Q(_source_stream_conv2d_16_source_6_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43450_ ( .CLK(CLK), .D(_02337_), .Q(_source_stream_conv2d_16_source_6_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43451_ ( .CLK(CLK), .D(_02338_), .Q(_source_stream_conv2d_16_source_6_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43452_ ( .CLK(CLK), .D(_02339_), .Q(_source_stream_conv2d_16_source_6_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43453_ ( .CLK(CLK), .D(_01400_), .Q(__variable_wdata_230) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43454_ ( .CLK(CLK), .D(_02344_), .Q(_source_stream_conv2d_16_source_8_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43455_ ( .CLK(CLK), .D(_02345_), .Q(_source_stream_conv2d_16_source_8_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43456_ ( .CLK(CLK), .D(_02346_), .Q(_source_stream_conv2d_16_source_8_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43457_ ( .CLK(CLK), .D(_02347_), .Q(_source_stream_conv2d_16_source_8_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43458_ ( .CLK(CLK), .D(_02348_), .Q(_source_stream_conv2d_16_source_8_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43459_ ( .CLK(CLK), .D(_02349_), .Q(_source_stream_conv2d_16_source_8_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43460_ ( .CLK(CLK), .D(_02350_), .Q(_source_stream_conv2d_16_source_8_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43461_ ( .CLK(CLK), .D(_02351_), .Q(_source_stream_conv2d_16_source_8_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43462_ ( .CLK(CLK), .D(_02356_), .Q(_source_stream_conv2d_16_source_8_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43463_ ( .CLK(CLK), .D(_02357_), .Q(_source_stream_conv2d_16_source_8_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43464_ ( .CLK(CLK), .D(_02358_), .Q(_source_stream_conv2d_16_source_8_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43465_ ( .CLK(CLK), .D(_02359_), .Q(_source_stream_conv2d_16_source_8_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43466_ ( .CLK(CLK), .D(_02340_), .Q(_source_stream_conv2d_16_source_8_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43467_ ( .CLK(CLK), .D(_02341_), .Q(_source_stream_conv2d_16_source_8_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43468_ ( .CLK(CLK), .D(_02342_), .Q(_source_stream_conv2d_16_source_8_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43469_ ( .CLK(CLK), .D(_02343_), .Q(_source_stream_conv2d_16_source_8_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43470_ ( .CLK(CLK), .D(_02352_), .Q(_source_stream_conv2d_16_source_8_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43471_ ( .CLK(CLK), .D(_02353_), .Q(_source_stream_conv2d_16_source_8_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43472_ ( .CLK(CLK), .D(_02354_), .Q(_source_stream_conv2d_16_source_8_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43473_ ( .CLK(CLK), .D(_02355_), .Q(_source_stream_conv2d_16_source_8_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43474_ ( .CLK(CLK), .D(_02360_), .Q(_source_stream_conv2d_16_source_8_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43475_ ( .CLK(CLK), .D(_02361_), .Q(_source_stream_conv2d_16_source_8_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43476_ ( .CLK(CLK), .D(_02362_), .Q(_source_stream_conv2d_16_source_8_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43477_ ( .CLK(CLK), .D(_02363_), .Q(_source_stream_conv2d_16_source_8_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43478_ ( .CLK(CLK), .D(_01401_), .Q(__variable_wdata_237) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43479_ ( .CLK(CLK), .D(_01402_), .Q(__variable_wdata_244) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43480_ ( .CLK(CLK), .D(_01404_), .Q(__variable_wdata_251) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43481_ ( .CLK(CLK), .D(_01405_), .Q(__variable_wdata_258) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __variable_wdata_264_reg  ( .CLK(CLK), .D(_01407_), .Q(__variable_wdata_264) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __variable_wdata_265_reg  ( .CLK(CLK), .D(_01408_), .Q(__variable_wdata_265) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43484_ ( .CLK(CLK), .D(_01409_), .Q(__variable_wdata_266) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43485_ ( .CLK(CLK), .D(_01888_), .Q(_source_stream_conv2d_16_source_19_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43486_ ( .CLK(CLK), .D(_01889_), .Q(_source_stream_conv2d_16_source_19_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43487_ ( .CLK(CLK), .D(_01890_), .Q(_source_stream_conv2d_16_source_19_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43488_ ( .CLK(CLK), .D(_01891_), .Q(_source_stream_conv2d_16_source_19_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43489_ ( .CLK(CLK), .D(_01892_), .Q(_source_stream_conv2d_16_source_19_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43490_ ( .CLK(CLK), .D(_01893_), .Q(_source_stream_conv2d_16_source_19_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43491_ ( .CLK(CLK), .D(_01894_), .Q(_source_stream_conv2d_16_source_19_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43492_ ( .CLK(CLK), .D(_01895_), .Q(_source_stream_conv2d_16_source_19_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43493_ ( .CLK(CLK), .D(_01900_), .Q(_source_stream_conv2d_16_source_19_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43494_ ( .CLK(CLK), .D(_01901_), .Q(_source_stream_conv2d_16_source_19_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43495_ ( .CLK(CLK), .D(_01902_), .Q(_source_stream_conv2d_16_source_19_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43496_ ( .CLK(CLK), .D(_01903_), .Q(_source_stream_conv2d_16_source_19_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43497_ ( .CLK(CLK), .D(_01884_), .Q(_source_stream_conv2d_16_source_19_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43498_ ( .CLK(CLK), .D(_01885_), .Q(_source_stream_conv2d_16_source_19_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43499_ ( .CLK(CLK), .D(_01886_), .Q(_source_stream_conv2d_16_source_19_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43500_ ( .CLK(CLK), .D(_01887_), .Q(_source_stream_conv2d_16_source_19_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43501_ ( .CLK(CLK), .D(_01896_), .Q(_source_stream_conv2d_16_source_19_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43502_ ( .CLK(CLK), .D(_01897_), .Q(_source_stream_conv2d_16_source_19_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43503_ ( .CLK(CLK), .D(_01898_), .Q(_source_stream_conv2d_16_source_19_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43504_ ( .CLK(CLK), .D(_01899_), .Q(_source_stream_conv2d_16_source_19_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43505_ ( .CLK(CLK), .D(_01904_), .Q(_source_stream_conv2d_16_source_19_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43506_ ( .CLK(CLK), .D(_01905_), .Q(_source_stream_conv2d_16_source_19_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43507_ ( .CLK(CLK), .D(_01906_), .Q(_source_stream_conv2d_16_source_19_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43508_ ( .CLK(CLK), .D(_01907_), .Q(_source_stream_conv2d_16_source_19_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43509_ ( .CLK(CLK), .D(_01410_), .Q(__variable_wdata_268) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43510_ ( .CLK(CLK), .D(_01912_), .Q(_source_stream_conv2d_16_source_20_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43511_ ( .CLK(CLK), .D(_01913_), .Q(_source_stream_conv2d_16_source_20_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43512_ ( .CLK(CLK), .D(_01914_), .Q(_source_stream_conv2d_16_source_20_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43513_ ( .CLK(CLK), .D(_01915_), .Q(_source_stream_conv2d_16_source_20_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43514_ ( .CLK(CLK), .D(_01916_), .Q(_source_stream_conv2d_16_source_20_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43515_ ( .CLK(CLK), .D(_01917_), .Q(_source_stream_conv2d_16_source_20_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43516_ ( .CLK(CLK), .D(_01918_), .Q(_source_stream_conv2d_16_source_20_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43517_ ( .CLK(CLK), .D(_01919_), .Q(_source_stream_conv2d_16_source_20_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43518_ ( .CLK(CLK), .D(_01924_), .Q(_source_stream_conv2d_16_source_20_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43519_ ( .CLK(CLK), .D(_01925_), .Q(_source_stream_conv2d_16_source_20_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43520_ ( .CLK(CLK), .D(_01926_), .Q(_source_stream_conv2d_16_source_20_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43521_ ( .CLK(CLK), .D(_01927_), .Q(_source_stream_conv2d_16_source_20_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43522_ ( .CLK(CLK), .D(_01908_), .Q(_source_stream_conv2d_16_source_20_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43523_ ( .CLK(CLK), .D(_01909_), .Q(_source_stream_conv2d_16_source_20_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43524_ ( .CLK(CLK), .D(_01910_), .Q(_source_stream_conv2d_16_source_20_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43525_ ( .CLK(CLK), .D(_01911_), .Q(_source_stream_conv2d_16_source_20_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43526_ ( .CLK(CLK), .D(_01920_), .Q(_source_stream_conv2d_16_source_20_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43527_ ( .CLK(CLK), .D(_01921_), .Q(_source_stream_conv2d_16_source_20_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43528_ ( .CLK(CLK), .D(_01922_), .Q(_source_stream_conv2d_16_source_20_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43529_ ( .CLK(CLK), .D(_01923_), .Q(_source_stream_conv2d_16_source_20_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43530_ ( .CLK(CLK), .D(_01928_), .Q(_source_stream_conv2d_16_source_20_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43531_ ( .CLK(CLK), .D(_01929_), .Q(_source_stream_conv2d_16_source_20_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43532_ ( .CLK(CLK), .D(_01930_), .Q(_source_stream_conv2d_16_source_20_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43533_ ( .CLK(CLK), .D(_01931_), .Q(_source_stream_conv2d_16_source_20_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43534_ ( .CLK(CLK), .D(_01411_), .Q(__variable_wdata_269) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43535_ ( .CLK(CLK), .D(_01936_), .Q(_source_stream_conv2d_16_source_21_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43536_ ( .CLK(CLK), .D(_01937_), .Q(_source_stream_conv2d_16_source_21_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43537_ ( .CLK(CLK), .D(_01938_), .Q(_source_stream_conv2d_16_source_21_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43538_ ( .CLK(CLK), .D(_01939_), .Q(_source_stream_conv2d_16_source_21_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43539_ ( .CLK(CLK), .D(_01940_), .Q(_source_stream_conv2d_16_source_21_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43540_ ( .CLK(CLK), .D(_01941_), .Q(_source_stream_conv2d_16_source_21_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43541_ ( .CLK(CLK), .D(_01942_), .Q(_source_stream_conv2d_16_source_21_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43542_ ( .CLK(CLK), .D(_01943_), .Q(_source_stream_conv2d_16_source_21_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43543_ ( .CLK(CLK), .D(_01948_), .Q(_source_stream_conv2d_16_source_21_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43544_ ( .CLK(CLK), .D(_01949_), .Q(_source_stream_conv2d_16_source_21_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43545_ ( .CLK(CLK), .D(_01950_), .Q(_source_stream_conv2d_16_source_21_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43546_ ( .CLK(CLK), .D(_01951_), .Q(_source_stream_conv2d_16_source_21_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43547_ ( .CLK(CLK), .D(_01932_), .Q(_source_stream_conv2d_16_source_21_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43548_ ( .CLK(CLK), .D(_01933_), .Q(_source_stream_conv2d_16_source_21_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43549_ ( .CLK(CLK), .D(_01934_), .Q(_source_stream_conv2d_16_source_21_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43550_ ( .CLK(CLK), .D(_01935_), .Q(_source_stream_conv2d_16_source_21_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43551_ ( .CLK(CLK), .D(_01944_), .Q(_source_stream_conv2d_16_source_21_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43552_ ( .CLK(CLK), .D(_01945_), .Q(_source_stream_conv2d_16_source_21_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43553_ ( .CLK(CLK), .D(_01946_), .Q(_source_stream_conv2d_16_source_21_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43554_ ( .CLK(CLK), .D(_01947_), .Q(_source_stream_conv2d_16_source_21_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43555_ ( .CLK(CLK), .D(_01952_), .Q(_source_stream_conv2d_16_source_21_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43556_ ( .CLK(CLK), .D(_01953_), .Q(_source_stream_conv2d_16_source_21_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43557_ ( .CLK(CLK), .D(_01954_), .Q(_source_stream_conv2d_16_source_21_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43558_ ( .CLK(CLK), .D(_01955_), .Q(_source_stream_conv2d_16_source_21_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43559_ ( .CLK(CLK), .D(_01413_), .Q(__variable_wdata_270) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43560_ ( .CLK(CLK), .D(_01960_), .Q(_source_stream_conv2d_16_source_22_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43561_ ( .CLK(CLK), .D(_01961_), .Q(_source_stream_conv2d_16_source_22_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43562_ ( .CLK(CLK), .D(_01962_), .Q(_source_stream_conv2d_16_source_22_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43563_ ( .CLK(CLK), .D(_01963_), .Q(_source_stream_conv2d_16_source_22_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43564_ ( .CLK(CLK), .D(_01964_), .Q(_source_stream_conv2d_16_source_22_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43565_ ( .CLK(CLK), .D(_01965_), .Q(_source_stream_conv2d_16_source_22_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43566_ ( .CLK(CLK), .D(_01966_), .Q(_source_stream_conv2d_16_source_22_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43567_ ( .CLK(CLK), .D(_01967_), .Q(_source_stream_conv2d_16_source_22_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43568_ ( .CLK(CLK), .D(_01972_), .Q(_source_stream_conv2d_16_source_22_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43569_ ( .CLK(CLK), .D(_01973_), .Q(_source_stream_conv2d_16_source_22_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43570_ ( .CLK(CLK), .D(_01974_), .Q(_source_stream_conv2d_16_source_22_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43571_ ( .CLK(CLK), .D(_01975_), .Q(_source_stream_conv2d_16_source_22_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43572_ ( .CLK(CLK), .D(_01956_), .Q(_source_stream_conv2d_16_source_22_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43573_ ( .CLK(CLK), .D(_01957_), .Q(_source_stream_conv2d_16_source_22_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43574_ ( .CLK(CLK), .D(_01958_), .Q(_source_stream_conv2d_16_source_22_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43575_ ( .CLK(CLK), .D(_01959_), .Q(_source_stream_conv2d_16_source_22_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43576_ ( .CLK(CLK), .D(_01968_), .Q(_source_stream_conv2d_16_source_22_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43577_ ( .CLK(CLK), .D(_01969_), .Q(_source_stream_conv2d_16_source_22_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43578_ ( .CLK(CLK), .D(_01970_), .Q(_source_stream_conv2d_16_source_22_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43579_ ( .CLK(CLK), .D(_01971_), .Q(_source_stream_conv2d_16_source_22_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43580_ ( .CLK(CLK), .D(_01976_), .Q(_source_stream_conv2d_16_source_22_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43581_ ( .CLK(CLK), .D(_01977_), .Q(_source_stream_conv2d_16_source_22_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43582_ ( .CLK(CLK), .D(_01978_), .Q(_source_stream_conv2d_16_source_22_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43583_ ( .CLK(CLK), .D(_01979_), .Q(_source_stream_conv2d_16_source_22_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43584_ ( .CLK(CLK), .D(_01414_), .Q(__variable_wdata_271) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43585_ ( .CLK(CLK), .D(_01984_), .Q(_source_stream_conv2d_16_source_23_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43586_ ( .CLK(CLK), .D(_01985_), .Q(_source_stream_conv2d_16_source_23_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43587_ ( .CLK(CLK), .D(_01986_), .Q(_source_stream_conv2d_16_source_23_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43588_ ( .CLK(CLK), .D(_01987_), .Q(_source_stream_conv2d_16_source_23_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43589_ ( .CLK(CLK), .D(_01988_), .Q(_source_stream_conv2d_16_source_23_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43590_ ( .CLK(CLK), .D(_01989_), .Q(_source_stream_conv2d_16_source_23_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43591_ ( .CLK(CLK), .D(_01990_), .Q(_source_stream_conv2d_16_source_23_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43592_ ( .CLK(CLK), .D(_01991_), .Q(_source_stream_conv2d_16_source_23_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43593_ ( .CLK(CLK), .D(_01996_), .Q(_source_stream_conv2d_16_source_23_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43594_ ( .CLK(CLK), .D(_01997_), .Q(_source_stream_conv2d_16_source_23_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43595_ ( .CLK(CLK), .D(_01998_), .Q(_source_stream_conv2d_16_source_23_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43596_ ( .CLK(CLK), .D(_01999_), .Q(_source_stream_conv2d_16_source_23_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43597_ ( .CLK(CLK), .D(_01980_), .Q(_source_stream_conv2d_16_source_23_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43598_ ( .CLK(CLK), .D(_01981_), .Q(_source_stream_conv2d_16_source_23_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43599_ ( .CLK(CLK), .D(_01982_), .Q(_source_stream_conv2d_16_source_23_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43600_ ( .CLK(CLK), .D(_01983_), .Q(_source_stream_conv2d_16_source_23_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43601_ ( .CLK(CLK), .D(_01992_), .Q(_source_stream_conv2d_16_source_23_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43602_ ( .CLK(CLK), .D(_01993_), .Q(_source_stream_conv2d_16_source_23_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43603_ ( .CLK(CLK), .D(_01994_), .Q(_source_stream_conv2d_16_source_23_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43604_ ( .CLK(CLK), .D(_01995_), .Q(_source_stream_conv2d_16_source_23_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43605_ ( .CLK(CLK), .D(_02000_), .Q(_source_stream_conv2d_16_source_23_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43606_ ( .CLK(CLK), .D(_02001_), .Q(_source_stream_conv2d_16_source_23_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43607_ ( .CLK(CLK), .D(_02002_), .Q(_source_stream_conv2d_16_source_23_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43608_ ( .CLK(CLK), .D(_02003_), .Q(_source_stream_conv2d_16_source_23_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43609_ ( .CLK(CLK), .D(_01415_), .Q(__variable_wdata_272) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43610_ ( .CLK(CLK), .D(_02008_), .Q(_source_stream_conv2d_16_source_24_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43611_ ( .CLK(CLK), .D(_02009_), .Q(_source_stream_conv2d_16_source_24_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43612_ ( .CLK(CLK), .D(_02010_), .Q(_source_stream_conv2d_16_source_24_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43613_ ( .CLK(CLK), .D(_02011_), .Q(_source_stream_conv2d_16_source_24_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43614_ ( .CLK(CLK), .D(_02012_), .Q(_source_stream_conv2d_16_source_24_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43615_ ( .CLK(CLK), .D(_02013_), .Q(_source_stream_conv2d_16_source_24_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43616_ ( .CLK(CLK), .D(_02014_), .Q(_source_stream_conv2d_16_source_24_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43617_ ( .CLK(CLK), .D(_02015_), .Q(_source_stream_conv2d_16_source_24_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43618_ ( .CLK(CLK), .D(_02020_), .Q(_source_stream_conv2d_16_source_24_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43619_ ( .CLK(CLK), .D(_02021_), .Q(_source_stream_conv2d_16_source_24_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43620_ ( .CLK(CLK), .D(_02022_), .Q(_source_stream_conv2d_16_source_24_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43621_ ( .CLK(CLK), .D(_02023_), .Q(_source_stream_conv2d_16_source_24_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43622_ ( .CLK(CLK), .D(_02004_), .Q(_source_stream_conv2d_16_source_24_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43623_ ( .CLK(CLK), .D(_02005_), .Q(_source_stream_conv2d_16_source_24_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43624_ ( .CLK(CLK), .D(_02006_), .Q(_source_stream_conv2d_16_source_24_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43625_ ( .CLK(CLK), .D(_02007_), .Q(_source_stream_conv2d_16_source_24_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43626_ ( .CLK(CLK), .D(_02016_), .Q(_source_stream_conv2d_16_source_24_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43627_ ( .CLK(CLK), .D(_02017_), .Q(_source_stream_conv2d_16_source_24_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43628_ ( .CLK(CLK), .D(_02018_), .Q(_source_stream_conv2d_16_source_24_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43629_ ( .CLK(CLK), .D(_02019_), .Q(_source_stream_conv2d_16_source_24_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43630_ ( .CLK(CLK), .D(_02024_), .Q(_source_stream_conv2d_16_source_24_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43631_ ( .CLK(CLK), .D(_02025_), .Q(_source_stream_conv2d_16_source_24_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43632_ ( .CLK(CLK), .D(_02026_), .Q(_source_stream_conv2d_16_source_24_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43633_ ( .CLK(CLK), .D(_02027_), .Q(_source_stream_conv2d_16_source_24_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43634_ ( .CLK(CLK), .D(_01416_), .Q(__variable_wdata_273) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43635_ ( .CLK(CLK), .D(_02032_), .Q(_source_stream_conv2d_16_source_25_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43636_ ( .CLK(CLK), .D(_02033_), .Q(_source_stream_conv2d_16_source_25_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43637_ ( .CLK(CLK), .D(_02034_), .Q(_source_stream_conv2d_16_source_25_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43638_ ( .CLK(CLK), .D(_02035_), .Q(_source_stream_conv2d_16_source_25_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43639_ ( .CLK(CLK), .D(_02036_), .Q(_source_stream_conv2d_16_source_25_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43640_ ( .CLK(CLK), .D(_02037_), .Q(_source_stream_conv2d_16_source_25_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43641_ ( .CLK(CLK), .D(_02038_), .Q(_source_stream_conv2d_16_source_25_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43642_ ( .CLK(CLK), .D(_02039_), .Q(_source_stream_conv2d_16_source_25_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43643_ ( .CLK(CLK), .D(_02044_), .Q(_source_stream_conv2d_16_source_25_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43644_ ( .CLK(CLK), .D(_02045_), .Q(_source_stream_conv2d_16_source_25_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43645_ ( .CLK(CLK), .D(_02046_), .Q(_source_stream_conv2d_16_source_25_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43646_ ( .CLK(CLK), .D(_02047_), .Q(_source_stream_conv2d_16_source_25_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43647_ ( .CLK(CLK), .D(_02028_), .Q(_source_stream_conv2d_16_source_25_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43648_ ( .CLK(CLK), .D(_02029_), .Q(_source_stream_conv2d_16_source_25_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43649_ ( .CLK(CLK), .D(_02030_), .Q(_source_stream_conv2d_16_source_25_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43650_ ( .CLK(CLK), .D(_02031_), .Q(_source_stream_conv2d_16_source_25_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43651_ ( .CLK(CLK), .D(_02040_), .Q(_source_stream_conv2d_16_source_25_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43652_ ( .CLK(CLK), .D(_02041_), .Q(_source_stream_conv2d_16_source_25_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43653_ ( .CLK(CLK), .D(_02042_), .Q(_source_stream_conv2d_16_source_25_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43654_ ( .CLK(CLK), .D(_02043_), .Q(_source_stream_conv2d_16_source_25_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43655_ ( .CLK(CLK), .D(_02048_), .Q(_source_stream_conv2d_16_source_25_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43656_ ( .CLK(CLK), .D(_02049_), .Q(_source_stream_conv2d_16_source_25_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43657_ ( .CLK(CLK), .D(_02050_), .Q(_source_stream_conv2d_16_source_25_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43658_ ( .CLK(CLK), .D(_02051_), .Q(_source_stream_conv2d_16_source_25_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43659_ ( .CLK(CLK), .D(_01417_), .Q(__variable_wdata_274) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43660_ ( .CLK(CLK), .D(_02056_), .Q(_source_stream_conv2d_16_source_26_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43661_ ( .CLK(CLK), .D(_02057_), .Q(_source_stream_conv2d_16_source_26_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43662_ ( .CLK(CLK), .D(_02058_), .Q(_source_stream_conv2d_16_source_26_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43663_ ( .CLK(CLK), .D(_02059_), .Q(_source_stream_conv2d_16_source_26_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43664_ ( .CLK(CLK), .D(_02060_), .Q(_source_stream_conv2d_16_source_26_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43665_ ( .CLK(CLK), .D(_02061_), .Q(_source_stream_conv2d_16_source_26_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43666_ ( .CLK(CLK), .D(_02062_), .Q(_source_stream_conv2d_16_source_26_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43667_ ( .CLK(CLK), .D(_02063_), .Q(_source_stream_conv2d_16_source_26_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43668_ ( .CLK(CLK), .D(_02068_), .Q(_source_stream_conv2d_16_source_26_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43669_ ( .CLK(CLK), .D(_02069_), .Q(_source_stream_conv2d_16_source_26_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43670_ ( .CLK(CLK), .D(_02070_), .Q(_source_stream_conv2d_16_source_26_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43671_ ( .CLK(CLK), .D(_02071_), .Q(_source_stream_conv2d_16_source_26_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43672_ ( .CLK(CLK), .D(_02052_), .Q(_source_stream_conv2d_16_source_26_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43673_ ( .CLK(CLK), .D(_02053_), .Q(_source_stream_conv2d_16_source_26_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43674_ ( .CLK(CLK), .D(_02054_), .Q(_source_stream_conv2d_16_source_26_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43675_ ( .CLK(CLK), .D(_02055_), .Q(_source_stream_conv2d_16_source_26_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43676_ ( .CLK(CLK), .D(_02064_), .Q(_source_stream_conv2d_16_source_26_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43677_ ( .CLK(CLK), .D(_02065_), .Q(_source_stream_conv2d_16_source_26_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43678_ ( .CLK(CLK), .D(_02066_), .Q(_source_stream_conv2d_16_source_26_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43679_ ( .CLK(CLK), .D(_02067_), .Q(_source_stream_conv2d_16_source_26_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43680_ ( .CLK(CLK), .D(_02072_), .Q(_source_stream_conv2d_16_source_26_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43681_ ( .CLK(CLK), .D(_02073_), .Q(_source_stream_conv2d_16_source_26_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43682_ ( .CLK(CLK), .D(_02074_), .Q(_source_stream_conv2d_16_source_26_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43683_ ( .CLK(CLK), .D(_02075_), .Q(_source_stream_conv2d_16_source_26_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43684_ ( .CLK(CLK), .D(_01418_), .Q(__variable_wdata_275) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43685_ ( .CLK(CLK), .D(_02080_), .Q(_source_stream_conv2d_16_source_27_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43686_ ( .CLK(CLK), .D(_02081_), .Q(_source_stream_conv2d_16_source_27_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43687_ ( .CLK(CLK), .D(_02082_), .Q(_source_stream_conv2d_16_source_27_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43688_ ( .CLK(CLK), .D(_02083_), .Q(_source_stream_conv2d_16_source_27_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43689_ ( .CLK(CLK), .D(_02084_), .Q(_source_stream_conv2d_16_source_27_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43690_ ( .CLK(CLK), .D(_02085_), .Q(_source_stream_conv2d_16_source_27_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43691_ ( .CLK(CLK), .D(_02086_), .Q(_source_stream_conv2d_16_source_27_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43692_ ( .CLK(CLK), .D(_02087_), .Q(_source_stream_conv2d_16_source_27_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43693_ ( .CLK(CLK), .D(_02092_), .Q(_source_stream_conv2d_16_source_27_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43694_ ( .CLK(CLK), .D(_02093_), .Q(_source_stream_conv2d_16_source_27_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43695_ ( .CLK(CLK), .D(_02094_), .Q(_source_stream_conv2d_16_source_27_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43696_ ( .CLK(CLK), .D(_02095_), .Q(_source_stream_conv2d_16_source_27_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43697_ ( .CLK(CLK), .D(_02076_), .Q(_source_stream_conv2d_16_source_27_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43698_ ( .CLK(CLK), .D(_02077_), .Q(_source_stream_conv2d_16_source_27_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43699_ ( .CLK(CLK), .D(_02078_), .Q(_source_stream_conv2d_16_source_27_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43700_ ( .CLK(CLK), .D(_02079_), .Q(_source_stream_conv2d_16_source_27_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43701_ ( .CLK(CLK), .D(_02088_), .Q(_source_stream_conv2d_16_source_27_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43702_ ( .CLK(CLK), .D(_02089_), .Q(_source_stream_conv2d_16_source_27_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43703_ ( .CLK(CLK), .D(_02090_), .Q(_source_stream_conv2d_16_source_27_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43704_ ( .CLK(CLK), .D(_02091_), .Q(_source_stream_conv2d_16_source_27_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43705_ ( .CLK(CLK), .D(_02096_), .Q(_source_stream_conv2d_16_source_27_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43706_ ( .CLK(CLK), .D(_02097_), .Q(_source_stream_conv2d_16_source_27_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43707_ ( .CLK(CLK), .D(_02098_), .Q(_source_stream_conv2d_16_source_27_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43708_ ( .CLK(CLK), .D(_02099_), .Q(_source_stream_conv2d_16_source_27_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _43709_ ( .CLK(CLK), .D(_01419_), .Q(__variable_wdata_276) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43710_ ( .CLK(CLK), .D(_02104_), .Q(_source_stream_conv2d_16_source_28_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43711_ ( .CLK(CLK), .D(_02105_), .Q(_source_stream_conv2d_16_source_28_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43712_ ( .CLK(CLK), .D(_02106_), .Q(_source_stream_conv2d_16_source_28_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43713_ ( .CLK(CLK), .D(_02107_), .Q(_source_stream_conv2d_16_source_28_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43714_ ( .CLK(CLK), .D(_02108_), .Q(_source_stream_conv2d_16_source_28_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43715_ ( .CLK(CLK), .D(_02109_), .Q(_source_stream_conv2d_16_source_28_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43716_ ( .CLK(CLK), .D(_02110_), .Q(_source_stream_conv2d_16_source_28_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43717_ ( .CLK(CLK), .D(_02111_), .Q(_source_stream_conv2d_16_source_28_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43718_ ( .CLK(CLK), .D(_02116_), .Q(_source_stream_conv2d_16_source_28_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43719_ ( .CLK(CLK), .D(_02117_), .Q(_source_stream_conv2d_16_source_28_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43720_ ( .CLK(CLK), .D(_02118_), .Q(_source_stream_conv2d_16_source_28_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43721_ ( .CLK(CLK), .D(_02119_), .Q(_source_stream_conv2d_16_source_28_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43722_ ( .CLK(CLK), .D(_02100_), .Q(_source_stream_conv2d_16_source_28_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43723_ ( .CLK(CLK), .D(_02101_), .Q(_source_stream_conv2d_16_source_28_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43724_ ( .CLK(CLK), .D(_02102_), .Q(_source_stream_conv2d_16_source_28_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43725_ ( .CLK(CLK), .D(_02103_), .Q(_source_stream_conv2d_16_source_28_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43726_ ( .CLK(CLK), .D(_02112_), .Q(_source_stream_conv2d_16_source_28_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43727_ ( .CLK(CLK), .D(_02113_), .Q(_source_stream_conv2d_16_source_28_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43728_ ( .CLK(CLK), .D(_02114_), .Q(_source_stream_conv2d_16_source_28_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43729_ ( .CLK(CLK), .D(_02115_), .Q(_source_stream_conv2d_16_source_28_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43730_ ( .CLK(CLK), .D(_02120_), .Q(_source_stream_conv2d_16_source_28_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43731_ ( .CLK(CLK), .D(_02121_), .Q(_source_stream_conv2d_16_source_28_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43732_ ( .CLK(CLK), .D(_02122_), .Q(_source_stream_conv2d_16_source_28_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43733_ ( .CLK(CLK), .D(_02123_), .Q(_source_stream_conv2d_16_source_28_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43734_ ( .CLK(CLK), .D(_01430_), .Q(__variable_wdata_502) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43735_ ( .CLK(CLK), .D(_02128_), .Q(_source_stream_conv2d_16_source_29_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43736_ ( .CLK(CLK), .D(_02129_), .Q(_source_stream_conv2d_16_source_29_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43737_ ( .CLK(CLK), .D(_02130_), .Q(_source_stream_conv2d_16_source_29_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43738_ ( .CLK(CLK), .D(_02131_), .Q(_source_stream_conv2d_16_source_29_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43739_ ( .CLK(CLK), .D(_02132_), .Q(_source_stream_conv2d_16_source_29_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43740_ ( .CLK(CLK), .D(_02133_), .Q(_source_stream_conv2d_16_source_29_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43741_ ( .CLK(CLK), .D(_02134_), .Q(_source_stream_conv2d_16_source_29_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43742_ ( .CLK(CLK), .D(_02135_), .Q(_source_stream_conv2d_16_source_29_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43743_ ( .CLK(CLK), .D(_02140_), .Q(_source_stream_conv2d_16_source_29_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43744_ ( .CLK(CLK), .D(_02141_), .Q(_source_stream_conv2d_16_source_29_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43745_ ( .CLK(CLK), .D(_02142_), .Q(_source_stream_conv2d_16_source_29_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43746_ ( .CLK(CLK), .D(_02143_), .Q(_source_stream_conv2d_16_source_29_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43747_ ( .CLK(CLK), .D(_02124_), .Q(_source_stream_conv2d_16_source_29_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43748_ ( .CLK(CLK), .D(_02125_), .Q(_source_stream_conv2d_16_source_29_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43749_ ( .CLK(CLK), .D(_02126_), .Q(_source_stream_conv2d_16_source_29_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43750_ ( .CLK(CLK), .D(_02127_), .Q(_source_stream_conv2d_16_source_29_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43751_ ( .CLK(CLK), .D(_02136_), .Q(_source_stream_conv2d_16_source_29_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43752_ ( .CLK(CLK), .D(_02137_), .Q(_source_stream_conv2d_16_source_29_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43753_ ( .CLK(CLK), .D(_02138_), .Q(_source_stream_conv2d_16_source_29_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43754_ ( .CLK(CLK), .D(_02139_), .Q(_source_stream_conv2d_16_source_29_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43755_ ( .CLK(CLK), .D(_02144_), .Q(_source_stream_conv2d_16_source_29_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43756_ ( .CLK(CLK), .D(_02145_), .Q(_source_stream_conv2d_16_source_29_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43757_ ( .CLK(CLK), .D(_02146_), .Q(_source_stream_conv2d_16_source_29_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43758_ ( .CLK(CLK), .D(_02147_), .Q(_source_stream_conv2d_16_source_29_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43759_ ( .CLK(CLK), .D(_01431_), .Q(__variable_wdata_503) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43760_ ( .CLK(CLK), .D(_02152_), .Q(_source_stream_conv2d_16_source_30_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43761_ ( .CLK(CLK), .D(_02153_), .Q(_source_stream_conv2d_16_source_30_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43762_ ( .CLK(CLK), .D(_02154_), .Q(_source_stream_conv2d_16_source_30_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43763_ ( .CLK(CLK), .D(_02155_), .Q(_source_stream_conv2d_16_source_30_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43764_ ( .CLK(CLK), .D(_02156_), .Q(_source_stream_conv2d_16_source_30_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43765_ ( .CLK(CLK), .D(_02157_), .Q(_source_stream_conv2d_16_source_30_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43766_ ( .CLK(CLK), .D(_02158_), .Q(_source_stream_conv2d_16_source_30_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43767_ ( .CLK(CLK), .D(_02159_), .Q(_source_stream_conv2d_16_source_30_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43768_ ( .CLK(CLK), .D(_02164_), .Q(_source_stream_conv2d_16_source_30_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43769_ ( .CLK(CLK), .D(_02165_), .Q(_source_stream_conv2d_16_source_30_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43770_ ( .CLK(CLK), .D(_02166_), .Q(_source_stream_conv2d_16_source_30_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43771_ ( .CLK(CLK), .D(_02167_), .Q(_source_stream_conv2d_16_source_30_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43772_ ( .CLK(CLK), .D(_02148_), .Q(_source_stream_conv2d_16_source_30_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43773_ ( .CLK(CLK), .D(_02149_), .Q(_source_stream_conv2d_16_source_30_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43774_ ( .CLK(CLK), .D(_02150_), .Q(_source_stream_conv2d_16_source_30_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43775_ ( .CLK(CLK), .D(_02151_), .Q(_source_stream_conv2d_16_source_30_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43776_ ( .CLK(CLK), .D(_02160_), .Q(_source_stream_conv2d_16_source_30_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43777_ ( .CLK(CLK), .D(_02161_), .Q(_source_stream_conv2d_16_source_30_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43778_ ( .CLK(CLK), .D(_02162_), .Q(_source_stream_conv2d_16_source_30_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43779_ ( .CLK(CLK), .D(_02163_), .Q(_source_stream_conv2d_16_source_30_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43780_ ( .CLK(CLK), .D(_02168_), .Q(_source_stream_conv2d_16_source_30_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43781_ ( .CLK(CLK), .D(_02169_), .Q(_source_stream_conv2d_16_source_30_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43782_ ( .CLK(CLK), .D(_02170_), .Q(_source_stream_conv2d_16_source_30_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43783_ ( .CLK(CLK), .D(_02171_), .Q(_source_stream_conv2d_16_source_30_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43784_ ( .CLK(CLK), .D(_01432_), .Q(__variable_wdata_504) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43785_ ( .CLK(CLK), .D(_02176_), .Q(_source_stream_conv2d_16_source_31_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43786_ ( .CLK(CLK), .D(_02177_), .Q(_source_stream_conv2d_16_source_31_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43787_ ( .CLK(CLK), .D(_02178_), .Q(_source_stream_conv2d_16_source_31_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43788_ ( .CLK(CLK), .D(_02179_), .Q(_source_stream_conv2d_16_source_31_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43789_ ( .CLK(CLK), .D(_02180_), .Q(_source_stream_conv2d_16_source_31_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43790_ ( .CLK(CLK), .D(_02181_), .Q(_source_stream_conv2d_16_source_31_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43791_ ( .CLK(CLK), .D(_02182_), .Q(_source_stream_conv2d_16_source_31_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43792_ ( .CLK(CLK), .D(_02183_), .Q(_source_stream_conv2d_16_source_31_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43793_ ( .CLK(CLK), .D(_02188_), .Q(_source_stream_conv2d_16_source_31_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43794_ ( .CLK(CLK), .D(_02189_), .Q(_source_stream_conv2d_16_source_31_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43795_ ( .CLK(CLK), .D(_02190_), .Q(_source_stream_conv2d_16_source_31_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43796_ ( .CLK(CLK), .D(_02191_), .Q(_source_stream_conv2d_16_source_31_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43797_ ( .CLK(CLK), .D(_02172_), .Q(_source_stream_conv2d_16_source_31_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43798_ ( .CLK(CLK), .D(_02173_), .Q(_source_stream_conv2d_16_source_31_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43799_ ( .CLK(CLK), .D(_02174_), .Q(_source_stream_conv2d_16_source_31_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43800_ ( .CLK(CLK), .D(_02175_), .Q(_source_stream_conv2d_16_source_31_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43801_ ( .CLK(CLK), .D(_02184_), .Q(_source_stream_conv2d_16_source_31_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43802_ ( .CLK(CLK), .D(_02185_), .Q(_source_stream_conv2d_16_source_31_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43803_ ( .CLK(CLK), .D(_02186_), .Q(_source_stream_conv2d_16_source_31_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43804_ ( .CLK(CLK), .D(_02187_), .Q(_source_stream_conv2d_16_source_31_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43805_ ( .CLK(CLK), .D(_02192_), .Q(_source_stream_conv2d_16_source_31_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43806_ ( .CLK(CLK), .D(_02193_), .Q(_source_stream_conv2d_16_source_31_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43807_ ( .CLK(CLK), .D(_02194_), .Q(_source_stream_conv2d_16_source_31_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43808_ ( .CLK(CLK), .D(_02195_), .Q(_source_stream_conv2d_16_source_31_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43809_ ( .CLK(CLK), .D(_01433_), .Q(__variable_wdata_505) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43810_ ( .CLK(CLK), .D(_02200_), .Q(_source_stream_conv2d_16_source_32_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43811_ ( .CLK(CLK), .D(_02201_), .Q(_source_stream_conv2d_16_source_32_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43812_ ( .CLK(CLK), .D(_02202_), .Q(_source_stream_conv2d_16_source_32_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43813_ ( .CLK(CLK), .D(_02203_), .Q(_source_stream_conv2d_16_source_32_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43814_ ( .CLK(CLK), .D(_02204_), .Q(_source_stream_conv2d_16_source_32_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43815_ ( .CLK(CLK), .D(_02205_), .Q(_source_stream_conv2d_16_source_32_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43816_ ( .CLK(CLK), .D(_02206_), .Q(_source_stream_conv2d_16_source_32_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43817_ ( .CLK(CLK), .D(_02207_), .Q(_source_stream_conv2d_16_source_32_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43818_ ( .CLK(CLK), .D(_02212_), .Q(_source_stream_conv2d_16_source_32_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43819_ ( .CLK(CLK), .D(_02213_), .Q(_source_stream_conv2d_16_source_32_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43820_ ( .CLK(CLK), .D(_02214_), .Q(_source_stream_conv2d_16_source_32_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43821_ ( .CLK(CLK), .D(_02215_), .Q(_source_stream_conv2d_16_source_32_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43822_ ( .CLK(CLK), .D(_02196_), .Q(_source_stream_conv2d_16_source_32_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43823_ ( .CLK(CLK), .D(_02197_), .Q(_source_stream_conv2d_16_source_32_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43824_ ( .CLK(CLK), .D(_02198_), .Q(_source_stream_conv2d_16_source_32_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43825_ ( .CLK(CLK), .D(_02199_), .Q(_source_stream_conv2d_16_source_32_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43826_ ( .CLK(CLK), .D(_02208_), .Q(_source_stream_conv2d_16_source_32_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43827_ ( .CLK(CLK), .D(_02209_), .Q(_source_stream_conv2d_16_source_32_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43828_ ( .CLK(CLK), .D(_02210_), .Q(_source_stream_conv2d_16_source_32_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43829_ ( .CLK(CLK), .D(_02211_), .Q(_source_stream_conv2d_16_source_32_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43830_ ( .CLK(CLK), .D(_02216_), .Q(_source_stream_conv2d_16_source_32_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43831_ ( .CLK(CLK), .D(_02217_), .Q(_source_stream_conv2d_16_source_32_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43832_ ( .CLK(CLK), .D(_02218_), .Q(_source_stream_conv2d_16_source_32_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43833_ ( .CLK(CLK), .D(_02219_), .Q(_source_stream_conv2d_16_source_32_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43834_ ( .CLK(CLK), .D(_01434_), .Q(__variable_wdata_506) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43835_ ( .CLK(CLK), .D(_02224_), .Q(_source_stream_conv2d_16_source_33_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43836_ ( .CLK(CLK), .D(_02225_), .Q(_source_stream_conv2d_16_source_33_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43837_ ( .CLK(CLK), .D(_02226_), .Q(_source_stream_conv2d_16_source_33_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43838_ ( .CLK(CLK), .D(_02227_), .Q(_source_stream_conv2d_16_source_33_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43839_ ( .CLK(CLK), .D(_02228_), .Q(_source_stream_conv2d_16_source_33_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43840_ ( .CLK(CLK), .D(_02229_), .Q(_source_stream_conv2d_16_source_33_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43841_ ( .CLK(CLK), .D(_02230_), .Q(_source_stream_conv2d_16_source_33_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43842_ ( .CLK(CLK), .D(_02231_), .Q(_source_stream_conv2d_16_source_33_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43843_ ( .CLK(CLK), .D(_02236_), .Q(_source_stream_conv2d_16_source_33_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43844_ ( .CLK(CLK), .D(_02237_), .Q(_source_stream_conv2d_16_source_33_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43845_ ( .CLK(CLK), .D(_02238_), .Q(_source_stream_conv2d_16_source_33_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43846_ ( .CLK(CLK), .D(_02239_), .Q(_source_stream_conv2d_16_source_33_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43847_ ( .CLK(CLK), .D(_02220_), .Q(_source_stream_conv2d_16_source_33_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43848_ ( .CLK(CLK), .D(_02221_), .Q(_source_stream_conv2d_16_source_33_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43849_ ( .CLK(CLK), .D(_02222_), .Q(_source_stream_conv2d_16_source_33_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43850_ ( .CLK(CLK), .D(_02223_), .Q(_source_stream_conv2d_16_source_33_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43851_ ( .CLK(CLK), .D(_02232_), .Q(_source_stream_conv2d_16_source_33_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43852_ ( .CLK(CLK), .D(_02233_), .Q(_source_stream_conv2d_16_source_33_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43853_ ( .CLK(CLK), .D(_02234_), .Q(_source_stream_conv2d_16_source_33_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43854_ ( .CLK(CLK), .D(_02235_), .Q(_source_stream_conv2d_16_source_33_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43855_ ( .CLK(CLK), .D(_02240_), .Q(_source_stream_conv2d_16_source_33_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43856_ ( .CLK(CLK), .D(_02241_), .Q(_source_stream_conv2d_16_source_33_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43857_ ( .CLK(CLK), .D(_02242_), .Q(_source_stream_conv2d_16_source_33_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43858_ ( .CLK(CLK), .D(_02243_), .Q(_source_stream_conv2d_16_source_33_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43859_ ( .CLK(CLK), .D(_01435_), .Q(__variable_wdata_507) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43860_ ( .CLK(CLK), .D(_02248_), .Q(_source_stream_conv2d_16_source_34_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43861_ ( .CLK(CLK), .D(_02249_), .Q(_source_stream_conv2d_16_source_34_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43862_ ( .CLK(CLK), .D(_02250_), .Q(_source_stream_conv2d_16_source_34_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43863_ ( .CLK(CLK), .D(_02251_), .Q(_source_stream_conv2d_16_source_34_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43864_ ( .CLK(CLK), .D(_02252_), .Q(_source_stream_conv2d_16_source_34_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43865_ ( .CLK(CLK), .D(_02253_), .Q(_source_stream_conv2d_16_source_34_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43866_ ( .CLK(CLK), .D(_02254_), .Q(_source_stream_conv2d_16_source_34_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43867_ ( .CLK(CLK), .D(_02255_), .Q(_source_stream_conv2d_16_source_34_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43868_ ( .CLK(CLK), .D(_02260_), .Q(_source_stream_conv2d_16_source_34_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43869_ ( .CLK(CLK), .D(_02261_), .Q(_source_stream_conv2d_16_source_34_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43870_ ( .CLK(CLK), .D(_02262_), .Q(_source_stream_conv2d_16_source_34_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43871_ ( .CLK(CLK), .D(_02263_), .Q(_source_stream_conv2d_16_source_34_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43872_ ( .CLK(CLK), .D(_02244_), .Q(_source_stream_conv2d_16_source_34_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43873_ ( .CLK(CLK), .D(_02245_), .Q(_source_stream_conv2d_16_source_34_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43874_ ( .CLK(CLK), .D(_02246_), .Q(_source_stream_conv2d_16_source_34_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43875_ ( .CLK(CLK), .D(_02247_), .Q(_source_stream_conv2d_16_source_34_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43876_ ( .CLK(CLK), .D(_02256_), .Q(_source_stream_conv2d_16_source_34_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43877_ ( .CLK(CLK), .D(_02257_), .Q(_source_stream_conv2d_16_source_34_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43878_ ( .CLK(CLK), .D(_02258_), .Q(_source_stream_conv2d_16_source_34_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43879_ ( .CLK(CLK), .D(_02259_), .Q(_source_stream_conv2d_16_source_34_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43880_ ( .CLK(CLK), .D(_02264_), .Q(_source_stream_conv2d_16_source_34_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43881_ ( .CLK(CLK), .D(_02265_), .Q(_source_stream_conv2d_16_source_34_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43882_ ( .CLK(CLK), .D(_02266_), .Q(_source_stream_conv2d_16_source_34_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43883_ ( .CLK(CLK), .D(_02267_), .Q(_source_stream_conv2d_16_source_34_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43884_ ( .CLK(CLK), .D(_01436_), .Q(__variable_wdata_508) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43885_ ( .CLK(CLK), .D(_02272_), .Q(_source_stream_conv2d_16_source_35_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43886_ ( .CLK(CLK), .D(_02273_), .Q(_source_stream_conv2d_16_source_35_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43887_ ( .CLK(CLK), .D(_02274_), .Q(_source_stream_conv2d_16_source_35_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43888_ ( .CLK(CLK), .D(_02275_), .Q(_source_stream_conv2d_16_source_35_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43889_ ( .CLK(CLK), .D(_02276_), .Q(_source_stream_conv2d_16_source_35_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43890_ ( .CLK(CLK), .D(_02277_), .Q(_source_stream_conv2d_16_source_35_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43891_ ( .CLK(CLK), .D(_02278_), .Q(_source_stream_conv2d_16_source_35_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43892_ ( .CLK(CLK), .D(_02279_), .Q(_source_stream_conv2d_16_source_35_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43893_ ( .CLK(CLK), .D(_02284_), .Q(_source_stream_conv2d_16_source_35_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43894_ ( .CLK(CLK), .D(_02285_), .Q(_source_stream_conv2d_16_source_35_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43895_ ( .CLK(CLK), .D(_02286_), .Q(_source_stream_conv2d_16_source_35_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43896_ ( .CLK(CLK), .D(_02287_), .Q(_source_stream_conv2d_16_source_35_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43897_ ( .CLK(CLK), .D(_02268_), .Q(_source_stream_conv2d_16_source_35_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43898_ ( .CLK(CLK), .D(_02269_), .Q(_source_stream_conv2d_16_source_35_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43899_ ( .CLK(CLK), .D(_02270_), .Q(_source_stream_conv2d_16_source_35_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43900_ ( .CLK(CLK), .D(_02271_), .Q(_source_stream_conv2d_16_source_35_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43901_ ( .CLK(CLK), .D(_02280_), .Q(_source_stream_conv2d_16_source_35_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43902_ ( .CLK(CLK), .D(_02281_), .Q(_source_stream_conv2d_16_source_35_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43903_ ( .CLK(CLK), .D(_02282_), .Q(_source_stream_conv2d_16_source_35_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43904_ ( .CLK(CLK), .D(_02283_), .Q(_source_stream_conv2d_16_source_35_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43905_ ( .CLK(CLK), .D(_02288_), .Q(_source_stream_conv2d_16_source_35_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43906_ ( .CLK(CLK), .D(_02289_), .Q(_source_stream_conv2d_16_source_35_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43907_ ( .CLK(CLK), .D(_02290_), .Q(_source_stream_conv2d_16_source_35_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43908_ ( .CLK(CLK), .D(_02291_), .Q(_source_stream_conv2d_16_source_35_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43909_ ( .CLK(CLK), .D(_01437_), .Q(__variable_wdata_509) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43910_ ( .CLK(CLK), .D(_02296_), .Q(_source_stream_conv2d_16_source_36_pat_cur_offset_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43911_ ( .CLK(CLK), .D(_02297_), .Q(_source_stream_conv2d_16_source_36_pat_cur_offset_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43912_ ( .CLK(CLK), .D(_02298_), .Q(_source_stream_conv2d_16_source_36_pat_cur_offset_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43913_ ( .CLK(CLK), .D(_02299_), .Q(_source_stream_conv2d_16_source_36_pat_cur_offset_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43914_ ( .CLK(CLK), .D(_02300_), .Q(_source_stream_conv2d_16_source_36_pat_size_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43915_ ( .CLK(CLK), .D(_02301_), .Q(_source_stream_conv2d_16_source_36_pat_size_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43916_ ( .CLK(CLK), .D(_02302_), .Q(_source_stream_conv2d_16_source_36_pat_size_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43917_ ( .CLK(CLK), .D(_02303_), .Q(_source_stream_conv2d_16_source_36_pat_size_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43918_ ( .CLK(CLK), .D(_02308_), .Q(_source_stream_conv2d_16_source_36_pat_stride_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43919_ ( .CLK(CLK), .D(_02309_), .Q(_source_stream_conv2d_16_source_36_pat_stride_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43920_ ( .CLK(CLK), .D(_02310_), .Q(_source_stream_conv2d_16_source_36_pat_stride_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43921_ ( .CLK(CLK), .D(_02311_), .Q(_source_stream_conv2d_16_source_36_pat_stride_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43922_ ( .CLK(CLK), .D(_02292_), .Q(_source_stream_conv2d_16_source_36_pat_count_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43923_ ( .CLK(CLK), .D(_02293_), .Q(_source_stream_conv2d_16_source_36_pat_count_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43924_ ( .CLK(CLK), .D(_02294_), .Q(_source_stream_conv2d_16_source_36_pat_count_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43925_ ( .CLK(CLK), .D(_02295_), .Q(_source_stream_conv2d_16_source_36_pat_count_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43926_ ( .CLK(CLK), .D(_02304_), .Q(_source_stream_conv2d_16_source_36_pat_size_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43927_ ( .CLK(CLK), .D(_02305_), .Q(_source_stream_conv2d_16_source_36_pat_size_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43928_ ( .CLK(CLK), .D(_02306_), .Q(_source_stream_conv2d_16_source_36_pat_size_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43929_ ( .CLK(CLK), .D(_02307_), .Q(_source_stream_conv2d_16_source_36_pat_size_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43930_ ( .CLK(CLK), .D(_02312_), .Q(_source_stream_conv2d_16_source_36_pat_stride_buf_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43931_ ( .CLK(CLK), .D(_02313_), .Q(_source_stream_conv2d_16_source_36_pat_stride_buf_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43932_ ( .CLK(CLK), .D(_02314_), .Q(_source_stream_conv2d_16_source_36_pat_stride_buf_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43933_ ( .CLK(CLK), .D(_02315_), .Q(_source_stream_conv2d_16_source_36_pat_stride_buf_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _43934_ ( .CLK(CLK), .D(_01438_), .Q(__variable_wdata_510) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _set_flag_710_reg  ( .CLK(CLK), .D(_01873_), .Q(_set_flag_710) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43936_ ( .CLK(CLK), .D(_00811_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43937_ ( .CLK(CLK), .D(_00822_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43938_ ( .CLK(CLK), .D(_00833_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43939_ ( .CLK(CLK), .D(_00840_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43940_ ( .CLK(CLK), .D(_00841_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43941_ ( .CLK(CLK), .D(_00842_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43942_ ( .CLK(CLK), .D(_00843_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43943_ ( .CLK(CLK), .D(_00844_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43944_ ( .CLK(CLK), .D(_00845_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43945_ ( .CLK(CLK), .D(_00801_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43946_ ( .CLK(CLK), .D(_00802_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43947_ ( .CLK(CLK), .D(_00803_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43948_ ( .CLK(CLK), .D(_00804_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43949_ ( .CLK(CLK), .D(_00805_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43950_ ( .CLK(CLK), .D(_00806_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43951_ ( .CLK(CLK), .D(_00807_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43952_ ( .CLK(CLK), .D(_00808_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43953_ ( .CLK(CLK), .D(_00809_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43954_ ( .CLK(CLK), .D(_00810_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43955_ ( .CLK(CLK), .D(_00812_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43956_ ( .CLK(CLK), .D(_00813_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43957_ ( .CLK(CLK), .D(_00814_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43958_ ( .CLK(CLK), .D(_00815_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43959_ ( .CLK(CLK), .D(_00816_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43960_ ( .CLK(CLK), .D(_00817_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43961_ ( .CLK(CLK), .D(_00818_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43962_ ( .CLK(CLK), .D(_00819_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43963_ ( .CLK(CLK), .D(_00820_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43964_ ( .CLK(CLK), .D(_00821_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43965_ ( .CLK(CLK), .D(_00823_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43966_ ( .CLK(CLK), .D(_00824_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43967_ ( .CLK(CLK), .D(_00825_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43968_ ( .CLK(CLK), .D(_00826_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43969_ ( .CLK(CLK), .D(_00827_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43970_ ( .CLK(CLK), .D(_00828_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43971_ ( .CLK(CLK), .D(_00829_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43972_ ( .CLK(CLK), .D(_00830_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43973_ ( .CLK(CLK), .D(_00831_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43974_ ( .CLK(CLK), .D(_00832_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43975_ ( .CLK(CLK), .D(_00834_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43976_ ( .CLK(CLK), .D(_00835_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43977_ ( .CLK(CLK), .D(_00836_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_42) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43978_ ( .CLK(CLK), .D(_00837_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_43) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43979_ ( .CLK(CLK), .D(_00838_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_44) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _43980_ ( .CLK(CLK), .D(_00839_), .Q(__stream_conv2d_16_sink_37_sink_offset_0_45) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43981_ ( .CLK(CLK), .D(_00856_), .Q(__stream_conv2d_16_sink_37_sink_size_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43982_ ( .CLK(CLK), .D(_00867_), .Q(__stream_conv2d_16_sink_37_sink_size_1_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43983_ ( .CLK(CLK), .D(_00878_), .Q(__stream_conv2d_16_sink_37_sink_size_1_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43984_ ( .CLK(CLK), .D(_00885_), .Q(__stream_conv2d_16_sink_37_sink_size_1_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43985_ ( .CLK(CLK), .D(_00886_), .Q(__stream_conv2d_16_sink_37_sink_size_1_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43986_ ( .CLK(CLK), .D(_00887_), .Q(__stream_conv2d_16_sink_37_sink_size_1_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43987_ ( .CLK(CLK), .D(_00888_), .Q(__stream_conv2d_16_sink_37_sink_size_1_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43988_ ( .CLK(CLK), .D(_00889_), .Q(__stream_conv2d_16_sink_37_sink_size_1_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43989_ ( .CLK(CLK), .D(_00890_), .Q(__stream_conv2d_16_sink_37_sink_size_1_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43990_ ( .CLK(CLK), .D(_00846_), .Q(__stream_conv2d_16_sink_37_sink_size_1_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43991_ ( .CLK(CLK), .D(_00847_), .Q(__stream_conv2d_16_sink_37_sink_size_1_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43992_ ( .CLK(CLK), .D(_00848_), .Q(__stream_conv2d_16_sink_37_sink_size_1_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43993_ ( .CLK(CLK), .D(_00849_), .Q(__stream_conv2d_16_sink_37_sink_size_1_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43994_ ( .CLK(CLK), .D(_00850_), .Q(__stream_conv2d_16_sink_37_sink_size_1_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43995_ ( .CLK(CLK), .D(_00851_), .Q(__stream_conv2d_16_sink_37_sink_size_1_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43996_ ( .CLK(CLK), .D(_00852_), .Q(__stream_conv2d_16_sink_37_sink_size_1_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43997_ ( .CLK(CLK), .D(_00853_), .Q(__stream_conv2d_16_sink_37_sink_size_1_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43998_ ( .CLK(CLK), .D(_00854_), .Q(__stream_conv2d_16_sink_37_sink_size_1_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _43999_ ( .CLK(CLK), .D(_00855_), .Q(__stream_conv2d_16_sink_37_sink_size_1_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44000_ ( .CLK(CLK), .D(_00857_), .Q(__stream_conv2d_16_sink_37_sink_size_1_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44001_ ( .CLK(CLK), .D(_00858_), .Q(__stream_conv2d_16_sink_37_sink_size_1_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44002_ ( .CLK(CLK), .D(_00859_), .Q(__stream_conv2d_16_sink_37_sink_size_1_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44003_ ( .CLK(CLK), .D(_00860_), .Q(__stream_conv2d_16_sink_37_sink_size_1_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44004_ ( .CLK(CLK), .D(_00861_), .Q(__stream_conv2d_16_sink_37_sink_size_1_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44005_ ( .CLK(CLK), .D(_00862_), .Q(__stream_conv2d_16_sink_37_sink_size_1_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44006_ ( .CLK(CLK), .D(_00863_), .Q(__stream_conv2d_16_sink_37_sink_size_1_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44007_ ( .CLK(CLK), .D(_00864_), .Q(__stream_conv2d_16_sink_37_sink_size_1_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44008_ ( .CLK(CLK), .D(_00865_), .Q(__stream_conv2d_16_sink_37_sink_size_1_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44009_ ( .CLK(CLK), .D(_00866_), .Q(__stream_conv2d_16_sink_37_sink_size_1_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44010_ ( .CLK(CLK), .D(_00868_), .Q(__stream_conv2d_16_sink_37_sink_size_1_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44011_ ( .CLK(CLK), .D(_00869_), .Q(__stream_conv2d_16_sink_37_sink_size_1_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44012_ ( .CLK(CLK), .D(_00870_), .Q(__stream_conv2d_16_sink_37_sink_size_1_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44013_ ( .CLK(CLK), .D(_00871_), .Q(__stream_conv2d_16_sink_37_sink_size_1_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44014_ ( .CLK(CLK), .D(_00872_), .Q(__stream_conv2d_16_sink_37_sink_size_1_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44015_ ( .CLK(CLK), .D(_00873_), .Q(__stream_conv2d_16_sink_37_sink_size_1_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44016_ ( .CLK(CLK), .D(_00874_), .Q(__stream_conv2d_16_sink_37_sink_size_1_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44017_ ( .CLK(CLK), .D(_00875_), .Q(__stream_conv2d_16_sink_37_sink_size_1_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44018_ ( .CLK(CLK), .D(_00876_), .Q(__stream_conv2d_16_sink_37_sink_size_1_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44019_ ( .CLK(CLK), .D(_00877_), .Q(__stream_conv2d_16_sink_37_sink_size_1_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44020_ ( .CLK(CLK), .D(_00879_), .Q(__stream_conv2d_16_sink_37_sink_size_1_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44021_ ( .CLK(CLK), .D(_00880_), .Q(__stream_conv2d_16_sink_37_sink_size_1_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44022_ ( .CLK(CLK), .D(_00881_), .Q(__stream_conv2d_16_sink_37_sink_size_1_42) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44023_ ( .CLK(CLK), .D(_00882_), .Q(__stream_conv2d_16_sink_37_sink_size_1_43) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44024_ ( .CLK(CLK), .D(_00883_), .Q(__stream_conv2d_16_sink_37_sink_size_1_44) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44025_ ( .CLK(CLK), .D(_00884_), .Q(__stream_conv2d_16_sink_37_sink_size_1_45) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_1_reg  ( .CLK(CLK), .D(_00766_), .Q(__set_flag_710_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_2_reg  ( .CLK(CLK), .D(_00777_), .Q(__set_flag_710_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_3_reg  ( .CLK(CLK), .D(_00788_), .Q(__set_flag_710_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_4_reg  ( .CLK(CLK), .D(_00795_), .Q(__set_flag_710_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_5_reg  ( .CLK(CLK), .D(_00796_), .Q(__set_flag_710_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_6_reg  ( .CLK(CLK), .D(_00797_), .Q(__set_flag_710_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_7_reg  ( .CLK(CLK), .D(_00798_), .Q(__set_flag_710_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_8_reg  ( .CLK(CLK), .D(_00799_), .Q(__set_flag_710_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_9_reg  ( .CLK(CLK), .D(_00800_), .Q(__set_flag_710_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_10_reg  ( .CLK(CLK), .D(_00756_), .Q(__set_flag_710_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_11_reg  ( .CLK(CLK), .D(_00757_), .Q(__set_flag_710_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_12_reg  ( .CLK(CLK), .D(_00758_), .Q(__set_flag_710_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_13_reg  ( .CLK(CLK), .D(_00759_), .Q(__set_flag_710_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_14_reg  ( .CLK(CLK), .D(_00760_), .Q(__set_flag_710_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_15_reg  ( .CLK(CLK), .D(_00761_), .Q(__set_flag_710_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_16_reg  ( .CLK(CLK), .D(_00762_), .Q(__set_flag_710_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_17_reg  ( .CLK(CLK), .D(_00763_), .Q(__set_flag_710_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_18_reg  ( .CLK(CLK), .D(_00764_), .Q(__set_flag_710_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_19_reg  ( .CLK(CLK), .D(_00765_), .Q(__set_flag_710_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_20_reg  ( .CLK(CLK), .D(_00767_), .Q(__set_flag_710_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_21_reg  ( .CLK(CLK), .D(_00768_), .Q(__set_flag_710_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_22_reg  ( .CLK(CLK), .D(_00769_), .Q(__set_flag_710_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_23_reg  ( .CLK(CLK), .D(_00770_), .Q(__set_flag_710_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_24_reg  ( .CLK(CLK), .D(_00771_), .Q(__set_flag_710_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_25_reg  ( .CLK(CLK), .D(_00772_), .Q(__set_flag_710_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_26_reg  ( .CLK(CLK), .D(_00773_), .Q(__set_flag_710_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_27_reg  ( .CLK(CLK), .D(_00774_), .Q(__set_flag_710_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_28_reg  ( .CLK(CLK), .D(_00775_), .Q(__set_flag_710_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_29_reg  ( .CLK(CLK), .D(_00776_), .Q(__set_flag_710_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_30_reg  ( .CLK(CLK), .D(_00778_), .Q(__set_flag_710_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_31_reg  ( .CLK(CLK), .D(_00779_), .Q(__set_flag_710_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_32_reg  ( .CLK(CLK), .D(_00780_), .Q(__set_flag_710_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_33_reg  ( .CLK(CLK), .D(_00781_), .Q(__set_flag_710_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_34_reg  ( .CLK(CLK), .D(_00782_), .Q(__set_flag_710_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_35_reg  ( .CLK(CLK), .D(_00783_), .Q(__set_flag_710_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_36_reg  ( .CLK(CLK), .D(_00784_), .Q(__set_flag_710_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_37_reg  ( .CLK(CLK), .D(_00785_), .Q(__set_flag_710_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_38_reg  ( .CLK(CLK), .D(_00786_), .Q(__set_flag_710_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_39_reg  ( .CLK(CLK), .D(_00787_), .Q(__set_flag_710_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_40_reg  ( .CLK(CLK), .D(_00789_), .Q(__set_flag_710_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_41_reg  ( .CLK(CLK), .D(_00790_), .Q(__set_flag_710_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_42_reg  ( .CLK(CLK), .D(_00791_), .Q(__set_flag_710_42) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_43_reg  ( .CLK(CLK), .D(_00792_), .Q(__set_flag_710_43) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_44_reg  ( .CLK(CLK), .D(_00793_), .Q(__set_flag_710_44) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __set_flag_710_45_reg  ( .CLK(CLK), .D(_00794_), .Q(__set_flag_710_45) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_1_reg  ( .CLK(CLK), .D(_00901_), .Q(__stream_conv2d_16_start_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_2_reg  ( .CLK(CLK), .D(_00912_), .Q(__stream_conv2d_16_start_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_3_reg  ( .CLK(CLK), .D(_00923_), .Q(__stream_conv2d_16_start_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_4_reg  ( .CLK(CLK), .D(_00931_), .Q(__stream_conv2d_16_start_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_5_reg  ( .CLK(CLK), .D(_00932_), .Q(__stream_conv2d_16_start_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_6_reg  ( .CLK(CLK), .D(_00933_), .Q(__stream_conv2d_16_start_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_7_reg  ( .CLK(CLK), .D(_00934_), .Q(__stream_conv2d_16_start_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_8_reg  ( .CLK(CLK), .D(_00935_), .Q(__stream_conv2d_16_start_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_9_reg  ( .CLK(CLK), .D(_00936_), .Q(__stream_conv2d_16_start_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_10_reg  ( .CLK(CLK), .D(_00891_), .Q(__stream_conv2d_16_start_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_11_reg  ( .CLK(CLK), .D(_00892_), .Q(__stream_conv2d_16_start_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_12_reg  ( .CLK(CLK), .D(_00893_), .Q(__stream_conv2d_16_start_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_13_reg  ( .CLK(CLK), .D(_00894_), .Q(__stream_conv2d_16_start_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_14_reg  ( .CLK(CLK), .D(_00895_), .Q(__stream_conv2d_16_start_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_15_reg  ( .CLK(CLK), .D(_00896_), .Q(__stream_conv2d_16_start_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_16_reg  ( .CLK(CLK), .D(_00897_), .Q(__stream_conv2d_16_start_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_17_reg  ( .CLK(CLK), .D(_00898_), .Q(__stream_conv2d_16_start_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_18_reg  ( .CLK(CLK), .D(_00899_), .Q(__stream_conv2d_16_start_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_19_reg  ( .CLK(CLK), .D(_00900_), .Q(__stream_conv2d_16_start_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_20_reg  ( .CLK(CLK), .D(_00902_), .Q(__stream_conv2d_16_start_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_21_reg  ( .CLK(CLK), .D(_00903_), .Q(__stream_conv2d_16_start_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_22_reg  ( .CLK(CLK), .D(_00904_), .Q(__stream_conv2d_16_start_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_23_reg  ( .CLK(CLK), .D(_00905_), .Q(__stream_conv2d_16_start_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_24_reg  ( .CLK(CLK), .D(_00906_), .Q(__stream_conv2d_16_start_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_25_reg  ( .CLK(CLK), .D(_00907_), .Q(__stream_conv2d_16_start_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_26_reg  ( .CLK(CLK), .D(_00908_), .Q(__stream_conv2d_16_start_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_27_reg  ( .CLK(CLK), .D(_00909_), .Q(__stream_conv2d_16_start_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_28_reg  ( .CLK(CLK), .D(_00910_), .Q(__stream_conv2d_16_start_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_29_reg  ( .CLK(CLK), .D(_00911_), .Q(__stream_conv2d_16_start_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_30_reg  ( .CLK(CLK), .D(_00913_), .Q(__stream_conv2d_16_start_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_31_reg  ( .CLK(CLK), .D(_00914_), .Q(__stream_conv2d_16_start_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_32_reg  ( .CLK(CLK), .D(_00915_), .Q(__stream_conv2d_16_start_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_33_reg  ( .CLK(CLK), .D(_00916_), .Q(__stream_conv2d_16_start_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_34_reg  ( .CLK(CLK), .D(_00917_), .Q(__stream_conv2d_16_start_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_35_reg  ( .CLK(CLK), .D(_00918_), .Q(__stream_conv2d_16_start_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_36_reg  ( .CLK(CLK), .D(_00919_), .Q(__stream_conv2d_16_start_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_37_reg  ( .CLK(CLK), .D(_00920_), .Q(__stream_conv2d_16_start_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_38_reg  ( .CLK(CLK), .D(_00921_), .Q(__stream_conv2d_16_start_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_39_reg  ( .CLK(CLK), .D(_00922_), .Q(__stream_conv2d_16_start_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_40_reg  ( .CLK(CLK), .D(_00924_), .Q(__stream_conv2d_16_start_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_41_reg  ( .CLK(CLK), .D(_00925_), .Q(__stream_conv2d_16_start_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_42_reg  ( .CLK(CLK), .D(_00926_), .Q(__stream_conv2d_16_start_42) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_43_reg  ( .CLK(CLK), .D(_00927_), .Q(__stream_conv2d_16_start_43) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_44_reg  ( .CLK(CLK), .D(_00928_), .Q(__stream_conv2d_16_start_44) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_45_reg  ( .CLK(CLK), .D(_00929_), .Q(__stream_conv2d_16_start_45) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __stream_conv2d_16_start_46_reg  ( .CLK(CLK), .D(_00930_), .Q(__stream_conv2d_16_start_46) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_1_reg  ( .CLK(CLK), .D(_01289_), .Q(__tmp_799_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_2_reg  ( .CLK(CLK), .D(_01290_), .Q(__tmp_799_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_3_reg  ( .CLK(CLK), .D(_01291_), .Q(__tmp_799_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_4_reg  ( .CLK(CLK), .D(_01292_), .Q(__tmp_799_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_5_reg  ( .CLK(CLK), .D(_01293_), .Q(__tmp_799_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_6_reg  ( .CLK(CLK), .D(_01297_), .Q(__tmp_799_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_7_reg  ( .CLK(CLK), .D(_01298_), .Q(__tmp_799_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_8_reg  ( .CLK(CLK), .D(_01299_), .Q(__tmp_799_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_9_reg  ( .CLK(CLK), .D(_01300_), .Q(__tmp_799_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_10_reg  ( .CLK(CLK), .D(_01294_), .Q(__tmp_799_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_11_reg  ( .CLK(CLK), .D(_01295_), .Q(__tmp_799_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_12_reg  ( .CLK(CLK), .D(_01296_), .Q(__tmp_799_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_13_reg  ( .CLK(CLK), .D(_01301_), .Q(__tmp_799_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_14_reg  ( .CLK(CLK), .D(_01302_), .Q(__tmp_799_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_15_reg  ( .CLK(CLK), .D(_01303_), .Q(__tmp_799_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_16_reg  ( .CLK(CLK), .D(_01304_), .Q(__tmp_799_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_17_reg  ( .CLK(CLK), .D(_01305_), .Q(__tmp_799_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_18_reg  ( .CLK(CLK), .D(_01306_), .Q(__tmp_799_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_19_reg  ( .CLK(CLK), .D(_01307_), .Q(__tmp_799_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_20_reg  ( .CLK(CLK), .D(_01308_), .Q(__tmp_799_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_21_reg  ( .CLK(CLK), .D(_01309_), .Q(__tmp_799_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_22_reg  ( .CLK(CLK), .D(_01310_), .Q(__tmp_799_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_23_reg  ( .CLK(CLK), .D(_01311_), .Q(__tmp_799_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_24_reg  ( .CLK(CLK), .D(_01312_), .Q(__tmp_799_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_25_reg  ( .CLK(CLK), .D(_01313_), .Q(__tmp_799_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_26_reg  ( .CLK(CLK), .D(_01314_), .Q(__tmp_799_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_27_reg  ( .CLK(CLK), .D(_01315_), .Q(__tmp_799_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_28_reg  ( .CLK(CLK), .D(_01316_), .Q(__tmp_799_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_29_reg  ( .CLK(CLK), .D(_01317_), .Q(__tmp_799_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_30_reg  ( .CLK(CLK), .D(_01318_), .Q(__tmp_799_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_31_reg  ( .CLK(CLK), .D(_01319_), .Q(__tmp_799_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_32_reg  ( .CLK(CLK), .D(_01320_), .Q(__tmp_799_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_33_reg  ( .CLK(CLK), .D(_01321_), .Q(__tmp_799_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_799_34_reg  ( .CLK(CLK), .D(_01322_), .Q(__tmp_799_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_967_43_reg  ( .CLK(CLK), .D(_01365_), .Q(__tmp_967_43) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_967_44_reg  ( .CLK(CLK), .D(_01366_), .Q(__tmp_967_44) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_967_45_reg  ( .CLK(CLK), .D(_01367_), .Q(__tmp_967_45) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_967_46_reg  ( .CLK(CLK), .D(_01368_), .Q(__tmp_967_46) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_13_reg  ( .CLK(CLK), .D(_01335_), .Q(__tmp_969_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_14_reg  ( .CLK(CLK), .D(_01336_), .Q(__tmp_969_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_15_reg  ( .CLK(CLK), .D(_01337_), .Q(__tmp_969_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_16_reg  ( .CLK(CLK), .D(_01338_), .Q(__tmp_969_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_17_reg  ( .CLK(CLK), .D(_01339_), .Q(__tmp_969_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_18_reg  ( .CLK(CLK), .D(_01340_), .Q(__tmp_969_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_19_reg  ( .CLK(CLK), .D(_01341_), .Q(__tmp_969_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_20_reg  ( .CLK(CLK), .D(_01342_), .Q(__tmp_969_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_21_reg  ( .CLK(CLK), .D(_01343_), .Q(__tmp_969_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_22_reg  ( .CLK(CLK), .D(_01344_), .Q(__tmp_969_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_23_reg  ( .CLK(CLK), .D(_01345_), .Q(__tmp_969_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_24_reg  ( .CLK(CLK), .D(_01346_), .Q(__tmp_969_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_25_reg  ( .CLK(CLK), .D(_01347_), .Q(__tmp_969_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_26_reg  ( .CLK(CLK), .D(_01348_), .Q(__tmp_969_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_27_reg  ( .CLK(CLK), .D(_01349_), .Q(__tmp_969_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_28_reg  ( .CLK(CLK), .D(_01350_), .Q(__tmp_969_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_29_reg  ( .CLK(CLK), .D(_01351_), .Q(__tmp_969_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_30_reg  ( .CLK(CLK), .D(_01352_), .Q(__tmp_969_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_31_reg  ( .CLK(CLK), .D(_01353_), .Q(__tmp_969_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_32_reg  ( .CLK(CLK), .D(_01354_), .Q(__tmp_969_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_33_reg  ( .CLK(CLK), .D(_01355_), .Q(__tmp_969_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_34_reg  ( .CLK(CLK), .D(_01356_), .Q(__tmp_969_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_35_reg  ( .CLK(CLK), .D(_01357_), .Q(__tmp_969_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_36_reg  ( .CLK(CLK), .D(_01358_), .Q(__tmp_969_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_37_reg  ( .CLK(CLK), .D(_01359_), .Q(__tmp_969_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_38_reg  ( .CLK(CLK), .D(_01360_), .Q(__tmp_969_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_39_reg  ( .CLK(CLK), .D(_01361_), .Q(__tmp_969_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_40_reg  ( .CLK(CLK), .D(_01362_), .Q(__tmp_969_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_41_reg  ( .CLK(CLK), .D(_01363_), .Q(__tmp_969_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_969_42_reg  ( .CLK(CLK), .D(_01364_), .Q(__tmp_969_42) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __reduce_max_13_reduce_reset_reg  ( .CLK(CLK), .D(_00705_), .Q(__reduce_max_13_reduce_reset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream__reduce_max_13_x_data_cond_792_42_reg  ( .CLK(CLK), .D(_02799_), .Q(_substream__reduce_max_13_x_data_cond_792_42) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream__reduce_max_13_size_data_cond_792_43_reg  ( .CLK(CLK), .D(_02798_), .Q(_substream__reduce_max_13_size_data_cond_792_43) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44188_ ( .CLK(CLK), .D(_01840_), .Q(_reducemax_data_211) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44189_ ( .CLK(CLK), .D(_01839_), .Q(_reducemax_count_211) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _pulse_data_213_reg  ( .CLK(CLK), .D(_01823_), .Q(_pulse_data_213) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44191_ ( .CLK(CLK), .D(_01821_), .Q(_pulse_count_213) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44192_ ( .CLK(CLK), .D(_01393_), .Q(__variable_wdata_207) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44193_ ( .CLK(CLK), .D(_01394_), .Q(__variable_wdata_208) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1060_1_reg  ( .CLK(CLK), .D(_01121_), .Q(__tmp_1060_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1060_2_reg  ( .CLK(CLK), .D(_01122_), .Q(__tmp_1060_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1060_3_reg  ( .CLK(CLK), .D(_01123_), .Q(__tmp_1060_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1060_4_reg  ( .CLK(CLK), .D(_01124_), .Q(__tmp_1060_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1060_5_reg  ( .CLK(CLK), .D(_01125_), .Q(__tmp_1060_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_12_x_data_cond_728_24_reg  ( .CLK(CLK), .D(_02823_), .Q(_substream_mul_12_x_data_cond_728_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_12_y_data_cond_728_25_reg  ( .CLK(CLK), .D(_02824_), .Q(_substream_mul_12_y_data_cond_728_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_12_rshift_data_cond_728_26_reg  ( .CLK(CLK), .D(_02822_), .Q(_substream_mul_12_rshift_data_cond_728_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greaterthan_data_193_reg  ( .CLK(CLK), .D(_01696_), .Q(_greaterthan_data_193) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44203_ ( .CLK(CLK), .D(_01805_), .Q(_minus_data_195) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44204_ ( .CLK(CLK), .D(_00597_), .Q(__delay_data_730) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44205_ ( .CLK(CLK), .D(_00600_), .Q(__delay_data_733) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44206_ ( .CLK(CLK), .D(_00603_), .Q(__delay_data_736) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(18) ) _44207_ ( .CLK(CLK), .D(_01879_), .Q(_sll_data_197) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_729_reg  ( .CLK(CLK), .D(_00596_), .Q(__delay_data_729) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44209_ ( .CLK(CLK), .D(_00598_), .Q(__delay_data_731) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44210_ ( .CLK(CLK), .D(_00601_), .Q(__delay_data_734) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44211_ ( .CLK(CLK), .D(_00604_), .Q(__delay_data_737) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44212_ ( .CLK(CLK), .D(_01474_), .Q(_cond_data_203) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44213_ ( .CLK(CLK), .D(_00599_), .Q(__delay_data_732) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44214_ ( .CLK(CLK), .D(_00602_), .Q(__delay_data_735) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44215_ ( .CLK(CLK), .D(_00605_), .Q(__delay_data_738) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44216_ ( .CLK(CLK), .D(_00698_), .Q(__muladd_madd_odata_reg_205) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44217_ ( .CLK(CLK), .D(_00606_), .Q(__delay_data_739) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44218_ ( .CLK(CLK), .D(_00607_), .Q(__delay_data_740) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44219_ ( .CLK(CLK), .D(_00608_), .Q(__delay_data_741) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44220_ ( .CLK(CLK), .D(_00609_), .Q(__delay_data_742) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44221_ ( .CLK(CLK), .D(_02490_), .Q(_sra_data_206) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44222_ ( .CLK(CLK), .D(_01389_), .Q(__variable_wdata_190) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44223_ ( .CLK(CLK), .D(_01390_), .Q(__variable_wdata_191) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44224_ ( .CLK(CLK), .D(_01391_), .Q(__variable_wdata_192) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_11_x_data_cond_711_21_reg  ( .CLK(CLK), .D(_02820_), .Q(_substream_mul_11_x_data_cond_711_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_11_y_data_cond_711_22_reg  ( .CLK(CLK), .D(_02821_), .Q(_substream_mul_11_y_data_cond_711_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_11_rshift_data_cond_711_23_reg  ( .CLK(CLK), .D(_02819_), .Q(_substream_mul_11_rshift_data_cond_711_23) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greaterthan_data_176_reg  ( .CLK(CLK), .D(_01695_), .Q(_greaterthan_data_176) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44229_ ( .CLK(CLK), .D(_01804_), .Q(_minus_data_178) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44230_ ( .CLK(CLK), .D(_00583_), .Q(__delay_data_713) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44231_ ( .CLK(CLK), .D(_00586_), .Q(__delay_data_716) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44232_ ( .CLK(CLK), .D(_00589_), .Q(__delay_data_719) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(18) ) _44233_ ( .CLK(CLK), .D(_01878_), .Q(_sll_data_180) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_712_reg  ( .CLK(CLK), .D(_00582_), .Q(__delay_data_712) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44235_ ( .CLK(CLK), .D(_00584_), .Q(__delay_data_714) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44236_ ( .CLK(CLK), .D(_00587_), .Q(__delay_data_717) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44237_ ( .CLK(CLK), .D(_00590_), .Q(__delay_data_720) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44238_ ( .CLK(CLK), .D(_01473_), .Q(_cond_data_186) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44239_ ( .CLK(CLK), .D(_00585_), .Q(__delay_data_715) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44240_ ( .CLK(CLK), .D(_00588_), .Q(__delay_data_718) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44241_ ( .CLK(CLK), .D(_00591_), .Q(__delay_data_721) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44242_ ( .CLK(CLK), .D(_00697_), .Q(__muladd_madd_odata_reg_188) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44243_ ( .CLK(CLK), .D(_00592_), .Q(__delay_data_722) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44244_ ( .CLK(CLK), .D(_00593_), .Q(__delay_data_723) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44245_ ( .CLK(CLK), .D(_00594_), .Q(__delay_data_724) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44246_ ( .CLK(CLK), .D(_00595_), .Q(__delay_data_725) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44247_ ( .CLK(CLK), .D(_02489_), .Q(_sra_data_189) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44248_ ( .CLK(CLK), .D(_01386_), .Q(__variable_wdata_173) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44249_ ( .CLK(CLK), .D(_01387_), .Q(__variable_wdata_174) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44250_ ( .CLK(CLK), .D(_01388_), .Q(__variable_wdata_175) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_10_x_data_cond_694_18_reg  ( .CLK(CLK), .D(_02817_), .Q(_substream_mul_10_x_data_cond_694_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_10_y_data_cond_694_19_reg  ( .CLK(CLK), .D(_02818_), .Q(_substream_mul_10_y_data_cond_694_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_10_rshift_data_cond_694_20_reg  ( .CLK(CLK), .D(_02816_), .Q(_substream_mul_10_rshift_data_cond_694_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greaterthan_data_159_reg  ( .CLK(CLK), .D(_01694_), .Q(_greaterthan_data_159) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44255_ ( .CLK(CLK), .D(_01803_), .Q(_minus_data_161) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44256_ ( .CLK(CLK), .D(_00569_), .Q(__delay_data_696) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44257_ ( .CLK(CLK), .D(_00572_), .Q(__delay_data_699) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44258_ ( .CLK(CLK), .D(_00575_), .Q(__delay_data_702) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(18) ) _44259_ ( .CLK(CLK), .D(_01877_), .Q(_sll_data_163) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_695_reg  ( .CLK(CLK), .D(_00568_), .Q(__delay_data_695) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44261_ ( .CLK(CLK), .D(_00570_), .Q(__delay_data_697) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44262_ ( .CLK(CLK), .D(_00573_), .Q(__delay_data_700) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44263_ ( .CLK(CLK), .D(_00576_), .Q(__delay_data_703) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44264_ ( .CLK(CLK), .D(_01472_), .Q(_cond_data_169) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44265_ ( .CLK(CLK), .D(_00571_), .Q(__delay_data_698) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44266_ ( .CLK(CLK), .D(_00574_), .Q(__delay_data_701) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44267_ ( .CLK(CLK), .D(_00577_), .Q(__delay_data_704) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44268_ ( .CLK(CLK), .D(_00696_), .Q(__muladd_madd_odata_reg_171) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44269_ ( .CLK(CLK), .D(_00578_), .Q(__delay_data_705) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44270_ ( .CLK(CLK), .D(_00579_), .Q(__delay_data_706) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44271_ ( .CLK(CLK), .D(_00580_), .Q(__delay_data_707) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44272_ ( .CLK(CLK), .D(_00581_), .Q(__delay_data_708) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44273_ ( .CLK(CLK), .D(_02488_), .Q(_sra_data_172) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44274_ ( .CLK(CLK), .D(_01383_), .Q(__variable_wdata_156) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44275_ ( .CLK(CLK), .D(_01384_), .Q(__variable_wdata_157) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44276_ ( .CLK(CLK), .D(_01385_), .Q(__variable_wdata_158) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_9_x_data_cond_677_15_reg  ( .CLK(CLK), .D(_02844_), .Q(_substream_mul_9_x_data_cond_677_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_9_y_data_cond_677_16_reg  ( .CLK(CLK), .D(_02845_), .Q(_substream_mul_9_y_data_cond_677_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_9_rshift_data_cond_677_17_reg  ( .CLK(CLK), .D(_02843_), .Q(_substream_mul_9_rshift_data_cond_677_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greaterthan_data_142_reg  ( .CLK(CLK), .D(_01693_), .Q(_greaterthan_data_142) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44281_ ( .CLK(CLK), .D(_01802_), .Q(_minus_data_144) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44282_ ( .CLK(CLK), .D(_00555_), .Q(__delay_data_679) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44283_ ( .CLK(CLK), .D(_00558_), .Q(__delay_data_682) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44284_ ( .CLK(CLK), .D(_00561_), .Q(__delay_data_685) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(18) ) _44285_ ( .CLK(CLK), .D(_01876_), .Q(_sll_data_146) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_678_reg  ( .CLK(CLK), .D(_00554_), .Q(__delay_data_678) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44287_ ( .CLK(CLK), .D(_00556_), .Q(__delay_data_680) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44288_ ( .CLK(CLK), .D(_00559_), .Q(__delay_data_683) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44289_ ( .CLK(CLK), .D(_00562_), .Q(__delay_data_686) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44290_ ( .CLK(CLK), .D(_01471_), .Q(_cond_data_152) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44291_ ( .CLK(CLK), .D(_00557_), .Q(__delay_data_681) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44292_ ( .CLK(CLK), .D(_00560_), .Q(__delay_data_684) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44293_ ( .CLK(CLK), .D(_00563_), .Q(__delay_data_687) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44294_ ( .CLK(CLK), .D(_00695_), .Q(__muladd_madd_odata_reg_154) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44295_ ( .CLK(CLK), .D(_00564_), .Q(__delay_data_688) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44296_ ( .CLK(CLK), .D(_00565_), .Q(__delay_data_689) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44297_ ( .CLK(CLK), .D(_00566_), .Q(__delay_data_690) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44298_ ( .CLK(CLK), .D(_00567_), .Q(__delay_data_691) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44299_ ( .CLK(CLK), .D(_02487_), .Q(_sra_data_155) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44300_ ( .CLK(CLK), .D(_01380_), .Q(__variable_wdata_139) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44301_ ( .CLK(CLK), .D(_01381_), .Q(__variable_wdata_140) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44302_ ( .CLK(CLK), .D(_01382_), .Q(__variable_wdata_141) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_8_x_data_cond_660_12_reg  ( .CLK(CLK), .D(_02841_), .Q(_substream_mul_8_x_data_cond_660_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_8_y_data_cond_660_13_reg  ( .CLK(CLK), .D(_02842_), .Q(_substream_mul_8_y_data_cond_660_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_8_rshift_data_cond_660_14_reg  ( .CLK(CLK), .D(_02840_), .Q(_substream_mul_8_rshift_data_cond_660_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greaterthan_data_125_reg  ( .CLK(CLK), .D(_01692_), .Q(_greaterthan_data_125) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44307_ ( .CLK(CLK), .D(_01801_), .Q(_minus_data_127) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44308_ ( .CLK(CLK), .D(_00541_), .Q(__delay_data_662) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44309_ ( .CLK(CLK), .D(_00544_), .Q(__delay_data_665) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44310_ ( .CLK(CLK), .D(_00547_), .Q(__delay_data_668) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(18) ) _44311_ ( .CLK(CLK), .D(_01875_), .Q(_sll_data_129) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_661_reg  ( .CLK(CLK), .D(_00540_), .Q(__delay_data_661) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44313_ ( .CLK(CLK), .D(_00542_), .Q(__delay_data_663) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44314_ ( .CLK(CLK), .D(_00545_), .Q(__delay_data_666) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44315_ ( .CLK(CLK), .D(_00548_), .Q(__delay_data_669) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44316_ ( .CLK(CLK), .D(_01469_), .Q(_cond_data_135) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44317_ ( .CLK(CLK), .D(_00543_), .Q(__delay_data_664) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44318_ ( .CLK(CLK), .D(_00546_), .Q(__delay_data_667) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44319_ ( .CLK(CLK), .D(_00549_), .Q(__delay_data_670) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44320_ ( .CLK(CLK), .D(_00694_), .Q(__muladd_madd_odata_reg_137) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44321_ ( .CLK(CLK), .D(_00550_), .Q(__delay_data_671) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44322_ ( .CLK(CLK), .D(_00551_), .Q(__delay_data_672) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44323_ ( .CLK(CLK), .D(_00552_), .Q(__delay_data_673) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44324_ ( .CLK(CLK), .D(_00553_), .Q(__delay_data_674) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44325_ ( .CLK(CLK), .D(_02486_), .Q(_sra_data_138) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44326_ ( .CLK(CLK), .D(_01377_), .Q(__variable_wdata_122) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44327_ ( .CLK(CLK), .D(_01378_), .Q(__variable_wdata_123) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44328_ ( .CLK(CLK), .D(_01379_), .Q(__variable_wdata_124) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_7_x_data_cond_643_9_reg  ( .CLK(CLK), .D(_02838_), .Q(_substream_mul_7_x_data_cond_643_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_7_y_data_cond_643_10_reg  ( .CLK(CLK), .D(_02839_), .Q(_substream_mul_7_y_data_cond_643_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_7_rshift_data_cond_643_11_reg  ( .CLK(CLK), .D(_02837_), .Q(_substream_mul_7_rshift_data_cond_643_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greaterthan_data_108_reg  ( .CLK(CLK), .D(_01691_), .Q(_greaterthan_data_108) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44333_ ( .CLK(CLK), .D(_01800_), .Q(_minus_data_110) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44334_ ( .CLK(CLK), .D(_00527_), .Q(__delay_data_645) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44335_ ( .CLK(CLK), .D(_00530_), .Q(__delay_data_648) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44336_ ( .CLK(CLK), .D(_00533_), .Q(__delay_data_651) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(18) ) _44337_ ( .CLK(CLK), .D(_01874_), .Q(_sll_data_112) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_644_reg  ( .CLK(CLK), .D(_00526_), .Q(__delay_data_644) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44339_ ( .CLK(CLK), .D(_00528_), .Q(__delay_data_646) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44340_ ( .CLK(CLK), .D(_00531_), .Q(__delay_data_649) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44341_ ( .CLK(CLK), .D(_00534_), .Q(__delay_data_652) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44342_ ( .CLK(CLK), .D(_01468_), .Q(_cond_data_118) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44343_ ( .CLK(CLK), .D(_00529_), .Q(__delay_data_647) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44344_ ( .CLK(CLK), .D(_00532_), .Q(__delay_data_650) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44345_ ( .CLK(CLK), .D(_00535_), .Q(__delay_data_653) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44346_ ( .CLK(CLK), .D(_00693_), .Q(__muladd_madd_odata_reg_120) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44347_ ( .CLK(CLK), .D(_00536_), .Q(__delay_data_654) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44348_ ( .CLK(CLK), .D(_00537_), .Q(__delay_data_655) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44349_ ( .CLK(CLK), .D(_00538_), .Q(__delay_data_656) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44350_ ( .CLK(CLK), .D(_00539_), .Q(__delay_data_657) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44351_ ( .CLK(CLK), .D(_02485_), .Q(_sra_data_121) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44352_ ( .CLK(CLK), .D(_01374_), .Q(__variable_wdata_105) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44353_ ( .CLK(CLK), .D(_01375_), .Q(__variable_wdata_106) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44354_ ( .CLK(CLK), .D(_01376_), .Q(__variable_wdata_107) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_6_x_data_cond_626_6_reg  ( .CLK(CLK), .D(_02835_), .Q(_substream_mul_6_x_data_cond_626_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_6_y_data_cond_626_7_reg  ( .CLK(CLK), .D(_02836_), .Q(_substream_mul_6_y_data_cond_626_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_6_rshift_data_cond_626_8_reg  ( .CLK(CLK), .D(_02834_), .Q(_substream_mul_6_rshift_data_cond_626_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greaterthan_data_91_reg  ( .CLK(CLK), .D(_01702_), .Q(_greaterthan_data_91) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44359_ ( .CLK(CLK), .D(_01809_), .Q(_minus_data_93) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44360_ ( .CLK(CLK), .D(_00513_), .Q(__delay_data_628) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44361_ ( .CLK(CLK), .D(_00516_), .Q(__delay_data_631) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44362_ ( .CLK(CLK), .D(_00519_), .Q(__delay_data_634) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(18) ) _44363_ ( .CLK(CLK), .D(_01883_), .Q(_sll_data_95) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_627_reg  ( .CLK(CLK), .D(_00512_), .Q(__delay_data_627) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44365_ ( .CLK(CLK), .D(_00514_), .Q(__delay_data_629) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44366_ ( .CLK(CLK), .D(_00517_), .Q(__delay_data_632) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44367_ ( .CLK(CLK), .D(_00520_), .Q(__delay_data_635) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44368_ ( .CLK(CLK), .D(_01467_), .Q(_cond_data_101) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44369_ ( .CLK(CLK), .D(_00515_), .Q(__delay_data_630) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44370_ ( .CLK(CLK), .D(_00518_), .Q(__delay_data_633) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44371_ ( .CLK(CLK), .D(_00521_), .Q(__delay_data_636) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44372_ ( .CLK(CLK), .D(_00692_), .Q(__muladd_madd_odata_reg_103) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44373_ ( .CLK(CLK), .D(_00522_), .Q(__delay_data_637) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44374_ ( .CLK(CLK), .D(_00523_), .Q(__delay_data_638) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44375_ ( .CLK(CLK), .D(_00524_), .Q(__delay_data_639) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44376_ ( .CLK(CLK), .D(_00525_), .Q(__delay_data_640) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44377_ ( .CLK(CLK), .D(_02484_), .Q(_sra_data_104) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44378_ ( .CLK(CLK), .D(_01463_), .Q(__variable_wdata_88) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44379_ ( .CLK(CLK), .D(_01464_), .Q(__variable_wdata_89) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44380_ ( .CLK(CLK), .D(_01465_), .Q(__variable_wdata_90) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_5_x_data_cond_609_3_reg  ( .CLK(CLK), .D(_02832_), .Q(_substream_mul_5_x_data_cond_609_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_5_y_data_cond_609_4_reg  ( .CLK(CLK), .D(_02833_), .Q(_substream_mul_5_y_data_cond_609_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_5_rshift_data_cond_609_5_reg  ( .CLK(CLK), .D(_02831_), .Q(_substream_mul_5_rshift_data_cond_609_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greaterthan_data_74_reg  ( .CLK(CLK), .D(_01700_), .Q(_greaterthan_data_74) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44385_ ( .CLK(CLK), .D(_01808_), .Q(_minus_data_76) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44386_ ( .CLK(CLK), .D(_00499_), .Q(__delay_data_611) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44387_ ( .CLK(CLK), .D(_00502_), .Q(__delay_data_614) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44388_ ( .CLK(CLK), .D(_00505_), .Q(__delay_data_617) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(18) ) _44389_ ( .CLK(CLK), .D(_01881_), .Q(_sll_data_78) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_610_reg  ( .CLK(CLK), .D(_00498_), .Q(__delay_data_610) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44391_ ( .CLK(CLK), .D(_00500_), .Q(__delay_data_612) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44392_ ( .CLK(CLK), .D(_00503_), .Q(__delay_data_615) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44393_ ( .CLK(CLK), .D(_00506_), .Q(__delay_data_618) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44394_ ( .CLK(CLK), .D(_01554_), .Q(_cond_data_84) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44395_ ( .CLK(CLK), .D(_00501_), .Q(__delay_data_613) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44396_ ( .CLK(CLK), .D(_00504_), .Q(__delay_data_616) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44397_ ( .CLK(CLK), .D(_00507_), .Q(__delay_data_619) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44398_ ( .CLK(CLK), .D(_00700_), .Q(__muladd_madd_odata_reg_86) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44399_ ( .CLK(CLK), .D(_00508_), .Q(__delay_data_620) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44400_ ( .CLK(CLK), .D(_00509_), .Q(__delay_data_621) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44401_ ( .CLK(CLK), .D(_00510_), .Q(__delay_data_622) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44402_ ( .CLK(CLK), .D(_00511_), .Q(__delay_data_623) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44403_ ( .CLK(CLK), .D(_02494_), .Q(_sra_data_87) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44404_ ( .CLK(CLK), .D(_01442_), .Q(__variable_wdata_71) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44405_ ( .CLK(CLK), .D(_01443_), .Q(__variable_wdata_72) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44406_ ( .CLK(CLK), .D(_01444_), .Q(__variable_wdata_73) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_4_x_data_cond_592_0_reg  ( .CLK(CLK), .D(_02827_), .Q(_substream_mul_4_x_data_cond_592_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_4_y_data_cond_592_1_reg  ( .CLK(CLK), .D(_02829_), .Q(_substream_mul_4_y_data_cond_592_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_4_rshift_data_cond_592_2_reg  ( .CLK(CLK), .D(_02825_), .Q(_substream_mul_4_rshift_data_cond_592_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_4_x_data_cond_874_44_reg  ( .CLK(CLK), .D(_02828_), .Q(_substream_mul_4_x_data_cond_874_44) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_4_y_data_cond_874_45_reg  ( .CLK(CLK), .D(_02830_), .Q(_substream_mul_4_y_data_cond_874_45) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_4_rshift_data_cond_874_46_reg  ( .CLK(CLK), .D(_02826_), .Q(_substream_mul_4_rshift_data_cond_874_46) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greaterthan_data_57_reg  ( .CLK(CLK), .D(_01699_), .Q(_greaterthan_data_57) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44414_ ( .CLK(CLK), .D(_01806_), .Q(_minus_data_59) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44415_ ( .CLK(CLK), .D(_00485_), .Q(__delay_data_594) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44416_ ( .CLK(CLK), .D(_00488_), .Q(__delay_data_597) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44417_ ( .CLK(CLK), .D(_00491_), .Q(__delay_data_600) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(18) ) _44418_ ( .CLK(CLK), .D(_01880_), .Q(_sll_data_61) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_593_reg  ( .CLK(CLK), .D(_00484_), .Q(__delay_data_593) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44420_ ( .CLK(CLK), .D(_00486_), .Q(__delay_data_595) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44421_ ( .CLK(CLK), .D(_00489_), .Q(__delay_data_598) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44422_ ( .CLK(CLK), .D(_00492_), .Q(__delay_data_601) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44423_ ( .CLK(CLK), .D(_01546_), .Q(_cond_data_67) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44424_ ( .CLK(CLK), .D(_00487_), .Q(__delay_data_596) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44425_ ( .CLK(CLK), .D(_00490_), .Q(__delay_data_599) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44426_ ( .CLK(CLK), .D(_00493_), .Q(__delay_data_602) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44427_ ( .CLK(CLK), .D(_00699_), .Q(__muladd_madd_odata_reg_69) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44428_ ( .CLK(CLK), .D(_00494_), .Q(__delay_data_603) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44429_ ( .CLK(CLK), .D(_00495_), .Q(__delay_data_604) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44430_ ( .CLK(CLK), .D(_00496_), .Q(__delay_data_605) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44431_ ( .CLK(CLK), .D(_00497_), .Q(__delay_data_606) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _44432_ ( .CLK(CLK), .D(_02493_), .Q(_sra_data_70) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44433_ ( .CLK(CLK), .D(_01439_), .Q(__variable_wdata_54) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44434_ ( .CLK(CLK), .D(_01440_), .Q(__variable_wdata_55) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44435_ ( .CLK(CLK), .D(_01441_), .Q(__variable_wdata_56) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_rshift_clip_3_x_data_cond_763_39_reg  ( .CLK(CLK), .D(_02848_), .Q(_substream_mul_rshift_clip_3_x_data_cond_763_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_rshift_clip_3_y_data_cond_763_40_reg  ( .CLK(CLK), .D(_02850_), .Q(_substream_mul_rshift_clip_3_y_data_cond_763_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_rshift_clip_3_rshift_data_cond_763_41_reg  ( .CLK(CLK), .D(_02846_), .Q(_substream_mul_rshift_clip_3_rshift_data_cond_763_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_rshift_clip_3_x_data_cond_884_51_reg  ( .CLK(CLK), .D(_02849_), .Q(_substream_mul_rshift_clip_3_x_data_cond_884_51) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_rshift_clip_3_y_data_cond_884_52_reg  ( .CLK(CLK), .D(_02851_), .Q(_substream_mul_rshift_clip_3_y_data_cond_884_52) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_mul_rshift_clip_3_rshift_data_cond_884_53_reg  ( .CLK(CLK), .D(_02847_), .Q(_substream_mul_rshift_clip_3_rshift_data_cond_884_53) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(40) ) _44442_ ( .CLK(CLK), .D(_02852_), .Q(_times_mul_odata_reg_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _44443_ ( .CLK(CLK), .D(_00621_), .Q(__delay_data_764) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _44444_ ( .CLK(CLK), .D(_00622_), .Q(__delay_data_765) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _44445_ ( .CLK(CLK), .D(_00623_), .Q(__delay_data_766) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _44446_ ( .CLK(CLK), .D(_00624_), .Q(__delay_data_767) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(40) ) _44447_ ( .CLK(CLK), .D(_02492_), .Q(_sra_data_42) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greaterthan_data_43_reg  ( .CLK(CLK), .D(_01698_), .Q(_greaterthan_data_43) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _lessthan_data_47_reg  ( .CLK(CLK), .D(_01703_), .Q(_lessthan_data_47) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greatereq_data_51_reg  ( .CLK(CLK), .D(_01690_), .Q(_greatereq_data_51) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(40) ) _44451_ ( .CLK(CLK), .D(_00625_), .Q(__delay_data_768) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(40) ) _44452_ ( .CLK(CLK), .D(_01534_), .Q(_cond_data_45) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(40) ) _44453_ ( .CLK(CLK), .D(_01535_), .Q(_cond_data_49) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_769_reg  ( .CLK(CLK), .D(_00626_), .Q(__delay_data_769) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44455_ ( .CLK(CLK), .D(_01536_), .Q(_cond_data_53) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44456_ ( .CLK(CLK), .D(_01427_), .Q(__variable_wdata_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44457_ ( .CLK(CLK), .D(_01428_), .Q(__variable_wdata_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _44458_ ( .CLK(CLK), .D(_01429_), .Q(__variable_wdata_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_959_10_reg  ( .CLK(CLK), .D(_01332_), .Q(__tmp_959_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_959_11_reg  ( .CLK(CLK), .D(_01333_), .Q(__tmp_959_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_959_12_reg  ( .CLK(CLK), .D(_01334_), .Q(__tmp_959_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_add_tree_2_var0_data_cond_745_27_reg  ( .CLK(CLK), .D(_02807_), .Q(_substream_add_tree_2_var0_data_cond_745_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_add_tree_2_var1_data_cond_745_28_reg  ( .CLK(CLK), .D(_02808_), .Q(_substream_add_tree_2_var1_data_cond_745_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_add_tree_2_var2_data_cond_745_29_reg  ( .CLK(CLK), .D(_02809_), .Q(_substream_add_tree_2_var2_data_cond_745_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_add_tree_2_var3_data_cond_745_30_reg  ( .CLK(CLK), .D(_02810_), .Q(_substream_add_tree_2_var3_data_cond_745_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_add_tree_2_var4_data_cond_745_31_reg  ( .CLK(CLK), .D(_02811_), .Q(_substream_add_tree_2_var4_data_cond_745_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_add_tree_2_var5_data_cond_745_32_reg  ( .CLK(CLK), .D(_02812_), .Q(_substream_add_tree_2_var5_data_cond_745_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_add_tree_2_var6_data_cond_745_33_reg  ( .CLK(CLK), .D(_02813_), .Q(_substream_add_tree_2_var6_data_cond_745_33) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_add_tree_2_var7_data_cond_745_34_reg  ( .CLK(CLK), .D(_02814_), .Q(_substream_add_tree_2_var7_data_cond_745_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_add_tree_2_var8_data_cond_745_35_reg  ( .CLK(CLK), .D(_02815_), .Q(_substream_add_tree_2_var8_data_cond_745_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44471_ ( .CLK(CLK), .D(_00701_), .Q(__plusn_data_34) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44472_ ( .CLK(CLK), .D(_00702_), .Q(__plusn_data_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44473_ ( .CLK(CLK), .D(_00703_), .Q(__plusn_data_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44474_ ( .CLK(CLK), .D(_00704_), .Q(__plusn_data_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44475_ ( .CLK(CLK), .D(_01403_), .Q(__variable_wdata_24) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44476_ ( .CLK(CLK), .D(_01406_), .Q(__variable_wdata_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44477_ ( .CLK(CLK), .D(_01412_), .Q(__variable_wdata_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44478_ ( .CLK(CLK), .D(_01420_), .Q(__variable_wdata_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44479_ ( .CLK(CLK), .D(_01421_), .Q(__variable_wdata_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44480_ ( .CLK(CLK), .D(_01422_), .Q(__variable_wdata_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44481_ ( .CLK(CLK), .D(_01424_), .Q(__variable_wdata_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44482_ ( .CLK(CLK), .D(_01425_), .Q(__variable_wdata_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44483_ ( .CLK(CLK), .D(_01426_), .Q(__variable_wdata_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_add_tree_1_var0_data_cond_877_47_reg  ( .CLK(CLK), .D(_02806_), .Q(_substream_add_tree_1_var0_data_cond_877_47) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44485_ ( .CLK(CLK), .D(_01399_), .Q(__variable_wdata_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _acc_0_reduce_reset_reg  ( .CLK(CLK), .D(_01466_), .Q(_acc_0_reduce_reset) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_acc_0_x_data_cond_747_36_reg  ( .CLK(CLK), .D(_02804_), .Q(_substream_acc_0_x_data_cond_747_36) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_acc_0_rshift_data_cond_747_37_reg  ( .CLK(CLK), .D(_02800_), .Q(_substream_acc_0_rshift_data_cond_747_37) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_acc_0_size_data_cond_747_38_reg  ( .CLK(CLK), .D(_02802_), .Q(_substream_acc_0_size_data_cond_747_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_acc_0_x_data_cond_879_48_reg  ( .CLK(CLK), .D(_02805_), .Q(_substream_acc_0_x_data_cond_879_48) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_acc_0_rshift_data_cond_879_49_reg  ( .CLK(CLK), .D(_02801_), .Q(_substream_acc_0_rshift_data_cond_879_49) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _substream_acc_0_size_data_cond_879_50_reg  ( .CLK(CLK), .D(_02803_), .Q(_substream_acc_0_size_data_cond_879_50) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _greaterthan_data_3_reg  ( .CLK(CLK), .D(_01697_), .Q(_greaterthan_data_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _44494_ ( .CLK(CLK), .D(_01807_), .Q(_minus_data_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44495_ ( .CLK(CLK), .D(_01838_), .Q(_reduceadd_data_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44496_ ( .CLK(CLK), .D(_01837_), .Q(_reduceadd_count_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _pulse_data_19_reg  ( .CLK(CLK), .D(_01822_), .Q(_pulse_data_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _44498_ ( .CLK(CLK), .D(_01820_), .Q(_pulse_count_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _44499_ ( .CLK(CLK), .D(_00613_), .Q(__delay_data_751) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(66) ) _44500_ ( .CLK(CLK), .D(_01882_), .Q(_sll_data_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_748_reg  ( .CLK(CLK), .D(_00610_), .Q(__delay_data_748) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44502_ ( .CLK(CLK), .D(_00611_), .Q(__delay_data_749) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _44503_ ( .CLK(CLK), .D(_00614_), .Q(__delay_data_752) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_755_reg  ( .CLK(CLK), .D(_00617_), .Q(__delay_data_755) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44505_ ( .CLK(CLK), .D(_01470_), .Q(_cond_data_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44506_ ( .CLK(CLK), .D(_00612_), .Q(__delay_data_750) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _44507_ ( .CLK(CLK), .D(_00615_), .Q(__delay_data_753) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_756_reg  ( .CLK(CLK), .D(_00618_), .Q(__delay_data_756) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44509_ ( .CLK(CLK), .D(_01810_), .Q(_plus_data_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _44510_ ( .CLK(CLK), .D(_00616_), .Q(__delay_data_754) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_757_reg  ( .CLK(CLK), .D(_00619_), .Q(__delay_data_757) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44512_ ( .CLK(CLK), .D(_02491_), .Q(_sra_data_21) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __delay_data_758_reg  ( .CLK(CLK), .D(_00620_), .Q(__delay_data_758) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44514_ ( .CLK(CLK), .D(_01373_), .Q(__variable_wdata_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _44515_ ( .CLK(CLK), .D(_01392_), .Q(__variable_wdata_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44516_ ( .CLK(CLK), .D(_01423_), .Q(__variable_wdata_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_947_1_reg  ( .CLK(CLK), .D(_01323_), .Q(__tmp_947_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_947_2_reg  ( .CLK(CLK), .D(_01324_), .Q(__tmp_947_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_947_3_reg  ( .CLK(CLK), .D(_01325_), .Q(__tmp_947_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_947_4_reg  ( .CLK(CLK), .D(_01326_), .Q(__tmp_947_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_947_5_reg  ( .CLK(CLK), .D(_01327_), .Q(__tmp_947_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_947_6_reg  ( .CLK(CLK), .D(_01328_), .Q(__tmp_947_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_947_7_reg  ( .CLK(CLK), .D(_01329_), .Q(__tmp_947_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_947_8_reg  ( .CLK(CLK), .D(_01330_), .Q(__tmp_947_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_947_9_reg  ( .CLK(CLK), .D(_01331_), .Q(__tmp_947_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44526_ ( .CLK(CLK), .D(_03713_), .Q(ram_w8_l2048_id11_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44527_ ( .CLK(CLK), .D(_03714_), .Q(ram_w8_l2048_id11_3_0_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id11_3_0_wenable_reg  ( .CLK(CLK), .D(_03715_), .Q(ram_w8_l2048_id11_3_0_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44529_ ( .CLK(CLK), .D(_03716_), .Q(ram_w8_l2048_id11_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id11_3_cond_0_1_reg  ( .CLK(CLK), .D(_01832_), .Q(_ram_w8_l2048_id11_3_cond_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1007_reg  ( .CLK(CLK), .D(_02859_), .Q(_tmp_1007) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1012_1_reg  ( .CLK(CLK), .D(_01107_), .Q(__tmp_1012_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44533_ ( .CLK(CLK), .D(_01108_), .Q(__tmp_1013_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1014_reg  ( .CLK(CLK), .D(_02861_), .Q(_tmp_1014) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1015_reg  ( .CLK(CLK), .D(_02862_), .Q(_tmp_1015) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1016_reg  ( .CLK(CLK), .D(_02863_), .Q(_tmp_1016) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1017_reg  ( .CLK(CLK), .D(_02864_), .Q(_tmp_1017) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44538_ ( .CLK(CLK), .D(_02865_), .Q(_tmp_1018) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44539_ ( .CLK(CLK), .D(_03709_), .Q(ram_w8_l2048_id11_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44540_ ( .CLK(CLK), .D(_03710_), .Q(ram_w8_l2048_id11_2_0_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id11_2_0_wenable_reg  ( .CLK(CLK), .D(_03711_), .Q(ram_w8_l2048_id11_2_0_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44542_ ( .CLK(CLK), .D(_03712_), .Q(ram_w8_l2048_id11_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id11_2_cond_0_1_reg  ( .CLK(CLK), .D(_01831_), .Q(_ram_w8_l2048_id11_2_cond_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_995_reg  ( .CLK(CLK), .D(_03170_), .Q(_tmp_995) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1000_1_reg  ( .CLK(CLK), .D(_01105_), .Q(__tmp_1000_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44546_ ( .CLK(CLK), .D(_01106_), .Q(__tmp_1001_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1002_reg  ( .CLK(CLK), .D(_02854_), .Q(_tmp_1002) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1003_reg  ( .CLK(CLK), .D(_02855_), .Q(_tmp_1003) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1004_reg  ( .CLK(CLK), .D(_02856_), .Q(_tmp_1004) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1005_reg  ( .CLK(CLK), .D(_02857_), .Q(_tmp_1005) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44551_ ( .CLK(CLK), .D(_02858_), .Q(_tmp_1006) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44552_ ( .CLK(CLK), .D(_03705_), .Q(ram_w8_l2048_id11_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44553_ ( .CLK(CLK), .D(_03706_), .Q(ram_w8_l2048_id11_1_0_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id11_1_0_wenable_reg  ( .CLK(CLK), .D(_03707_), .Q(ram_w8_l2048_id11_1_0_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44555_ ( .CLK(CLK), .D(_03708_), .Q(ram_w8_l2048_id11_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id11_1_cond_0_1_reg  ( .CLK(CLK), .D(_01830_), .Q(_ram_w8_l2048_id11_1_cond_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_983_reg  ( .CLK(CLK), .D(_03164_), .Q(_tmp_983) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_988_1_reg  ( .CLK(CLK), .D(_01371_), .Q(__tmp_988_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44559_ ( .CLK(CLK), .D(_01372_), .Q(__tmp_989_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_990_reg  ( .CLK(CLK), .D(_03165_), .Q(_tmp_990) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_991_reg  ( .CLK(CLK), .D(_03166_), .Q(_tmp_991) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_992_reg  ( .CLK(CLK), .D(_03167_), .Q(_tmp_992) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_993_reg  ( .CLK(CLK), .D(_03168_), .Q(_tmp_993) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44564_ ( .CLK(CLK), .D(_03169_), .Q(_tmp_994) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44565_ ( .CLK(CLK), .D(_01588_), .Q(_dataflow_cat_data_98) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_cat_valid_98_reg  ( .CLK(CLK), .D(_01591_), .Q(_dataflow_cat_valid_98) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44567_ ( .CLK(CLK), .D(_03701_), .Q(ram_w8_l2048_id11_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44568_ ( .CLK(CLK), .D(_03702_), .Q(ram_w8_l2048_id11_0_0_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id11_0_0_wenable_reg  ( .CLK(CLK), .D(_03703_), .Q(ram_w8_l2048_id11_0_0_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44570_ ( .CLK(CLK), .D(_03704_), .Q(ram_w8_l2048_id11_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id11_0_cond_0_1_reg  ( .CLK(CLK), .D(_01829_), .Q(_ram_w8_l2048_id11_0_cond_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_971_reg  ( .CLK(CLK), .D(_03158_), .Q(_tmp_971) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_976_1_reg  ( .CLK(CLK), .D(_01369_), .Q(__tmp_976_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44574_ ( .CLK(CLK), .D(_01370_), .Q(__tmp_977_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_978_reg  ( .CLK(CLK), .D(_03159_), .Q(_tmp_978) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_979_reg  ( .CLK(CLK), .D(_03160_), .Q(_tmp_979) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_980_reg  ( .CLK(CLK), .D(_03161_), .Q(_tmp_980) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_981_reg  ( .CLK(CLK), .D(_03162_), .Q(_tmp_981) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44579_ ( .CLK(CLK), .D(_03163_), .Q(_tmp_982) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44580_ ( .CLK(CLK), .D(_03697_), .Q(ram_w8_l2048_id10_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44581_ ( .CLK(CLK), .D(_03698_), .Q(ram_w8_l2048_id10_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44582_ ( .CLK(CLK), .D(_03699_), .Q(ram_w8_l2048_id10_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id10_3_1_wenable_reg  ( .CLK(CLK), .D(_03700_), .Q(ram_w8_l2048_id10_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44584_ ( .CLK(CLK), .D(_03693_), .Q(ram_w8_l2048_id10_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44585_ ( .CLK(CLK), .D(_03694_), .Q(ram_w8_l2048_id10_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44586_ ( .CLK(CLK), .D(_03695_), .Q(ram_w8_l2048_id10_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id10_2_1_wenable_reg  ( .CLK(CLK), .D(_03696_), .Q(ram_w8_l2048_id10_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44588_ ( .CLK(CLK), .D(_03689_), .Q(ram_w8_l2048_id10_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44589_ ( .CLK(CLK), .D(_03690_), .Q(ram_w8_l2048_id10_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44590_ ( .CLK(CLK), .D(_03691_), .Q(ram_w8_l2048_id10_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id10_1_1_wenable_reg  ( .CLK(CLK), .D(_03692_), .Q(ram_w8_l2048_id10_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44592_ ( .CLK(CLK), .D(_03685_), .Q(ram_w8_l2048_id10_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44593_ ( .CLK(CLK), .D(_03686_), .Q(ram_w8_l2048_id10_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44594_ ( .CLK(CLK), .D(_03687_), .Q(ram_w8_l2048_id10_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id10_0_1_wenable_reg  ( .CLK(CLK), .D(_03688_), .Q(ram_w8_l2048_id10_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id10_0_cond_2_1_reg  ( .CLK(CLK), .D(_01261_), .Q(_ram_w8_l2048_id10_0_cond_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44597_ ( .CLK(CLK), .D(_03865_), .Q(ram_w8_l2048_id9_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44598_ ( .CLK(CLK), .D(_03866_), .Q(ram_w8_l2048_id9_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44599_ ( .CLK(CLK), .D(_03867_), .Q(ram_w8_l2048_id9_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id9_3_1_wenable_reg  ( .CLK(CLK), .D(_03868_), .Q(ram_w8_l2048_id9_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44601_ ( .CLK(CLK), .D(_03861_), .Q(ram_w8_l2048_id9_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44602_ ( .CLK(CLK), .D(_03862_), .Q(ram_w8_l2048_id9_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44603_ ( .CLK(CLK), .D(_03863_), .Q(ram_w8_l2048_id9_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id9_2_1_wenable_reg  ( .CLK(CLK), .D(_03864_), .Q(ram_w8_l2048_id9_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44605_ ( .CLK(CLK), .D(_03857_), .Q(ram_w8_l2048_id9_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44606_ ( .CLK(CLK), .D(_03858_), .Q(ram_w8_l2048_id9_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44607_ ( .CLK(CLK), .D(_03859_), .Q(ram_w8_l2048_id9_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id9_1_1_wenable_reg  ( .CLK(CLK), .D(_03860_), .Q(ram_w8_l2048_id9_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44609_ ( .CLK(CLK), .D(_03853_), .Q(ram_w8_l2048_id9_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44610_ ( .CLK(CLK), .D(_03854_), .Q(ram_w8_l2048_id9_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44611_ ( .CLK(CLK), .D(_03855_), .Q(ram_w8_l2048_id9_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id9_0_1_wenable_reg  ( .CLK(CLK), .D(_03856_), .Q(ram_w8_l2048_id9_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id9_0_cond_2_1_reg  ( .CLK(CLK), .D(_01258_), .Q(_ram_w8_l2048_id9_0_cond_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44614_ ( .CLK(CLK), .D(_03849_), .Q(ram_w8_l2048_id8_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44615_ ( .CLK(CLK), .D(_03850_), .Q(ram_w8_l2048_id8_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44616_ ( .CLK(CLK), .D(_03851_), .Q(ram_w8_l2048_id8_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id8_3_1_wenable_reg  ( .CLK(CLK), .D(_03852_), .Q(ram_w8_l2048_id8_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44618_ ( .CLK(CLK), .D(_03130_), .Q(_tmp_444) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44619_ ( .CLK(CLK), .D(_03131_), .Q(_tmp_445) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_446_reg  ( .CLK(CLK), .D(_03132_), .Q(_tmp_446) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44621_ ( .CLK(CLK), .D(_03133_), .Q(_tmp_447) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44622_ ( .CLK(CLK), .D(_03134_), .Q(_tmp_448) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44623_ ( .CLK(CLK), .D(_03135_), .Q(_tmp_449) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _44624_ ( .CLK(CLK), .D(_03137_), .Q(_tmp_456) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44625_ ( .CLK(CLK), .D(_03845_), .Q(ram_w8_l2048_id8_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44626_ ( .CLK(CLK), .D(_03846_), .Q(ram_w8_l2048_id8_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44627_ ( .CLK(CLK), .D(_03847_), .Q(ram_w8_l2048_id8_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id8_2_1_wenable_reg  ( .CLK(CLK), .D(_03848_), .Q(ram_w8_l2048_id8_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44629_ ( .CLK(CLK), .D(_03122_), .Q(_tmp_431) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44630_ ( .CLK(CLK), .D(_03123_), .Q(_tmp_432) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_433_reg  ( .CLK(CLK), .D(_03124_), .Q(_tmp_433) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44632_ ( .CLK(CLK), .D(_03125_), .Q(_tmp_434) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44633_ ( .CLK(CLK), .D(_03126_), .Q(_tmp_435) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44634_ ( .CLK(CLK), .D(_03127_), .Q(_tmp_436) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _44635_ ( .CLK(CLK), .D(_03129_), .Q(_tmp_443) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44636_ ( .CLK(CLK), .D(_03841_), .Q(ram_w8_l2048_id8_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44637_ ( .CLK(CLK), .D(_03842_), .Q(ram_w8_l2048_id8_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44638_ ( .CLK(CLK), .D(_03843_), .Q(ram_w8_l2048_id8_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id8_1_1_wenable_reg  ( .CLK(CLK), .D(_03844_), .Q(ram_w8_l2048_id8_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44640_ ( .CLK(CLK), .D(_03113_), .Q(_tmp_418) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44641_ ( .CLK(CLK), .D(_03114_), .Q(_tmp_419) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_420_reg  ( .CLK(CLK), .D(_03116_), .Q(_tmp_420) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44643_ ( .CLK(CLK), .D(_03117_), .Q(_tmp_421) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44644_ ( .CLK(CLK), .D(_03118_), .Q(_tmp_422) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44645_ ( .CLK(CLK), .D(_03119_), .Q(_tmp_423) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _44646_ ( .CLK(CLK), .D(_03121_), .Q(_tmp_430) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44647_ ( .CLK(CLK), .D(_03837_), .Q(ram_w8_l2048_id8_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44648_ ( .CLK(CLK), .D(_03838_), .Q(ram_w8_l2048_id8_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44649_ ( .CLK(CLK), .D(_03839_), .Q(ram_w8_l2048_id8_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id8_0_1_wenable_reg  ( .CLK(CLK), .D(_03840_), .Q(ram_w8_l2048_id8_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44651_ ( .CLK(CLK), .D(_03105_), .Q(_tmp_405) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44652_ ( .CLK(CLK), .D(_03106_), .Q(_tmp_406) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_407_reg  ( .CLK(CLK), .D(_03107_), .Q(_tmp_407) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44654_ ( .CLK(CLK), .D(_03108_), .Q(_tmp_408) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44655_ ( .CLK(CLK), .D(_03109_), .Q(_tmp_409) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44656_ ( .CLK(CLK), .D(_03111_), .Q(_tmp_410) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _44657_ ( .CLK(CLK), .D(_03112_), .Q(_tmp_417) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id8_0_cond_3_1_reg  ( .CLK(CLK), .D(_01255_), .Q(_ram_w8_l2048_id8_0_cond_3_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44659_ ( .CLK(CLK), .D(_03833_), .Q(ram_w8_l2048_id7_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44660_ ( .CLK(CLK), .D(_03834_), .Q(ram_w8_l2048_id7_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44661_ ( .CLK(CLK), .D(_03835_), .Q(ram_w8_l2048_id7_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id7_3_1_wenable_reg  ( .CLK(CLK), .D(_03836_), .Q(ram_w8_l2048_id7_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44663_ ( .CLK(CLK), .D(_03829_), .Q(ram_w8_l2048_id7_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44664_ ( .CLK(CLK), .D(_03830_), .Q(ram_w8_l2048_id7_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44665_ ( .CLK(CLK), .D(_03831_), .Q(ram_w8_l2048_id7_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id7_2_1_wenable_reg  ( .CLK(CLK), .D(_03832_), .Q(ram_w8_l2048_id7_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44667_ ( .CLK(CLK), .D(_03825_), .Q(ram_w8_l2048_id7_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44668_ ( .CLK(CLK), .D(_03826_), .Q(ram_w8_l2048_id7_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44669_ ( .CLK(CLK), .D(_03827_), .Q(ram_w8_l2048_id7_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id7_1_1_wenable_reg  ( .CLK(CLK), .D(_03828_), .Q(ram_w8_l2048_id7_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44671_ ( .CLK(CLK), .D(_03821_), .Q(ram_w8_l2048_id7_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44672_ ( .CLK(CLK), .D(_03822_), .Q(ram_w8_l2048_id7_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44673_ ( .CLK(CLK), .D(_03823_), .Q(ram_w8_l2048_id7_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id7_0_1_wenable_reg  ( .CLK(CLK), .D(_03824_), .Q(ram_w8_l2048_id7_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id7_0_cond_2_1_reg  ( .CLK(CLK), .D(_01252_), .Q(_ram_w8_l2048_id7_0_cond_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44676_ ( .CLK(CLK), .D(_03817_), .Q(ram_w8_l2048_id6_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44677_ ( .CLK(CLK), .D(_03818_), .Q(ram_w8_l2048_id6_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44678_ ( .CLK(CLK), .D(_03819_), .Q(ram_w8_l2048_id6_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id6_3_1_wenable_reg  ( .CLK(CLK), .D(_03820_), .Q(ram_w8_l2048_id6_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44680_ ( .CLK(CLK), .D(_03813_), .Q(ram_w8_l2048_id6_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44681_ ( .CLK(CLK), .D(_03814_), .Q(ram_w8_l2048_id6_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44682_ ( .CLK(CLK), .D(_03815_), .Q(ram_w8_l2048_id6_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id6_2_1_wenable_reg  ( .CLK(CLK), .D(_03816_), .Q(ram_w8_l2048_id6_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44684_ ( .CLK(CLK), .D(_03809_), .Q(ram_w8_l2048_id6_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44685_ ( .CLK(CLK), .D(_03810_), .Q(ram_w8_l2048_id6_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44686_ ( .CLK(CLK), .D(_03811_), .Q(ram_w8_l2048_id6_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id6_1_1_wenable_reg  ( .CLK(CLK), .D(_03812_), .Q(ram_w8_l2048_id6_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44688_ ( .CLK(CLK), .D(_03805_), .Q(ram_w8_l2048_id6_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44689_ ( .CLK(CLK), .D(_03806_), .Q(ram_w8_l2048_id6_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44690_ ( .CLK(CLK), .D(_03807_), .Q(ram_w8_l2048_id6_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id6_0_1_wenable_reg  ( .CLK(CLK), .D(_03808_), .Q(ram_w8_l2048_id6_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id6_0_cond_2_1_reg  ( .CLK(CLK), .D(_01249_), .Q(_ram_w8_l2048_id6_0_cond_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44693_ ( .CLK(CLK), .D(_03801_), .Q(ram_w8_l2048_id5_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44694_ ( .CLK(CLK), .D(_03802_), .Q(ram_w8_l2048_id5_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44695_ ( .CLK(CLK), .D(_03803_), .Q(ram_w8_l2048_id5_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id5_3_1_wenable_reg  ( .CLK(CLK), .D(_03804_), .Q(ram_w8_l2048_id5_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44697_ ( .CLK(CLK), .D(_03095_), .Q(_tmp_387) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44698_ ( .CLK(CLK), .D(_03096_), .Q(_tmp_388) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_389_reg  ( .CLK(CLK), .D(_03097_), .Q(_tmp_389) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44700_ ( .CLK(CLK), .D(_03099_), .Q(_tmp_390) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44701_ ( .CLK(CLK), .D(_03100_), .Q(_tmp_391) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44702_ ( .CLK(CLK), .D(_03101_), .Q(_tmp_392) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _44703_ ( .CLK(CLK), .D(_03102_), .Q(_tmp_399) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44704_ ( .CLK(CLK), .D(_03797_), .Q(ram_w8_l2048_id5_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44705_ ( .CLK(CLK), .D(_03798_), .Q(ram_w8_l2048_id5_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44706_ ( .CLK(CLK), .D(_03799_), .Q(ram_w8_l2048_id5_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id5_2_1_wenable_reg  ( .CLK(CLK), .D(_03800_), .Q(ram_w8_l2048_id5_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44708_ ( .CLK(CLK), .D(_03088_), .Q(_tmp_374) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44709_ ( .CLK(CLK), .D(_03089_), .Q(_tmp_375) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_376_reg  ( .CLK(CLK), .D(_03090_), .Q(_tmp_376) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44711_ ( .CLK(CLK), .D(_03091_), .Q(_tmp_377) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44712_ ( .CLK(CLK), .D(_03092_), .Q(_tmp_378) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44713_ ( .CLK(CLK), .D(_03093_), .Q(_tmp_379) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _44714_ ( .CLK(CLK), .D(_03094_), .Q(_tmp_386) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44715_ ( .CLK(CLK), .D(_03793_), .Q(ram_w8_l2048_id5_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44716_ ( .CLK(CLK), .D(_03794_), .Q(ram_w8_l2048_id5_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44717_ ( .CLK(CLK), .D(_03795_), .Q(ram_w8_l2048_id5_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id5_1_1_wenable_reg  ( .CLK(CLK), .D(_03796_), .Q(ram_w8_l2048_id5_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44719_ ( .CLK(CLK), .D(_03081_), .Q(_tmp_361) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44720_ ( .CLK(CLK), .D(_03082_), .Q(_tmp_362) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_363_reg  ( .CLK(CLK), .D(_03083_), .Q(_tmp_363) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44722_ ( .CLK(CLK), .D(_03084_), .Q(_tmp_364) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44723_ ( .CLK(CLK), .D(_03085_), .Q(_tmp_365) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44724_ ( .CLK(CLK), .D(_03086_), .Q(_tmp_366) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _44725_ ( .CLK(CLK), .D(_03087_), .Q(_tmp_373) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44726_ ( .CLK(CLK), .D(_03789_), .Q(ram_w8_l2048_id5_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44727_ ( .CLK(CLK), .D(_03790_), .Q(ram_w8_l2048_id5_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44728_ ( .CLK(CLK), .D(_03791_), .Q(ram_w8_l2048_id5_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id5_0_1_wenable_reg  ( .CLK(CLK), .D(_03792_), .Q(ram_w8_l2048_id5_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44730_ ( .CLK(CLK), .D(_03074_), .Q(_tmp_348) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44731_ ( .CLK(CLK), .D(_03075_), .Q(_tmp_349) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_350_reg  ( .CLK(CLK), .D(_03076_), .Q(_tmp_350) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44733_ ( .CLK(CLK), .D(_03077_), .Q(_tmp_351) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44734_ ( .CLK(CLK), .D(_03078_), .Q(_tmp_352) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44735_ ( .CLK(CLK), .D(_03079_), .Q(_tmp_353) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _44736_ ( .CLK(CLK), .D(_03080_), .Q(_tmp_360) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id5_0_cond_3_1_reg  ( .CLK(CLK), .D(_01246_), .Q(_ram_w8_l2048_id5_0_cond_3_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44738_ ( .CLK(CLK), .D(_03785_), .Q(ram_w8_l2048_id4_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44739_ ( .CLK(CLK), .D(_03786_), .Q(ram_w8_l2048_id4_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44740_ ( .CLK(CLK), .D(_03787_), .Q(ram_w8_l2048_id4_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id4_3_1_wenable_reg  ( .CLK(CLK), .D(_03788_), .Q(ram_w8_l2048_id4_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44742_ ( .CLK(CLK), .D(_03781_), .Q(ram_w8_l2048_id4_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44743_ ( .CLK(CLK), .D(_03782_), .Q(ram_w8_l2048_id4_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44744_ ( .CLK(CLK), .D(_03783_), .Q(ram_w8_l2048_id4_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id4_2_1_wenable_reg  ( .CLK(CLK), .D(_03784_), .Q(ram_w8_l2048_id4_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44746_ ( .CLK(CLK), .D(_03777_), .Q(ram_w8_l2048_id4_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44747_ ( .CLK(CLK), .D(_03778_), .Q(ram_w8_l2048_id4_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44748_ ( .CLK(CLK), .D(_03779_), .Q(ram_w8_l2048_id4_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id4_1_1_wenable_reg  ( .CLK(CLK), .D(_03780_), .Q(ram_w8_l2048_id4_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44750_ ( .CLK(CLK), .D(_03773_), .Q(ram_w8_l2048_id4_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44751_ ( .CLK(CLK), .D(_03774_), .Q(ram_w8_l2048_id4_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44752_ ( .CLK(CLK), .D(_03775_), .Q(ram_w8_l2048_id4_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id4_0_1_wenable_reg  ( .CLK(CLK), .D(_03776_), .Q(ram_w8_l2048_id4_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id4_0_cond_2_1_reg  ( .CLK(CLK), .D(_01243_), .Q(_ram_w8_l2048_id4_0_cond_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44755_ ( .CLK(CLK), .D(_03769_), .Q(ram_w8_l2048_id3_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44756_ ( .CLK(CLK), .D(_03770_), .Q(ram_w8_l2048_id3_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44757_ ( .CLK(CLK), .D(_03771_), .Q(ram_w8_l2048_id3_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id3_3_1_wenable_reg  ( .CLK(CLK), .D(_03772_), .Q(ram_w8_l2048_id3_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44759_ ( .CLK(CLK), .D(_02934_), .Q(_tmp_1161) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1162_reg  ( .CLK(CLK), .D(_02935_), .Q(_tmp_1162) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44761_ ( .CLK(CLK), .D(_03765_), .Q(ram_w8_l2048_id3_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44762_ ( .CLK(CLK), .D(_03766_), .Q(ram_w8_l2048_id3_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44763_ ( .CLK(CLK), .D(_03767_), .Q(ram_w8_l2048_id3_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id3_2_1_wenable_reg  ( .CLK(CLK), .D(_03768_), .Q(ram_w8_l2048_id3_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44765_ ( .CLK(CLK), .D(_02932_), .Q(_tmp_1159) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1160_reg  ( .CLK(CLK), .D(_02933_), .Q(_tmp_1160) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44767_ ( .CLK(CLK), .D(_03761_), .Q(ram_w8_l2048_id3_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44768_ ( .CLK(CLK), .D(_03762_), .Q(ram_w8_l2048_id3_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44769_ ( .CLK(CLK), .D(_03763_), .Q(ram_w8_l2048_id3_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id3_1_1_wenable_reg  ( .CLK(CLK), .D(_03764_), .Q(ram_w8_l2048_id3_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44771_ ( .CLK(CLK), .D(_02930_), .Q(_tmp_1157) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1158_reg  ( .CLK(CLK), .D(_02931_), .Q(_tmp_1158) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44773_ ( .CLK(CLK), .D(_03757_), .Q(ram_w8_l2048_id3_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44774_ ( .CLK(CLK), .D(_03758_), .Q(ram_w8_l2048_id3_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44775_ ( .CLK(CLK), .D(_03759_), .Q(ram_w8_l2048_id3_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id3_0_1_wenable_reg  ( .CLK(CLK), .D(_03760_), .Q(ram_w8_l2048_id3_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id3_0_cond_2_1_reg  ( .CLK(CLK), .D(_01240_), .Q(_ram_w8_l2048_id3_0_cond_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44778_ ( .CLK(CLK), .D(_02928_), .Q(_tmp_1155) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1156_reg  ( .CLK(CLK), .D(_02929_), .Q(_tmp_1156) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id3_0_cond_5_1_reg  ( .CLK(CLK), .D(_01147_), .Q(_ram_w8_l2048_id3_0_cond_5_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44781_ ( .CLK(CLK), .D(_03753_), .Q(ram_w8_l2048_id2_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44782_ ( .CLK(CLK), .D(_03754_), .Q(ram_w8_l2048_id2_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44783_ ( .CLK(CLK), .D(_03755_), .Q(ram_w8_l2048_id2_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id2_3_1_wenable_reg  ( .CLK(CLK), .D(_03756_), .Q(ram_w8_l2048_id2_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44785_ ( .CLK(CLK), .D(_03067_), .Q(_tmp_330) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44786_ ( .CLK(CLK), .D(_03068_), .Q(_tmp_331) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_332_reg  ( .CLK(CLK), .D(_03069_), .Q(_tmp_332) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44788_ ( .CLK(CLK), .D(_03070_), .Q(_tmp_333) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44789_ ( .CLK(CLK), .D(_03071_), .Q(_tmp_334) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44790_ ( .CLK(CLK), .D(_03072_), .Q(_tmp_335) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _44791_ ( .CLK(CLK), .D(_03073_), .Q(_tmp_342) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44792_ ( .CLK(CLK), .D(_02910_), .Q(_tmp_1130) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1131_reg  ( .CLK(CLK), .D(_02911_), .Q(_tmp_1131) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44794_ ( .CLK(CLK), .D(_03749_), .Q(ram_w8_l2048_id2_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44795_ ( .CLK(CLK), .D(_03750_), .Q(ram_w8_l2048_id2_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44796_ ( .CLK(CLK), .D(_03751_), .Q(ram_w8_l2048_id2_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id2_2_1_wenable_reg  ( .CLK(CLK), .D(_03752_), .Q(ram_w8_l2048_id2_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44798_ ( .CLK(CLK), .D(_03058_), .Q(_tmp_317) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44799_ ( .CLK(CLK), .D(_03059_), .Q(_tmp_318) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_319_reg  ( .CLK(CLK), .D(_03060_), .Q(_tmp_319) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44801_ ( .CLK(CLK), .D(_03062_), .Q(_tmp_320) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44802_ ( .CLK(CLK), .D(_03063_), .Q(_tmp_321) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44803_ ( .CLK(CLK), .D(_03064_), .Q(_tmp_322) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _44804_ ( .CLK(CLK), .D(_03065_), .Q(_tmp_329) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44805_ ( .CLK(CLK), .D(_02908_), .Q(_tmp_1128) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1129_reg  ( .CLK(CLK), .D(_02909_), .Q(_tmp_1129) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44807_ ( .CLK(CLK), .D(_03745_), .Q(ram_w8_l2048_id2_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44808_ ( .CLK(CLK), .D(_03746_), .Q(ram_w8_l2048_id2_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44809_ ( .CLK(CLK), .D(_03747_), .Q(ram_w8_l2048_id2_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id2_1_1_wenable_reg  ( .CLK(CLK), .D(_03748_), .Q(ram_w8_l2048_id2_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44811_ ( .CLK(CLK), .D(_03050_), .Q(_tmp_304) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44812_ ( .CLK(CLK), .D(_03051_), .Q(_tmp_305) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_306_reg  ( .CLK(CLK), .D(_03052_), .Q(_tmp_306) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44814_ ( .CLK(CLK), .D(_03053_), .Q(_tmp_307) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44815_ ( .CLK(CLK), .D(_03054_), .Q(_tmp_308) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44816_ ( .CLK(CLK), .D(_03055_), .Q(_tmp_309) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _44817_ ( .CLK(CLK), .D(_03057_), .Q(_tmp_316) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44818_ ( .CLK(CLK), .D(_02906_), .Q(_tmp_1126) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1127_reg  ( .CLK(CLK), .D(_02907_), .Q(_tmp_1127) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44820_ ( .CLK(CLK), .D(_03741_), .Q(ram_w8_l2048_id2_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44821_ ( .CLK(CLK), .D(_03742_), .Q(ram_w8_l2048_id2_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44822_ ( .CLK(CLK), .D(_03743_), .Q(ram_w8_l2048_id2_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id2_0_1_wenable_reg  ( .CLK(CLK), .D(_03744_), .Q(ram_w8_l2048_id2_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44824_ ( .CLK(CLK), .D(_03041_), .Q(_tmp_291) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44825_ ( .CLK(CLK), .D(_03042_), .Q(_tmp_292) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_293_reg  ( .CLK(CLK), .D(_03043_), .Q(_tmp_293) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44827_ ( .CLK(CLK), .D(_03044_), .Q(_tmp_294) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44828_ ( .CLK(CLK), .D(_03045_), .Q(_tmp_295) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44829_ ( .CLK(CLK), .D(_03046_), .Q(_tmp_296) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(2) ) _44830_ ( .CLK(CLK), .D(_03049_), .Q(_tmp_303) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id2_0_cond_3_1_reg  ( .CLK(CLK), .D(_01237_), .Q(_ram_w8_l2048_id2_0_cond_3_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44832_ ( .CLK(CLK), .D(_02904_), .Q(_tmp_1124) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1125_reg  ( .CLK(CLK), .D(_02905_), .Q(_tmp_1125) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id2_0_cond_6_1_reg  ( .CLK(CLK), .D(_01141_), .Q(_ram_w8_l2048_id2_0_cond_6_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44835_ ( .CLK(CLK), .D(_03735_), .Q(ram_w8_l2048_id1_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44836_ ( .CLK(CLK), .D(_03736_), .Q(ram_w8_l2048_id1_3_0_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id1_3_0_wenable_reg  ( .CLK(CLK), .D(_03737_), .Q(ram_w8_l2048_id1_3_0_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44838_ ( .CLK(CLK), .D(_03738_), .Q(ram_w8_l2048_id1_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44839_ ( .CLK(CLK), .D(_03739_), .Q(ram_w8_l2048_id1_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id1_3_1_wenable_reg  ( .CLK(CLK), .D(_03740_), .Q(ram_w8_l2048_id1_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44841_ ( .CLK(CLK), .D(_02993_), .Q(_tmp_18) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_19_reg  ( .CLK(CLK), .D(_03002_), .Q(_tmp_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id1_3_cond_5_1_reg  ( .CLK(CLK), .D(_01836_), .Q(_ram_w8_l2048_id1_3_cond_5_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1345_reg  ( .CLK(CLK), .D(_02959_), .Q(_tmp_1345) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1350_1_reg  ( .CLK(CLK), .D(_01227_), .Q(__tmp_1350_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44846_ ( .CLK(CLK), .D(_01228_), .Q(__tmp_1351_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1352_reg  ( .CLK(CLK), .D(_02961_), .Q(_tmp_1352) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1353_reg  ( .CLK(CLK), .D(_02962_), .Q(_tmp_1353) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1354_reg  ( .CLK(CLK), .D(_02963_), .Q(_tmp_1354) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1355_reg  ( .CLK(CLK), .D(_02964_), .Q(_tmp_1355) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44851_ ( .CLK(CLK), .D(_02965_), .Q(_tmp_1356) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44852_ ( .CLK(CLK), .D(_03729_), .Q(ram_w8_l2048_id1_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44853_ ( .CLK(CLK), .D(_03730_), .Q(ram_w8_l2048_id1_2_0_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id1_2_0_wenable_reg  ( .CLK(CLK), .D(_03731_), .Q(ram_w8_l2048_id1_2_0_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44855_ ( .CLK(CLK), .D(_03732_), .Q(ram_w8_l2048_id1_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44856_ ( .CLK(CLK), .D(_03733_), .Q(ram_w8_l2048_id1_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id1_2_1_wenable_reg  ( .CLK(CLK), .D(_03734_), .Q(ram_w8_l2048_id1_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44858_ ( .CLK(CLK), .D(_02987_), .Q(_tmp_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_17_reg  ( .CLK(CLK), .D(_02992_), .Q(_tmp_17) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id1_2_cond_5_1_reg  ( .CLK(CLK), .D(_01835_), .Q(_ram_w8_l2048_id1_2_cond_5_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1333_reg  ( .CLK(CLK), .D(_02952_), .Q(_tmp_1333) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1338_1_reg  ( .CLK(CLK), .D(_01225_), .Q(__tmp_1338_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44863_ ( .CLK(CLK), .D(_01226_), .Q(__tmp_1339_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1340_reg  ( .CLK(CLK), .D(_02954_), .Q(_tmp_1340) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1341_reg  ( .CLK(CLK), .D(_02955_), .Q(_tmp_1341) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1342_reg  ( .CLK(CLK), .D(_02956_), .Q(_tmp_1342) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1343_reg  ( .CLK(CLK), .D(_02957_), .Q(_tmp_1343) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44868_ ( .CLK(CLK), .D(_02958_), .Q(_tmp_1344) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44869_ ( .CLK(CLK), .D(_03723_), .Q(ram_w8_l2048_id1_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44870_ ( .CLK(CLK), .D(_03724_), .Q(ram_w8_l2048_id1_1_0_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id1_1_0_wenable_reg  ( .CLK(CLK), .D(_03725_), .Q(ram_w8_l2048_id1_1_0_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44872_ ( .CLK(CLK), .D(_03726_), .Q(ram_w8_l2048_id1_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44873_ ( .CLK(CLK), .D(_03727_), .Q(ram_w8_l2048_id1_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id1_1_1_wenable_reg  ( .CLK(CLK), .D(_03728_), .Q(ram_w8_l2048_id1_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44875_ ( .CLK(CLK), .D(_02976_), .Q(_tmp_14) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_15_reg  ( .CLK(CLK), .D(_02977_), .Q(_tmp_15) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id1_1_cond_5_1_reg  ( .CLK(CLK), .D(_01834_), .Q(_ram_w8_l2048_id1_1_cond_5_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1321_reg  ( .CLK(CLK), .D(_02945_), .Q(_tmp_1321) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1326_1_reg  ( .CLK(CLK), .D(_01223_), .Q(__tmp_1326_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44880_ ( .CLK(CLK), .D(_01224_), .Q(__tmp_1327_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1328_reg  ( .CLK(CLK), .D(_02946_), .Q(_tmp_1328) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1329_reg  ( .CLK(CLK), .D(_02947_), .Q(_tmp_1329) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1330_reg  ( .CLK(CLK), .D(_02949_), .Q(_tmp_1330) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1331_reg  ( .CLK(CLK), .D(_02950_), .Q(_tmp_1331) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44885_ ( .CLK(CLK), .D(_02951_), .Q(_tmp_1332) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44886_ ( .CLK(CLK), .D(_01587_), .Q(_dataflow_cat_data_167) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_cat_valid_167_reg  ( .CLK(CLK), .D(_01590_), .Q(_dataflow_cat_valid_167) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44888_ ( .CLK(CLK), .D(_03717_), .Q(ram_w8_l2048_id1_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44889_ ( .CLK(CLK), .D(_03718_), .Q(ram_w8_l2048_id1_0_0_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id1_0_0_wenable_reg  ( .CLK(CLK), .D(_03719_), .Q(ram_w8_l2048_id1_0_0_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44891_ ( .CLK(CLK), .D(_03720_), .Q(ram_w8_l2048_id1_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44892_ ( .CLK(CLK), .D(_03721_), .Q(ram_w8_l2048_id1_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id1_0_1_wenable_reg  ( .CLK(CLK), .D(_03722_), .Q(ram_w8_l2048_id1_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44894_ ( .CLK(CLK), .D(_02936_), .Q(_tmp_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_13_reg  ( .CLK(CLK), .D(_02972_), .Q(_tmp_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id1_0_cond_2_1_reg  ( .CLK(CLK), .D(_01231_), .Q(_ram_w8_l2048_id1_0_cond_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id1_0_cond_4_1_reg  ( .CLK(CLK), .D(_01111_), .Q(_ram_w8_l2048_id1_0_cond_4_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id1_0_cond_5_1_reg  ( .CLK(CLK), .D(_01833_), .Q(_ram_w8_l2048_id1_0_cond_5_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1309_reg  ( .CLK(CLK), .D(_02937_), .Q(_tmp_1309) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1314_1_reg  ( .CLK(CLK), .D(_01221_), .Q(__tmp_1314_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44901_ ( .CLK(CLK), .D(_01222_), .Q(__tmp_1315_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1316_reg  ( .CLK(CLK), .D(_02939_), .Q(_tmp_1316) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1317_reg  ( .CLK(CLK), .D(_02940_), .Q(_tmp_1317) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1318_reg  ( .CLK(CLK), .D(_02941_), .Q(_tmp_1318) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1319_reg  ( .CLK(CLK), .D(_02942_), .Q(_tmp_1319) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44906_ ( .CLK(CLK), .D(_02944_), .Q(_tmp_1320) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44907_ ( .CLK(CLK), .D(_03679_), .Q(ram_w8_l2048_id0_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44908_ ( .CLK(CLK), .D(_03680_), .Q(ram_w8_l2048_id0_3_0_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id0_3_0_wenable_reg  ( .CLK(CLK), .D(_03681_), .Q(ram_w8_l2048_id0_3_0_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44910_ ( .CLK(CLK), .D(_03682_), .Q(ram_w8_l2048_id0_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44911_ ( .CLK(CLK), .D(_03683_), .Q(ram_w8_l2048_id0_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id0_3_1_wenable_reg  ( .CLK(CLK), .D(_03684_), .Q(ram_w8_l2048_id0_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44913_ ( .CLK(CLK), .D(_03061_), .Q(_tmp_31) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_32_reg  ( .CLK(CLK), .D(_03066_), .Q(_tmp_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id0_3_cond_0_1_reg  ( .CLK(CLK), .D(_01824_), .Q(_ram_w8_l2048_id0_3_cond_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id0_3_cond_2_1_reg  ( .CLK(CLK), .D(_01234_), .Q(_ram_w8_l2048_id0_3_cond_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id0_3_cond_3_1_reg  ( .CLK(CLK), .D(_01828_), .Q(_ram_w8_l2048_id0_3_cond_3_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1108_reg  ( .CLK(CLK), .D(_02895_), .Q(_tmp_1108) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1113_1_reg  ( .CLK(CLK), .D(_01137_), .Q(__tmp_1113_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44920_ ( .CLK(CLK), .D(_01138_), .Q(__tmp_1114_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1115_reg  ( .CLK(CLK), .D(_02897_), .Q(_tmp_1115) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1116_reg  ( .CLK(CLK), .D(_02898_), .Q(_tmp_1116) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1117_reg  ( .CLK(CLK), .D(_02899_), .Q(_tmp_1117) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1118_reg  ( .CLK(CLK), .D(_02900_), .Q(_tmp_1118) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44925_ ( .CLK(CLK), .D(_02901_), .Q(_tmp_1119) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id0_3_cond_5_1_reg  ( .CLK(CLK), .D(_01144_), .Q(_ram_w8_l2048_id0_3_cond_5_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44927_ ( .CLK(CLK), .D(_03673_), .Q(ram_w8_l2048_id0_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44928_ ( .CLK(CLK), .D(_03674_), .Q(ram_w8_l2048_id0_2_0_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id0_2_0_wenable_reg  ( .CLK(CLK), .D(_03675_), .Q(ram_w8_l2048_id0_2_0_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44930_ ( .CLK(CLK), .D(_03676_), .Q(ram_w8_l2048_id0_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44931_ ( .CLK(CLK), .D(_03677_), .Q(ram_w8_l2048_id0_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id0_2_1_wenable_reg  ( .CLK(CLK), .D(_03678_), .Q(ram_w8_l2048_id0_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44933_ ( .CLK(CLK), .D(_03047_), .Q(_tmp_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_30_reg  ( .CLK(CLK), .D(_03056_), .Q(_tmp_30) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id0_2_cond_3_1_reg  ( .CLK(CLK), .D(_01827_), .Q(_ram_w8_l2048_id0_2_cond_3_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1096_reg  ( .CLK(CLK), .D(_02888_), .Q(_tmp_1096) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1101_1_reg  ( .CLK(CLK), .D(_01135_), .Q(__tmp_1101_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44938_ ( .CLK(CLK), .D(_01136_), .Q(__tmp_1102_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1103_reg  ( .CLK(CLK), .D(_02890_), .Q(_tmp_1103) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1104_reg  ( .CLK(CLK), .D(_02891_), .Q(_tmp_1104) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1105_reg  ( .CLK(CLK), .D(_02892_), .Q(_tmp_1105) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1106_reg  ( .CLK(CLK), .D(_02893_), .Q(_tmp_1106) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44943_ ( .CLK(CLK), .D(_02894_), .Q(_tmp_1107) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44944_ ( .CLK(CLK), .D(_03667_), .Q(ram_w8_l2048_id0_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44945_ ( .CLK(CLK), .D(_03668_), .Q(ram_w8_l2048_id0_1_0_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id0_1_0_wenable_reg  ( .CLK(CLK), .D(_03669_), .Q(ram_w8_l2048_id0_1_0_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44947_ ( .CLK(CLK), .D(_03670_), .Q(ram_w8_l2048_id0_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44948_ ( .CLK(CLK), .D(_03671_), .Q(ram_w8_l2048_id0_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id0_1_1_wenable_reg  ( .CLK(CLK), .D(_03672_), .Q(ram_w8_l2048_id0_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44950_ ( .CLK(CLK), .D(_03038_), .Q(_tmp_27) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_28_reg  ( .CLK(CLK), .D(_03040_), .Q(_tmp_28) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id0_1_cond_3_1_reg  ( .CLK(CLK), .D(_01826_), .Q(_ram_w8_l2048_id0_1_cond_3_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1084_reg  ( .CLK(CLK), .D(_02881_), .Q(_tmp_1084) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1089_1_reg  ( .CLK(CLK), .D(_01133_), .Q(__tmp_1089_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44955_ ( .CLK(CLK), .D(_01134_), .Q(__tmp_1090_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1091_reg  ( .CLK(CLK), .D(_02883_), .Q(_tmp_1091) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1092_reg  ( .CLK(CLK), .D(_02884_), .Q(_tmp_1092) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1093_reg  ( .CLK(CLK), .D(_02885_), .Q(_tmp_1093) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1094_reg  ( .CLK(CLK), .D(_02886_), .Q(_tmp_1094) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44960_ ( .CLK(CLK), .D(_02887_), .Q(_tmp_1095) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _44961_ ( .CLK(CLK), .D(_01586_), .Q(_dataflow_cat_data_107) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_cat_valid_107_reg  ( .CLK(CLK), .D(_01589_), .Q(_dataflow_cat_valid_107) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44963_ ( .CLK(CLK), .D(_03661_), .Q(ram_w8_l2048_id0_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44964_ ( .CLK(CLK), .D(_03662_), .Q(ram_w8_l2048_id0_0_0_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id0_0_0_wenable_reg  ( .CLK(CLK), .D(_03663_), .Q(ram_w8_l2048_id0_0_0_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _44966_ ( .CLK(CLK), .D(_03664_), .Q(ram_w8_l2048_id0_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44967_ ( .CLK(CLK), .D(_03665_), .Q(ram_w8_l2048_id0_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w8_l2048_id0_0_1_wenable_reg  ( .CLK(CLK), .D(_03666_), .Q(ram_w8_l2048_id0_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44969_ ( .CLK(CLK), .D(_03029_), .Q(_tmp_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_26_reg  ( .CLK(CLK), .D(_03037_), .Q(_tmp_26) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w8_l2048_id0_0_cond_3_1_reg  ( .CLK(CLK), .D(_01825_), .Q(_ram_w8_l2048_id0_0_cond_3_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1072_reg  ( .CLK(CLK), .D(_02874_), .Q(_tmp_1072) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) __tmp_1077_1_reg  ( .CLK(CLK), .D(_01131_), .Q(__tmp_1077_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _44974_ ( .CLK(CLK), .D(_01132_), .Q(__tmp_1078_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1079_reg  ( .CLK(CLK), .D(_02875_), .Q(_tmp_1079) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1080_reg  ( .CLK(CLK), .D(_02877_), .Q(_tmp_1080) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1081_reg  ( .CLK(CLK), .D(_02878_), .Q(_tmp_1081) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1082_reg  ( .CLK(CLK), .D(_02879_), .Q(_tmp_1082) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _44979_ ( .CLK(CLK), .D(_02880_), .Q(_tmp_1083) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44980_ ( .CLK(CLK), .D(_03657_), .Q(ram_w4_l8192_id8_7_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44981_ ( .CLK(CLK), .D(_03658_), .Q(ram_w4_l8192_id8_7_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44982_ ( .CLK(CLK), .D(_03659_), .Q(ram_w4_l8192_id8_7_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id8_7_1_wenable_reg  ( .CLK(CLK), .D(_03660_), .Q(ram_w4_l8192_id8_7_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44984_ ( .CLK(CLK), .D(_03653_), .Q(ram_w4_l8192_id8_6_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44985_ ( .CLK(CLK), .D(_03654_), .Q(ram_w4_l8192_id8_6_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44986_ ( .CLK(CLK), .D(_03655_), .Q(ram_w4_l8192_id8_6_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id8_6_1_wenable_reg  ( .CLK(CLK), .D(_03656_), .Q(ram_w4_l8192_id8_6_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44988_ ( .CLK(CLK), .D(_03649_), .Q(ram_w4_l8192_id8_5_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44989_ ( .CLK(CLK), .D(_03650_), .Q(ram_w4_l8192_id8_5_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44990_ ( .CLK(CLK), .D(_03651_), .Q(ram_w4_l8192_id8_5_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id8_5_1_wenable_reg  ( .CLK(CLK), .D(_03652_), .Q(ram_w4_l8192_id8_5_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44992_ ( .CLK(CLK), .D(_03645_), .Q(ram_w4_l8192_id8_4_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44993_ ( .CLK(CLK), .D(_03646_), .Q(ram_w4_l8192_id8_4_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44994_ ( .CLK(CLK), .D(_03647_), .Q(ram_w4_l8192_id8_4_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id8_4_1_wenable_reg  ( .CLK(CLK), .D(_03648_), .Q(ram_w4_l8192_id8_4_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44996_ ( .CLK(CLK), .D(_03641_), .Q(ram_w4_l8192_id8_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _44997_ ( .CLK(CLK), .D(_03642_), .Q(ram_w4_l8192_id8_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _44998_ ( .CLK(CLK), .D(_03643_), .Q(ram_w4_l8192_id8_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id8_3_1_wenable_reg  ( .CLK(CLK), .D(_03644_), .Q(ram_w4_l8192_id8_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45000_ ( .CLK(CLK), .D(_03637_), .Q(ram_w4_l8192_id8_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45001_ ( .CLK(CLK), .D(_03638_), .Q(ram_w4_l8192_id8_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45002_ ( .CLK(CLK), .D(_03639_), .Q(ram_w4_l8192_id8_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id8_2_1_wenable_reg  ( .CLK(CLK), .D(_03640_), .Q(ram_w4_l8192_id8_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45004_ ( .CLK(CLK), .D(_03633_), .Q(ram_w4_l8192_id8_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45005_ ( .CLK(CLK), .D(_03634_), .Q(ram_w4_l8192_id8_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45006_ ( .CLK(CLK), .D(_03635_), .Q(ram_w4_l8192_id8_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id8_1_1_wenable_reg  ( .CLK(CLK), .D(_03636_), .Q(ram_w4_l8192_id8_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45008_ ( .CLK(CLK), .D(_03629_), .Q(ram_w4_l8192_id8_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45009_ ( .CLK(CLK), .D(_03630_), .Q(ram_w4_l8192_id8_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45010_ ( .CLK(CLK), .D(_03631_), .Q(ram_w4_l8192_id8_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id8_0_1_wenable_reg  ( .CLK(CLK), .D(_03632_), .Q(ram_w4_l8192_id8_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w4_l8192_id8_0_cond_1_1_reg  ( .CLK(CLK), .D(_01288_), .Q(_ram_w4_l8192_id8_0_cond_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45013_ ( .CLK(CLK), .D(_03625_), .Q(ram_w4_l8192_id7_7_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45014_ ( .CLK(CLK), .D(_03626_), .Q(ram_w4_l8192_id7_7_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45015_ ( .CLK(CLK), .D(_03627_), .Q(ram_w4_l8192_id7_7_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id7_7_1_wenable_reg  ( .CLK(CLK), .D(_03628_), .Q(ram_w4_l8192_id7_7_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w4_l8192_id7_7_cond_1_1_reg  ( .CLK(CLK), .D(_01285_), .Q(_ram_w4_l8192_id7_7_cond_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45018_ ( .CLK(CLK), .D(_03621_), .Q(ram_w4_l8192_id7_6_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45019_ ( .CLK(CLK), .D(_03622_), .Q(ram_w4_l8192_id7_6_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45020_ ( .CLK(CLK), .D(_03623_), .Q(ram_w4_l8192_id7_6_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id7_6_1_wenable_reg  ( .CLK(CLK), .D(_03624_), .Q(ram_w4_l8192_id7_6_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45022_ ( .CLK(CLK), .D(_03617_), .Q(ram_w4_l8192_id7_5_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45023_ ( .CLK(CLK), .D(_03618_), .Q(ram_w4_l8192_id7_5_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45024_ ( .CLK(CLK), .D(_03619_), .Q(ram_w4_l8192_id7_5_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id7_5_1_wenable_reg  ( .CLK(CLK), .D(_03620_), .Q(ram_w4_l8192_id7_5_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45026_ ( .CLK(CLK), .D(_03613_), .Q(ram_w4_l8192_id7_4_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45027_ ( .CLK(CLK), .D(_03614_), .Q(ram_w4_l8192_id7_4_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45028_ ( .CLK(CLK), .D(_03615_), .Q(ram_w4_l8192_id7_4_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id7_4_1_wenable_reg  ( .CLK(CLK), .D(_03616_), .Q(ram_w4_l8192_id7_4_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45030_ ( .CLK(CLK), .D(_03609_), .Q(ram_w4_l8192_id7_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45031_ ( .CLK(CLK), .D(_03610_), .Q(ram_w4_l8192_id7_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45032_ ( .CLK(CLK), .D(_03611_), .Q(ram_w4_l8192_id7_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id7_3_1_wenable_reg  ( .CLK(CLK), .D(_03612_), .Q(ram_w4_l8192_id7_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45034_ ( .CLK(CLK), .D(_03605_), .Q(ram_w4_l8192_id7_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45035_ ( .CLK(CLK), .D(_03606_), .Q(ram_w4_l8192_id7_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45036_ ( .CLK(CLK), .D(_03607_), .Q(ram_w4_l8192_id7_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id7_2_1_wenable_reg  ( .CLK(CLK), .D(_03608_), .Q(ram_w4_l8192_id7_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45038_ ( .CLK(CLK), .D(_03601_), .Q(ram_w4_l8192_id7_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45039_ ( .CLK(CLK), .D(_03602_), .Q(ram_w4_l8192_id7_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45040_ ( .CLK(CLK), .D(_03603_), .Q(ram_w4_l8192_id7_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id7_1_1_wenable_reg  ( .CLK(CLK), .D(_03604_), .Q(ram_w4_l8192_id7_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45042_ ( .CLK(CLK), .D(_03597_), .Q(ram_w4_l8192_id7_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45043_ ( .CLK(CLK), .D(_03598_), .Q(ram_w4_l8192_id7_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45044_ ( .CLK(CLK), .D(_03599_), .Q(ram_w4_l8192_id7_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id7_0_1_wenable_reg  ( .CLK(CLK), .D(_03600_), .Q(ram_w4_l8192_id7_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45046_ ( .CLK(CLK), .D(_03593_), .Q(ram_w4_l8192_id6_7_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45047_ ( .CLK(CLK), .D(_03594_), .Q(ram_w4_l8192_id6_7_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45048_ ( .CLK(CLK), .D(_03595_), .Q(ram_w4_l8192_id6_7_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id6_7_1_wenable_reg  ( .CLK(CLK), .D(_03596_), .Q(ram_w4_l8192_id6_7_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45050_ ( .CLK(CLK), .D(_03589_), .Q(ram_w4_l8192_id6_6_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45051_ ( .CLK(CLK), .D(_03590_), .Q(ram_w4_l8192_id6_6_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45052_ ( .CLK(CLK), .D(_03591_), .Q(ram_w4_l8192_id6_6_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id6_6_1_wenable_reg  ( .CLK(CLK), .D(_03592_), .Q(ram_w4_l8192_id6_6_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45054_ ( .CLK(CLK), .D(_03585_), .Q(ram_w4_l8192_id6_5_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45055_ ( .CLK(CLK), .D(_03586_), .Q(ram_w4_l8192_id6_5_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45056_ ( .CLK(CLK), .D(_03587_), .Q(ram_w4_l8192_id6_5_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id6_5_1_wenable_reg  ( .CLK(CLK), .D(_03588_), .Q(ram_w4_l8192_id6_5_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45058_ ( .CLK(CLK), .D(_03581_), .Q(ram_w4_l8192_id6_4_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45059_ ( .CLK(CLK), .D(_03582_), .Q(ram_w4_l8192_id6_4_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45060_ ( .CLK(CLK), .D(_03583_), .Q(ram_w4_l8192_id6_4_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id6_4_1_wenable_reg  ( .CLK(CLK), .D(_03584_), .Q(ram_w4_l8192_id6_4_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45062_ ( .CLK(CLK), .D(_03577_), .Q(ram_w4_l8192_id6_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45063_ ( .CLK(CLK), .D(_03578_), .Q(ram_w4_l8192_id6_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45064_ ( .CLK(CLK), .D(_03579_), .Q(ram_w4_l8192_id6_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id6_3_1_wenable_reg  ( .CLK(CLK), .D(_03580_), .Q(ram_w4_l8192_id6_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45066_ ( .CLK(CLK), .D(_03573_), .Q(ram_w4_l8192_id6_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45067_ ( .CLK(CLK), .D(_03574_), .Q(ram_w4_l8192_id6_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45068_ ( .CLK(CLK), .D(_03575_), .Q(ram_w4_l8192_id6_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id6_2_1_wenable_reg  ( .CLK(CLK), .D(_03576_), .Q(ram_w4_l8192_id6_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w4_l8192_id6_2_cond_1_1_reg  ( .CLK(CLK), .D(_01282_), .Q(_ram_w4_l8192_id6_2_cond_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45071_ ( .CLK(CLK), .D(_03569_), .Q(ram_w4_l8192_id6_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45072_ ( .CLK(CLK), .D(_03570_), .Q(ram_w4_l8192_id6_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45073_ ( .CLK(CLK), .D(_03571_), .Q(ram_w4_l8192_id6_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id6_1_1_wenable_reg  ( .CLK(CLK), .D(_03572_), .Q(ram_w4_l8192_id6_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45075_ ( .CLK(CLK), .D(_03565_), .Q(ram_w4_l8192_id6_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45076_ ( .CLK(CLK), .D(_03566_), .Q(ram_w4_l8192_id6_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45077_ ( .CLK(CLK), .D(_03567_), .Q(ram_w4_l8192_id6_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id6_0_1_wenable_reg  ( .CLK(CLK), .D(_03568_), .Q(ram_w4_l8192_id6_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45079_ ( .CLK(CLK), .D(_03561_), .Q(ram_w4_l8192_id5_7_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45080_ ( .CLK(CLK), .D(_03562_), .Q(ram_w4_l8192_id5_7_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45081_ ( .CLK(CLK), .D(_03563_), .Q(ram_w4_l8192_id5_7_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id5_7_1_wenable_reg  ( .CLK(CLK), .D(_03564_), .Q(ram_w4_l8192_id5_7_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w4_l8192_id5_7_cond_2_1_reg  ( .CLK(CLK), .D(_01279_), .Q(_ram_w4_l8192_id5_7_cond_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45084_ ( .CLK(CLK), .D(_03557_), .Q(ram_w4_l8192_id5_6_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45085_ ( .CLK(CLK), .D(_03558_), .Q(ram_w4_l8192_id5_6_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45086_ ( .CLK(CLK), .D(_03559_), .Q(ram_w4_l8192_id5_6_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id5_6_1_wenable_reg  ( .CLK(CLK), .D(_03560_), .Q(ram_w4_l8192_id5_6_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45088_ ( .CLK(CLK), .D(_03553_), .Q(ram_w4_l8192_id5_5_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45089_ ( .CLK(CLK), .D(_03554_), .Q(ram_w4_l8192_id5_5_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45090_ ( .CLK(CLK), .D(_03555_), .Q(ram_w4_l8192_id5_5_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id5_5_1_wenable_reg  ( .CLK(CLK), .D(_03556_), .Q(ram_w4_l8192_id5_5_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45092_ ( .CLK(CLK), .D(_03549_), .Q(ram_w4_l8192_id5_4_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45093_ ( .CLK(CLK), .D(_03550_), .Q(ram_w4_l8192_id5_4_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45094_ ( .CLK(CLK), .D(_03551_), .Q(ram_w4_l8192_id5_4_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id5_4_1_wenable_reg  ( .CLK(CLK), .D(_03552_), .Q(ram_w4_l8192_id5_4_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45096_ ( .CLK(CLK), .D(_03545_), .Q(ram_w4_l8192_id5_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45097_ ( .CLK(CLK), .D(_03546_), .Q(ram_w4_l8192_id5_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45098_ ( .CLK(CLK), .D(_03547_), .Q(ram_w4_l8192_id5_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id5_3_1_wenable_reg  ( .CLK(CLK), .D(_03548_), .Q(ram_w4_l8192_id5_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45100_ ( .CLK(CLK), .D(_03541_), .Q(ram_w4_l8192_id5_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45101_ ( .CLK(CLK), .D(_03542_), .Q(ram_w4_l8192_id5_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45102_ ( .CLK(CLK), .D(_03543_), .Q(ram_w4_l8192_id5_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id5_2_1_wenable_reg  ( .CLK(CLK), .D(_03544_), .Q(ram_w4_l8192_id5_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45104_ ( .CLK(CLK), .D(_03537_), .Q(ram_w4_l8192_id5_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45105_ ( .CLK(CLK), .D(_03538_), .Q(ram_w4_l8192_id5_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45106_ ( .CLK(CLK), .D(_03539_), .Q(ram_w4_l8192_id5_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id5_1_1_wenable_reg  ( .CLK(CLK), .D(_03540_), .Q(ram_w4_l8192_id5_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45108_ ( .CLK(CLK), .D(_03533_), .Q(ram_w4_l8192_id5_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45109_ ( .CLK(CLK), .D(_03534_), .Q(ram_w4_l8192_id5_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45110_ ( .CLK(CLK), .D(_03535_), .Q(ram_w4_l8192_id5_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id5_0_1_wenable_reg  ( .CLK(CLK), .D(_03536_), .Q(ram_w4_l8192_id5_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45112_ ( .CLK(CLK), .D(_03529_), .Q(ram_w4_l8192_id4_7_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45113_ ( .CLK(CLK), .D(_03530_), .Q(ram_w4_l8192_id4_7_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45114_ ( .CLK(CLK), .D(_03531_), .Q(ram_w4_l8192_id4_7_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id4_7_1_wenable_reg  ( .CLK(CLK), .D(_03532_), .Q(ram_w4_l8192_id4_7_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w4_l8192_id4_7_cond_1_1_reg  ( .CLK(CLK), .D(_01276_), .Q(_ram_w4_l8192_id4_7_cond_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45117_ ( .CLK(CLK), .D(_03525_), .Q(ram_w4_l8192_id4_6_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45118_ ( .CLK(CLK), .D(_03526_), .Q(ram_w4_l8192_id4_6_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45119_ ( .CLK(CLK), .D(_03527_), .Q(ram_w4_l8192_id4_6_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id4_6_1_wenable_reg  ( .CLK(CLK), .D(_03528_), .Q(ram_w4_l8192_id4_6_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45121_ ( .CLK(CLK), .D(_03521_), .Q(ram_w4_l8192_id4_5_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45122_ ( .CLK(CLK), .D(_03522_), .Q(ram_w4_l8192_id4_5_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45123_ ( .CLK(CLK), .D(_03523_), .Q(ram_w4_l8192_id4_5_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id4_5_1_wenable_reg  ( .CLK(CLK), .D(_03524_), .Q(ram_w4_l8192_id4_5_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45125_ ( .CLK(CLK), .D(_03517_), .Q(ram_w4_l8192_id4_4_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45126_ ( .CLK(CLK), .D(_03518_), .Q(ram_w4_l8192_id4_4_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45127_ ( .CLK(CLK), .D(_03519_), .Q(ram_w4_l8192_id4_4_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id4_4_1_wenable_reg  ( .CLK(CLK), .D(_03520_), .Q(ram_w4_l8192_id4_4_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45129_ ( .CLK(CLK), .D(_03513_), .Q(ram_w4_l8192_id4_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45130_ ( .CLK(CLK), .D(_03514_), .Q(ram_w4_l8192_id4_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45131_ ( .CLK(CLK), .D(_03515_), .Q(ram_w4_l8192_id4_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id4_3_1_wenable_reg  ( .CLK(CLK), .D(_03516_), .Q(ram_w4_l8192_id4_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45133_ ( .CLK(CLK), .D(_03509_), .Q(ram_w4_l8192_id4_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45134_ ( .CLK(CLK), .D(_03510_), .Q(ram_w4_l8192_id4_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45135_ ( .CLK(CLK), .D(_03511_), .Q(ram_w4_l8192_id4_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id4_2_1_wenable_reg  ( .CLK(CLK), .D(_03512_), .Q(ram_w4_l8192_id4_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45137_ ( .CLK(CLK), .D(_03505_), .Q(ram_w4_l8192_id4_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45138_ ( .CLK(CLK), .D(_03506_), .Q(ram_w4_l8192_id4_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45139_ ( .CLK(CLK), .D(_03507_), .Q(ram_w4_l8192_id4_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id4_1_1_wenable_reg  ( .CLK(CLK), .D(_03508_), .Q(ram_w4_l8192_id4_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45141_ ( .CLK(CLK), .D(_03501_), .Q(ram_w4_l8192_id4_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45142_ ( .CLK(CLK), .D(_03502_), .Q(ram_w4_l8192_id4_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45143_ ( .CLK(CLK), .D(_03503_), .Q(ram_w4_l8192_id4_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id4_0_1_wenable_reg  ( .CLK(CLK), .D(_03504_), .Q(ram_w4_l8192_id4_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45145_ ( .CLK(CLK), .D(_03497_), .Q(ram_w4_l8192_id3_7_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45146_ ( .CLK(CLK), .D(_03498_), .Q(ram_w4_l8192_id3_7_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45147_ ( .CLK(CLK), .D(_03499_), .Q(ram_w4_l8192_id3_7_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id3_7_1_wenable_reg  ( .CLK(CLK), .D(_03500_), .Q(ram_w4_l8192_id3_7_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w4_l8192_id3_7_cond_1_1_reg  ( .CLK(CLK), .D(_01273_), .Q(_ram_w4_l8192_id3_7_cond_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45150_ ( .CLK(CLK), .D(_03493_), .Q(ram_w4_l8192_id3_6_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45151_ ( .CLK(CLK), .D(_03494_), .Q(ram_w4_l8192_id3_6_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45152_ ( .CLK(CLK), .D(_03495_), .Q(ram_w4_l8192_id3_6_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id3_6_1_wenable_reg  ( .CLK(CLK), .D(_03496_), .Q(ram_w4_l8192_id3_6_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45154_ ( .CLK(CLK), .D(_03489_), .Q(ram_w4_l8192_id3_5_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45155_ ( .CLK(CLK), .D(_03490_), .Q(ram_w4_l8192_id3_5_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45156_ ( .CLK(CLK), .D(_03491_), .Q(ram_w4_l8192_id3_5_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id3_5_1_wenable_reg  ( .CLK(CLK), .D(_03492_), .Q(ram_w4_l8192_id3_5_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45158_ ( .CLK(CLK), .D(_03485_), .Q(ram_w4_l8192_id3_4_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45159_ ( .CLK(CLK), .D(_03486_), .Q(ram_w4_l8192_id3_4_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45160_ ( .CLK(CLK), .D(_03487_), .Q(ram_w4_l8192_id3_4_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id3_4_1_wenable_reg  ( .CLK(CLK), .D(_03488_), .Q(ram_w4_l8192_id3_4_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45162_ ( .CLK(CLK), .D(_03481_), .Q(ram_w4_l8192_id3_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45163_ ( .CLK(CLK), .D(_03482_), .Q(ram_w4_l8192_id3_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45164_ ( .CLK(CLK), .D(_03483_), .Q(ram_w4_l8192_id3_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id3_3_1_wenable_reg  ( .CLK(CLK), .D(_03484_), .Q(ram_w4_l8192_id3_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45166_ ( .CLK(CLK), .D(_03477_), .Q(ram_w4_l8192_id3_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45167_ ( .CLK(CLK), .D(_03478_), .Q(ram_w4_l8192_id3_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45168_ ( .CLK(CLK), .D(_03479_), .Q(ram_w4_l8192_id3_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id3_2_1_wenable_reg  ( .CLK(CLK), .D(_03480_), .Q(ram_w4_l8192_id3_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45170_ ( .CLK(CLK), .D(_03473_), .Q(ram_w4_l8192_id3_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45171_ ( .CLK(CLK), .D(_03474_), .Q(ram_w4_l8192_id3_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45172_ ( .CLK(CLK), .D(_03475_), .Q(ram_w4_l8192_id3_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id3_1_1_wenable_reg  ( .CLK(CLK), .D(_03476_), .Q(ram_w4_l8192_id3_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45174_ ( .CLK(CLK), .D(_03469_), .Q(ram_w4_l8192_id3_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45175_ ( .CLK(CLK), .D(_03470_), .Q(ram_w4_l8192_id3_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45176_ ( .CLK(CLK), .D(_03471_), .Q(ram_w4_l8192_id3_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id3_0_1_wenable_reg  ( .CLK(CLK), .D(_03472_), .Q(ram_w4_l8192_id3_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45178_ ( .CLK(CLK), .D(_03465_), .Q(ram_w4_l8192_id2_7_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45179_ ( .CLK(CLK), .D(_03466_), .Q(ram_w4_l8192_id2_7_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45180_ ( .CLK(CLK), .D(_03467_), .Q(ram_w4_l8192_id2_7_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id2_7_1_wenable_reg  ( .CLK(CLK), .D(_03468_), .Q(ram_w4_l8192_id2_7_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w4_l8192_id2_7_cond_1_1_reg  ( .CLK(CLK), .D(_01270_), .Q(_ram_w4_l8192_id2_7_cond_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45183_ ( .CLK(CLK), .D(_03461_), .Q(ram_w4_l8192_id2_6_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45184_ ( .CLK(CLK), .D(_03462_), .Q(ram_w4_l8192_id2_6_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45185_ ( .CLK(CLK), .D(_03463_), .Q(ram_w4_l8192_id2_6_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id2_6_1_wenable_reg  ( .CLK(CLK), .D(_03464_), .Q(ram_w4_l8192_id2_6_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45187_ ( .CLK(CLK), .D(_03457_), .Q(ram_w4_l8192_id2_5_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45188_ ( .CLK(CLK), .D(_03458_), .Q(ram_w4_l8192_id2_5_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45189_ ( .CLK(CLK), .D(_03459_), .Q(ram_w4_l8192_id2_5_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id2_5_1_wenable_reg  ( .CLK(CLK), .D(_03460_), .Q(ram_w4_l8192_id2_5_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45191_ ( .CLK(CLK), .D(_03453_), .Q(ram_w4_l8192_id2_4_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45192_ ( .CLK(CLK), .D(_03454_), .Q(ram_w4_l8192_id2_4_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45193_ ( .CLK(CLK), .D(_03455_), .Q(ram_w4_l8192_id2_4_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id2_4_1_wenable_reg  ( .CLK(CLK), .D(_03456_), .Q(ram_w4_l8192_id2_4_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45195_ ( .CLK(CLK), .D(_03449_), .Q(ram_w4_l8192_id2_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45196_ ( .CLK(CLK), .D(_03450_), .Q(ram_w4_l8192_id2_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45197_ ( .CLK(CLK), .D(_03451_), .Q(ram_w4_l8192_id2_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id2_3_1_wenable_reg  ( .CLK(CLK), .D(_03452_), .Q(ram_w4_l8192_id2_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45199_ ( .CLK(CLK), .D(_03445_), .Q(ram_w4_l8192_id2_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45200_ ( .CLK(CLK), .D(_03446_), .Q(ram_w4_l8192_id2_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45201_ ( .CLK(CLK), .D(_03447_), .Q(ram_w4_l8192_id2_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id2_2_1_wenable_reg  ( .CLK(CLK), .D(_03448_), .Q(ram_w4_l8192_id2_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45203_ ( .CLK(CLK), .D(_03441_), .Q(ram_w4_l8192_id2_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45204_ ( .CLK(CLK), .D(_03442_), .Q(ram_w4_l8192_id2_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45205_ ( .CLK(CLK), .D(_03443_), .Q(ram_w4_l8192_id2_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id2_1_1_wenable_reg  ( .CLK(CLK), .D(_03444_), .Q(ram_w4_l8192_id2_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45207_ ( .CLK(CLK), .D(_03437_), .Q(ram_w4_l8192_id2_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45208_ ( .CLK(CLK), .D(_03438_), .Q(ram_w4_l8192_id2_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45209_ ( .CLK(CLK), .D(_03439_), .Q(ram_w4_l8192_id2_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id2_0_1_wenable_reg  ( .CLK(CLK), .D(_03440_), .Q(ram_w4_l8192_id2_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45211_ ( .CLK(CLK), .D(_03433_), .Q(ram_w4_l8192_id1_7_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45212_ ( .CLK(CLK), .D(_03434_), .Q(ram_w4_l8192_id1_7_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45213_ ( .CLK(CLK), .D(_03435_), .Q(ram_w4_l8192_id1_7_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id1_7_1_wenable_reg  ( .CLK(CLK), .D(_03436_), .Q(ram_w4_l8192_id1_7_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w4_l8192_id1_7_cond_1_1_reg  ( .CLK(CLK), .D(_01267_), .Q(_ram_w4_l8192_id1_7_cond_1_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45216_ ( .CLK(CLK), .D(_03429_), .Q(ram_w4_l8192_id1_6_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45217_ ( .CLK(CLK), .D(_03430_), .Q(ram_w4_l8192_id1_6_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45218_ ( .CLK(CLK), .D(_03431_), .Q(ram_w4_l8192_id1_6_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id1_6_1_wenable_reg  ( .CLK(CLK), .D(_03432_), .Q(ram_w4_l8192_id1_6_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45220_ ( .CLK(CLK), .D(_03425_), .Q(ram_w4_l8192_id1_5_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45221_ ( .CLK(CLK), .D(_03426_), .Q(ram_w4_l8192_id1_5_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45222_ ( .CLK(CLK), .D(_03427_), .Q(ram_w4_l8192_id1_5_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id1_5_1_wenable_reg  ( .CLK(CLK), .D(_03428_), .Q(ram_w4_l8192_id1_5_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45224_ ( .CLK(CLK), .D(_03421_), .Q(ram_w4_l8192_id1_4_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45225_ ( .CLK(CLK), .D(_03422_), .Q(ram_w4_l8192_id1_4_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45226_ ( .CLK(CLK), .D(_03423_), .Q(ram_w4_l8192_id1_4_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id1_4_1_wenable_reg  ( .CLK(CLK), .D(_03424_), .Q(ram_w4_l8192_id1_4_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45228_ ( .CLK(CLK), .D(_03417_), .Q(ram_w4_l8192_id1_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45229_ ( .CLK(CLK), .D(_03418_), .Q(ram_w4_l8192_id1_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45230_ ( .CLK(CLK), .D(_03419_), .Q(ram_w4_l8192_id1_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id1_3_1_wenable_reg  ( .CLK(CLK), .D(_03420_), .Q(ram_w4_l8192_id1_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45232_ ( .CLK(CLK), .D(_03413_), .Q(ram_w4_l8192_id1_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45233_ ( .CLK(CLK), .D(_03414_), .Q(ram_w4_l8192_id1_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45234_ ( .CLK(CLK), .D(_03415_), .Q(ram_w4_l8192_id1_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id1_2_1_wenable_reg  ( .CLK(CLK), .D(_03416_), .Q(ram_w4_l8192_id1_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45236_ ( .CLK(CLK), .D(_03409_), .Q(ram_w4_l8192_id1_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45237_ ( .CLK(CLK), .D(_03410_), .Q(ram_w4_l8192_id1_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45238_ ( .CLK(CLK), .D(_03411_), .Q(ram_w4_l8192_id1_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id1_1_1_wenable_reg  ( .CLK(CLK), .D(_03412_), .Q(ram_w4_l8192_id1_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45240_ ( .CLK(CLK), .D(_03405_), .Q(ram_w4_l8192_id1_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45241_ ( .CLK(CLK), .D(_03406_), .Q(ram_w4_l8192_id1_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45242_ ( .CLK(CLK), .D(_03407_), .Q(ram_w4_l8192_id1_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id1_0_1_wenable_reg  ( .CLK(CLK), .D(_03408_), .Q(ram_w4_l8192_id1_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45244_ ( .CLK(CLK), .D(_03401_), .Q(ram_w4_l8192_id0_7_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45245_ ( .CLK(CLK), .D(_03402_), .Q(ram_w4_l8192_id0_7_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45246_ ( .CLK(CLK), .D(_03403_), .Q(ram_w4_l8192_id0_7_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id0_7_1_wenable_reg  ( .CLK(CLK), .D(_03404_), .Q(ram_w4_l8192_id0_7_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _45248_ ( .CLK(CLK), .D(_03024_), .Q(_tmp_255) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45249_ ( .CLK(CLK), .D(_03025_), .Q(_tmp_256) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_257_reg  ( .CLK(CLK), .D(_03026_), .Q(_tmp_257) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45251_ ( .CLK(CLK), .D(_03027_), .Q(_tmp_258) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45252_ ( .CLK(CLK), .D(_03028_), .Q(_tmp_259) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45253_ ( .CLK(CLK), .D(_03030_), .Q(_tmp_260) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45254_ ( .CLK(CLK), .D(_03031_), .Q(_tmp_261) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45255_ ( .CLK(CLK), .D(_03032_), .Q(_tmp_262) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45256_ ( .CLK(CLK), .D(_03033_), .Q(_tmp_263) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45257_ ( .CLK(CLK), .D(_03034_), .Q(_tmp_264) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45258_ ( .CLK(CLK), .D(_03035_), .Q(_tmp_265) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45259_ ( .CLK(CLK), .D(_03036_), .Q(_tmp_266) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45260_ ( .CLK(CLK), .D(_03039_), .Q(_tmp_285) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _ram_w4_l8192_id0_7_cond_2_1_reg  ( .CLK(CLK), .D(_01264_), .Q(_ram_w4_l8192_id0_7_cond_2_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45262_ ( .CLK(CLK), .D(_02926_), .Q(_tmp_1150) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1151_reg  ( .CLK(CLK), .D(_02927_), .Q(_tmp_1151) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45264_ ( .CLK(CLK), .D(_03397_), .Q(ram_w4_l8192_id0_6_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45265_ ( .CLK(CLK), .D(_03398_), .Q(ram_w4_l8192_id0_6_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45266_ ( .CLK(CLK), .D(_03399_), .Q(ram_w4_l8192_id0_6_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id0_6_1_wenable_reg  ( .CLK(CLK), .D(_03400_), .Q(ram_w4_l8192_id0_6_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _45268_ ( .CLK(CLK), .D(_03011_), .Q(_tmp_224) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45269_ ( .CLK(CLK), .D(_03012_), .Q(_tmp_225) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_226_reg  ( .CLK(CLK), .D(_03013_), .Q(_tmp_226) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45271_ ( .CLK(CLK), .D(_03014_), .Q(_tmp_227) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45272_ ( .CLK(CLK), .D(_03015_), .Q(_tmp_228) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45273_ ( .CLK(CLK), .D(_03016_), .Q(_tmp_229) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45274_ ( .CLK(CLK), .D(_03017_), .Q(_tmp_230) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45275_ ( .CLK(CLK), .D(_03018_), .Q(_tmp_231) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45276_ ( .CLK(CLK), .D(_03019_), .Q(_tmp_232) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45277_ ( .CLK(CLK), .D(_03020_), .Q(_tmp_233) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45278_ ( .CLK(CLK), .D(_03021_), .Q(_tmp_234) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45279_ ( .CLK(CLK), .D(_03022_), .Q(_tmp_235) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45280_ ( .CLK(CLK), .D(_03023_), .Q(_tmp_254) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45281_ ( .CLK(CLK), .D(_02924_), .Q(_tmp_1148) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1149_reg  ( .CLK(CLK), .D(_02925_), .Q(_tmp_1149) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45283_ ( .CLK(CLK), .D(_03393_), .Q(ram_w4_l8192_id0_5_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45284_ ( .CLK(CLK), .D(_03394_), .Q(ram_w4_l8192_id0_5_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45285_ ( .CLK(CLK), .D(_03395_), .Q(ram_w4_l8192_id0_5_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id0_5_1_wenable_reg  ( .CLK(CLK), .D(_03396_), .Q(ram_w4_l8192_id0_5_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _45287_ ( .CLK(CLK), .D(_02995_), .Q(_tmp_193) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45288_ ( .CLK(CLK), .D(_02996_), .Q(_tmp_194) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_195_reg  ( .CLK(CLK), .D(_02997_), .Q(_tmp_195) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45290_ ( .CLK(CLK), .D(_02998_), .Q(_tmp_196) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45291_ ( .CLK(CLK), .D(_02999_), .Q(_tmp_197) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45292_ ( .CLK(CLK), .D(_03000_), .Q(_tmp_198) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45293_ ( .CLK(CLK), .D(_03001_), .Q(_tmp_199) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45294_ ( .CLK(CLK), .D(_03004_), .Q(_tmp_200) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45295_ ( .CLK(CLK), .D(_03005_), .Q(_tmp_201) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45296_ ( .CLK(CLK), .D(_03006_), .Q(_tmp_202) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45297_ ( .CLK(CLK), .D(_03007_), .Q(_tmp_203) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45298_ ( .CLK(CLK), .D(_03008_), .Q(_tmp_204) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45299_ ( .CLK(CLK), .D(_03010_), .Q(_tmp_223) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45300_ ( .CLK(CLK), .D(_02922_), .Q(_tmp_1146) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1147_reg  ( .CLK(CLK), .D(_02923_), .Q(_tmp_1147) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45302_ ( .CLK(CLK), .D(_03389_), .Q(ram_w4_l8192_id0_4_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45303_ ( .CLK(CLK), .D(_03390_), .Q(ram_w4_l8192_id0_4_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45304_ ( .CLK(CLK), .D(_03391_), .Q(ram_w4_l8192_id0_4_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id0_4_1_wenable_reg  ( .CLK(CLK), .D(_03392_), .Q(ram_w4_l8192_id0_4_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _45306_ ( .CLK(CLK), .D(_02979_), .Q(_tmp_162) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45307_ ( .CLK(CLK), .D(_02980_), .Q(_tmp_163) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_164_reg  ( .CLK(CLK), .D(_02981_), .Q(_tmp_164) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45309_ ( .CLK(CLK), .D(_02982_), .Q(_tmp_165) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45310_ ( .CLK(CLK), .D(_02983_), .Q(_tmp_166) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45311_ ( .CLK(CLK), .D(_02984_), .Q(_tmp_167) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45312_ ( .CLK(CLK), .D(_02985_), .Q(_tmp_168) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45313_ ( .CLK(CLK), .D(_02986_), .Q(_tmp_169) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45314_ ( .CLK(CLK), .D(_02988_), .Q(_tmp_170) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45315_ ( .CLK(CLK), .D(_02989_), .Q(_tmp_171) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45316_ ( .CLK(CLK), .D(_02990_), .Q(_tmp_172) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45317_ ( .CLK(CLK), .D(_02991_), .Q(_tmp_173) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45318_ ( .CLK(CLK), .D(_02994_), .Q(_tmp_192) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45319_ ( .CLK(CLK), .D(_02920_), .Q(_tmp_1144) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1145_reg  ( .CLK(CLK), .D(_02921_), .Q(_tmp_1145) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45321_ ( .CLK(CLK), .D(_03385_), .Q(ram_w4_l8192_id0_3_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45322_ ( .CLK(CLK), .D(_03386_), .Q(ram_w4_l8192_id0_3_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45323_ ( .CLK(CLK), .D(_03387_), .Q(ram_w4_l8192_id0_3_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id0_3_1_wenable_reg  ( .CLK(CLK), .D(_03388_), .Q(ram_w4_l8192_id0_3_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _45325_ ( .CLK(CLK), .D(_02943_), .Q(_tmp_131) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45326_ ( .CLK(CLK), .D(_02948_), .Q(_tmp_132) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_133_reg  ( .CLK(CLK), .D(_02953_), .Q(_tmp_133) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45328_ ( .CLK(CLK), .D(_02960_), .Q(_tmp_134) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45329_ ( .CLK(CLK), .D(_02967_), .Q(_tmp_135) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45330_ ( .CLK(CLK), .D(_02968_), .Q(_tmp_136) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45331_ ( .CLK(CLK), .D(_02969_), .Q(_tmp_137) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45332_ ( .CLK(CLK), .D(_02970_), .Q(_tmp_138) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45333_ ( .CLK(CLK), .D(_02971_), .Q(_tmp_139) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45334_ ( .CLK(CLK), .D(_02973_), .Q(_tmp_140) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45335_ ( .CLK(CLK), .D(_02974_), .Q(_tmp_141) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45336_ ( .CLK(CLK), .D(_02975_), .Q(_tmp_142) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45337_ ( .CLK(CLK), .D(_02978_), .Q(_tmp_161) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45338_ ( .CLK(CLK), .D(_02918_), .Q(_tmp_1142) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1143_reg  ( .CLK(CLK), .D(_02919_), .Q(_tmp_1143) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45340_ ( .CLK(CLK), .D(_03381_), .Q(ram_w4_l8192_id0_2_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45341_ ( .CLK(CLK), .D(_03382_), .Q(ram_w4_l8192_id0_2_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45342_ ( .CLK(CLK), .D(_03383_), .Q(ram_w4_l8192_id0_2_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id0_2_1_wenable_reg  ( .CLK(CLK), .D(_03384_), .Q(ram_w4_l8192_id0_2_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _45344_ ( .CLK(CLK), .D(_02860_), .Q(_tmp_100) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45345_ ( .CLK(CLK), .D(_02867_), .Q(_tmp_101) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_102_reg  ( .CLK(CLK), .D(_02869_), .Q(_tmp_102) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45347_ ( .CLK(CLK), .D(_02870_), .Q(_tmp_103) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45348_ ( .CLK(CLK), .D(_02871_), .Q(_tmp_104) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45349_ ( .CLK(CLK), .D(_02872_), .Q(_tmp_105) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45350_ ( .CLK(CLK), .D(_02873_), .Q(_tmp_106) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45351_ ( .CLK(CLK), .D(_02876_), .Q(_tmp_107) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45352_ ( .CLK(CLK), .D(_02882_), .Q(_tmp_108) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45353_ ( .CLK(CLK), .D(_02889_), .Q(_tmp_109) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45354_ ( .CLK(CLK), .D(_02896_), .Q(_tmp_110) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45355_ ( .CLK(CLK), .D(_02902_), .Q(_tmp_111) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45356_ ( .CLK(CLK), .D(_02938_), .Q(_tmp_130) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45357_ ( .CLK(CLK), .D(_02916_), .Q(_tmp_1140) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1141_reg  ( .CLK(CLK), .D(_02917_), .Q(_tmp_1141) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45359_ ( .CLK(CLK), .D(_03377_), .Q(ram_w4_l8192_id0_1_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45360_ ( .CLK(CLK), .D(_03378_), .Q(ram_w4_l8192_id0_1_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45361_ ( .CLK(CLK), .D(_03379_), .Q(ram_w4_l8192_id0_1_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id0_1_1_wenable_reg  ( .CLK(CLK), .D(_03380_), .Q(ram_w4_l8192_id0_1_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _45363_ ( .CLK(CLK), .D(_03146_), .Q(_tmp_69) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45364_ ( .CLK(CLK), .D(_03147_), .Q(_tmp_70) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_71_reg  ( .CLK(CLK), .D(_03148_), .Q(_tmp_71) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45366_ ( .CLK(CLK), .D(_03149_), .Q(_tmp_72) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45367_ ( .CLK(CLK), .D(_03150_), .Q(_tmp_73) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45368_ ( .CLK(CLK), .D(_03151_), .Q(_tmp_74) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45369_ ( .CLK(CLK), .D(_03152_), .Q(_tmp_75) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45370_ ( .CLK(CLK), .D(_03153_), .Q(_tmp_76) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45371_ ( .CLK(CLK), .D(_03154_), .Q(_tmp_77) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45372_ ( .CLK(CLK), .D(_03155_), .Q(_tmp_78) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45373_ ( .CLK(CLK), .D(_03156_), .Q(_tmp_79) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45374_ ( .CLK(CLK), .D(_03157_), .Q(_tmp_80) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45375_ ( .CLK(CLK), .D(_03171_), .Q(_tmp_99) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45376_ ( .CLK(CLK), .D(_02914_), .Q(_tmp_1138) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1139_reg  ( .CLK(CLK), .D(_02915_), .Q(_tmp_1139) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45378_ ( .CLK(CLK), .D(_03373_), .Q(ram_w4_l8192_id0_0_0_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45379_ ( .CLK(CLK), .D(_03374_), .Q(ram_w4_l8192_id0_0_1_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45380_ ( .CLK(CLK), .D(_03375_), .Q(ram_w4_l8192_id0_0_1_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) ram_w4_l8192_id0_0_1_wenable_reg  ( .CLK(CLK), .D(_03376_), .Q(ram_w4_l8192_id0_0_1_wenable) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(11) ) _45382_ ( .CLK(CLK), .D(_03098_), .Q(_tmp_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45383_ ( .CLK(CLK), .D(_03103_), .Q(_tmp_39) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_40_reg  ( .CLK(CLK), .D(_03110_), .Q(_tmp_40) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45385_ ( .CLK(CLK), .D(_03115_), .Q(_tmp_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45386_ ( .CLK(CLK), .D(_03120_), .Q(_tmp_42) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45387_ ( .CLK(CLK), .D(_03128_), .Q(_tmp_43) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45388_ ( .CLK(CLK), .D(_03136_), .Q(_tmp_44) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45389_ ( .CLK(CLK), .D(_03138_), .Q(_tmp_45) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45390_ ( .CLK(CLK), .D(_03139_), .Q(_tmp_46) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45391_ ( .CLK(CLK), .D(_03140_), .Q(_tmp_47) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45392_ ( .CLK(CLK), .D(_03141_), .Q(_tmp_48) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(10) ) _45393_ ( .CLK(CLK), .D(_03142_), .Q(_tmp_49) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45394_ ( .CLK(CLK), .D(_03145_), .Q(_tmp_68) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(34) ) _45395_ ( .CLK(CLK), .D(_02912_), .Q(_tmp_1136) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1137_reg  ( .CLK(CLK), .D(_02913_), .Q(_tmp_1137) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) RST_reg  ( .CLK(CLK), .D(_00000_), .Q(RST) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _rst_logic_1_reg  ( .CLK(CLK), .D(rst_logic), .Q(_rst_logic_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _rst_logic_2_reg  ( .CLK(CLK), .D(_rst_logic_1), .Q(_rst_logic_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45400_ ( .CLK(CLK), .D(_01869_), .Q(_saxi_register_fsm) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45401_ ( .CLK(CLK), .D(_03144_), .Q(_tmp_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) saxi_bvalid_reg  ( .CLK(CLK), .D(_03873_), .Q(saxi_bvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45403_ ( .CLK(CLK), .D(_03874_), .Q(saxi_rdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) saxi_rvalid_reg  ( .CLK(CLK), .D(_03875_), .Q(saxi_rvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45405_ ( .CLK(CLK), .D(_01855_), .Q(_saxi_register_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45406_ ( .CLK(CLK), .D(_01860_), .Q(_saxi_register_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45407_ ( .CLK(CLK), .D(_01861_), .Q(_saxi_register_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45408_ ( .CLK(CLK), .D(_01862_), .Q(_saxi_register_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45409_ ( .CLK(CLK), .D(_01863_), .Q(_saxi_register_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45410_ ( .CLK(CLK), .D(_01864_), .Q(_saxi_register_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45411_ ( .CLK(CLK), .D(_01865_), .Q(_saxi_register_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45412_ ( .CLK(CLK), .D(_01866_), .Q(_saxi_register_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45413_ ( .CLK(CLK), .D(_01867_), .Q(_saxi_register_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45414_ ( .CLK(CLK), .D(_01868_), .Q(_saxi_register_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45415_ ( .CLK(CLK), .D(_01856_), .Q(_saxi_register_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45416_ ( .CLK(CLK), .D(_01857_), .Q(_saxi_register_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45417_ ( .CLK(CLK), .D(_01858_), .Q(_saxi_register_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45418_ ( .CLK(CLK), .D(_01859_), .Q(_saxi_register_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_0_reg  ( .CLK(CLK), .D(_01841_), .Q(_saxi_flag_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_1_reg  ( .CLK(CLK), .D(_01846_), .Q(_saxi_flag_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_2_reg  ( .CLK(CLK), .D(_01847_), .Q(_saxi_flag_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_3_reg  ( .CLK(CLK), .D(_01848_), .Q(_saxi_flag_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_4_reg  ( .CLK(CLK), .D(_01849_), .Q(_saxi_flag_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_5_reg  ( .CLK(CLK), .D(_01850_), .Q(_saxi_flag_5) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_6_reg  ( .CLK(CLK), .D(_01851_), .Q(_saxi_flag_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_7_reg  ( .CLK(CLK), .D(_01852_), .Q(_saxi_flag_7) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_8_reg  ( .CLK(CLK), .D(_01853_), .Q(_saxi_flag_8) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_9_reg  ( .CLK(CLK), .D(_01854_), .Q(_saxi_flag_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_10_reg  ( .CLK(CLK), .D(_01842_), .Q(_saxi_flag_10) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_11_reg  ( .CLK(CLK), .D(_01843_), .Q(_saxi_flag_11) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_12_reg  ( .CLK(CLK), .D(_01844_), .Q(_saxi_flag_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_flag_13_reg  ( .CLK(CLK), .D(_01845_), .Q(_saxi_flag_13) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(6) ) _45433_ ( .CLK(CLK), .D(_02853_), .Q(_tmp_0) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1_reg  ( .CLK(CLK), .D(_03003_), .Q(_tmp_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_2_reg  ( .CLK(CLK), .D(_03048_), .Q(_tmp_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_3_reg  ( .CLK(CLK), .D(_03104_), .Q(_tmp_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_4_reg  ( .CLK(CLK), .D(_03143_), .Q(_tmp_4) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _saxi_cond_0_1_reg  ( .CLK(CLK), .D(_01704_), .Q(_saxi_cond_0_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45439_ ( .CLK(CLK), .D(_01617_), .Q(_dataflow_slice_data_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_3_reg  ( .CLK(CLK), .D(_01661_), .Q(_dataflow_slice_valid_3) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45441_ ( .CLK(CLK), .D(_01627_), .Q(_dataflow_slice_data_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_6_reg  ( .CLK(CLK), .D(_01671_), .Q(_dataflow_slice_valid_6) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45443_ ( .CLK(CLK), .D(_01635_), .Q(_dataflow_slice_data_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_9_reg  ( .CLK(CLK), .D(_01679_), .Q(_dataflow_slice_valid_9) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45445_ ( .CLK(CLK), .D(_01598_), .Q(_dataflow_slice_data_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_12_reg  ( .CLK(CLK), .D(_01642_), .Q(_dataflow_slice_valid_12) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45447_ ( .CLK(CLK), .D(_01609_), .Q(_dataflow_slice_data_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_16_reg  ( .CLK(CLK), .D(_01653_), .Q(_dataflow_slice_valid_16) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45449_ ( .CLK(CLK), .D(_01610_), .Q(_dataflow_slice_data_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_19_reg  ( .CLK(CLK), .D(_01654_), .Q(_dataflow_slice_valid_19) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45451_ ( .CLK(CLK), .D(_01611_), .Q(_dataflow_slice_data_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_22_reg  ( .CLK(CLK), .D(_01655_), .Q(_dataflow_slice_valid_22) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45453_ ( .CLK(CLK), .D(_01612_), .Q(_dataflow_slice_data_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_25_reg  ( .CLK(CLK), .D(_01656_), .Q(_dataflow_slice_valid_25) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45455_ ( .CLK(CLK), .D(_01613_), .Q(_dataflow_slice_data_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_29_reg  ( .CLK(CLK), .D(_01657_), .Q(_dataflow_slice_valid_29) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45457_ ( .CLK(CLK), .D(_01614_), .Q(_dataflow_slice_data_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_32_reg  ( .CLK(CLK), .D(_01658_), .Q(_dataflow_slice_valid_32) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45459_ ( .CLK(CLK), .D(_01615_), .Q(_dataflow_slice_data_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_35_reg  ( .CLK(CLK), .D(_01659_), .Q(_dataflow_slice_valid_35) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45461_ ( .CLK(CLK), .D(_01616_), .Q(_dataflow_slice_data_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_38_reg  ( .CLK(CLK), .D(_01660_), .Q(_dataflow_slice_valid_38) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45463_ ( .CLK(CLK), .D(_01618_), .Q(_dataflow_slice_data_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_41_reg  ( .CLK(CLK), .D(_01662_), .Q(_dataflow_slice_valid_41) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45465_ ( .CLK(CLK), .D(_01619_), .Q(_dataflow_slice_data_44) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_44_reg  ( .CLK(CLK), .D(_01663_), .Q(_dataflow_slice_valid_44) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45467_ ( .CLK(CLK), .D(_01620_), .Q(_dataflow_slice_data_47) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_47_reg  ( .CLK(CLK), .D(_01664_), .Q(_dataflow_slice_valid_47) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45469_ ( .CLK(CLK), .D(_01621_), .Q(_dataflow_slice_data_50) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_50_reg  ( .CLK(CLK), .D(_01665_), .Q(_dataflow_slice_valid_50) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45471_ ( .CLK(CLK), .D(_01622_), .Q(_dataflow_slice_data_54) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_54_reg  ( .CLK(CLK), .D(_01666_), .Q(_dataflow_slice_valid_54) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45473_ ( .CLK(CLK), .D(_01623_), .Q(_dataflow_slice_data_57) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_57_reg  ( .CLK(CLK), .D(_01667_), .Q(_dataflow_slice_valid_57) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45475_ ( .CLK(CLK), .D(_01624_), .Q(_dataflow_slice_data_60) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_60_reg  ( .CLK(CLK), .D(_01668_), .Q(_dataflow_slice_valid_60) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45477_ ( .CLK(CLK), .D(_01625_), .Q(_dataflow_slice_data_63) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_63_reg  ( .CLK(CLK), .D(_01669_), .Q(_dataflow_slice_valid_63) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45479_ ( .CLK(CLK), .D(_01626_), .Q(_dataflow_slice_data_67) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_67_reg  ( .CLK(CLK), .D(_01670_), .Q(_dataflow_slice_valid_67) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45481_ ( .CLK(CLK), .D(_01628_), .Q(_dataflow_slice_data_70) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_70_reg  ( .CLK(CLK), .D(_01672_), .Q(_dataflow_slice_valid_70) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45483_ ( .CLK(CLK), .D(_01629_), .Q(_dataflow_slice_data_73) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_73_reg  ( .CLK(CLK), .D(_01673_), .Q(_dataflow_slice_valid_73) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45485_ ( .CLK(CLK), .D(_01630_), .Q(_dataflow_slice_data_76) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_76_reg  ( .CLK(CLK), .D(_01674_), .Q(_dataflow_slice_valid_76) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45487_ ( .CLK(CLK), .D(_01631_), .Q(_dataflow_slice_data_80) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_80_reg  ( .CLK(CLK), .D(_01675_), .Q(_dataflow_slice_valid_80) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45489_ ( .CLK(CLK), .D(_01632_), .Q(_dataflow_slice_data_83) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_83_reg  ( .CLK(CLK), .D(_01676_), .Q(_dataflow_slice_valid_83) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45491_ ( .CLK(CLK), .D(_01633_), .Q(_dataflow_slice_data_86) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_86_reg  ( .CLK(CLK), .D(_01677_), .Q(_dataflow_slice_valid_86) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45493_ ( .CLK(CLK), .D(_01634_), .Q(_dataflow_slice_data_89) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_89_reg  ( .CLK(CLK), .D(_01678_), .Q(_dataflow_slice_valid_89) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45495_ ( .CLK(CLK), .D(_01592_), .Q(_dataflow_slice_data_111) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_111_reg  ( .CLK(CLK), .D(_01636_), .Q(_dataflow_slice_valid_111) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45497_ ( .CLK(CLK), .D(_01593_), .Q(_dataflow_slice_data_114) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_114_reg  ( .CLK(CLK), .D(_01637_), .Q(_dataflow_slice_valid_114) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45499_ ( .CLK(CLK), .D(_01594_), .Q(_dataflow_slice_data_117) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_117_reg  ( .CLK(CLK), .D(_01638_), .Q(_dataflow_slice_valid_117) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45501_ ( .CLK(CLK), .D(_01595_), .Q(_dataflow_slice_data_120) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_120_reg  ( .CLK(CLK), .D(_01639_), .Q(_dataflow_slice_valid_120) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45503_ ( .CLK(CLK), .D(_01596_), .Q(_dataflow_slice_data_124) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_124_reg  ( .CLK(CLK), .D(_01640_), .Q(_dataflow_slice_valid_124) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45505_ ( .CLK(CLK), .D(_01597_), .Q(_dataflow_slice_data_127) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_127_reg  ( .CLK(CLK), .D(_01641_), .Q(_dataflow_slice_valid_127) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45507_ ( .CLK(CLK), .D(_01599_), .Q(_dataflow_slice_data_130) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_130_reg  ( .CLK(CLK), .D(_01643_), .Q(_dataflow_slice_valid_130) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45509_ ( .CLK(CLK), .D(_01600_), .Q(_dataflow_slice_data_133) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_133_reg  ( .CLK(CLK), .D(_01644_), .Q(_dataflow_slice_valid_133) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45511_ ( .CLK(CLK), .D(_01601_), .Q(_dataflow_slice_data_136) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_136_reg  ( .CLK(CLK), .D(_01645_), .Q(_dataflow_slice_valid_136) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45513_ ( .CLK(CLK), .D(_01602_), .Q(_dataflow_slice_data_139) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_139_reg  ( .CLK(CLK), .D(_01646_), .Q(_dataflow_slice_valid_139) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45515_ ( .CLK(CLK), .D(_01603_), .Q(_dataflow_slice_data_142) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_142_reg  ( .CLK(CLK), .D(_01647_), .Q(_dataflow_slice_valid_142) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45517_ ( .CLK(CLK), .D(_01604_), .Q(_dataflow_slice_data_145) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_145_reg  ( .CLK(CLK), .D(_01648_), .Q(_dataflow_slice_valid_145) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45519_ ( .CLK(CLK), .D(_01605_), .Q(_dataflow_slice_data_149) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_149_reg  ( .CLK(CLK), .D(_01649_), .Q(_dataflow_slice_valid_149) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45521_ ( .CLK(CLK), .D(_01606_), .Q(_dataflow_slice_data_152) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_152_reg  ( .CLK(CLK), .D(_01650_), .Q(_dataflow_slice_valid_152) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45523_ ( .CLK(CLK), .D(_01607_), .Q(_dataflow_slice_data_155) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_155_reg  ( .CLK(CLK), .D(_01651_), .Q(_dataflow_slice_valid_155) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45525_ ( .CLK(CLK), .D(_01608_), .Q(_dataflow_slice_data_158) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _dataflow_slice_valid_158_reg  ( .CLK(CLK), .D(_01652_), .Q(_dataflow_slice_valid_158) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45527_ ( .CLK(CLK), .D(_03366_), .Q(maxi_awaddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45528_ ( .CLK(CLK), .D(_03367_), .Q(maxi_awlen) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) maxi_awvalid_reg  ( .CLK(CLK), .D(_03368_), .Q(maxi_awvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45530_ ( .CLK(CLK), .D(_03369_), .Q(maxi_wdata) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _45531_ ( .CLK(CLK), .D(_03371_), .Q(maxi_wstrb) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) maxi_wlast_reg  ( .CLK(CLK), .D(_03370_), .Q(maxi_wlast) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) maxi_wvalid_reg  ( .CLK(CLK), .D(_03372_), .Q(maxi_wvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45534_ ( .CLK(CLK), .D(_03363_), .Q(maxi_araddr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45535_ ( .CLK(CLK), .D(_03364_), .Q(maxi_arlen) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) maxi_arvalid_reg  ( .CLK(CLK), .D(_03365_), .Q(maxi_arvalid) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_read_start_reg  ( .CLK(CLK), .D(_01788_), .Q(_maxi_read_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45538_ ( .CLK(CLK), .D(_01785_), .Q(_maxi_read_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45539_ ( .CLK(CLK), .D(_01783_), .Q(_maxi_read_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45540_ ( .CLK(CLK), .D(_01781_), .Q(_maxi_read_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45541_ ( .CLK(CLK), .D(_01787_), .Q(_maxi_read_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45542_ ( .CLK(CLK), .D(_01784_), .Q(_maxi_read_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_read_idle_reg  ( .CLK(CLK), .D(_01782_), .Q(_maxi_read_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_write_start_reg  ( .CLK(CLK), .D(_01799_), .Q(_maxi_write_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45545_ ( .CLK(CLK), .D(_01796_), .Q(_maxi_write_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45546_ ( .CLK(CLK), .D(_01794_), .Q(_maxi_write_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45547_ ( .CLK(CLK), .D(_01792_), .Q(_maxi_write_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45548_ ( .CLK(CLK), .D(_01798_), .Q(_maxi_write_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45549_ ( .CLK(CLK), .D(_01795_), .Q(_maxi_write_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_write_idle_reg  ( .CLK(CLK), .D(_01793_), .Q(_maxi_write_idle) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45551_ ( .CLK(CLK), .D(_01705_), .Q(_maxi_global_base_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_ram_w8_l2048_id1_1_read_start_reg  ( .CLK(CLK), .D(_01741_), .Q(_maxi_ram_w8_l2048_id1_1_read_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45553_ ( .CLK(CLK), .D(_01739_), .Q(_maxi_ram_w8_l2048_id1_1_read_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45554_ ( .CLK(CLK), .D(_01737_), .Q(_maxi_ram_w8_l2048_id1_1_read_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45555_ ( .CLK(CLK), .D(_01736_), .Q(_maxi_ram_w8_l2048_id1_1_read_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45556_ ( .CLK(CLK), .D(_01740_), .Q(_maxi_ram_w8_l2048_id1_1_read_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45557_ ( .CLK(CLK), .D(_01738_), .Q(_maxi_ram_w8_l2048_id1_1_read_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _45558_ ( .CLK(CLK), .D(_03009_), .Q(_tmp_20) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_ram_w8_l2048_id0_1_read_start_reg  ( .CLK(CLK), .D(_01723_), .Q(_maxi_ram_w8_l2048_id0_1_read_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45560_ ( .CLK(CLK), .D(_01721_), .Q(_maxi_ram_w8_l2048_id0_1_read_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45561_ ( .CLK(CLK), .D(_01719_), .Q(_maxi_ram_w8_l2048_id0_1_read_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45562_ ( .CLK(CLK), .D(_01718_), .Q(_maxi_ram_w8_l2048_id0_1_read_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45563_ ( .CLK(CLK), .D(_01722_), .Q(_maxi_ram_w8_l2048_id0_1_read_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45564_ ( .CLK(CLK), .D(_01720_), .Q(_maxi_ram_w8_l2048_id0_1_read_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start_reg  ( .CLK(CLK), .D(_01717_), .Q(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45566_ ( .CLK(CLK), .D(_01715_), .Q(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45567_ ( .CLK(CLK), .D(_01713_), .Q(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45568_ ( .CLK(CLK), .D(_01712_), .Q(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45569_ ( .CLK(CLK), .D(_01716_), .Q(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45570_ ( .CLK(CLK), .D(_01714_), .Q(_maxi_ram_w4_l8192_id0_ram_w4_l8192_id1_ram_w4_l8192_id2_ram_w4_l8192_id3_ram_w4_l8192_id4_ram_w4_l8192_id5_ram_w4_l8192_id6_ram_w4_l8192_id7_ram_w4_l8192_id8_1_read_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start_reg  ( .CLK(CLK), .D(_01759_), .Q(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45572_ ( .CLK(CLK), .D(_01757_), .Q(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45573_ ( .CLK(CLK), .D(_01755_), .Q(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45574_ ( .CLK(CLK), .D(_01754_), .Q(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45575_ ( .CLK(CLK), .D(_01758_), .Q(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45576_ ( .CLK(CLK), .D(_01756_), .Q(_maxi_ram_w8_l2048_id2_ram_w8_l2048_id3_ram_w8_l2048_id4_1_read_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start_reg  ( .CLK(CLK), .D(_01771_), .Q(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45578_ ( .CLK(CLK), .D(_01769_), .Q(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45579_ ( .CLK(CLK), .D(_01767_), .Q(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45580_ ( .CLK(CLK), .D(_01766_), .Q(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45581_ ( .CLK(CLK), .D(_01770_), .Q(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45582_ ( .CLK(CLK), .D(_01768_), .Q(_maxi_ram_w8_l2048_id5_ram_w8_l2048_id6_ram_w8_l2048_id7_1_read_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start_reg  ( .CLK(CLK), .D(_01777_), .Q(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45584_ ( .CLK(CLK), .D(_01775_), .Q(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45585_ ( .CLK(CLK), .D(_01773_), .Q(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45586_ ( .CLK(CLK), .D(_01772_), .Q(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45587_ ( .CLK(CLK), .D(_01776_), .Q(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45588_ ( .CLK(CLK), .D(_01774_), .Q(_maxi_ram_w8_l2048_id8_ram_w8_l2048_id9_ram_w8_l2048_id10_1_read_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_ram_w8_l2048_id11_1_write_start_reg  ( .CLK(CLK), .D(_01735_), .Q(_maxi_ram_w8_l2048_id11_1_write_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45590_ ( .CLK(CLK), .D(_01733_), .Q(_maxi_ram_w8_l2048_id11_1_write_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45591_ ( .CLK(CLK), .D(_01731_), .Q(_maxi_ram_w8_l2048_id11_1_write_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45592_ ( .CLK(CLK), .D(_01730_), .Q(_maxi_ram_w8_l2048_id11_1_write_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45593_ ( .CLK(CLK), .D(_01734_), .Q(_maxi_ram_w8_l2048_id11_1_write_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45594_ ( .CLK(CLK), .D(_01732_), .Q(_maxi_ram_w8_l2048_id11_1_write_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(9) ) _45595_ ( .CLK(CLK), .D(_02866_), .Q(_tmp_1019) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1020_reg  ( .CLK(CLK), .D(_02868_), .Q(_tmp_1020) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_ram_w8_l2048_id0_1_write_start_reg  ( .CLK(CLK), .D(_01729_), .Q(_maxi_ram_w8_l2048_id0_1_write_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45598_ ( .CLK(CLK), .D(_01727_), .Q(_maxi_ram_w8_l2048_id0_1_write_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45599_ ( .CLK(CLK), .D(_01725_), .Q(_maxi_ram_w8_l2048_id0_1_write_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45600_ ( .CLK(CLK), .D(_01724_), .Q(_maxi_ram_w8_l2048_id0_1_write_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45601_ ( .CLK(CLK), .D(_01728_), .Q(_maxi_ram_w8_l2048_id0_1_write_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45602_ ( .CLK(CLK), .D(_01726_), .Q(_maxi_ram_w8_l2048_id0_1_write_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1120_reg  ( .CLK(CLK), .D(_02903_), .Q(_tmp_1120) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_ram_w8_l2048_id2_1_read_start_reg  ( .CLK(CLK), .D(_01753_), .Q(_maxi_ram_w8_l2048_id2_1_read_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45605_ ( .CLK(CLK), .D(_01751_), .Q(_maxi_ram_w8_l2048_id2_1_read_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45606_ ( .CLK(CLK), .D(_01749_), .Q(_maxi_ram_w8_l2048_id2_1_read_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45607_ ( .CLK(CLK), .D(_01748_), .Q(_maxi_ram_w8_l2048_id2_1_read_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45608_ ( .CLK(CLK), .D(_01752_), .Q(_maxi_ram_w8_l2048_id2_1_read_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45609_ ( .CLK(CLK), .D(_01750_), .Q(_maxi_ram_w8_l2048_id2_1_read_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_ram_w4_l8192_id0_1_read_start_reg  ( .CLK(CLK), .D(_01711_), .Q(_maxi_ram_w4_l8192_id0_1_read_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45611_ ( .CLK(CLK), .D(_01709_), .Q(_maxi_ram_w4_l8192_id0_1_read_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45612_ ( .CLK(CLK), .D(_01707_), .Q(_maxi_ram_w4_l8192_id0_1_read_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45613_ ( .CLK(CLK), .D(_01706_), .Q(_maxi_ram_w4_l8192_id0_1_read_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45614_ ( .CLK(CLK), .D(_01710_), .Q(_maxi_ram_w4_l8192_id0_1_read_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45615_ ( .CLK(CLK), .D(_01708_), .Q(_maxi_ram_w4_l8192_id0_1_read_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_ram_w8_l2048_id3_1_read_start_reg  ( .CLK(CLK), .D(_01765_), .Q(_maxi_ram_w8_l2048_id3_1_read_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45617_ ( .CLK(CLK), .D(_01763_), .Q(_maxi_ram_w8_l2048_id3_1_read_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45618_ ( .CLK(CLK), .D(_01761_), .Q(_maxi_ram_w8_l2048_id3_1_read_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45619_ ( .CLK(CLK), .D(_01760_), .Q(_maxi_ram_w8_l2048_id3_1_read_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45620_ ( .CLK(CLK), .D(_01764_), .Q(_maxi_ram_w8_l2048_id3_1_read_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45621_ ( .CLK(CLK), .D(_01762_), .Q(_maxi_ram_w8_l2048_id3_1_read_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _maxi_ram_w8_l2048_id1_1_write_start_reg  ( .CLK(CLK), .D(_01747_), .Q(_maxi_ram_w8_l2048_id1_1_write_start) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _45623_ ( .CLK(CLK), .D(_01745_), .Q(_maxi_ram_w8_l2048_id1_1_write_op_sel) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45624_ ( .CLK(CLK), .D(_01743_), .Q(_maxi_ram_w8_l2048_id1_1_write_local_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45625_ ( .CLK(CLK), .D(_01742_), .Q(_maxi_ram_w8_l2048_id1_1_write_global_addr) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(33) ) _45626_ ( .CLK(CLK), .D(_01746_), .Q(_maxi_ram_w8_l2048_id1_1_write_size) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _45627_ ( .CLK(CLK), .D(_01744_), .Q(_maxi_ram_w8_l2048_id1_1_write_local_stride) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _tmp_1357_reg  ( .CLK(CLK), .D(_02966_), .Q(_tmp_1357) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _RESETN_inv_1_reg  ( .CLK(CLK), .D(RESETN_inv), .Q(_RESETN_inv_1) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(1) ) _RESETN_inv_2_reg  ( .CLK(CLK), .D(_RESETN_inv_1), .Q(_RESETN_inv_2) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54134_ ( .CLK(CLK), .D(_cond_data_101), .Q(\__muladd_madd_103.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _54135_ ( .CLK(CLK), .D(__delay_data_633), .Q(\__muladd_madd_103.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54136_ ( .CLK(CLK), .D(\__muladd_madd_103.madd._madd ), .Q(\__muladd_madd_103.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _54137_ ( .CLK(CLK), .D(__delay_data_630), .Q(\__muladd_madd_103.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54138_ ( .CLK(CLK), .D(\__muladd_madd_103.madd._pipe_madd0 ), .Q(\__muladd_madd_103.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54141_ ( .CLK(CLK), .D(_cond_data_118), .Q(\__muladd_madd_120.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _54142_ ( .CLK(CLK), .D(__delay_data_650), .Q(\__muladd_madd_120.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54143_ ( .CLK(CLK), .D(\__muladd_madd_120.madd._madd ), .Q(\__muladd_madd_120.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _54144_ ( .CLK(CLK), .D(__delay_data_647), .Q(\__muladd_madd_120.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54145_ ( .CLK(CLK), .D(\__muladd_madd_120.madd._pipe_madd0 ), .Q(\__muladd_madd_120.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54148_ ( .CLK(CLK), .D(_cond_data_135), .Q(\__muladd_madd_137.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _54149_ ( .CLK(CLK), .D(__delay_data_667), .Q(\__muladd_madd_137.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54150_ ( .CLK(CLK), .D(\__muladd_madd_137.madd._madd ), .Q(\__muladd_madd_137.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _54151_ ( .CLK(CLK), .D(__delay_data_664), .Q(\__muladd_madd_137.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54152_ ( .CLK(CLK), .D(\__muladd_madd_137.madd._pipe_madd0 ), .Q(\__muladd_madd_137.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54155_ ( .CLK(CLK), .D(_cond_data_152), .Q(\__muladd_madd_154.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _54156_ ( .CLK(CLK), .D(__delay_data_684), .Q(\__muladd_madd_154.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54157_ ( .CLK(CLK), .D(\__muladd_madd_154.madd._madd ), .Q(\__muladd_madd_154.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _54158_ ( .CLK(CLK), .D(__delay_data_681), .Q(\__muladd_madd_154.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54159_ ( .CLK(CLK), .D(\__muladd_madd_154.madd._pipe_madd0 ), .Q(\__muladd_madd_154.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54162_ ( .CLK(CLK), .D(_cond_data_169), .Q(\__muladd_madd_171.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _54163_ ( .CLK(CLK), .D(__delay_data_701), .Q(\__muladd_madd_171.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54164_ ( .CLK(CLK), .D(\__muladd_madd_171.madd._madd ), .Q(\__muladd_madd_171.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _54165_ ( .CLK(CLK), .D(__delay_data_698), .Q(\__muladd_madd_171.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54166_ ( .CLK(CLK), .D(\__muladd_madd_171.madd._pipe_madd0 ), .Q(\__muladd_madd_171.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54169_ ( .CLK(CLK), .D(_cond_data_186), .Q(\__muladd_madd_188.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _54170_ ( .CLK(CLK), .D(__delay_data_718), .Q(\__muladd_madd_188.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54171_ ( .CLK(CLK), .D(\__muladd_madd_188.madd._madd ), .Q(\__muladd_madd_188.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _54172_ ( .CLK(CLK), .D(__delay_data_715), .Q(\__muladd_madd_188.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54173_ ( .CLK(CLK), .D(\__muladd_madd_188.madd._pipe_madd0 ), .Q(\__muladd_madd_188.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54176_ ( .CLK(CLK), .D(_cond_data_203), .Q(\__muladd_madd_205.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _54177_ ( .CLK(CLK), .D(__delay_data_735), .Q(\__muladd_madd_205.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54178_ ( .CLK(CLK), .D(\__muladd_madd_205.madd._madd ), .Q(\__muladd_madd_205.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _54179_ ( .CLK(CLK), .D(__delay_data_732), .Q(\__muladd_madd_205.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54180_ ( .CLK(CLK), .D(\__muladd_madd_205.madd._pipe_madd0 ), .Q(\__muladd_madd_205.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54183_ ( .CLK(CLK), .D(_cond_data_67), .Q(\__muladd_madd_69.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _54184_ ( .CLK(CLK), .D(__delay_data_599), .Q(\__muladd_madd_69.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54185_ ( .CLK(CLK), .D(\__muladd_madd_69.madd._madd ), .Q(\__muladd_madd_69.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _54186_ ( .CLK(CLK), .D(__delay_data_596), .Q(\__muladd_madd_69.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54187_ ( .CLK(CLK), .D(\__muladd_madd_69.madd._pipe_madd0 ), .Q(\__muladd_madd_69.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54190_ ( .CLK(CLK), .D(_cond_data_84), .Q(\__muladd_madd_86.madd._c ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(4) ) _54191_ ( .CLK(CLK), .D(__delay_data_616), .Q(\__muladd_madd_86.madd._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54192_ ( .CLK(CLK), .D(\__muladd_madd_86.madd._madd ), .Q(\__muladd_madd_86.madd._pipe_madd0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _54193_ ( .CLK(CLK), .D(__delay_data_613), .Q(\__muladd_madd_86.madd._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(12) ) _54194_ ( .CLK(CLK), .D(\__muladd_madd_86.madd._pipe_madd0 ), .Q(\__muladd_madd_86.madd._pipe_madd1 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(8) ) _54196_ ( .CLK(CLK), .D(__variable_wdata_39), .Q(\_times_mul_41.mult._b ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(32) ) _54197_ ( .CLK(CLK), .D(__variable_wdata_38), .Q(\_times_mul_41.mult._a ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(40) ) _54198_ ( .CLK(CLK), .D(\_times_mul_41.mult._mul ), .Q(\_times_mul_41.mult._pipe_mul0 ) );
  \$dff  #( .CLK_POLARITY(1'h1), .WIDTH(40) ) _54199_ ( .CLK(CLK), .D(\_times_mul_41.mult._pipe_mul0 ), .Q(\_times_mul_41.mult._pipe_mul1 ) );
  ram_w4_l8192_id0_0 inst_ram_w4_l8192_id0_0 ( .CLK(CLK), .ram_w4_l8192_id0_0_0_addr(ram_w4_l8192_id0_0_0_addr), .ram_w4_l8192_id0_0_0_rdata(ram_w4_l8192_id0_0_0_rdata), .ram_w4_l8192_id0_0_0_wdata(4'h0), .ram_w4_l8192_id0_0_0_wenable(1'h0), .ram_w4_l8192_id0_0_1_addr(ram_w4_l8192_id0_0_1_addr), .ram_w4_l8192_id0_0_1_rdata(ram_w4_l8192_id0_0_1_rdata), .ram_w4_l8192_id0_0_1_wdata(ram_w4_l8192_id0_0_1_wdata), .ram_w4_l8192_id0_0_1_wenable(ram_w4_l8192_id0_0_1_wenable) );
  ram_w4_l8192_id0_1 inst_ram_w4_l8192_id0_1 ( .CLK(CLK), .ram_w4_l8192_id0_1_0_addr(ram_w4_l8192_id0_1_0_addr), .ram_w4_l8192_id0_1_0_rdata(ram_w4_l8192_id0_1_0_rdata), .ram_w4_l8192_id0_1_0_wdata(4'h0), .ram_w4_l8192_id0_1_0_wenable(1'h0), .ram_w4_l8192_id0_1_1_addr(ram_w4_l8192_id0_1_1_addr), .ram_w4_l8192_id0_1_1_rdata(ram_w4_l8192_id0_1_1_rdata), .ram_w4_l8192_id0_1_1_wdata(ram_w4_l8192_id0_1_1_wdata), .ram_w4_l8192_id0_1_1_wenable(ram_w4_l8192_id0_1_1_wenable) );
  ram_w4_l8192_id0_2 inst_ram_w4_l8192_id0_2 ( .CLK(CLK), .ram_w4_l8192_id0_2_0_addr(ram_w4_l8192_id0_2_0_addr), .ram_w4_l8192_id0_2_0_rdata(ram_w4_l8192_id0_2_0_rdata), .ram_w4_l8192_id0_2_0_wdata(4'h0), .ram_w4_l8192_id0_2_0_wenable(1'h0), .ram_w4_l8192_id0_2_1_addr(ram_w4_l8192_id0_2_1_addr), .ram_w4_l8192_id0_2_1_rdata(ram_w4_l8192_id0_2_1_rdata), .ram_w4_l8192_id0_2_1_wdata(ram_w4_l8192_id0_2_1_wdata), .ram_w4_l8192_id0_2_1_wenable(ram_w4_l8192_id0_2_1_wenable) );
  ram_w4_l8192_id0_3 inst_ram_w4_l8192_id0_3 ( .CLK(CLK), .ram_w4_l8192_id0_3_0_addr(ram_w4_l8192_id0_3_0_addr), .ram_w4_l8192_id0_3_0_rdata(ram_w4_l8192_id0_3_0_rdata), .ram_w4_l8192_id0_3_0_wdata(4'h0), .ram_w4_l8192_id0_3_0_wenable(1'h0), .ram_w4_l8192_id0_3_1_addr(ram_w4_l8192_id0_3_1_addr), .ram_w4_l8192_id0_3_1_rdata(ram_w4_l8192_id0_3_1_rdata), .ram_w4_l8192_id0_3_1_wdata(ram_w4_l8192_id0_3_1_wdata), .ram_w4_l8192_id0_3_1_wenable(ram_w4_l8192_id0_3_1_wenable) );
  ram_w4_l8192_id0_4 inst_ram_w4_l8192_id0_4 ( .CLK(CLK), .ram_w4_l8192_id0_4_0_addr(ram_w4_l8192_id0_4_0_addr), .ram_w4_l8192_id0_4_0_rdata(ram_w4_l8192_id0_4_0_rdata), .ram_w4_l8192_id0_4_0_wdata(4'h0), .ram_w4_l8192_id0_4_0_wenable(1'h0), .ram_w4_l8192_id0_4_1_addr(ram_w4_l8192_id0_4_1_addr), .ram_w4_l8192_id0_4_1_rdata(ram_w4_l8192_id0_4_1_rdata), .ram_w4_l8192_id0_4_1_wdata(ram_w4_l8192_id0_4_1_wdata), .ram_w4_l8192_id0_4_1_wenable(ram_w4_l8192_id0_4_1_wenable) );
  ram_w4_l8192_id0_5 inst_ram_w4_l8192_id0_5 ( .CLK(CLK), .ram_w4_l8192_id0_5_0_addr(ram_w4_l8192_id0_5_0_addr), .ram_w4_l8192_id0_5_0_rdata(ram_w4_l8192_id0_5_0_rdata), .ram_w4_l8192_id0_5_0_wdata(4'h0), .ram_w4_l8192_id0_5_0_wenable(1'h0), .ram_w4_l8192_id0_5_1_addr(ram_w4_l8192_id0_5_1_addr), .ram_w4_l8192_id0_5_1_rdata(ram_w4_l8192_id0_5_1_rdata), .ram_w4_l8192_id0_5_1_wdata(ram_w4_l8192_id0_5_1_wdata), .ram_w4_l8192_id0_5_1_wenable(ram_w4_l8192_id0_5_1_wenable) );
  ram_w4_l8192_id0_6 inst_ram_w4_l8192_id0_6 ( .CLK(CLK), .ram_w4_l8192_id0_6_0_addr(ram_w4_l8192_id0_6_0_addr), .ram_w4_l8192_id0_6_0_rdata(ram_w4_l8192_id0_6_0_rdata), .ram_w4_l8192_id0_6_0_wdata(4'h0), .ram_w4_l8192_id0_6_0_wenable(1'h0), .ram_w4_l8192_id0_6_1_addr(ram_w4_l8192_id0_6_1_addr), .ram_w4_l8192_id0_6_1_rdata(ram_w4_l8192_id0_6_1_rdata), .ram_w4_l8192_id0_6_1_wdata(ram_w4_l8192_id0_6_1_wdata), .ram_w4_l8192_id0_6_1_wenable(ram_w4_l8192_id0_6_1_wenable) );
  ram_w4_l8192_id0_7 inst_ram_w4_l8192_id0_7 ( .CLK(CLK), .ram_w4_l8192_id0_7_0_addr(ram_w4_l8192_id0_7_0_addr), .ram_w4_l8192_id0_7_0_rdata(ram_w4_l8192_id0_7_0_rdata), .ram_w4_l8192_id0_7_0_wdata(4'h0), .ram_w4_l8192_id0_7_0_wenable(1'h0), .ram_w4_l8192_id0_7_1_addr(ram_w4_l8192_id0_7_1_addr), .ram_w4_l8192_id0_7_1_rdata(ram_w4_l8192_id0_7_1_rdata), .ram_w4_l8192_id0_7_1_wdata(ram_w4_l8192_id0_7_1_wdata), .ram_w4_l8192_id0_7_1_wenable(ram_w4_l8192_id0_7_1_wenable) );
  ram_w4_l8192_id1_0 inst_ram_w4_l8192_id1_0 ( .CLK(CLK), .ram_w4_l8192_id1_0_0_addr(ram_w4_l8192_id1_0_0_addr), .ram_w4_l8192_id1_0_0_rdata(ram_w4_l8192_id1_0_0_rdata), .ram_w4_l8192_id1_0_0_wdata(4'h0), .ram_w4_l8192_id1_0_0_wenable(1'h0), .ram_w4_l8192_id1_0_1_addr(ram_w4_l8192_id1_0_1_addr), .ram_w4_l8192_id1_0_1_rdata(ram_w4_l8192_id1_0_1_rdata), .ram_w4_l8192_id1_0_1_wdata(ram_w4_l8192_id1_0_1_wdata), .ram_w4_l8192_id1_0_1_wenable(ram_w4_l8192_id1_0_1_wenable) );
  ram_w4_l8192_id1_1 inst_ram_w4_l8192_id1_1 ( .CLK(CLK), .ram_w4_l8192_id1_1_0_addr(ram_w4_l8192_id1_1_0_addr), .ram_w4_l8192_id1_1_0_rdata(ram_w4_l8192_id1_1_0_rdata), .ram_w4_l8192_id1_1_0_wdata(4'h0), .ram_w4_l8192_id1_1_0_wenable(1'h0), .ram_w4_l8192_id1_1_1_addr(ram_w4_l8192_id1_1_1_addr), .ram_w4_l8192_id1_1_1_rdata(ram_w4_l8192_id1_1_1_rdata), .ram_w4_l8192_id1_1_1_wdata(ram_w4_l8192_id1_1_1_wdata), .ram_w4_l8192_id1_1_1_wenable(ram_w4_l8192_id1_1_1_wenable) );
  ram_w4_l8192_id1_2 inst_ram_w4_l8192_id1_2 ( .CLK(CLK), .ram_w4_l8192_id1_2_0_addr(ram_w4_l8192_id1_2_0_addr), .ram_w4_l8192_id1_2_0_rdata(ram_w4_l8192_id1_2_0_rdata), .ram_w4_l8192_id1_2_0_wdata(4'h0), .ram_w4_l8192_id1_2_0_wenable(1'h0), .ram_w4_l8192_id1_2_1_addr(ram_w4_l8192_id1_2_1_addr), .ram_w4_l8192_id1_2_1_rdata(ram_w4_l8192_id1_2_1_rdata), .ram_w4_l8192_id1_2_1_wdata(ram_w4_l8192_id1_2_1_wdata), .ram_w4_l8192_id1_2_1_wenable(ram_w4_l8192_id1_2_1_wenable) );
  ram_w4_l8192_id1_3 inst_ram_w4_l8192_id1_3 ( .CLK(CLK), .ram_w4_l8192_id1_3_0_addr(ram_w4_l8192_id1_3_0_addr), .ram_w4_l8192_id1_3_0_rdata(ram_w4_l8192_id1_3_0_rdata), .ram_w4_l8192_id1_3_0_wdata(4'h0), .ram_w4_l8192_id1_3_0_wenable(1'h0), .ram_w4_l8192_id1_3_1_addr(ram_w4_l8192_id1_3_1_addr), .ram_w4_l8192_id1_3_1_rdata(ram_w4_l8192_id1_3_1_rdata), .ram_w4_l8192_id1_3_1_wdata(ram_w4_l8192_id1_3_1_wdata), .ram_w4_l8192_id1_3_1_wenable(ram_w4_l8192_id1_3_1_wenable) );
  ram_w4_l8192_id1_4 inst_ram_w4_l8192_id1_4 ( .CLK(CLK), .ram_w4_l8192_id1_4_0_addr(ram_w4_l8192_id1_4_0_addr), .ram_w4_l8192_id1_4_0_rdata(ram_w4_l8192_id1_4_0_rdata), .ram_w4_l8192_id1_4_0_wdata(4'h0), .ram_w4_l8192_id1_4_0_wenable(1'h0), .ram_w4_l8192_id1_4_1_addr(ram_w4_l8192_id1_4_1_addr), .ram_w4_l8192_id1_4_1_rdata(ram_w4_l8192_id1_4_1_rdata), .ram_w4_l8192_id1_4_1_wdata(ram_w4_l8192_id1_4_1_wdata), .ram_w4_l8192_id1_4_1_wenable(ram_w4_l8192_id1_4_1_wenable) );
  ram_w4_l8192_id1_5 inst_ram_w4_l8192_id1_5 ( .CLK(CLK), .ram_w4_l8192_id1_5_0_addr(ram_w4_l8192_id1_5_0_addr), .ram_w4_l8192_id1_5_0_rdata(ram_w4_l8192_id1_5_0_rdata), .ram_w4_l8192_id1_5_0_wdata(4'h0), .ram_w4_l8192_id1_5_0_wenable(1'h0), .ram_w4_l8192_id1_5_1_addr(ram_w4_l8192_id1_5_1_addr), .ram_w4_l8192_id1_5_1_rdata(ram_w4_l8192_id1_5_1_rdata), .ram_w4_l8192_id1_5_1_wdata(ram_w4_l8192_id1_5_1_wdata), .ram_w4_l8192_id1_5_1_wenable(ram_w4_l8192_id1_5_1_wenable) );
  ram_w4_l8192_id1_6 inst_ram_w4_l8192_id1_6 ( .CLK(CLK), .ram_w4_l8192_id1_6_0_addr(ram_w4_l8192_id1_6_0_addr), .ram_w4_l8192_id1_6_0_rdata(ram_w4_l8192_id1_6_0_rdata), .ram_w4_l8192_id1_6_0_wdata(4'h0), .ram_w4_l8192_id1_6_0_wenable(1'h0), .ram_w4_l8192_id1_6_1_addr(ram_w4_l8192_id1_6_1_addr), .ram_w4_l8192_id1_6_1_rdata(ram_w4_l8192_id1_6_1_rdata), .ram_w4_l8192_id1_6_1_wdata(ram_w4_l8192_id1_6_1_wdata), .ram_w4_l8192_id1_6_1_wenable(ram_w4_l8192_id1_6_1_wenable) );
  ram_w4_l8192_id1_7 inst_ram_w4_l8192_id1_7 ( .CLK(CLK), .ram_w4_l8192_id1_7_0_addr(ram_w4_l8192_id1_7_0_addr), .ram_w4_l8192_id1_7_0_rdata(ram_w4_l8192_id1_7_0_rdata), .ram_w4_l8192_id1_7_0_wdata(4'h0), .ram_w4_l8192_id1_7_0_wenable(1'h0), .ram_w4_l8192_id1_7_1_addr(ram_w4_l8192_id1_7_1_addr), .ram_w4_l8192_id1_7_1_rdata(ram_w4_l8192_id1_7_1_rdata), .ram_w4_l8192_id1_7_1_wdata(ram_w4_l8192_id1_7_1_wdata), .ram_w4_l8192_id1_7_1_wenable(ram_w4_l8192_id1_7_1_wenable) );
  ram_w4_l8192_id2_0 inst_ram_w4_l8192_id2_0 ( .CLK(CLK), .ram_w4_l8192_id2_0_0_addr(ram_w4_l8192_id2_0_0_addr), .ram_w4_l8192_id2_0_0_rdata(ram_w4_l8192_id2_0_0_rdata), .ram_w4_l8192_id2_0_0_wdata(4'h0), .ram_w4_l8192_id2_0_0_wenable(1'h0), .ram_w4_l8192_id2_0_1_addr(ram_w4_l8192_id2_0_1_addr), .ram_w4_l8192_id2_0_1_rdata(ram_w4_l8192_id2_0_1_rdata), .ram_w4_l8192_id2_0_1_wdata(ram_w4_l8192_id2_0_1_wdata), .ram_w4_l8192_id2_0_1_wenable(ram_w4_l8192_id2_0_1_wenable) );
  ram_w4_l8192_id2_1 inst_ram_w4_l8192_id2_1 ( .CLK(CLK), .ram_w4_l8192_id2_1_0_addr(ram_w4_l8192_id2_1_0_addr), .ram_w4_l8192_id2_1_0_rdata(ram_w4_l8192_id2_1_0_rdata), .ram_w4_l8192_id2_1_0_wdata(4'h0), .ram_w4_l8192_id2_1_0_wenable(1'h0), .ram_w4_l8192_id2_1_1_addr(ram_w4_l8192_id2_1_1_addr), .ram_w4_l8192_id2_1_1_rdata(ram_w4_l8192_id2_1_1_rdata), .ram_w4_l8192_id2_1_1_wdata(ram_w4_l8192_id2_1_1_wdata), .ram_w4_l8192_id2_1_1_wenable(ram_w4_l8192_id2_1_1_wenable) );
  ram_w4_l8192_id2_2 inst_ram_w4_l8192_id2_2 ( .CLK(CLK), .ram_w4_l8192_id2_2_0_addr(ram_w4_l8192_id2_2_0_addr), .ram_w4_l8192_id2_2_0_rdata(ram_w4_l8192_id2_2_0_rdata), .ram_w4_l8192_id2_2_0_wdata(4'h0), .ram_w4_l8192_id2_2_0_wenable(1'h0), .ram_w4_l8192_id2_2_1_addr(ram_w4_l8192_id2_2_1_addr), .ram_w4_l8192_id2_2_1_rdata(ram_w4_l8192_id2_2_1_rdata), .ram_w4_l8192_id2_2_1_wdata(ram_w4_l8192_id2_2_1_wdata), .ram_w4_l8192_id2_2_1_wenable(ram_w4_l8192_id2_2_1_wenable) );
  ram_w4_l8192_id2_3 inst_ram_w4_l8192_id2_3 ( .CLK(CLK), .ram_w4_l8192_id2_3_0_addr(ram_w4_l8192_id2_3_0_addr), .ram_w4_l8192_id2_3_0_rdata(ram_w4_l8192_id2_3_0_rdata), .ram_w4_l8192_id2_3_0_wdata(4'h0), .ram_w4_l8192_id2_3_0_wenable(1'h0), .ram_w4_l8192_id2_3_1_addr(ram_w4_l8192_id2_3_1_addr), .ram_w4_l8192_id2_3_1_rdata(ram_w4_l8192_id2_3_1_rdata), .ram_w4_l8192_id2_3_1_wdata(ram_w4_l8192_id2_3_1_wdata), .ram_w4_l8192_id2_3_1_wenable(ram_w4_l8192_id2_3_1_wenable) );
  ram_w4_l8192_id2_4 inst_ram_w4_l8192_id2_4 ( .CLK(CLK), .ram_w4_l8192_id2_4_0_addr(ram_w4_l8192_id2_4_0_addr), .ram_w4_l8192_id2_4_0_rdata(ram_w4_l8192_id2_4_0_rdata), .ram_w4_l8192_id2_4_0_wdata(4'h0), .ram_w4_l8192_id2_4_0_wenable(1'h0), .ram_w4_l8192_id2_4_1_addr(ram_w4_l8192_id2_4_1_addr), .ram_w4_l8192_id2_4_1_rdata(ram_w4_l8192_id2_4_1_rdata), .ram_w4_l8192_id2_4_1_wdata(ram_w4_l8192_id2_4_1_wdata), .ram_w4_l8192_id2_4_1_wenable(ram_w4_l8192_id2_4_1_wenable) );
  ram_w4_l8192_id2_5 inst_ram_w4_l8192_id2_5 ( .CLK(CLK), .ram_w4_l8192_id2_5_0_addr(ram_w4_l8192_id2_5_0_addr), .ram_w4_l8192_id2_5_0_rdata(ram_w4_l8192_id2_5_0_rdata), .ram_w4_l8192_id2_5_0_wdata(4'h0), .ram_w4_l8192_id2_5_0_wenable(1'h0), .ram_w4_l8192_id2_5_1_addr(ram_w4_l8192_id2_5_1_addr), .ram_w4_l8192_id2_5_1_rdata(ram_w4_l8192_id2_5_1_rdata), .ram_w4_l8192_id2_5_1_wdata(ram_w4_l8192_id2_5_1_wdata), .ram_w4_l8192_id2_5_1_wenable(ram_w4_l8192_id2_5_1_wenable) );
  ram_w4_l8192_id2_6 inst_ram_w4_l8192_id2_6 ( .CLK(CLK), .ram_w4_l8192_id2_6_0_addr(ram_w4_l8192_id2_6_0_addr), .ram_w4_l8192_id2_6_0_rdata(ram_w4_l8192_id2_6_0_rdata), .ram_w4_l8192_id2_6_0_wdata(4'h0), .ram_w4_l8192_id2_6_0_wenable(1'h0), .ram_w4_l8192_id2_6_1_addr(ram_w4_l8192_id2_6_1_addr), .ram_w4_l8192_id2_6_1_rdata(ram_w4_l8192_id2_6_1_rdata), .ram_w4_l8192_id2_6_1_wdata(ram_w4_l8192_id2_6_1_wdata), .ram_w4_l8192_id2_6_1_wenable(ram_w4_l8192_id2_6_1_wenable) );
  ram_w4_l8192_id2_7 inst_ram_w4_l8192_id2_7 ( .CLK(CLK), .ram_w4_l8192_id2_7_0_addr(ram_w4_l8192_id2_7_0_addr), .ram_w4_l8192_id2_7_0_rdata(ram_w4_l8192_id2_7_0_rdata), .ram_w4_l8192_id2_7_0_wdata(4'h0), .ram_w4_l8192_id2_7_0_wenable(1'h0), .ram_w4_l8192_id2_7_1_addr(ram_w4_l8192_id2_7_1_addr), .ram_w4_l8192_id2_7_1_rdata(ram_w4_l8192_id2_7_1_rdata), .ram_w4_l8192_id2_7_1_wdata(ram_w4_l8192_id2_7_1_wdata), .ram_w4_l8192_id2_7_1_wenable(ram_w4_l8192_id2_7_1_wenable) );
  ram_w4_l8192_id3_0 inst_ram_w4_l8192_id3_0 ( .CLK(CLK), .ram_w4_l8192_id3_0_0_addr(ram_w4_l8192_id3_0_0_addr), .ram_w4_l8192_id3_0_0_rdata(ram_w4_l8192_id3_0_0_rdata), .ram_w4_l8192_id3_0_0_wdata(4'h0), .ram_w4_l8192_id3_0_0_wenable(1'h0), .ram_w4_l8192_id3_0_1_addr(ram_w4_l8192_id3_0_1_addr), .ram_w4_l8192_id3_0_1_rdata(ram_w4_l8192_id3_0_1_rdata), .ram_w4_l8192_id3_0_1_wdata(ram_w4_l8192_id3_0_1_wdata), .ram_w4_l8192_id3_0_1_wenable(ram_w4_l8192_id3_0_1_wenable) );
  ram_w4_l8192_id3_1 inst_ram_w4_l8192_id3_1 ( .CLK(CLK), .ram_w4_l8192_id3_1_0_addr(ram_w4_l8192_id3_1_0_addr), .ram_w4_l8192_id3_1_0_rdata(ram_w4_l8192_id3_1_0_rdata), .ram_w4_l8192_id3_1_0_wdata(4'h0), .ram_w4_l8192_id3_1_0_wenable(1'h0), .ram_w4_l8192_id3_1_1_addr(ram_w4_l8192_id3_1_1_addr), .ram_w4_l8192_id3_1_1_rdata(ram_w4_l8192_id3_1_1_rdata), .ram_w4_l8192_id3_1_1_wdata(ram_w4_l8192_id3_1_1_wdata), .ram_w4_l8192_id3_1_1_wenable(ram_w4_l8192_id3_1_1_wenable) );
  ram_w4_l8192_id3_2 inst_ram_w4_l8192_id3_2 ( .CLK(CLK), .ram_w4_l8192_id3_2_0_addr(ram_w4_l8192_id3_2_0_addr), .ram_w4_l8192_id3_2_0_rdata(ram_w4_l8192_id3_2_0_rdata), .ram_w4_l8192_id3_2_0_wdata(4'h0), .ram_w4_l8192_id3_2_0_wenable(1'h0), .ram_w4_l8192_id3_2_1_addr(ram_w4_l8192_id3_2_1_addr), .ram_w4_l8192_id3_2_1_rdata(ram_w4_l8192_id3_2_1_rdata), .ram_w4_l8192_id3_2_1_wdata(ram_w4_l8192_id3_2_1_wdata), .ram_w4_l8192_id3_2_1_wenable(ram_w4_l8192_id3_2_1_wenable) );
  ram_w4_l8192_id3_3 inst_ram_w4_l8192_id3_3 ( .CLK(CLK), .ram_w4_l8192_id3_3_0_addr(ram_w4_l8192_id3_3_0_addr), .ram_w4_l8192_id3_3_0_rdata(ram_w4_l8192_id3_3_0_rdata), .ram_w4_l8192_id3_3_0_wdata(4'h0), .ram_w4_l8192_id3_3_0_wenable(1'h0), .ram_w4_l8192_id3_3_1_addr(ram_w4_l8192_id3_3_1_addr), .ram_w4_l8192_id3_3_1_rdata(ram_w4_l8192_id3_3_1_rdata), .ram_w4_l8192_id3_3_1_wdata(ram_w4_l8192_id3_3_1_wdata), .ram_w4_l8192_id3_3_1_wenable(ram_w4_l8192_id3_3_1_wenable) );
  ram_w4_l8192_id3_4 inst_ram_w4_l8192_id3_4 ( .CLK(CLK), .ram_w4_l8192_id3_4_0_addr(ram_w4_l8192_id3_4_0_addr), .ram_w4_l8192_id3_4_0_rdata(ram_w4_l8192_id3_4_0_rdata), .ram_w4_l8192_id3_4_0_wdata(4'h0), .ram_w4_l8192_id3_4_0_wenable(1'h0), .ram_w4_l8192_id3_4_1_addr(ram_w4_l8192_id3_4_1_addr), .ram_w4_l8192_id3_4_1_rdata(ram_w4_l8192_id3_4_1_rdata), .ram_w4_l8192_id3_4_1_wdata(ram_w4_l8192_id3_4_1_wdata), .ram_w4_l8192_id3_4_1_wenable(ram_w4_l8192_id3_4_1_wenable) );
  ram_w4_l8192_id3_5 inst_ram_w4_l8192_id3_5 ( .CLK(CLK), .ram_w4_l8192_id3_5_0_addr(ram_w4_l8192_id3_5_0_addr), .ram_w4_l8192_id3_5_0_rdata(ram_w4_l8192_id3_5_0_rdata), .ram_w4_l8192_id3_5_0_wdata(4'h0), .ram_w4_l8192_id3_5_0_wenable(1'h0), .ram_w4_l8192_id3_5_1_addr(ram_w4_l8192_id3_5_1_addr), .ram_w4_l8192_id3_5_1_rdata(ram_w4_l8192_id3_5_1_rdata), .ram_w4_l8192_id3_5_1_wdata(ram_w4_l8192_id3_5_1_wdata), .ram_w4_l8192_id3_5_1_wenable(ram_w4_l8192_id3_5_1_wenable) );
  ram_w4_l8192_id3_6 inst_ram_w4_l8192_id3_6 ( .CLK(CLK), .ram_w4_l8192_id3_6_0_addr(ram_w4_l8192_id3_6_0_addr), .ram_w4_l8192_id3_6_0_rdata(ram_w4_l8192_id3_6_0_rdata), .ram_w4_l8192_id3_6_0_wdata(4'h0), .ram_w4_l8192_id3_6_0_wenable(1'h0), .ram_w4_l8192_id3_6_1_addr(ram_w4_l8192_id3_6_1_addr), .ram_w4_l8192_id3_6_1_rdata(ram_w4_l8192_id3_6_1_rdata), .ram_w4_l8192_id3_6_1_wdata(ram_w4_l8192_id3_6_1_wdata), .ram_w4_l8192_id3_6_1_wenable(ram_w4_l8192_id3_6_1_wenable) );
  ram_w4_l8192_id3_7 inst_ram_w4_l8192_id3_7 ( .CLK(CLK), .ram_w4_l8192_id3_7_0_addr(ram_w4_l8192_id3_7_0_addr), .ram_w4_l8192_id3_7_0_rdata(ram_w4_l8192_id3_7_0_rdata), .ram_w4_l8192_id3_7_0_wdata(4'h0), .ram_w4_l8192_id3_7_0_wenable(1'h0), .ram_w4_l8192_id3_7_1_addr(ram_w4_l8192_id3_7_1_addr), .ram_w4_l8192_id3_7_1_rdata(ram_w4_l8192_id3_7_1_rdata), .ram_w4_l8192_id3_7_1_wdata(ram_w4_l8192_id3_7_1_wdata), .ram_w4_l8192_id3_7_1_wenable(ram_w4_l8192_id3_7_1_wenable) );
  ram_w4_l8192_id4_0 inst_ram_w4_l8192_id4_0 ( .CLK(CLK), .ram_w4_l8192_id4_0_0_addr(ram_w4_l8192_id4_0_0_addr), .ram_w4_l8192_id4_0_0_rdata(ram_w4_l8192_id4_0_0_rdata), .ram_w4_l8192_id4_0_0_wdata(4'h0), .ram_w4_l8192_id4_0_0_wenable(1'h0), .ram_w4_l8192_id4_0_1_addr(ram_w4_l8192_id4_0_1_addr), .ram_w4_l8192_id4_0_1_rdata(ram_w4_l8192_id4_0_1_rdata), .ram_w4_l8192_id4_0_1_wdata(ram_w4_l8192_id4_0_1_wdata), .ram_w4_l8192_id4_0_1_wenable(ram_w4_l8192_id4_0_1_wenable) );
  ram_w4_l8192_id4_1 inst_ram_w4_l8192_id4_1 ( .CLK(CLK), .ram_w4_l8192_id4_1_0_addr(ram_w4_l8192_id4_1_0_addr), .ram_w4_l8192_id4_1_0_rdata(ram_w4_l8192_id4_1_0_rdata), .ram_w4_l8192_id4_1_0_wdata(4'h0), .ram_w4_l8192_id4_1_0_wenable(1'h0), .ram_w4_l8192_id4_1_1_addr(ram_w4_l8192_id4_1_1_addr), .ram_w4_l8192_id4_1_1_rdata(ram_w4_l8192_id4_1_1_rdata), .ram_w4_l8192_id4_1_1_wdata(ram_w4_l8192_id4_1_1_wdata), .ram_w4_l8192_id4_1_1_wenable(ram_w4_l8192_id4_1_1_wenable) );
  ram_w4_l8192_id4_2 inst_ram_w4_l8192_id4_2 ( .CLK(CLK), .ram_w4_l8192_id4_2_0_addr(ram_w4_l8192_id4_2_0_addr), .ram_w4_l8192_id4_2_0_rdata(ram_w4_l8192_id4_2_0_rdata), .ram_w4_l8192_id4_2_0_wdata(4'h0), .ram_w4_l8192_id4_2_0_wenable(1'h0), .ram_w4_l8192_id4_2_1_addr(ram_w4_l8192_id4_2_1_addr), .ram_w4_l8192_id4_2_1_rdata(ram_w4_l8192_id4_2_1_rdata), .ram_w4_l8192_id4_2_1_wdata(ram_w4_l8192_id4_2_1_wdata), .ram_w4_l8192_id4_2_1_wenable(ram_w4_l8192_id4_2_1_wenable) );
  ram_w4_l8192_id4_3 inst_ram_w4_l8192_id4_3 ( .CLK(CLK), .ram_w4_l8192_id4_3_0_addr(ram_w4_l8192_id4_3_0_addr), .ram_w4_l8192_id4_3_0_rdata(ram_w4_l8192_id4_3_0_rdata), .ram_w4_l8192_id4_3_0_wdata(4'h0), .ram_w4_l8192_id4_3_0_wenable(1'h0), .ram_w4_l8192_id4_3_1_addr(ram_w4_l8192_id4_3_1_addr), .ram_w4_l8192_id4_3_1_rdata(ram_w4_l8192_id4_3_1_rdata), .ram_w4_l8192_id4_3_1_wdata(ram_w4_l8192_id4_3_1_wdata), .ram_w4_l8192_id4_3_1_wenable(ram_w4_l8192_id4_3_1_wenable) );
  ram_w4_l8192_id4_4 inst_ram_w4_l8192_id4_4 ( .CLK(CLK), .ram_w4_l8192_id4_4_0_addr(ram_w4_l8192_id4_4_0_addr), .ram_w4_l8192_id4_4_0_rdata(ram_w4_l8192_id4_4_0_rdata), .ram_w4_l8192_id4_4_0_wdata(4'h0), .ram_w4_l8192_id4_4_0_wenable(1'h0), .ram_w4_l8192_id4_4_1_addr(ram_w4_l8192_id4_4_1_addr), .ram_w4_l8192_id4_4_1_rdata(ram_w4_l8192_id4_4_1_rdata), .ram_w4_l8192_id4_4_1_wdata(ram_w4_l8192_id4_4_1_wdata), .ram_w4_l8192_id4_4_1_wenable(ram_w4_l8192_id4_4_1_wenable) );
  ram_w4_l8192_id4_5 inst_ram_w4_l8192_id4_5 ( .CLK(CLK), .ram_w4_l8192_id4_5_0_addr(ram_w4_l8192_id4_5_0_addr), .ram_w4_l8192_id4_5_0_rdata(ram_w4_l8192_id4_5_0_rdata), .ram_w4_l8192_id4_5_0_wdata(4'h0), .ram_w4_l8192_id4_5_0_wenable(1'h0), .ram_w4_l8192_id4_5_1_addr(ram_w4_l8192_id4_5_1_addr), .ram_w4_l8192_id4_5_1_rdata(ram_w4_l8192_id4_5_1_rdata), .ram_w4_l8192_id4_5_1_wdata(ram_w4_l8192_id4_5_1_wdata), .ram_w4_l8192_id4_5_1_wenable(ram_w4_l8192_id4_5_1_wenable) );
  ram_w4_l8192_id4_6 inst_ram_w4_l8192_id4_6 ( .CLK(CLK), .ram_w4_l8192_id4_6_0_addr(ram_w4_l8192_id4_6_0_addr), .ram_w4_l8192_id4_6_0_rdata(ram_w4_l8192_id4_6_0_rdata), .ram_w4_l8192_id4_6_0_wdata(4'h0), .ram_w4_l8192_id4_6_0_wenable(1'h0), .ram_w4_l8192_id4_6_1_addr(ram_w4_l8192_id4_6_1_addr), .ram_w4_l8192_id4_6_1_rdata(ram_w4_l8192_id4_6_1_rdata), .ram_w4_l8192_id4_6_1_wdata(ram_w4_l8192_id4_6_1_wdata), .ram_w4_l8192_id4_6_1_wenable(ram_w4_l8192_id4_6_1_wenable) );
  ram_w4_l8192_id4_7 inst_ram_w4_l8192_id4_7 ( .CLK(CLK), .ram_w4_l8192_id4_7_0_addr(ram_w4_l8192_id4_7_0_addr), .ram_w4_l8192_id4_7_0_rdata(ram_w4_l8192_id4_7_0_rdata), .ram_w4_l8192_id4_7_0_wdata(4'h0), .ram_w4_l8192_id4_7_0_wenable(1'h0), .ram_w4_l8192_id4_7_1_addr(ram_w4_l8192_id4_7_1_addr), .ram_w4_l8192_id4_7_1_rdata(ram_w4_l8192_id4_7_1_rdata), .ram_w4_l8192_id4_7_1_wdata(ram_w4_l8192_id4_7_1_wdata), .ram_w4_l8192_id4_7_1_wenable(ram_w4_l8192_id4_7_1_wenable) );
  ram_w4_l8192_id5_0 inst_ram_w4_l8192_id5_0 ( .CLK(CLK), .ram_w4_l8192_id5_0_0_addr(ram_w4_l8192_id5_0_0_addr), .ram_w4_l8192_id5_0_0_rdata(ram_w4_l8192_id5_0_0_rdata), .ram_w4_l8192_id5_0_0_wdata(4'h0), .ram_w4_l8192_id5_0_0_wenable(1'h0), .ram_w4_l8192_id5_0_1_addr(ram_w4_l8192_id5_0_1_addr), .ram_w4_l8192_id5_0_1_rdata(ram_w4_l8192_id5_0_1_rdata), .ram_w4_l8192_id5_0_1_wdata(ram_w4_l8192_id5_0_1_wdata), .ram_w4_l8192_id5_0_1_wenable(ram_w4_l8192_id5_0_1_wenable) );
  ram_w4_l8192_id5_1 inst_ram_w4_l8192_id5_1 ( .CLK(CLK), .ram_w4_l8192_id5_1_0_addr(ram_w4_l8192_id5_1_0_addr), .ram_w4_l8192_id5_1_0_rdata(ram_w4_l8192_id5_1_0_rdata), .ram_w4_l8192_id5_1_0_wdata(4'h0), .ram_w4_l8192_id5_1_0_wenable(1'h0), .ram_w4_l8192_id5_1_1_addr(ram_w4_l8192_id5_1_1_addr), .ram_w4_l8192_id5_1_1_rdata(ram_w4_l8192_id5_1_1_rdata), .ram_w4_l8192_id5_1_1_wdata(ram_w4_l8192_id5_1_1_wdata), .ram_w4_l8192_id5_1_1_wenable(ram_w4_l8192_id5_1_1_wenable) );
  ram_w4_l8192_id5_2 inst_ram_w4_l8192_id5_2 ( .CLK(CLK), .ram_w4_l8192_id5_2_0_addr(ram_w4_l8192_id5_2_0_addr), .ram_w4_l8192_id5_2_0_rdata(ram_w4_l8192_id5_2_0_rdata), .ram_w4_l8192_id5_2_0_wdata(4'h0), .ram_w4_l8192_id5_2_0_wenable(1'h0), .ram_w4_l8192_id5_2_1_addr(ram_w4_l8192_id5_2_1_addr), .ram_w4_l8192_id5_2_1_rdata(ram_w4_l8192_id5_2_1_rdata), .ram_w4_l8192_id5_2_1_wdata(ram_w4_l8192_id5_2_1_wdata), .ram_w4_l8192_id5_2_1_wenable(ram_w4_l8192_id5_2_1_wenable) );
  ram_w4_l8192_id5_3 inst_ram_w4_l8192_id5_3 ( .CLK(CLK), .ram_w4_l8192_id5_3_0_addr(ram_w4_l8192_id5_3_0_addr), .ram_w4_l8192_id5_3_0_rdata(ram_w4_l8192_id5_3_0_rdata), .ram_w4_l8192_id5_3_0_wdata(4'h0), .ram_w4_l8192_id5_3_0_wenable(1'h0), .ram_w4_l8192_id5_3_1_addr(ram_w4_l8192_id5_3_1_addr), .ram_w4_l8192_id5_3_1_rdata(ram_w4_l8192_id5_3_1_rdata), .ram_w4_l8192_id5_3_1_wdata(ram_w4_l8192_id5_3_1_wdata), .ram_w4_l8192_id5_3_1_wenable(ram_w4_l8192_id5_3_1_wenable) );
  ram_w4_l8192_id5_4 inst_ram_w4_l8192_id5_4 ( .CLK(CLK), .ram_w4_l8192_id5_4_0_addr(ram_w4_l8192_id5_4_0_addr), .ram_w4_l8192_id5_4_0_rdata(ram_w4_l8192_id5_4_0_rdata), .ram_w4_l8192_id5_4_0_wdata(4'h0), .ram_w4_l8192_id5_4_0_wenable(1'h0), .ram_w4_l8192_id5_4_1_addr(ram_w4_l8192_id5_4_1_addr), .ram_w4_l8192_id5_4_1_rdata(ram_w4_l8192_id5_4_1_rdata), .ram_w4_l8192_id5_4_1_wdata(ram_w4_l8192_id5_4_1_wdata), .ram_w4_l8192_id5_4_1_wenable(ram_w4_l8192_id5_4_1_wenable) );
  ram_w4_l8192_id5_5 inst_ram_w4_l8192_id5_5 ( .CLK(CLK), .ram_w4_l8192_id5_5_0_addr(ram_w4_l8192_id5_5_0_addr), .ram_w4_l8192_id5_5_0_rdata(ram_w4_l8192_id5_5_0_rdata), .ram_w4_l8192_id5_5_0_wdata(4'h0), .ram_w4_l8192_id5_5_0_wenable(1'h0), .ram_w4_l8192_id5_5_1_addr(ram_w4_l8192_id5_5_1_addr), .ram_w4_l8192_id5_5_1_rdata(ram_w4_l8192_id5_5_1_rdata), .ram_w4_l8192_id5_5_1_wdata(ram_w4_l8192_id5_5_1_wdata), .ram_w4_l8192_id5_5_1_wenable(ram_w4_l8192_id5_5_1_wenable) );
  ram_w4_l8192_id5_6 inst_ram_w4_l8192_id5_6 ( .CLK(CLK), .ram_w4_l8192_id5_6_0_addr(ram_w4_l8192_id5_6_0_addr), .ram_w4_l8192_id5_6_0_rdata(ram_w4_l8192_id5_6_0_rdata), .ram_w4_l8192_id5_6_0_wdata(4'h0), .ram_w4_l8192_id5_6_0_wenable(1'h0), .ram_w4_l8192_id5_6_1_addr(ram_w4_l8192_id5_6_1_addr), .ram_w4_l8192_id5_6_1_rdata(ram_w4_l8192_id5_6_1_rdata), .ram_w4_l8192_id5_6_1_wdata(ram_w4_l8192_id5_6_1_wdata), .ram_w4_l8192_id5_6_1_wenable(ram_w4_l8192_id5_6_1_wenable) );
  ram_w4_l8192_id5_7 inst_ram_w4_l8192_id5_7 ( .CLK(CLK), .ram_w4_l8192_id5_7_0_addr(ram_w4_l8192_id5_7_0_addr), .ram_w4_l8192_id5_7_0_rdata(ram_w4_l8192_id5_7_0_rdata), .ram_w4_l8192_id5_7_0_wdata(4'h0), .ram_w4_l8192_id5_7_0_wenable(1'h0), .ram_w4_l8192_id5_7_1_addr(ram_w4_l8192_id5_7_1_addr), .ram_w4_l8192_id5_7_1_rdata(ram_w4_l8192_id5_7_1_rdata), .ram_w4_l8192_id5_7_1_wdata(ram_w4_l8192_id5_7_1_wdata), .ram_w4_l8192_id5_7_1_wenable(ram_w4_l8192_id5_7_1_wenable) );
  ram_w4_l8192_id6_0 inst_ram_w4_l8192_id6_0 ( .CLK(CLK), .ram_w4_l8192_id6_0_0_addr(ram_w4_l8192_id6_0_0_addr), .ram_w4_l8192_id6_0_0_rdata(ram_w4_l8192_id6_0_0_rdata), .ram_w4_l8192_id6_0_0_wdata(4'h0), .ram_w4_l8192_id6_0_0_wenable(1'h0), .ram_w4_l8192_id6_0_1_addr(ram_w4_l8192_id6_0_1_addr), .ram_w4_l8192_id6_0_1_rdata(ram_w4_l8192_id6_0_1_rdata), .ram_w4_l8192_id6_0_1_wdata(ram_w4_l8192_id6_0_1_wdata), .ram_w4_l8192_id6_0_1_wenable(ram_w4_l8192_id6_0_1_wenable) );
  ram_w4_l8192_id6_1 inst_ram_w4_l8192_id6_1 ( .CLK(CLK), .ram_w4_l8192_id6_1_0_addr(ram_w4_l8192_id6_1_0_addr), .ram_w4_l8192_id6_1_0_rdata(ram_w4_l8192_id6_1_0_rdata), .ram_w4_l8192_id6_1_0_wdata(4'h0), .ram_w4_l8192_id6_1_0_wenable(1'h0), .ram_w4_l8192_id6_1_1_addr(ram_w4_l8192_id6_1_1_addr), .ram_w4_l8192_id6_1_1_rdata(ram_w4_l8192_id6_1_1_rdata), .ram_w4_l8192_id6_1_1_wdata(ram_w4_l8192_id6_1_1_wdata), .ram_w4_l8192_id6_1_1_wenable(ram_w4_l8192_id6_1_1_wenable) );
  ram_w4_l8192_id6_2 inst_ram_w4_l8192_id6_2 ( .CLK(CLK), .ram_w4_l8192_id6_2_0_addr(ram_w4_l8192_id6_2_0_addr), .ram_w4_l8192_id6_2_0_rdata(ram_w4_l8192_id6_2_0_rdata), .ram_w4_l8192_id6_2_0_wdata(4'h0), .ram_w4_l8192_id6_2_0_wenable(1'h0), .ram_w4_l8192_id6_2_1_addr(ram_w4_l8192_id6_2_1_addr), .ram_w4_l8192_id6_2_1_rdata(ram_w4_l8192_id6_2_1_rdata), .ram_w4_l8192_id6_2_1_wdata(ram_w4_l8192_id6_2_1_wdata), .ram_w4_l8192_id6_2_1_wenable(ram_w4_l8192_id6_2_1_wenable) );
  ram_w4_l8192_id6_3 inst_ram_w4_l8192_id6_3 ( .CLK(CLK), .ram_w4_l8192_id6_3_0_addr(ram_w4_l8192_id6_3_0_addr), .ram_w4_l8192_id6_3_0_rdata(ram_w4_l8192_id6_3_0_rdata), .ram_w4_l8192_id6_3_0_wdata(4'h0), .ram_w4_l8192_id6_3_0_wenable(1'h0), .ram_w4_l8192_id6_3_1_addr(ram_w4_l8192_id6_3_1_addr), .ram_w4_l8192_id6_3_1_rdata(ram_w4_l8192_id6_3_1_rdata), .ram_w4_l8192_id6_3_1_wdata(ram_w4_l8192_id6_3_1_wdata), .ram_w4_l8192_id6_3_1_wenable(ram_w4_l8192_id6_3_1_wenable) );
  ram_w4_l8192_id6_4 inst_ram_w4_l8192_id6_4 ( .CLK(CLK), .ram_w4_l8192_id6_4_0_addr(ram_w4_l8192_id6_4_0_addr), .ram_w4_l8192_id6_4_0_rdata(ram_w4_l8192_id6_4_0_rdata), .ram_w4_l8192_id6_4_0_wdata(4'h0), .ram_w4_l8192_id6_4_0_wenable(1'h0), .ram_w4_l8192_id6_4_1_addr(ram_w4_l8192_id6_4_1_addr), .ram_w4_l8192_id6_4_1_rdata(ram_w4_l8192_id6_4_1_rdata), .ram_w4_l8192_id6_4_1_wdata(ram_w4_l8192_id6_4_1_wdata), .ram_w4_l8192_id6_4_1_wenable(ram_w4_l8192_id6_4_1_wenable) );
  ram_w4_l8192_id6_5 inst_ram_w4_l8192_id6_5 ( .CLK(CLK), .ram_w4_l8192_id6_5_0_addr(ram_w4_l8192_id6_5_0_addr), .ram_w4_l8192_id6_5_0_rdata(ram_w4_l8192_id6_5_0_rdata), .ram_w4_l8192_id6_5_0_wdata(4'h0), .ram_w4_l8192_id6_5_0_wenable(1'h0), .ram_w4_l8192_id6_5_1_addr(ram_w4_l8192_id6_5_1_addr), .ram_w4_l8192_id6_5_1_rdata(ram_w4_l8192_id6_5_1_rdata), .ram_w4_l8192_id6_5_1_wdata(ram_w4_l8192_id6_5_1_wdata), .ram_w4_l8192_id6_5_1_wenable(ram_w4_l8192_id6_5_1_wenable) );
  ram_w4_l8192_id6_6 inst_ram_w4_l8192_id6_6 ( .CLK(CLK), .ram_w4_l8192_id6_6_0_addr(ram_w4_l8192_id6_6_0_addr), .ram_w4_l8192_id6_6_0_rdata(ram_w4_l8192_id6_6_0_rdata), .ram_w4_l8192_id6_6_0_wdata(4'h0), .ram_w4_l8192_id6_6_0_wenable(1'h0), .ram_w4_l8192_id6_6_1_addr(ram_w4_l8192_id6_6_1_addr), .ram_w4_l8192_id6_6_1_rdata(ram_w4_l8192_id6_6_1_rdata), .ram_w4_l8192_id6_6_1_wdata(ram_w4_l8192_id6_6_1_wdata), .ram_w4_l8192_id6_6_1_wenable(ram_w4_l8192_id6_6_1_wenable) );
  ram_w4_l8192_id6_7 inst_ram_w4_l8192_id6_7 ( .CLK(CLK), .ram_w4_l8192_id6_7_0_addr(ram_w4_l8192_id6_7_0_addr), .ram_w4_l8192_id6_7_0_rdata(ram_w4_l8192_id6_7_0_rdata), .ram_w4_l8192_id6_7_0_wdata(4'h0), .ram_w4_l8192_id6_7_0_wenable(1'h0), .ram_w4_l8192_id6_7_1_addr(ram_w4_l8192_id6_7_1_addr), .ram_w4_l8192_id6_7_1_rdata(ram_w4_l8192_id6_7_1_rdata), .ram_w4_l8192_id6_7_1_wdata(ram_w4_l8192_id6_7_1_wdata), .ram_w4_l8192_id6_7_1_wenable(ram_w4_l8192_id6_7_1_wenable) );
  ram_w4_l8192_id7_0 inst_ram_w4_l8192_id7_0 ( .CLK(CLK), .ram_w4_l8192_id7_0_0_addr(ram_w4_l8192_id7_0_0_addr), .ram_w4_l8192_id7_0_0_rdata(ram_w4_l8192_id7_0_0_rdata), .ram_w4_l8192_id7_0_0_wdata(4'h0), .ram_w4_l8192_id7_0_0_wenable(1'h0), .ram_w4_l8192_id7_0_1_addr(ram_w4_l8192_id7_0_1_addr), .ram_w4_l8192_id7_0_1_rdata(ram_w4_l8192_id7_0_1_rdata), .ram_w4_l8192_id7_0_1_wdata(ram_w4_l8192_id7_0_1_wdata), .ram_w4_l8192_id7_0_1_wenable(ram_w4_l8192_id7_0_1_wenable) );
  ram_w4_l8192_id7_1 inst_ram_w4_l8192_id7_1 ( .CLK(CLK), .ram_w4_l8192_id7_1_0_addr(ram_w4_l8192_id7_1_0_addr), .ram_w4_l8192_id7_1_0_rdata(ram_w4_l8192_id7_1_0_rdata), .ram_w4_l8192_id7_1_0_wdata(4'h0), .ram_w4_l8192_id7_1_0_wenable(1'h0), .ram_w4_l8192_id7_1_1_addr(ram_w4_l8192_id7_1_1_addr), .ram_w4_l8192_id7_1_1_rdata(ram_w4_l8192_id7_1_1_rdata), .ram_w4_l8192_id7_1_1_wdata(ram_w4_l8192_id7_1_1_wdata), .ram_w4_l8192_id7_1_1_wenable(ram_w4_l8192_id7_1_1_wenable) );
  ram_w4_l8192_id7_2 inst_ram_w4_l8192_id7_2 ( .CLK(CLK), .ram_w4_l8192_id7_2_0_addr(ram_w4_l8192_id7_2_0_addr), .ram_w4_l8192_id7_2_0_rdata(ram_w4_l8192_id7_2_0_rdata), .ram_w4_l8192_id7_2_0_wdata(4'h0), .ram_w4_l8192_id7_2_0_wenable(1'h0), .ram_w4_l8192_id7_2_1_addr(ram_w4_l8192_id7_2_1_addr), .ram_w4_l8192_id7_2_1_rdata(ram_w4_l8192_id7_2_1_rdata), .ram_w4_l8192_id7_2_1_wdata(ram_w4_l8192_id7_2_1_wdata), .ram_w4_l8192_id7_2_1_wenable(ram_w4_l8192_id7_2_1_wenable) );
  ram_w4_l8192_id7_3 inst_ram_w4_l8192_id7_3 ( .CLK(CLK), .ram_w4_l8192_id7_3_0_addr(ram_w4_l8192_id7_3_0_addr), .ram_w4_l8192_id7_3_0_rdata(ram_w4_l8192_id7_3_0_rdata), .ram_w4_l8192_id7_3_0_wdata(4'h0), .ram_w4_l8192_id7_3_0_wenable(1'h0), .ram_w4_l8192_id7_3_1_addr(ram_w4_l8192_id7_3_1_addr), .ram_w4_l8192_id7_3_1_rdata(ram_w4_l8192_id7_3_1_rdata), .ram_w4_l8192_id7_3_1_wdata(ram_w4_l8192_id7_3_1_wdata), .ram_w4_l8192_id7_3_1_wenable(ram_w4_l8192_id7_3_1_wenable) );
  ram_w4_l8192_id7_4 inst_ram_w4_l8192_id7_4 ( .CLK(CLK), .ram_w4_l8192_id7_4_0_addr(ram_w4_l8192_id7_4_0_addr), .ram_w4_l8192_id7_4_0_rdata(ram_w4_l8192_id7_4_0_rdata), .ram_w4_l8192_id7_4_0_wdata(4'h0), .ram_w4_l8192_id7_4_0_wenable(1'h0), .ram_w4_l8192_id7_4_1_addr(ram_w4_l8192_id7_4_1_addr), .ram_w4_l8192_id7_4_1_rdata(ram_w4_l8192_id7_4_1_rdata), .ram_w4_l8192_id7_4_1_wdata(ram_w4_l8192_id7_4_1_wdata), .ram_w4_l8192_id7_4_1_wenable(ram_w4_l8192_id7_4_1_wenable) );
  ram_w4_l8192_id7_5 inst_ram_w4_l8192_id7_5 ( .CLK(CLK), .ram_w4_l8192_id7_5_0_addr(ram_w4_l8192_id7_5_0_addr), .ram_w4_l8192_id7_5_0_rdata(ram_w4_l8192_id7_5_0_rdata), .ram_w4_l8192_id7_5_0_wdata(4'h0), .ram_w4_l8192_id7_5_0_wenable(1'h0), .ram_w4_l8192_id7_5_1_addr(ram_w4_l8192_id7_5_1_addr), .ram_w4_l8192_id7_5_1_rdata(ram_w4_l8192_id7_5_1_rdata), .ram_w4_l8192_id7_5_1_wdata(ram_w4_l8192_id7_5_1_wdata), .ram_w4_l8192_id7_5_1_wenable(ram_w4_l8192_id7_5_1_wenable) );
  ram_w4_l8192_id7_6 inst_ram_w4_l8192_id7_6 ( .CLK(CLK), .ram_w4_l8192_id7_6_0_addr(ram_w4_l8192_id7_6_0_addr), .ram_w4_l8192_id7_6_0_rdata(ram_w4_l8192_id7_6_0_rdata), .ram_w4_l8192_id7_6_0_wdata(4'h0), .ram_w4_l8192_id7_6_0_wenable(1'h0), .ram_w4_l8192_id7_6_1_addr(ram_w4_l8192_id7_6_1_addr), .ram_w4_l8192_id7_6_1_rdata(ram_w4_l8192_id7_6_1_rdata), .ram_w4_l8192_id7_6_1_wdata(ram_w4_l8192_id7_6_1_wdata), .ram_w4_l8192_id7_6_1_wenable(ram_w4_l8192_id7_6_1_wenable) );
  ram_w4_l8192_id7_7 inst_ram_w4_l8192_id7_7 ( .CLK(CLK), .ram_w4_l8192_id7_7_0_addr(ram_w4_l8192_id7_7_0_addr), .ram_w4_l8192_id7_7_0_rdata(ram_w4_l8192_id7_7_0_rdata), .ram_w4_l8192_id7_7_0_wdata(4'h0), .ram_w4_l8192_id7_7_0_wenable(1'h0), .ram_w4_l8192_id7_7_1_addr(ram_w4_l8192_id7_7_1_addr), .ram_w4_l8192_id7_7_1_rdata(ram_w4_l8192_id7_7_1_rdata), .ram_w4_l8192_id7_7_1_wdata(ram_w4_l8192_id7_7_1_wdata), .ram_w4_l8192_id7_7_1_wenable(ram_w4_l8192_id7_7_1_wenable) );
  ram_w4_l8192_id8_0 inst_ram_w4_l8192_id8_0 ( .CLK(CLK), .ram_w4_l8192_id8_0_0_addr(ram_w4_l8192_id8_0_0_addr), .ram_w4_l8192_id8_0_0_rdata(ram_w4_l8192_id8_0_0_rdata), .ram_w4_l8192_id8_0_0_wdata(4'h0), .ram_w4_l8192_id8_0_0_wenable(1'h0), .ram_w4_l8192_id8_0_1_addr(ram_w4_l8192_id8_0_1_addr), .ram_w4_l8192_id8_0_1_rdata(ram_w4_l8192_id8_0_1_rdata), .ram_w4_l8192_id8_0_1_wdata(ram_w4_l8192_id8_0_1_wdata), .ram_w4_l8192_id8_0_1_wenable(ram_w4_l8192_id8_0_1_wenable) );
  ram_w4_l8192_id8_1 inst_ram_w4_l8192_id8_1 ( .CLK(CLK), .ram_w4_l8192_id8_1_0_addr(ram_w4_l8192_id8_1_0_addr), .ram_w4_l8192_id8_1_0_rdata(ram_w4_l8192_id8_1_0_rdata), .ram_w4_l8192_id8_1_0_wdata(4'h0), .ram_w4_l8192_id8_1_0_wenable(1'h0), .ram_w4_l8192_id8_1_1_addr(ram_w4_l8192_id8_1_1_addr), .ram_w4_l8192_id8_1_1_rdata(ram_w4_l8192_id8_1_1_rdata), .ram_w4_l8192_id8_1_1_wdata(ram_w4_l8192_id8_1_1_wdata), .ram_w4_l8192_id8_1_1_wenable(ram_w4_l8192_id8_1_1_wenable) );
  ram_w4_l8192_id8_2 inst_ram_w4_l8192_id8_2 ( .CLK(CLK), .ram_w4_l8192_id8_2_0_addr(ram_w4_l8192_id8_2_0_addr), .ram_w4_l8192_id8_2_0_rdata(ram_w4_l8192_id8_2_0_rdata), .ram_w4_l8192_id8_2_0_wdata(4'h0), .ram_w4_l8192_id8_2_0_wenable(1'h0), .ram_w4_l8192_id8_2_1_addr(ram_w4_l8192_id8_2_1_addr), .ram_w4_l8192_id8_2_1_rdata(ram_w4_l8192_id8_2_1_rdata), .ram_w4_l8192_id8_2_1_wdata(ram_w4_l8192_id8_2_1_wdata), .ram_w4_l8192_id8_2_1_wenable(ram_w4_l8192_id8_2_1_wenable) );
  ram_w4_l8192_id8_3 inst_ram_w4_l8192_id8_3 ( .CLK(CLK), .ram_w4_l8192_id8_3_0_addr(ram_w4_l8192_id8_3_0_addr), .ram_w4_l8192_id8_3_0_rdata(ram_w4_l8192_id8_3_0_rdata), .ram_w4_l8192_id8_3_0_wdata(4'h0), .ram_w4_l8192_id8_3_0_wenable(1'h0), .ram_w4_l8192_id8_3_1_addr(ram_w4_l8192_id8_3_1_addr), .ram_w4_l8192_id8_3_1_rdata(ram_w4_l8192_id8_3_1_rdata), .ram_w4_l8192_id8_3_1_wdata(ram_w4_l8192_id8_3_1_wdata), .ram_w4_l8192_id8_3_1_wenable(ram_w4_l8192_id8_3_1_wenable) );
  ram_w4_l8192_id8_4 inst_ram_w4_l8192_id8_4 ( .CLK(CLK), .ram_w4_l8192_id8_4_0_addr(ram_w4_l8192_id8_4_0_addr), .ram_w4_l8192_id8_4_0_rdata(ram_w4_l8192_id8_4_0_rdata), .ram_w4_l8192_id8_4_0_wdata(4'h0), .ram_w4_l8192_id8_4_0_wenable(1'h0), .ram_w4_l8192_id8_4_1_addr(ram_w4_l8192_id8_4_1_addr), .ram_w4_l8192_id8_4_1_rdata(ram_w4_l8192_id8_4_1_rdata), .ram_w4_l8192_id8_4_1_wdata(ram_w4_l8192_id8_4_1_wdata), .ram_w4_l8192_id8_4_1_wenable(ram_w4_l8192_id8_4_1_wenable) );
  ram_w4_l8192_id8_5 inst_ram_w4_l8192_id8_5 ( .CLK(CLK), .ram_w4_l8192_id8_5_0_addr(ram_w4_l8192_id8_5_0_addr), .ram_w4_l8192_id8_5_0_rdata(ram_w4_l8192_id8_5_0_rdata), .ram_w4_l8192_id8_5_0_wdata(4'h0), .ram_w4_l8192_id8_5_0_wenable(1'h0), .ram_w4_l8192_id8_5_1_addr(ram_w4_l8192_id8_5_1_addr), .ram_w4_l8192_id8_5_1_rdata(ram_w4_l8192_id8_5_1_rdata), .ram_w4_l8192_id8_5_1_wdata(ram_w4_l8192_id8_5_1_wdata), .ram_w4_l8192_id8_5_1_wenable(ram_w4_l8192_id8_5_1_wenable) );
  ram_w4_l8192_id8_6 inst_ram_w4_l8192_id8_6 ( .CLK(CLK), .ram_w4_l8192_id8_6_0_addr(ram_w4_l8192_id8_6_0_addr), .ram_w4_l8192_id8_6_0_rdata(ram_w4_l8192_id8_6_0_rdata), .ram_w4_l8192_id8_6_0_wdata(4'h0), .ram_w4_l8192_id8_6_0_wenable(1'h0), .ram_w4_l8192_id8_6_1_addr(ram_w4_l8192_id8_6_1_addr), .ram_w4_l8192_id8_6_1_rdata(ram_w4_l8192_id8_6_1_rdata), .ram_w4_l8192_id8_6_1_wdata(ram_w4_l8192_id8_6_1_wdata), .ram_w4_l8192_id8_6_1_wenable(ram_w4_l8192_id8_6_1_wenable) );
  ram_w4_l8192_id8_7 inst_ram_w4_l8192_id8_7 ( .CLK(CLK), .ram_w4_l8192_id8_7_0_addr(ram_w4_l8192_id8_7_0_addr), .ram_w4_l8192_id8_7_0_rdata(ram_w4_l8192_id8_7_0_rdata), .ram_w4_l8192_id8_7_0_wdata(4'h0), .ram_w4_l8192_id8_7_0_wenable(1'h0), .ram_w4_l8192_id8_7_1_addr(ram_w4_l8192_id8_7_1_addr), .ram_w4_l8192_id8_7_1_rdata(ram_w4_l8192_id8_7_1_rdata), .ram_w4_l8192_id8_7_1_wdata(ram_w4_l8192_id8_7_1_wdata), .ram_w4_l8192_id8_7_1_wenable(ram_w4_l8192_id8_7_1_wenable) );
  ram_w8_l2048_id0_0 inst_ram_w8_l2048_id0_0 ( .CLK(CLK), .ram_w8_l2048_id0_0_0_addr(ram_w8_l2048_id0_0_0_addr), .ram_w8_l2048_id0_0_0_rdata(ram_w8_l2048_id0_0_0_rdata), .ram_w8_l2048_id0_0_0_wdata(ram_w8_l2048_id0_0_0_wdata), .ram_w8_l2048_id0_0_0_wenable(ram_w8_l2048_id0_0_0_wenable), .ram_w8_l2048_id0_0_1_addr(ram_w8_l2048_id0_0_1_addr), .ram_w8_l2048_id0_0_1_rdata(ram_w8_l2048_id0_0_1_rdata), .ram_w8_l2048_id0_0_1_wdata(ram_w8_l2048_id0_0_1_wdata), .ram_w8_l2048_id0_0_1_wenable(ram_w8_l2048_id0_0_1_wenable) );
  ram_w8_l2048_id0_1 inst_ram_w8_l2048_id0_1 ( .CLK(CLK), .ram_w8_l2048_id0_1_0_addr(ram_w8_l2048_id0_1_0_addr), .ram_w8_l2048_id0_1_0_rdata(ram_w8_l2048_id0_1_0_rdata), .ram_w8_l2048_id0_1_0_wdata(ram_w8_l2048_id0_1_0_wdata), .ram_w8_l2048_id0_1_0_wenable(ram_w8_l2048_id0_1_0_wenable), .ram_w8_l2048_id0_1_1_addr(ram_w8_l2048_id0_1_1_addr), .ram_w8_l2048_id0_1_1_rdata(ram_w8_l2048_id0_1_1_rdata), .ram_w8_l2048_id0_1_1_wdata(ram_w8_l2048_id0_1_1_wdata), .ram_w8_l2048_id0_1_1_wenable(ram_w8_l2048_id0_1_1_wenable) );
  ram_w8_l2048_id0_2 inst_ram_w8_l2048_id0_2 ( .CLK(CLK), .ram_w8_l2048_id0_2_0_addr(ram_w8_l2048_id0_2_0_addr), .ram_w8_l2048_id0_2_0_rdata(ram_w8_l2048_id0_2_0_rdata), .ram_w8_l2048_id0_2_0_wdata(ram_w8_l2048_id0_2_0_wdata), .ram_w8_l2048_id0_2_0_wenable(ram_w8_l2048_id0_2_0_wenable), .ram_w8_l2048_id0_2_1_addr(ram_w8_l2048_id0_2_1_addr), .ram_w8_l2048_id0_2_1_rdata(ram_w8_l2048_id0_2_1_rdata), .ram_w8_l2048_id0_2_1_wdata(ram_w8_l2048_id0_2_1_wdata), .ram_w8_l2048_id0_2_1_wenable(ram_w8_l2048_id0_2_1_wenable) );
  ram_w8_l2048_id0_3 inst_ram_w8_l2048_id0_3 ( .CLK(CLK), .ram_w8_l2048_id0_3_0_addr(ram_w8_l2048_id0_3_0_addr), .ram_w8_l2048_id0_3_0_rdata(ram_w8_l2048_id0_3_0_rdata), .ram_w8_l2048_id0_3_0_wdata(ram_w8_l2048_id0_3_0_wdata), .ram_w8_l2048_id0_3_0_wenable(ram_w8_l2048_id0_3_0_wenable), .ram_w8_l2048_id0_3_1_addr(ram_w8_l2048_id0_3_1_addr), .ram_w8_l2048_id0_3_1_rdata(ram_w8_l2048_id0_3_1_rdata), .ram_w8_l2048_id0_3_1_wdata(ram_w8_l2048_id0_3_1_wdata), .ram_w8_l2048_id0_3_1_wenable(ram_w8_l2048_id0_3_1_wenable) );
  ram_w8_l2048_id10_0 inst_ram_w8_l2048_id10_0 ( .CLK(CLK), .ram_w8_l2048_id10_0_0_addr(ram_w8_l2048_id10_0_0_addr), .ram_w8_l2048_id10_0_0_rdata(ram_w8_l2048_id10_0_0_rdata), .ram_w8_l2048_id10_0_0_wdata(8'h00), .ram_w8_l2048_id10_0_0_wenable(1'h0), .ram_w8_l2048_id10_0_1_addr(ram_w8_l2048_id10_0_1_addr), .ram_w8_l2048_id10_0_1_rdata(ram_w8_l2048_id10_0_1_rdata), .ram_w8_l2048_id10_0_1_wdata(ram_w8_l2048_id10_0_1_wdata), .ram_w8_l2048_id10_0_1_wenable(ram_w8_l2048_id10_0_1_wenable) );
  ram_w8_l2048_id10_1 inst_ram_w8_l2048_id10_1 ( .CLK(CLK), .ram_w8_l2048_id10_1_0_addr(ram_w8_l2048_id10_1_0_addr), .ram_w8_l2048_id10_1_0_rdata(ram_w8_l2048_id10_1_0_rdata), .ram_w8_l2048_id10_1_0_wdata(8'h00), .ram_w8_l2048_id10_1_0_wenable(1'h0), .ram_w8_l2048_id10_1_1_addr(ram_w8_l2048_id10_1_1_addr), .ram_w8_l2048_id10_1_1_rdata(ram_w8_l2048_id10_1_1_rdata), .ram_w8_l2048_id10_1_1_wdata(ram_w8_l2048_id10_1_1_wdata), .ram_w8_l2048_id10_1_1_wenable(ram_w8_l2048_id10_1_1_wenable) );
  ram_w8_l2048_id10_2 inst_ram_w8_l2048_id10_2 ( .CLK(CLK), .ram_w8_l2048_id10_2_0_addr(ram_w8_l2048_id10_2_0_addr), .ram_w8_l2048_id10_2_0_rdata(ram_w8_l2048_id10_2_0_rdata), .ram_w8_l2048_id10_2_0_wdata(8'h00), .ram_w8_l2048_id10_2_0_wenable(1'h0), .ram_w8_l2048_id10_2_1_addr(ram_w8_l2048_id10_2_1_addr), .ram_w8_l2048_id10_2_1_rdata(ram_w8_l2048_id10_2_1_rdata), .ram_w8_l2048_id10_2_1_wdata(ram_w8_l2048_id10_2_1_wdata), .ram_w8_l2048_id10_2_1_wenable(ram_w8_l2048_id10_2_1_wenable) );
  ram_w8_l2048_id10_3 inst_ram_w8_l2048_id10_3 ( .CLK(CLK), .ram_w8_l2048_id10_3_0_addr(ram_w8_l2048_id10_3_0_addr), .ram_w8_l2048_id10_3_0_rdata(ram_w8_l2048_id10_3_0_rdata), .ram_w8_l2048_id10_3_0_wdata(8'h00), .ram_w8_l2048_id10_3_0_wenable(1'h0), .ram_w8_l2048_id10_3_1_addr(ram_w8_l2048_id10_3_1_addr), .ram_w8_l2048_id10_3_1_rdata(ram_w8_l2048_id10_3_1_rdata), .ram_w8_l2048_id10_3_1_wdata(ram_w8_l2048_id10_3_1_wdata), .ram_w8_l2048_id10_3_1_wenable(ram_w8_l2048_id10_3_1_wenable) );
  ram_w8_l2048_id11_0 inst_ram_w8_l2048_id11_0 ( .CLK(CLK), .ram_w8_l2048_id11_0_0_addr(ram_w8_l2048_id11_0_0_addr), .ram_w8_l2048_id11_0_0_rdata(ram_w8_l2048_id11_0_0_rdata), .ram_w8_l2048_id11_0_0_wdata(ram_w8_l2048_id11_0_0_wdata), .ram_w8_l2048_id11_0_0_wenable(ram_w8_l2048_id11_0_0_wenable), .ram_w8_l2048_id11_0_1_addr(ram_w8_l2048_id11_0_1_addr), .ram_w8_l2048_id11_0_1_rdata(ram_w8_l2048_id11_0_1_rdata), .ram_w8_l2048_id11_0_1_wdata(8'h00), .ram_w8_l2048_id11_0_1_wenable(1'h0) );
  ram_w8_l2048_id11_1 inst_ram_w8_l2048_id11_1 ( .CLK(CLK), .ram_w8_l2048_id11_1_0_addr(ram_w8_l2048_id11_1_0_addr), .ram_w8_l2048_id11_1_0_rdata(ram_w8_l2048_id11_1_0_rdata), .ram_w8_l2048_id11_1_0_wdata(ram_w8_l2048_id11_1_0_wdata), .ram_w8_l2048_id11_1_0_wenable(ram_w8_l2048_id11_1_0_wenable), .ram_w8_l2048_id11_1_1_addr(ram_w8_l2048_id11_1_1_addr), .ram_w8_l2048_id11_1_1_rdata(ram_w8_l2048_id11_1_1_rdata), .ram_w8_l2048_id11_1_1_wdata(8'h00), .ram_w8_l2048_id11_1_1_wenable(1'h0) );
  ram_w8_l2048_id11_2 inst_ram_w8_l2048_id11_2 ( .CLK(CLK), .ram_w8_l2048_id11_2_0_addr(ram_w8_l2048_id11_2_0_addr), .ram_w8_l2048_id11_2_0_rdata(ram_w8_l2048_id11_2_0_rdata), .ram_w8_l2048_id11_2_0_wdata(ram_w8_l2048_id11_2_0_wdata), .ram_w8_l2048_id11_2_0_wenable(ram_w8_l2048_id11_2_0_wenable), .ram_w8_l2048_id11_2_1_addr(ram_w8_l2048_id11_2_1_addr), .ram_w8_l2048_id11_2_1_rdata(ram_w8_l2048_id11_2_1_rdata), .ram_w8_l2048_id11_2_1_wdata(8'h00), .ram_w8_l2048_id11_2_1_wenable(1'h0) );
  ram_w8_l2048_id11_3 inst_ram_w8_l2048_id11_3 ( .CLK(CLK), .ram_w8_l2048_id11_3_0_addr(ram_w8_l2048_id11_3_0_addr), .ram_w8_l2048_id11_3_0_rdata(ram_w8_l2048_id11_3_0_rdata), .ram_w8_l2048_id11_3_0_wdata(ram_w8_l2048_id11_3_0_wdata), .ram_w8_l2048_id11_3_0_wenable(ram_w8_l2048_id11_3_0_wenable), .ram_w8_l2048_id11_3_1_addr(ram_w8_l2048_id11_3_1_addr), .ram_w8_l2048_id11_3_1_rdata(ram_w8_l2048_id11_3_1_rdata), .ram_w8_l2048_id11_3_1_wdata(8'h00), .ram_w8_l2048_id11_3_1_wenable(1'h0) );
  ram_w8_l2048_id1_0 inst_ram_w8_l2048_id1_0 ( .CLK(CLK), .ram_w8_l2048_id1_0_0_addr(ram_w8_l2048_id1_0_0_addr), .ram_w8_l2048_id1_0_0_rdata(ram_w8_l2048_id1_0_0_rdata), .ram_w8_l2048_id1_0_0_wdata(ram_w8_l2048_id1_0_0_wdata), .ram_w8_l2048_id1_0_0_wenable(ram_w8_l2048_id1_0_0_wenable), .ram_w8_l2048_id1_0_1_addr(ram_w8_l2048_id1_0_1_addr), .ram_w8_l2048_id1_0_1_rdata(ram_w8_l2048_id1_0_1_rdata), .ram_w8_l2048_id1_0_1_wdata(ram_w8_l2048_id1_0_1_wdata), .ram_w8_l2048_id1_0_1_wenable(ram_w8_l2048_id1_0_1_wenable) );
  ram_w8_l2048_id1_1 inst_ram_w8_l2048_id1_1 ( .CLK(CLK), .ram_w8_l2048_id1_1_0_addr(ram_w8_l2048_id1_1_0_addr), .ram_w8_l2048_id1_1_0_rdata(ram_w8_l2048_id1_1_0_rdata), .ram_w8_l2048_id1_1_0_wdata(ram_w8_l2048_id1_1_0_wdata), .ram_w8_l2048_id1_1_0_wenable(ram_w8_l2048_id1_1_0_wenable), .ram_w8_l2048_id1_1_1_addr(ram_w8_l2048_id1_1_1_addr), .ram_w8_l2048_id1_1_1_rdata(ram_w8_l2048_id1_1_1_rdata), .ram_w8_l2048_id1_1_1_wdata(ram_w8_l2048_id1_1_1_wdata), .ram_w8_l2048_id1_1_1_wenable(ram_w8_l2048_id1_1_1_wenable) );
  ram_w8_l2048_id1_2 inst_ram_w8_l2048_id1_2 ( .CLK(CLK), .ram_w8_l2048_id1_2_0_addr(ram_w8_l2048_id1_2_0_addr), .ram_w8_l2048_id1_2_0_rdata(ram_w8_l2048_id1_2_0_rdata), .ram_w8_l2048_id1_2_0_wdata(ram_w8_l2048_id1_2_0_wdata), .ram_w8_l2048_id1_2_0_wenable(ram_w8_l2048_id1_2_0_wenable), .ram_w8_l2048_id1_2_1_addr(ram_w8_l2048_id1_2_1_addr), .ram_w8_l2048_id1_2_1_rdata(ram_w8_l2048_id1_2_1_rdata), .ram_w8_l2048_id1_2_1_wdata(ram_w8_l2048_id1_2_1_wdata), .ram_w8_l2048_id1_2_1_wenable(ram_w8_l2048_id1_2_1_wenable) );
  ram_w8_l2048_id1_3 inst_ram_w8_l2048_id1_3 ( .CLK(CLK), .ram_w8_l2048_id1_3_0_addr(ram_w8_l2048_id1_3_0_addr), .ram_w8_l2048_id1_3_0_rdata(ram_w8_l2048_id1_3_0_rdata), .ram_w8_l2048_id1_3_0_wdata(ram_w8_l2048_id1_3_0_wdata), .ram_w8_l2048_id1_3_0_wenable(ram_w8_l2048_id1_3_0_wenable), .ram_w8_l2048_id1_3_1_addr(ram_w8_l2048_id1_3_1_addr), .ram_w8_l2048_id1_3_1_rdata(ram_w8_l2048_id1_3_1_rdata), .ram_w8_l2048_id1_3_1_wdata(ram_w8_l2048_id1_3_1_wdata), .ram_w8_l2048_id1_3_1_wenable(ram_w8_l2048_id1_3_1_wenable) );
  ram_w8_l2048_id2_0 inst_ram_w8_l2048_id2_0 ( .CLK(CLK), .ram_w8_l2048_id2_0_0_addr(ram_w8_l2048_id2_0_0_addr), .ram_w8_l2048_id2_0_0_rdata(ram_w8_l2048_id2_0_0_rdata), .ram_w8_l2048_id2_0_0_wdata(8'h00), .ram_w8_l2048_id2_0_0_wenable(1'h0), .ram_w8_l2048_id2_0_1_addr(ram_w8_l2048_id2_0_1_addr), .ram_w8_l2048_id2_0_1_rdata(ram_w8_l2048_id2_0_1_rdata), .ram_w8_l2048_id2_0_1_wdata(ram_w8_l2048_id2_0_1_wdata), .ram_w8_l2048_id2_0_1_wenable(ram_w8_l2048_id2_0_1_wenable) );
  ram_w8_l2048_id2_1 inst_ram_w8_l2048_id2_1 ( .CLK(CLK), .ram_w8_l2048_id2_1_0_addr(ram_w8_l2048_id2_1_0_addr), .ram_w8_l2048_id2_1_0_rdata(ram_w8_l2048_id2_1_0_rdata), .ram_w8_l2048_id2_1_0_wdata(8'h00), .ram_w8_l2048_id2_1_0_wenable(1'h0), .ram_w8_l2048_id2_1_1_addr(ram_w8_l2048_id2_1_1_addr), .ram_w8_l2048_id2_1_1_rdata(ram_w8_l2048_id2_1_1_rdata), .ram_w8_l2048_id2_1_1_wdata(ram_w8_l2048_id2_1_1_wdata), .ram_w8_l2048_id2_1_1_wenable(ram_w8_l2048_id2_1_1_wenable) );
  ram_w8_l2048_id2_2 inst_ram_w8_l2048_id2_2 ( .CLK(CLK), .ram_w8_l2048_id2_2_0_addr(ram_w8_l2048_id2_2_0_addr), .ram_w8_l2048_id2_2_0_rdata(ram_w8_l2048_id2_2_0_rdata), .ram_w8_l2048_id2_2_0_wdata(8'h00), .ram_w8_l2048_id2_2_0_wenable(1'h0), .ram_w8_l2048_id2_2_1_addr(ram_w8_l2048_id2_2_1_addr), .ram_w8_l2048_id2_2_1_rdata(ram_w8_l2048_id2_2_1_rdata), .ram_w8_l2048_id2_2_1_wdata(ram_w8_l2048_id2_2_1_wdata), .ram_w8_l2048_id2_2_1_wenable(ram_w8_l2048_id2_2_1_wenable) );
  ram_w8_l2048_id2_3 inst_ram_w8_l2048_id2_3 ( .CLK(CLK), .ram_w8_l2048_id2_3_0_addr(ram_w8_l2048_id2_3_0_addr), .ram_w8_l2048_id2_3_0_rdata(ram_w8_l2048_id2_3_0_rdata), .ram_w8_l2048_id2_3_0_wdata(8'h00), .ram_w8_l2048_id2_3_0_wenable(1'h0), .ram_w8_l2048_id2_3_1_addr(ram_w8_l2048_id2_3_1_addr), .ram_w8_l2048_id2_3_1_rdata(ram_w8_l2048_id2_3_1_rdata), .ram_w8_l2048_id2_3_1_wdata(ram_w8_l2048_id2_3_1_wdata), .ram_w8_l2048_id2_3_1_wenable(ram_w8_l2048_id2_3_1_wenable) );
  ram_w8_l2048_id3_0 inst_ram_w8_l2048_id3_0 ( .CLK(CLK), .ram_w8_l2048_id3_0_0_addr(ram_w8_l2048_id3_0_0_addr), .ram_w8_l2048_id3_0_0_rdata(ram_w8_l2048_id3_0_0_rdata), .ram_w8_l2048_id3_0_0_wdata(8'h00), .ram_w8_l2048_id3_0_0_wenable(1'h0), .ram_w8_l2048_id3_0_1_addr(ram_w8_l2048_id3_0_1_addr), .ram_w8_l2048_id3_0_1_rdata(ram_w8_l2048_id3_0_1_rdata), .ram_w8_l2048_id3_0_1_wdata(ram_w8_l2048_id3_0_1_wdata), .ram_w8_l2048_id3_0_1_wenable(ram_w8_l2048_id3_0_1_wenable) );
  ram_w8_l2048_id3_1 inst_ram_w8_l2048_id3_1 ( .CLK(CLK), .ram_w8_l2048_id3_1_0_addr(ram_w8_l2048_id3_1_0_addr), .ram_w8_l2048_id3_1_0_rdata(ram_w8_l2048_id3_1_0_rdata), .ram_w8_l2048_id3_1_0_wdata(8'h00), .ram_w8_l2048_id3_1_0_wenable(1'h0), .ram_w8_l2048_id3_1_1_addr(ram_w8_l2048_id3_1_1_addr), .ram_w8_l2048_id3_1_1_rdata(ram_w8_l2048_id3_1_1_rdata), .ram_w8_l2048_id3_1_1_wdata(ram_w8_l2048_id3_1_1_wdata), .ram_w8_l2048_id3_1_1_wenable(ram_w8_l2048_id3_1_1_wenable) );
  ram_w8_l2048_id3_2 inst_ram_w8_l2048_id3_2 ( .CLK(CLK), .ram_w8_l2048_id3_2_0_addr(ram_w8_l2048_id3_2_0_addr), .ram_w8_l2048_id3_2_0_rdata(ram_w8_l2048_id3_2_0_rdata), .ram_w8_l2048_id3_2_0_wdata(8'h00), .ram_w8_l2048_id3_2_0_wenable(1'h0), .ram_w8_l2048_id3_2_1_addr(ram_w8_l2048_id3_2_1_addr), .ram_w8_l2048_id3_2_1_rdata(ram_w8_l2048_id3_2_1_rdata), .ram_w8_l2048_id3_2_1_wdata(ram_w8_l2048_id3_2_1_wdata), .ram_w8_l2048_id3_2_1_wenable(ram_w8_l2048_id3_2_1_wenable) );
  ram_w8_l2048_id3_3 inst_ram_w8_l2048_id3_3 ( .CLK(CLK), .ram_w8_l2048_id3_3_0_addr(ram_w8_l2048_id3_3_0_addr), .ram_w8_l2048_id3_3_0_rdata(ram_w8_l2048_id3_3_0_rdata), .ram_w8_l2048_id3_3_0_wdata(8'h00), .ram_w8_l2048_id3_3_0_wenable(1'h0), .ram_w8_l2048_id3_3_1_addr(ram_w8_l2048_id3_3_1_addr), .ram_w8_l2048_id3_3_1_rdata(ram_w8_l2048_id3_3_1_rdata), .ram_w8_l2048_id3_3_1_wdata(ram_w8_l2048_id3_3_1_wdata), .ram_w8_l2048_id3_3_1_wenable(ram_w8_l2048_id3_3_1_wenable) );
  ram_w8_l2048_id4_0 inst_ram_w8_l2048_id4_0 ( .CLK(CLK), .ram_w8_l2048_id4_0_0_addr(ram_w8_l2048_id4_0_0_addr), .ram_w8_l2048_id4_0_0_rdata(ram_w8_l2048_id4_0_0_rdata), .ram_w8_l2048_id4_0_0_wdata(8'h00), .ram_w8_l2048_id4_0_0_wenable(1'h0), .ram_w8_l2048_id4_0_1_addr(ram_w8_l2048_id4_0_1_addr), .ram_w8_l2048_id4_0_1_rdata(ram_w8_l2048_id4_0_1_rdata), .ram_w8_l2048_id4_0_1_wdata(ram_w8_l2048_id4_0_1_wdata), .ram_w8_l2048_id4_0_1_wenable(ram_w8_l2048_id4_0_1_wenable) );
  ram_w8_l2048_id4_1 inst_ram_w8_l2048_id4_1 ( .CLK(CLK), .ram_w8_l2048_id4_1_0_addr(ram_w8_l2048_id4_1_0_addr), .ram_w8_l2048_id4_1_0_rdata(ram_w8_l2048_id4_1_0_rdata), .ram_w8_l2048_id4_1_0_wdata(8'h00), .ram_w8_l2048_id4_1_0_wenable(1'h0), .ram_w8_l2048_id4_1_1_addr(ram_w8_l2048_id4_1_1_addr), .ram_w8_l2048_id4_1_1_rdata(ram_w8_l2048_id4_1_1_rdata), .ram_w8_l2048_id4_1_1_wdata(ram_w8_l2048_id4_1_1_wdata), .ram_w8_l2048_id4_1_1_wenable(ram_w8_l2048_id4_1_1_wenable) );
  ram_w8_l2048_id4_2 inst_ram_w8_l2048_id4_2 ( .CLK(CLK), .ram_w8_l2048_id4_2_0_addr(ram_w8_l2048_id4_2_0_addr), .ram_w8_l2048_id4_2_0_rdata(ram_w8_l2048_id4_2_0_rdata), .ram_w8_l2048_id4_2_0_wdata(8'h00), .ram_w8_l2048_id4_2_0_wenable(1'h0), .ram_w8_l2048_id4_2_1_addr(ram_w8_l2048_id4_2_1_addr), .ram_w8_l2048_id4_2_1_rdata(ram_w8_l2048_id4_2_1_rdata), .ram_w8_l2048_id4_2_1_wdata(ram_w8_l2048_id4_2_1_wdata), .ram_w8_l2048_id4_2_1_wenable(ram_w8_l2048_id4_2_1_wenable) );
  ram_w8_l2048_id4_3 inst_ram_w8_l2048_id4_3 ( .CLK(CLK), .ram_w8_l2048_id4_3_0_addr(ram_w8_l2048_id4_3_0_addr), .ram_w8_l2048_id4_3_0_rdata(ram_w8_l2048_id4_3_0_rdata), .ram_w8_l2048_id4_3_0_wdata(8'h00), .ram_w8_l2048_id4_3_0_wenable(1'h0), .ram_w8_l2048_id4_3_1_addr(ram_w8_l2048_id4_3_1_addr), .ram_w8_l2048_id4_3_1_rdata(ram_w8_l2048_id4_3_1_rdata), .ram_w8_l2048_id4_3_1_wdata(ram_w8_l2048_id4_3_1_wdata), .ram_w8_l2048_id4_3_1_wenable(ram_w8_l2048_id4_3_1_wenable) );
  ram_w8_l2048_id5_0 inst_ram_w8_l2048_id5_0 ( .CLK(CLK), .ram_w8_l2048_id5_0_0_addr(ram_w8_l2048_id5_0_0_addr), .ram_w8_l2048_id5_0_0_rdata(ram_w8_l2048_id5_0_0_rdata), .ram_w8_l2048_id5_0_0_wdata(8'h00), .ram_w8_l2048_id5_0_0_wenable(1'h0), .ram_w8_l2048_id5_0_1_addr(ram_w8_l2048_id5_0_1_addr), .ram_w8_l2048_id5_0_1_rdata(ram_w8_l2048_id5_0_1_rdata), .ram_w8_l2048_id5_0_1_wdata(ram_w8_l2048_id5_0_1_wdata), .ram_w8_l2048_id5_0_1_wenable(ram_w8_l2048_id5_0_1_wenable) );
  ram_w8_l2048_id5_1 inst_ram_w8_l2048_id5_1 ( .CLK(CLK), .ram_w8_l2048_id5_1_0_addr(ram_w8_l2048_id5_1_0_addr), .ram_w8_l2048_id5_1_0_rdata(ram_w8_l2048_id5_1_0_rdata), .ram_w8_l2048_id5_1_0_wdata(8'h00), .ram_w8_l2048_id5_1_0_wenable(1'h0), .ram_w8_l2048_id5_1_1_addr(ram_w8_l2048_id5_1_1_addr), .ram_w8_l2048_id5_1_1_rdata(ram_w8_l2048_id5_1_1_rdata), .ram_w8_l2048_id5_1_1_wdata(ram_w8_l2048_id5_1_1_wdata), .ram_w8_l2048_id5_1_1_wenable(ram_w8_l2048_id5_1_1_wenable) );
  ram_w8_l2048_id5_2 inst_ram_w8_l2048_id5_2 ( .CLK(CLK), .ram_w8_l2048_id5_2_0_addr(ram_w8_l2048_id5_2_0_addr), .ram_w8_l2048_id5_2_0_rdata(ram_w8_l2048_id5_2_0_rdata), .ram_w8_l2048_id5_2_0_wdata(8'h00), .ram_w8_l2048_id5_2_0_wenable(1'h0), .ram_w8_l2048_id5_2_1_addr(ram_w8_l2048_id5_2_1_addr), .ram_w8_l2048_id5_2_1_rdata(ram_w8_l2048_id5_2_1_rdata), .ram_w8_l2048_id5_2_1_wdata(ram_w8_l2048_id5_2_1_wdata), .ram_w8_l2048_id5_2_1_wenable(ram_w8_l2048_id5_2_1_wenable) );
  ram_w8_l2048_id5_3 inst_ram_w8_l2048_id5_3 ( .CLK(CLK), .ram_w8_l2048_id5_3_0_addr(ram_w8_l2048_id5_3_0_addr), .ram_w8_l2048_id5_3_0_rdata(ram_w8_l2048_id5_3_0_rdata), .ram_w8_l2048_id5_3_0_wdata(8'h00), .ram_w8_l2048_id5_3_0_wenable(1'h0), .ram_w8_l2048_id5_3_1_addr(ram_w8_l2048_id5_3_1_addr), .ram_w8_l2048_id5_3_1_rdata(ram_w8_l2048_id5_3_1_rdata), .ram_w8_l2048_id5_3_1_wdata(ram_w8_l2048_id5_3_1_wdata), .ram_w8_l2048_id5_3_1_wenable(ram_w8_l2048_id5_3_1_wenable) );
  ram_w8_l2048_id6_0 inst_ram_w8_l2048_id6_0 ( .CLK(CLK), .ram_w8_l2048_id6_0_0_addr(ram_w8_l2048_id6_0_0_addr), .ram_w8_l2048_id6_0_0_rdata(ram_w8_l2048_id6_0_0_rdata), .ram_w8_l2048_id6_0_0_wdata(8'h00), .ram_w8_l2048_id6_0_0_wenable(1'h0), .ram_w8_l2048_id6_0_1_addr(ram_w8_l2048_id6_0_1_addr), .ram_w8_l2048_id6_0_1_rdata(ram_w8_l2048_id6_0_1_rdata), .ram_w8_l2048_id6_0_1_wdata(ram_w8_l2048_id6_0_1_wdata), .ram_w8_l2048_id6_0_1_wenable(ram_w8_l2048_id6_0_1_wenable) );
  ram_w8_l2048_id6_1 inst_ram_w8_l2048_id6_1 ( .CLK(CLK), .ram_w8_l2048_id6_1_0_addr(ram_w8_l2048_id6_1_0_addr), .ram_w8_l2048_id6_1_0_rdata(ram_w8_l2048_id6_1_0_rdata), .ram_w8_l2048_id6_1_0_wdata(8'h00), .ram_w8_l2048_id6_1_0_wenable(1'h0), .ram_w8_l2048_id6_1_1_addr(ram_w8_l2048_id6_1_1_addr), .ram_w8_l2048_id6_1_1_rdata(ram_w8_l2048_id6_1_1_rdata), .ram_w8_l2048_id6_1_1_wdata(ram_w8_l2048_id6_1_1_wdata), .ram_w8_l2048_id6_1_1_wenable(ram_w8_l2048_id6_1_1_wenable) );
  ram_w8_l2048_id6_2 inst_ram_w8_l2048_id6_2 ( .CLK(CLK), .ram_w8_l2048_id6_2_0_addr(ram_w8_l2048_id6_2_0_addr), .ram_w8_l2048_id6_2_0_rdata(ram_w8_l2048_id6_2_0_rdata), .ram_w8_l2048_id6_2_0_wdata(8'h00), .ram_w8_l2048_id6_2_0_wenable(1'h0), .ram_w8_l2048_id6_2_1_addr(ram_w8_l2048_id6_2_1_addr), .ram_w8_l2048_id6_2_1_rdata(ram_w8_l2048_id6_2_1_rdata), .ram_w8_l2048_id6_2_1_wdata(ram_w8_l2048_id6_2_1_wdata), .ram_w8_l2048_id6_2_1_wenable(ram_w8_l2048_id6_2_1_wenable) );
  ram_w8_l2048_id6_3 inst_ram_w8_l2048_id6_3 ( .CLK(CLK), .ram_w8_l2048_id6_3_0_addr(ram_w8_l2048_id6_3_0_addr), .ram_w8_l2048_id6_3_0_rdata(ram_w8_l2048_id6_3_0_rdata), .ram_w8_l2048_id6_3_0_wdata(8'h00), .ram_w8_l2048_id6_3_0_wenable(1'h0), .ram_w8_l2048_id6_3_1_addr(ram_w8_l2048_id6_3_1_addr), .ram_w8_l2048_id6_3_1_rdata(ram_w8_l2048_id6_3_1_rdata), .ram_w8_l2048_id6_3_1_wdata(ram_w8_l2048_id6_3_1_wdata), .ram_w8_l2048_id6_3_1_wenable(ram_w8_l2048_id6_3_1_wenable) );
  ram_w8_l2048_id7_0 inst_ram_w8_l2048_id7_0 ( .CLK(CLK), .ram_w8_l2048_id7_0_0_addr(ram_w8_l2048_id7_0_0_addr), .ram_w8_l2048_id7_0_0_rdata(ram_w8_l2048_id7_0_0_rdata), .ram_w8_l2048_id7_0_0_wdata(8'h00), .ram_w8_l2048_id7_0_0_wenable(1'h0), .ram_w8_l2048_id7_0_1_addr(ram_w8_l2048_id7_0_1_addr), .ram_w8_l2048_id7_0_1_rdata(ram_w8_l2048_id7_0_1_rdata), .ram_w8_l2048_id7_0_1_wdata(ram_w8_l2048_id7_0_1_wdata), .ram_w8_l2048_id7_0_1_wenable(ram_w8_l2048_id7_0_1_wenable) );
  ram_w8_l2048_id7_1 inst_ram_w8_l2048_id7_1 ( .CLK(CLK), .ram_w8_l2048_id7_1_0_addr(ram_w8_l2048_id7_1_0_addr), .ram_w8_l2048_id7_1_0_rdata(ram_w8_l2048_id7_1_0_rdata), .ram_w8_l2048_id7_1_0_wdata(8'h00), .ram_w8_l2048_id7_1_0_wenable(1'h0), .ram_w8_l2048_id7_1_1_addr(ram_w8_l2048_id7_1_1_addr), .ram_w8_l2048_id7_1_1_rdata(ram_w8_l2048_id7_1_1_rdata), .ram_w8_l2048_id7_1_1_wdata(ram_w8_l2048_id7_1_1_wdata), .ram_w8_l2048_id7_1_1_wenable(ram_w8_l2048_id7_1_1_wenable) );
  ram_w8_l2048_id7_2 inst_ram_w8_l2048_id7_2 ( .CLK(CLK), .ram_w8_l2048_id7_2_0_addr(ram_w8_l2048_id7_2_0_addr), .ram_w8_l2048_id7_2_0_rdata(ram_w8_l2048_id7_2_0_rdata), .ram_w8_l2048_id7_2_0_wdata(8'h00), .ram_w8_l2048_id7_2_0_wenable(1'h0), .ram_w8_l2048_id7_2_1_addr(ram_w8_l2048_id7_2_1_addr), .ram_w8_l2048_id7_2_1_rdata(ram_w8_l2048_id7_2_1_rdata), .ram_w8_l2048_id7_2_1_wdata(ram_w8_l2048_id7_2_1_wdata), .ram_w8_l2048_id7_2_1_wenable(ram_w8_l2048_id7_2_1_wenable) );
  ram_w8_l2048_id7_3 inst_ram_w8_l2048_id7_3 ( .CLK(CLK), .ram_w8_l2048_id7_3_0_addr(ram_w8_l2048_id7_3_0_addr), .ram_w8_l2048_id7_3_0_rdata(ram_w8_l2048_id7_3_0_rdata), .ram_w8_l2048_id7_3_0_wdata(8'h00), .ram_w8_l2048_id7_3_0_wenable(1'h0), .ram_w8_l2048_id7_3_1_addr(ram_w8_l2048_id7_3_1_addr), .ram_w8_l2048_id7_3_1_rdata(ram_w8_l2048_id7_3_1_rdata), .ram_w8_l2048_id7_3_1_wdata(ram_w8_l2048_id7_3_1_wdata), .ram_w8_l2048_id7_3_1_wenable(ram_w8_l2048_id7_3_1_wenable) );
  ram_w8_l2048_id8_0 inst_ram_w8_l2048_id8_0 ( .CLK(CLK), .ram_w8_l2048_id8_0_0_addr(ram_w8_l2048_id8_0_0_addr), .ram_w8_l2048_id8_0_0_rdata(ram_w8_l2048_id8_0_0_rdata), .ram_w8_l2048_id8_0_0_wdata(8'h00), .ram_w8_l2048_id8_0_0_wenable(1'h0), .ram_w8_l2048_id8_0_1_addr(ram_w8_l2048_id8_0_1_addr), .ram_w8_l2048_id8_0_1_rdata(ram_w8_l2048_id8_0_1_rdata), .ram_w8_l2048_id8_0_1_wdata(ram_w8_l2048_id8_0_1_wdata), .ram_w8_l2048_id8_0_1_wenable(ram_w8_l2048_id8_0_1_wenable) );
  ram_w8_l2048_id8_1 inst_ram_w8_l2048_id8_1 ( .CLK(CLK), .ram_w8_l2048_id8_1_0_addr(ram_w8_l2048_id8_1_0_addr), .ram_w8_l2048_id8_1_0_rdata(ram_w8_l2048_id8_1_0_rdata), .ram_w8_l2048_id8_1_0_wdata(8'h00), .ram_w8_l2048_id8_1_0_wenable(1'h0), .ram_w8_l2048_id8_1_1_addr(ram_w8_l2048_id8_1_1_addr), .ram_w8_l2048_id8_1_1_rdata(ram_w8_l2048_id8_1_1_rdata), .ram_w8_l2048_id8_1_1_wdata(ram_w8_l2048_id8_1_1_wdata), .ram_w8_l2048_id8_1_1_wenable(ram_w8_l2048_id8_1_1_wenable) );
  ram_w8_l2048_id8_2 inst_ram_w8_l2048_id8_2 ( .CLK(CLK), .ram_w8_l2048_id8_2_0_addr(ram_w8_l2048_id8_2_0_addr), .ram_w8_l2048_id8_2_0_rdata(ram_w8_l2048_id8_2_0_rdata), .ram_w8_l2048_id8_2_0_wdata(8'h00), .ram_w8_l2048_id8_2_0_wenable(1'h0), .ram_w8_l2048_id8_2_1_addr(ram_w8_l2048_id8_2_1_addr), .ram_w8_l2048_id8_2_1_rdata(ram_w8_l2048_id8_2_1_rdata), .ram_w8_l2048_id8_2_1_wdata(ram_w8_l2048_id8_2_1_wdata), .ram_w8_l2048_id8_2_1_wenable(ram_w8_l2048_id8_2_1_wenable) );
  ram_w8_l2048_id8_3 inst_ram_w8_l2048_id8_3 ( .CLK(CLK), .ram_w8_l2048_id8_3_0_addr(ram_w8_l2048_id8_3_0_addr), .ram_w8_l2048_id8_3_0_rdata(ram_w8_l2048_id8_3_0_rdata), .ram_w8_l2048_id8_3_0_wdata(8'h00), .ram_w8_l2048_id8_3_0_wenable(1'h0), .ram_w8_l2048_id8_3_1_addr(ram_w8_l2048_id8_3_1_addr), .ram_w8_l2048_id8_3_1_rdata(ram_w8_l2048_id8_3_1_rdata), .ram_w8_l2048_id8_3_1_wdata(ram_w8_l2048_id8_3_1_wdata), .ram_w8_l2048_id8_3_1_wenable(ram_w8_l2048_id8_3_1_wenable) );
  ram_w8_l2048_id9_0 inst_ram_w8_l2048_id9_0 ( .CLK(CLK), .ram_w8_l2048_id9_0_0_addr(ram_w8_l2048_id9_0_0_addr), .ram_w8_l2048_id9_0_0_rdata(ram_w8_l2048_id9_0_0_rdata), .ram_w8_l2048_id9_0_0_wdata(8'h00), .ram_w8_l2048_id9_0_0_wenable(1'h0), .ram_w8_l2048_id9_0_1_addr(ram_w8_l2048_id9_0_1_addr), .ram_w8_l2048_id9_0_1_rdata(ram_w8_l2048_id9_0_1_rdata), .ram_w8_l2048_id9_0_1_wdata(ram_w8_l2048_id9_0_1_wdata), .ram_w8_l2048_id9_0_1_wenable(ram_w8_l2048_id9_0_1_wenable) );
  ram_w8_l2048_id9_1 inst_ram_w8_l2048_id9_1 ( .CLK(CLK), .ram_w8_l2048_id9_1_0_addr(ram_w8_l2048_id9_1_0_addr), .ram_w8_l2048_id9_1_0_rdata(ram_w8_l2048_id9_1_0_rdata), .ram_w8_l2048_id9_1_0_wdata(8'h00), .ram_w8_l2048_id9_1_0_wenable(1'h0), .ram_w8_l2048_id9_1_1_addr(ram_w8_l2048_id9_1_1_addr), .ram_w8_l2048_id9_1_1_rdata(ram_w8_l2048_id9_1_1_rdata), .ram_w8_l2048_id9_1_1_wdata(ram_w8_l2048_id9_1_1_wdata), .ram_w8_l2048_id9_1_1_wenable(ram_w8_l2048_id9_1_1_wenable) );
  ram_w8_l2048_id9_2 inst_ram_w8_l2048_id9_2 ( .CLK(CLK), .ram_w8_l2048_id9_2_0_addr(ram_w8_l2048_id9_2_0_addr), .ram_w8_l2048_id9_2_0_rdata(ram_w8_l2048_id9_2_0_rdata), .ram_w8_l2048_id9_2_0_wdata(8'h00), .ram_w8_l2048_id9_2_0_wenable(1'h0), .ram_w8_l2048_id9_2_1_addr(ram_w8_l2048_id9_2_1_addr), .ram_w8_l2048_id9_2_1_rdata(ram_w8_l2048_id9_2_1_rdata), .ram_w8_l2048_id9_2_1_wdata(ram_w8_l2048_id9_2_1_wdata), .ram_w8_l2048_id9_2_1_wenable(ram_w8_l2048_id9_2_1_wenable) );
  ram_w8_l2048_id9_3 inst_ram_w8_l2048_id9_3 ( .CLK(CLK), .ram_w8_l2048_id9_3_0_addr(ram_w8_l2048_id9_3_0_addr), .ram_w8_l2048_id9_3_0_rdata(ram_w8_l2048_id9_3_0_rdata), .ram_w8_l2048_id9_3_0_wdata(8'h00), .ram_w8_l2048_id9_3_0_wenable(1'h0), .ram_w8_l2048_id9_3_1_addr(ram_w8_l2048_id9_3_1_addr), .ram_w8_l2048_id9_3_1_rdata(ram_w8_l2048_id9_3_1_rdata), .ram_w8_l2048_id9_3_1_wdata(ram_w8_l2048_id9_3_1_wdata), .ram_w8_l2048_id9_3_1_wenable(ram_w8_l2048_id9_3_1_wenable) );
endmodule
